BZh91AY&SYJX2�?_�px����������ai� �Q�2U� �y"��   �h    �   P   ���J@ ��   �   AB� @Q!))T )@�   P (
 U.   m�:��( P��`���r޲�&�#vr� Ό]:so6w���� t��ׇ��� ���� X ҨY`(b i� D�*�
0Ц!�S�t8�����*�(   ,:��(   �1�R��F6WӖ���m=5��]7�VM{5ŕV=β�� Ҭ���}㺞��=:���/x ����-ͧ�9k�K�S�x� ��_mn;��;����Ԯ�]Q{��� �@ ,` o}J��w���;��Ū{o�n�\ ��n�J�;�Vm*�5�n�+ޥ7n�W_ twW��˕U��:�d�e\��rj�wx��� �yS�]*�W�^ZWN]R��ϐ) �JP PP� �>����^��}�x�]�st�` 'Qc�*sj�q�9��]. ���y����u�i�  ����\��� �S�6ꛟ{�K���}�'�J� 'Jd�ŏ^�ON����O�z�( PP P�(� :>�K�2���^#ݫ��[n k��J��4��ʼ=�^R� �����|����  �9omz�}�W� /g���6�{���oZy=;���m7 �=Jǻ���f�iɡY5/x          �S�&)�*J�4 ��a14"��h��U)       E?���04� #&F� 4i����U*�&��     ?BI���J4�0��L�0��F�@)�	��1Ojh���4zh�)�'Ꟁ����߿���]?����}]{���������7�QU� �*��U�H�����U��((��`�(�������P�(����/�� J�rj�?������'󾏧����17���11�3�LL��1��LLL�8���1���q���A���$ę��.1111�LI���c9�`�Øa�Xi�ΌLL���1��bc�&$Ġ�	���8���Ę�����2��i��h�N1[�112�q�8�q����8�11�L�p��3���=��Za���_!`����&1�Lg�c8�7ah��,Zi�9�
�D�4�0�F&1�Lc�1�c���&7bc�M4�Ni�H�)�D��11������}}?H���Y��z�OXee4��(:สD�D�����YWmSJ"AR�WJ��+j��T�˺���"+�ҡ$v�_{\p卪�����H�*�WQSvժA��Ծ']�R��@�Ҋ�vR*��O�*��+O�+����U$gh���C�-��P�3�Ra�S���5s���Z6��S�v��죩8U'EH�].�*u��,u�D���r��}���Y����ev/�8�N��t�K�V40A�'#(Ƭ�3�H�BP�hc
�d��LLؔ�塋!(p2t�.9	��IƘX(XyO\�,��(MC�����[�1�t��Z�L`he_�W�\���s����}�o�[�"����z�8�`Pf�2�A�a�����}��|·2	�A՜w������5a�e�y�{�ٲ;9.9�2vrLp�q5	[#�f���L��T�	K�F�Ӭɚpw���"u��*����e�E3�����.QIC����˷��L�yćz��A�kF�����ĖP�I�F�4D�FF8�o�E��Vu.�>�\aC��T��n�n8����F��}�u������|g%_)���R�"��;����f{����ov�y�<޻;�����=��n�\�d��9z��tF�k'4�A�4%b8�Y�sZl��M��Z�utu����t��LZ�͐��h3`�M�:\���s��ѐa�%�
�cѢt�5DV;�F�޷��7���he�X�f���,�������a���)$%�l5hĞkD8%`��%b�F:e��d%	��B��&!P�a����8霒58kS�{��5BV�%�t�A�P��L���`h��M�Da5I$b�a)6k5Kp'*�3v"��ܨ���EA(fL�߽�`��U3|��,���w~K�W�
��#�R��Y��.��r���f�ՠ3pd��8�k�]��t!!�=��:S�-�����~g�t.t~K��ʠ���r�[�v�%�v:��]��e,�{;-I�gtyٺ!�8N�%X���1d.>�J���J\J$K�O�����O��m��%���!T����s��uw�P�3�>��Z�K�����V�r�������o�rt�k����y�s��ݼ	�ڥ�v�}��{�,����8T�QH�&�'L����3CM��,f�d�FI�e�t1p'IBQ�C��S.9.�B=�t�&&P0$Д%&40c�i0J�Врd%.<��3,C�f�r�N.N����I�Ը�2�I�X:��.BrM%m�Q�3I�����Q�M&���'�98��11M�g ��dK 4d�w�Nf���d`l5	F:n�㐖B{�p0r�#c�P�:���49.9h6��s�(JLMF��BTI��	N����dv��t�����rFKP��Cm15���q�@P��r0xk1�%�A�L�Ʌ&�Z�̝.N�X�`勣R�2�:�2��:\%Ɲ.lp3:+����(O3C���S��12C2M�`�`�A��L��պݖ�ZM�53g �ѵ�8�(0�j\u��`K�c	��A��hZ���<��ġ�Vtp#�1��A��:6n5�0���0�1Ջ8�3Q��K�$�8&f8�P����F��1ӣa�a�n�X�T��:��j0Д�c�e��Z���t!�X�����N͑��I(��ka����g 0�9�Zݎ�����mkIV-����ճ!.V�'Z�2̝Nd�`�Li�5�K��wz��w�����x莧7���p�'pc�fN3�\8x�r�35�����q����6�]����T�NRh�yIݭ����ê��'y�x�kBzf#�I5ì�s4Q���>��[�R����~tv��FǇ�㘘�����0�5:6k��,&�����l��1�m����0(Ѿtgzv�g{S�HUC+�Q7m�U>U�L<�f�,H2ă'$�Ýw�4o8��֟mԘǚ���Z�.�zM1��2��N��������C��KPl���2p���	�w��;��a�f	Į��ȝ���E�:�@���v��k ɨ�2C2g�����ѽ<z��$��G�kXYgeZ�C��Ө�֥��BX�K��nu:\�hJP�����٬�83�V!�!�%X�	LI������(0y�`���=w�!͉Bu	F��a�.d%	��Ӑ�%	BH�@Kz�7	J�z٣:����(J`(O3�\��,\J�k���������a���s~k~FZ��\���Z�p���[5�4A��y���1���	O�:�u�Q�9%�ߘz��OM�:8��4�0ٚ�����:�r0�\�����6l����Ƃ�.h6�Z�����]s�GRi2C2!)d�7�o�<c7�uٳ���sN�21l���WGY���[��[�f�j3Vh-�N��������2E8�I�L��%��<��	��Ԓu��$ZC��7�A��5	�:	�\��' 6u	�KBw�������	G���ݷ�����CߒP��>.`mǻ��5&�(a�6@h�C26�u�	�6>��'pG�p;������:ֶq{�	N�؝BrC�X<��v�����i��X�g��Gq��0�l:�۝$w�%�0-N:a��{�78i9���/�F�`�=�O61���f��n8��h'�e���Y����IZ���\wWIO"}\�P���e_(��8j��3t�nrċZM\w�l��{ѣda�l�є�9a�b�Hd��)�4ƒ���b�`�%!�!��C�bY������.KE8�	X2	����(JLL�\��(J"��@dc�I�8I���d8�e���%C����a%���@1f]&�$a)�
��t��f	BQ���&�5	I,�uK@Le$��H�89N|󽡒���4��BX:�4c�t�`Bo1�8l�N��"�%	K�!(0r'�K�#`d8��2�\ \�`�&@a���V!�������L�i�N�1�:ؔ<��J������Q���b����ti��CӨ5[0�:ބ�L�Q��4j"���������F�8�4m#5ӳul ��$���0Ѭ�*p3E��Z{���t�o��f�4s7!��j�DД�;�Q��8q{�a��4����f:s}��E�5�u�*#Zc5�0����6xf6Xt�gfa�kHe��(�2��::�&�ӹ�=����n�͜�a�a��7�᎓PoO-�6d�������\�I��L�:�ِ�2\r0 �X�r0�pڊ��ӥT���]QlT�9uLI�O}�5䛵��]D�I$.��2\r���# �4ề�)�X�����XN:6s<�|Ѿ��9G;����0�1�'�t���Ġ0��8BV!�����'N�Pt�Ոd`N�:\�aí����̵�]v�I�Lh6p5�Zp6W{ �A�o^=�����Z-����,Og���# �KI�Ȑ�5h �S�Ө{u����GF��Z� ��I�1[C0�[3���p6p���f��;��m�k�����.�~����7�JLjqr@�G[�WV�<ނ޶o��f�0�y��1#�-9��sM�̌1��0�uhN�	N0d`A��lf��#7���u6Zv���2՚�:�o|N�V���8f���5;F��
��LB�I��Bhu���U�f�0vJe
I��`��Np�h�tj�яzݣ	&04j4A�sfkz���tbqi!�,{|ѳpa�$�HŏK޳N�SDc9BV�vѳ^w��u�u��2�u8�27!���і�N�$$�I�V�L�ͺ�4i%�`��K�����3%�c���9�^9�:�5�%0M!���)��c!�3���bh���˿F�2ќ뽇$�{��^uθw����Hd��L�w�{���J����9u��w|\�[�x�f�5�]wێ�X�;u���v�>����W�;ϲ�*>5Mҡ��$/h�n<�n4��*U�n@��ԃ�.;��s.��� g��m۫) �l*S��⮂�j�r�')�I�B��~��it좚��0t�q��q�:MV+����N&s�U�:�~������=��Z��$�I$�� )@A��P805l  �ro.����f���yi�5!D75��m�Aں�gMņ�ӫ�Wf|���n�+u��;^�t�-�vx�l�t'Eܕ�lH'��s:�j��J�IN��-ΖUt;h�+�d���ͅ�^��[y�  m[ ��6�6  Im 2D�m���p   [@ m�v�M��  	    �Ѷ� 8p��`6�   Gꇠ    � n�� ����m@[@ �J v�m�h"@ �ZlH Ԁ   H	  �6�k[@86��M�`�m�m��     $��p��qm6ٶ�8ʶ�   I�  m��4�l�Z��A���v�x�9݋Y~��NKE�ڶ  ��e�Ml	Cm� -���  [%��HޫI6ԅ���-�mm�a � ���[\նޭ�� m�@ �-� � ���` v�lp ���) I�*@�c[�[��&�  �� � m  ���A%�$m� ��vn�i�m��]��*p� ��[m��H�@#�lm��mp ��ܓ�n���mհ��|ds�e [D��-�mjG [@   � h� �@		   �� Hl 8��v apm�  [���ؐ��}zh � �r@[vؓm�h 8�B����m� ְ�J.�� ���u�e� 9�m�N-��h [@��i"۝l�     m �c�    h �� H��kn  N�  ����[F�	�� l�f�q�i���$    l�(!�� [m�	h� � m��[@9���mÁ��-�l[V�X�K'J�:��N���Ͷ�$l �6�   �mm�  �i�	�-� E  � �$  � �������m6�����UEP(��bq$k��m��-��M����lHz����� m���h��TQҭV�O+@HMt�5آ�XH�V��*�U@R�+�#�E�G���r������f��m ��˵�t�.�.ۘ�����j� 5��$�7F��Ͷ��   �d�i �`��  �i� $m�U�F�  +Yx��^۞����Ic�nV�UV�]1���vP��wb:�1E� 2=v�f�j���QʛK���
^kh
��e���[:7�H�$����	m�����f��J���([\ m� ����� �|���{O6�� -��p 9��0m����֎,��� �H川 �j��`m ��WU[RnQ�5 �v 	zP����Hp $��   ���n�l 0�$p-�Xש�:��s����n�^�@ ��  � ��� �   p� ���l�L���m�����H   �l-��a��   6�;l�G8��pb��m�O���$6��m&����V�� �%�@�%�;`[@ �m���p@  ��Ҥ��$	  I�� �l��m� ��-��H8z{o�m��  �   �` �p m  9���m�m� -�l۶���p[@   -��h8�g6ͤ�U�Wʁ�2�U*�rC�H�  m�hlH �趶ۍ�� 	 mÜ   �t��[g@ �.�-�e�$[M�8�`6�p�Yѻi) Im&� �r@�-�&K��`�]��v����v����B�J�U�=�Јj`ճ{���a�l_}�t���6�T
��{F�A��u�#�h��À܂��v�8]�v)� 
��r�l@J�K��ͷd���mNT��� �8l�ڐ [Wl�G[yj��ZA%�[B��M��[M�p -��;� p��m&��ܬ9bʯ0msmGe%m� �m-�m�Ƶ�  ඉ
P�m�`  �=����-���v*��S�(�Z�h( ll�   ���   �Ͷ k�6�'$  l�4P$6�/Z�   -�[@qi��J��]�s:�����v-���  ��H    H�� ��hl��[�� ��l6�ڶ�  -������� ��� �����f���Z�[���U��b�U��yKNkt 	 � 6[���� ��m   H     ��m-��   88   ���`�  �Ԁ6ضJ	  im  8-� �    l �� p h���spX�n�V6ī��J�VSj�l�=`櫫�]�g�և8[%��� V�m� �	��L6�"@-�m  ��=��]� m� �� �Sb�0Z��sm� ��l` :ْە�t�WX�����T�6��h 	m� m�m� m�֕&���fٶ�%�H 	uT2��UyyCf؇k���
�U*�U��qC+ڶ�v��vi�c���M��ImI��. ,��q%��[!U��r��m<����C	i���q�T9�y�f����,n%v"��U��U��m$ l���k���9@��̶��` ���h�vb����A{m&D� �  -[@�`(jׯ����Z������γP ��m�3�8HڢP�����p@K�A�*�^P�h ٵlp$m�r1e��@*�Us� [UK�Ĥ�Щ�� 	�m����i�0p$ �m[%��ju l S^%���l�l����E�M��,�֛lM�	 =����� �d� ź�p���l5�!l�,['�t�6ؐ�� H -��L���Jm�� m�f�m��-�����p7UuU@.(J�у�mz  @     ڳM�
�UU@�Xv�>-%��[m� r&�Cm� i-��d�J Z�m���.^�� m[@  6����A͔�`K$�[&�9��8m���i1;UH	ҭ@$  m�$�	�   �6� 6�m�  6���   �  8� m �  	 �m�H 8l��#�@8  ���l �#]���M�m�|m����e�K�d�� �d�l�8 ��Ě��m  �c8�v�g� �P�n�$m��e��q*�6��v�0m��q mۤ� 6�mr� m��  p6�6ض�I��$I7n�K��m��פ͆� !oP� 6�m�   �@�A��l� h  m��c� ��$6��6�B@ ���m�   �m  hА    ۰p���  �hH �m��� -� m��VŴ �8�� �Á:$/6�  @ 6ض�"Kn�����o$�lS uS�����m��rY@8kmٕ����n�P�<��6�y���"��HG=��մm�m    9��  ��p    �b� � -��H�p ��ށm -� -�۶�	�i �H �`��8 6��@ -�   8�h  ��mm�0ٶl` m&�t�bI�p �ٺi�"�*Kh�a�Xq��줜�*�Uҭ���[&k��!m ��[@��   [A�H@  6�I��  � H��pB@[@����� H ��m$H�mR��UU����@� t�o��Sn�:t����eu����@ �{o�m��w��p>�m��m�  $���q"��� �`�e�M�'[\�6vZ�#j�&  K)im� ��@ @  -�� �%�&�9�  +a��kZ)�j�(�T��2t�F��F�p8G7[$[(�5�1tF�Noh�,�v �:��᷾�E�4po%�CǄ�$���]�3�wh$���KI�_�QE��8�*��؂��~� �����v��"���I(&�ぐf��d�S��Da��a��"bC�t�#��㳰8$�A���ꢪ���*��������������*��������B��D*��J������������~O��z@��?���t+��;�����*UWB�zjOب^b 2<^��PM�L� �ب�tG��_bUڈ.�q1P��������Dl OPC�C^����
=zz��v���t#����B)�qC���. "c &�L<^��x0���/�,����Hc���b����e�6&��X=v�&m;I���8���x���UN�@��(����pD`�����Xv� JJA}W�a�HAOW���m� i<4q!�T��*����Q�` ��u7��
�	���dR�*���P�&�SAG�wঁ8���d��V;P!�@uЯ�A�#ӱ#�����U�^U�^U�^PW�yW�yW�y�yW�yW�yW�yW�yݷm�vݷm�^wm�{+��^UU�_����������y��������ϩ�>���w����|�&�kd��w� �?��I(����ŷ�Y��_�O�'+�W-+��ӄ�bv���N��;U/ uߞy�7|�� �NW�m��Lh5�g��gi�Mr7glԫ�
��걻����Z���KZ�F�r�8.۷k0���+�E]�vst&S��׾�||ogZ�m��9:uN;&WBq�O�mu�n�v�*�� 3��,BM�)���(lYvϱ�ܝ.Z��Ivꫫ��!dUT��]��
is��D���	-���݄��([b�' �\���Y5Ƈ%\:E����yu��\E�ƫ�e�A���T�-͐ 1��+r��ѱ\��I�K��L�=qՌ���-X�:0�vU�v��i����:���غ��k��fU۱F�����mgWl�kr-��tӫF��Iy��e�u݂mzEXئ6*�.�B��e�n7�Tݣ����%����z�; +/0UtqUm�M��nt�4�d^Tܝ�-%��)6 6j�獩ʹ�V�hN��XCpU�[n���Lhz��ۖ���Uɲ��m������bɩ�[�9���XP%%Nd;�e3�RT�m�[e�N�Xm$��b��m��m8���|�[\lZKS���nD�RZڶ���W���$΅V�Ďup�4PS�*���X�.�m���T�r=e��9�u;r���ݦ��U��f;����X�kQ�;v�nۋ'�=vm��@�ѹU�jD��]$]�<�Rt�2�Z��N��5�J��p"����MR�X7$D�Kk��$t��2�(�Umm��a�v�SG�Kr
�˶7c����ʒgi��;b�6A��z�(��=���c�[�K��kj^�W
RJK��G�D��(`�L�IR�H|�F��y���-�X8
Q{ �ǀ���>�I��!5.\�&����[�)<a��\7j��rf�dz�C�.�v4��y^Y�6�v�q2���4ϩ�3nd��gp�d�^�i�h��$�Y5�߻�.u�6ٔܗl;"14�:Cb���%��}p��MEJ8�6��R�7��������3}����}�(<^����O�< H}��@�E�pQ�h�K�df��W0�� ݴh��:��u�zѮ���qą��`&vdiȸ�ݷ,&
��޶%�2�~>���-�ö��V��[���3[��ϋ��E�w;	z�(�z��Y�k%*�l�=f;-b�h�;L���oi#rBh�k��`ۇ;L$�ص�S-��մ�<��H��`�%�vu��[r���u�Om�;v��;��w{��s���\��ԛN�T:n�i�/*�vrq��Ǳ�`��9^ANw�p2������q�D�e�����%ˀy�qڀC�KY�6�Li�Q�X/{�9I�6Xy�>�����,�$�n%�iR�����m2ʘ��L�2wZ�36�T�D�J����=�L�m2���jâ"&{_U���L���QJT��U6ͦX�ޜmX�u`f/b�>�>3$�Ԓ�S�	
#m7Z������񦐰��Ҙn�\�qLP<J��Fх�#�I!`v�َ�����R>oج�L�7E���IR��UJ�s���u�*I"�@g� /�^�}�G���?���~���e�KZ�X���ƪ4�HКn;=酁�zaf�Z���^�v�ʱb*&�D�S2%E�6�m����`9�j�{�� �*X̡��cNR�����c��W�T��X��STED�K�F]m�������Wh�#����u�xsL�g�����
,Ś~�~�����v�jdy��ζ�͇��|EITM$�RT���L�m2�s��َ����>��¥%��R8X�q`cZ�X�#���DTDX��Հ�i�{~�ED�I)*�UUUT|��f6�y��=����	T�I*U4�Uǜ��s��Gk\|����Q2�VF׫�)�Y�)J�;U� >�ɰ�x:��yæ�Ż��vʛN� s&�߿�775C>z۸fk_n�×$T�355����gD�Ϭ8������dhpRHJRUBIQ�Ǯ᙭|��y�3���"M��J8�亘��>g����ױ�g����"��u�}w�N��PEITM$�UR���n��|���f��N�PM5PT�}�[�5������4^�-�4Ţ����s+�Z`)T��*�1T���|��6����Ƿ��&*IIR���UG�3]�1��&��g���_� ��*�������{���ݧqf��*ffR�JT��>;7��\|�5�3A^�ʌ���IBTiˬ��ڮUs��<���<��>�߾낼^�C�A��v{�/{Ƿ�߻~�x�[2��*��v�;.�v �nѳl���E����vn�1�dR���Y'{Z[1�۱d�S�Lی������vҟ�_��s]aλdے-�(&����W`q��,u���K�ю<��t6��6r�	����OWV���'�\�7��9��v�F8�յD���
�s�N��+�6	��ە���+�r&N�T*�ݷ���۱�J������������d����x�����ۮm������5��u�[�X�y�UՍ�~���,)J��D�B����:�������L���.�JR��UJ�Up�mi6��=�3��]{�VrD�Q
6����7p�]D<���f6��q��EA4�hUUp�]D<�����cw�7�D�I)**��R���݃1���n��3�߽��.���]��HK�t��9T�3�Ţ)7���uY���[[[w�l^��l�R��q������u�u��f���e��赚����{�^��^*�����_�O��J��{��3_ndL�Tʙ�*)L�U��u��f6�c~��0ـ�bi�RNms��۷Z{u����\=�Q��8��*���Q*����>��{��TC�n.-�b�:�TB�����vУ�m��	�2i8vs�2�����s��>6D�"T�5n>}�f]g���;���������_Q3DLR*����C�Is����3u��y�K���%B���bN�d���J���E�۽V�MrwRIq5�sk�������U���g"Ӄ�G*������wu�E�7a���B\S$�)@�*_{ۮ���n�ڍF�����n��ͯ�]U�p.r*j�ʮU���̊m��M+�vm�i���5WD=�Q�n�����w=&"4��))%W}���}�,��{.��Y+j����iOiF��I#i9|�n�w��]g��*��.���9)��
�D)"����מ{��<�a�����O@�@� |ET�H��=�˿4G���"b�UUJ���v����w~����kD��[�v�i��)=��d�Bp۶�SWk�Q��޻�[�m�n�%j%UD^cw����{u�=�Q��DT�R�R*UU�<n�>��3�o�"��F���\S$J�*�K���p�]Q��ǌm}��aJT�T)�SUp�\W�{u������w��a�rI5(JD�UD^cw�����Z�{����&�K�`5�@\f�[g�J�xd�ݔ�C�t�W�"�El0M
Zq�C�7�۶6�p��,KM�.,T�����V�ۛAl ��X� ;0����.�̆�V�ݥ{S�=�aXmv &��۶���l��&j짞:����LY�%qE�{/d֐M	�,��x��nxQW[>ݜN\��������v�Ϗ@m/�ewH�]R�o�x�{�{�ݷ���^�=��Y�%��AŇ��=q���.�v�u�ln���GZ�ƹ��j�\�(��Q������7a���`��&eU*��{u�=�Q���n���YK�%
u)���{%S����3����u�V�����4��%UD{u���u����먌�6�*A)R�*�_�3';���9�y{7���9�}�Y���D�lє6�����XW[OAa�q�R�F,G=vٳ�6��
QQ"���4�|�}��͔��6Z�8�3�72� ���V���Y����=��/j��Y�BN.)I$�����Z}��]�msVB�R��TLMUD^cw�����먏k�6��)UP��R��ڋ=;���˨��n�$9�&*��J��K�fl��{��=���1��DG���]4�e%Y�6ت�e'te�ec���]�p���u����:`�Q�MJ\�Q0��v�3eU��w�1���������ADʚHU
�"��w����u�먋�ؘ"�M8��tb�1�������yw-��I���7���'��Ns�UH�W��� v��a�
	]A�HP	�U?FkP����J�h�R��D��G^�a6��D �(JU
��E7���� ����|k� ��Ҁ��V��I� ���P��zGl�v�؂~�;�hC���r�o�qJ�������ԥ ��g��|��#4F�f��qJ���=��R�����)JRu�}��R��<��qJR��o0���͖�o{�+�����)Jg��ÊR��}���r���g�k�R����pz��r��\�*���5��)�� lR�3n��<,����u��6�l���q�۞��vs�9�,��խkz3{�Ҕ�'~�}����%>�>�\R���}��ԥ)���Àa�s���i�J4�r��rIuΜ�J}�}���)I�w�pz��d����)JP��g���O�rS��z�̋�,խ���\R���Ͼ��� R�{��8��d���~��)J}�}���)I��|c���hޮs��.R��O���)JRy�����R���^}���	!�C�g����$}�?��߮�Ӝ��+k�j*�@N!��nKR���Ͻ��ԥ!?y���}�����9\��粝���(aB�0�TF����f�����ۡ)�j -4��ȁ�7��s��j�k�U\�/}����)N���q�%)>���s�9A�Q���Q"���4�|R��r��pz��>�߹�)JN���=JR�g���)@�����Q�l�F��淮s�ԥ)����/�d�'~��\{�)O�߹�)JR���}�R�����Y�ְֵ����)JN���pz��>�=�\R��<��~��!��O���pR��=���{�z�ozٚٚ�o�ԥ)�����R�=��g�
(���qJR�����R�ʤW�*��~�o��ԉK� �M�9ޜ�����Ek��1v6���m��&`���8l�)�Ds���l���o)��J��۲�m�q�m��F˻Fp������`姶��Xw �/fCǉU�ʝ�۶
�5Z"��n,���{aۮ��ݜ4u����콶������aw<�c�*�U��-���	uM�q7WV����y��l�qg�1��5�ݷi����{����|��곙�& ��I��c�e�b��O%u^N!#����QJ�?���ﳻM���j��e����(~�����S�=���):�Ͼ�r�R�R��3]��+��+��IA�e����s�S�=���)=�!��~�ԥ)�y��┥ w߾����&Jy����q	ԃrU��+��ۮt��R�g���)MC�~���J�}۫�(9�W�ب��D�����\�}	g�}�)OP޽��/P�)���ÊP4�y��pz��#���3������Y�o\R��r��pz��>�߸pZR��<��4�)J|�����(9ZF�5�#��ӎ	+,;;�����%CQ�|8��<���v�U���}�\%Њ�$���wuΜ�+��۫�
R��<��P)�y���~Ȁ˒�>y�ߛ�JR�g�}~�f��fkY��ַ��)JϾ��D~�~y����߿5�)JS�?>��)@r~�ߺ8�������/�~�f����l�f���R��~k߿5�iJ<�߸=H~,d��~p�f)I�~u��R��+jjT�"��r�w�Ps���{~���Jg��ÊP��'�{�\�
S��ߵ�)L�N���s��f���\�7�pz��>�߸qJR�����	�<�#Rk�~��(|�߾�JR��w����_�K�у�m,-�z�����sĥ;�q*��Gb��cM��\<f�f�����5��)JRy�����iK�>�|R�({��~��)J}�p�)I�{��a���kYf�[�o}p4������JD}����(���R����>��ԥ){y��f|E���,�Zַ�)JP��pz������)O���0��ߺ����)J_��}�)JP��y^�YխZ��9����)J}�p�{JRw�u��R�����)J^��߸=JP6�-���m&Ԓ�%_9A�Pr��n�s�J���N������R��;���ԥ)����R����|G�~f�{ܐ�Mu�ۛ�������n�.�M׵���h,�F�7;�p�n$j��#~;ߙJR�����JR��<��ps��H}�tqJR��=��R�������3-�,���k{���iJ���=JR�{��8�)I�}��JR�Ͼ��):��=όw��ц�p���pz��>�߸qJR��<��/R����}�Rd�z��=JR�z}��խ�ٽ淳�P��'���\�)K�>�|R�������C �!���~���.�9���)I����G�ճk,��f�[��J'>���)J;��=Hҟ{��8�'���O}�pz��?>?}��6��v�ї��4�sԢ��bn��B�l�Ls���Cͬ���ݠַٚ�)KAC�}��ZS�}���)<��~��	�@�y��┤W=X�Q�ӑ+rK��Nr�����ÊR��y��k�ԥ)}��o�R�W3ۚ�Ӝ��R3e����m$��ַ��R�����pz��/���R�����ԥ)���ÊR��y�����N29����Nr����n��R�=���pz��>�߸qJ�k3?~�s�9A�V�~�?��"#�8�R��￾��ԥ)����┥�y���)K�>�|S��R~��W��8O��K"6�t�^�{5ȅ�6ƃvݔk[�1�G[���v�TY�N4���7Q8M�dB�7n=H�`�L;b��|�%��E�����Ƌ�ļ�qG1�������۸ѝr��۷M�v�¡�J)�J�'Y�;��P�-�u��N6݀�Ժun	ݓK�{dz�	�/N��FfN�!�n#+����YT���1�I؏�ID�� s������Wk�uɋi��j��e��;F��<��cE��c����^�a�Gn̹C�EǠs�������R�����)JRy�}��R�����+�L��}���)O=>���u���[7���qJR��<��R�<�>���)J<�߸=JR�{��8�s�¼����D�89.�Ӝ��_y��┥*w��}��R���~��)JO<��=C�d�{y����Dj�՛�fkZ���)K�}��JS�}���)<�Ͼ��)J_y��┥W>��fЈ4��Nܒ���9H����R����~��ԥ)}��o�RwC�����)N��>�3Y���7����J��04sn���؀�z�Dw{]��m�ٺ�LU�+��2��3]���{ݷ�������,��>�_o�R��w��pz��>�߸qJR��>2���oY���f�f��R����}���� �;^��{|���R��w��R��}��)O(9^���s�W���{ǭ�"��No7��JR�����R����}���S���d�{�����R��?7�)@�w�m.D���Wq˺�Nr�������)<��~��)J_y��┤s��sn�Ӝ��+ٻJ�uI1HD�{��)Os�>��R�}��^�~o�P9�>�����9.J}�p┥'�[w�=���]�iVR)lS�Z���W���ʉ�;J�s�\XOc;uθ�Y��f�{��R��~��rR�;��=JR�y��8�)Iߞ}��JR|����"7f�kZֵ��┥}���ܝG਒)��ߗ)JR6�꓊�q8�����������3y���j�o{��JS�}���)<�Ͼ��.G����,��+����?7�)J|���ԥ)����Dm��)��(9�W��ۮt�(����)J^���=KAJ}�p┥'�|e���,��37�ek{��)J_y���K������ԥ)���ÊR��y��pz��/~�֏����@<܆��:헰I�N^P�n�^�ˆ(gkNp�g'>d��mQW�����A￾��ԥ)���ÊS�I����JR��~��):��=�|i����4k����R���{�)JRy�}��R���߷�)J�N����)\�{h�'D��i�nJ�r����{�>��ԥ)}�o�S��u������?�)���ÊR������f�F�淾R������)JP���}��R���~���\��!�'BB �D� ��=<}�}~��ԥ)~^�}~�#u��zՖ���R�?|ۥ�9�	/�	s��j��	p8�wޤ�!���{���)C�^{��k7��RC��3L:�ns�z�� Wn�gp����u���G%�v�J&���}�wޏR���{�)JRy�}���%/����ZR�����R���^�j�F�m))�%_+
�9�
�fon�Ҵ�2R�=�|R��￾����%>�5]_9\r�����fЅ"�$9,z��/����JR�����P!J}�p��)I����JS�u|���f[��[�oy��R�K�}��J~����R����>���x&��콗�|r��Pr���V��"IB0wn]�z��>�߸qJR�O<�ﹹ:��/�>�|��H��}���)M�^m��m$��ۻ������QG?qW�<"Y��
JKs(7������н�c8���ky����\"
gFBc�����X`�111�%��������F�8ȽAY�a�oB��`�%fKX�$*eCV��A�c�QAI�I�F9�H�P��KkRf8@nZ�*�����Z3Y���L)�e����,qM��(JX�rT-������`�$.by�'%�vD!�a��6��5.HD��HC����+��v��4ᬳI	c�ƌL���KAf9�2�̳��5�%()���'�;�QM���3LI�t�3)��$4Д'`�$���H�K��)"Hz`�j�`��Ԃ�!���@�t��@H$�@��W-h� �qs�ǐ@2̡$�	pf�L��!(�ʲ"�(\L,ɰ&�R$L���(����3+=����4�7үdl�1#	�5M%S,I�i���e�fR41�%$�h��*��򲢩J$�>nK�E���7�qɷ�߇V����y�p[N1�ڔ4�7+�)'���d�S���V\��U��U��Z�n�A�Tʪ�9���F׵���l�C�m`�N��
V�V�C��gs���q	����[�tr
L��H9�����P�X�m��:]����3n�eܒ=k�{d�jW��kf�լm��P6mS��,Q��nvi6�L��;]&��N���q��F��������lv]"�[9M��=�Nۻh4�t����nZV�:槬�JZ��j�U�z��*q8�[,]F�Æi�^ln��a�T��sIfS#۰`��`�m�������v0�e.U��[�f۝f��c���5T��@M]�N�/7+B�r�M"���W*���X�3O�� �Z�S��*mU�/.��ڊ���ؖj�e��H8E��krsRp/;XۛGYk=i���jҌ.�%gcv^�P��5�ѭݜ�t��zn���Ӵc�m����hZ�؋�,��ӎ��*�8;���̭.��]UC�m��{uTP&l���:%b��ګ�۲l/ 5[^A���Ӄu��$����e��W�׷����$T6e�\(l�'ql��í�:�Z6³S��cl�!�Y�j�lQ�q��[NPʹU��;>lb`1���6���{v�$<}�p�A�-�X�6�ĸ{ƒ�o[�����u���@��9ű�F �F#�(6��)�طJ�8u�a7�v�iV꺶���i��v}E)U�)XM8Dlrp�"�R�nU��j8���Cg:�.��w��vkf�Ù^,���tU��������f]��Ҭ�x7j�\pqeR[�S���@�`8
'O9-v�Uj��9M�E���kfq=\����q�]��W�t��G����&�c2�Y�L�0���U�P�ñ����f�ljj�v�+i�l8��3enZ\��݌h�q;X��NAU�F��� V6Q.KsïXwb�r�YujlU�	~?_��w{ޱ�v8w�t<GGj���⿲�w۶�����fq��Pt��rj�{�"]n�{aM͙Ŭ�B�]<� !� �m\��[�r�nJ0*Ln��Ӛ{5C�:z�=��u���99�7f�
Gie���^�؂������|v��}%��5�s�sA��R�`�׭�]��ϳ��=Kj�}�T��[������3)f��<�a�w%�0��q��e뉞��\��y�{��{����:��oc���rF��B]�H�M�u���m�uG*�������_w���������Z��[��(�Hd�~�oۮR����}�)JP���}�N��)���ÊR��w����f�F�淾R��x��K�#�Pg��<ߩP�ݗ�<yQ���P�Q4��X�n����Pp31�� ��4�Z�`��*Gs����u`ff�z�ݖ��`^:>^ƕ%iҐm�V�v �m���J���7�u-i�AHB[�n��`�gl�pc��k�z�@@F�vs�Xõ��t�O����� [nf�73iy.r�~�ށ����)"E$�:��%��Kx�.�8��t�����7;��������R�I).�$��]Xb�ͫ� �m�y�B)uL�ٔ7$���oWP��}H��=캰;�`V�"
lh�s�i�vXwse���]_R<��ށ��l�8�De8��-s!��Γ��8�\Z ����P�F��l婸��ѻ[��'e�� ?nh��T}�ݠ�� fhhu�jF5%�䓠^�ok�g�w� �n� ��l���A��fĩ(�lNSnJ�77޻ x��Ư����9�,�/�����6��u`{�%Y�Q�GMȢ$�B��/ gwU�ɸ�ņķ�� �&��E
�JBG�w1��}�<n-�@���`g��m�En��M�CC�2�	c�Nծ��'�h������Nݗ#R��REF�q��rN��ݺ�}^�<�w���r��`�QR*nJ�IVfn��ynk�Iwwe��.��
d@�% ԓ�IZ�X�������,��{��?}l�V����J2��ľٲZ}�ue����uf~���,�R�w����`��0Т�$hN�w:{v���݁���h�sUb�[��L٘3��h�Q��^�o=����B����k3Nώ��Ɗ"�m��$���ݻ!�� +m��}�J��q�A�	ʎ����%繮�s��A�~��XZ�n������Ǵ��*�DR*V��.gq�� }��<�XA�f�Z�.D�jS]��g�n�{۽�<s5���,�g����1TrWc�ٙT�7vC�ڸ�Pۚ76����u�W���1�nI 'I��RS��nmʯ3�l��挲�ђ ��ihv����Y��fE�Ю���<����\�;3��G��'I�+�t���{3�A�苊%����bq���\'�I�1�=�e]��v(��x��;���V�=Y�oF5 Z��m���@�"�՛�������nG�8d�� �;�gNɌ��˙��۱ۭ���s�u�n7��s�K�rF�l��JP��Xn]� ���utl��X���h���N�	L�gn���7 ԓz���]�WwvYi{=�_�9Ĺ�p�z����{������w�� ��ג�\�5�@n�������a���(�$�N�w/�3sn����9�����:�!δI2�L�rJ�=���@�y��+��ܖ{���]_�3b\�m
&�bn)$�@��q@{��!}�9�5�F�n���~����U��X�EI�%u�<�"\��]6�磣�ں�P���SsF�u��J7�WwrX�eՁ�noN��y��3�m�R�IF�5��:n����_���\�I�~�}V���v�-�5�s�K�ks4T]:�LN(��J�7w����z�A���������n�
% �5 2I���-�v�ݖ��ua����zu�=��kQ�uv{@ۚ �͕@fcw`l=}T��1�ܕ'�D��7HI����`ld;C�˞.��[��u�w�����g��8���r;����V����[��������$�l�rJ�33\�bI �z�@6� �ͥ\��֩�6�RTME���1n۰���~��?��0�4"d�������J��y��w�K�`D)���w���m���J�������\IC��`}���Q�MtrN���u`fcw`l=}�m˸��nf{�=����vVGb����d힀�8�۱��2����p�X�sфY��������?�v��� �q��p�Ҡ1���(
����$�@Ź��U]��`{�˫���z���V��pM!N&㰸�m��nҠ31��FC�� ���u��I��Q���۫1,���~��n�A�����]%�\\��{�@-Xe6�m�
A�%X��oz����s@g۴���\��o����w��8���]{[Q��p��Q�m�;u�7cbgf+j�m@1�(�&�?�����ҰwuX�w��77��Z;��*b]J�$�7�wv_��]Ձ�{w��s]��*�ٳ�%>D�jS]��=��P������������՞�Qt��jH�$�`Q]^�����|���Ws&�w�"�bRUJ�����O��>��q��6e��}�ܩ�Ϫ�er�r�H�?���nI�6�kW.�k��B�qcb6�u��!XZ:�n0q�GQ�E�?˻��\�f.U<���*��+�R��c�z��v���m�(��k�F\���8�J�8��W��v�J���l;Z��3z�e�9ŝ��X�v��\e��#�����Ǆv�kd-틞��j�u�aW�r�q�QH���m����B�cy��݊��>�́�u[�nӓ<����)�;WZ-ނ׋�nsQ�&�H��Y^:wG�����Z�o��`{�˫=��{�Չ� ��0m%RA�n;�>K�8�����(����`�Q�m:JAI",���@�^j�6��vX�2����%Z��FӄME����(�s@f�ҠFf7vDG۲>9B�%%4�
�wvX���t��_u���\O�tG��LO{M�)����z�!�7]g!丝6@��!�JE��2
�$��+�u})�$�R����??Tf7v�����m�LA��
����I#rIV}������W �VUv�Y}���3�G�y��΀�{w���s�>�h5�&���\�>� ��?q.$qq.r��;�����@<f:+YQq&"18�
��s@V}�j������8�ŏ��P������$����t��ՀUs�����7���.� �.�MM �=m�Ql���ͺ��b5����͕�IV�vnS����w��9���U�Vj� o�v>� ���I..$q.X�۫?��+�(�p�������� ?��϶6��8dF�N='RJJi�a�}�e�{��Vb��#` ��www}�ώ�ꢹʢC�_�_S����&І�-�8X�@ĮhS�d�e�k�;2�V��٘�P��S$�@�(%(��!��|���`�d�ڝX�a"	�������⪽
�Ȁ����Ҡ��j��
LU_��� �"���]�(i@����^]ϋ������7߾�v���MZ��"J5�)'@��mmՁ�{w�ې�a\����
��CP�GS5T��n��\��p6�Ϸj�{�X��*!�L�N�m����/��qh�{����%��ճ<�ߏwã��T��JI}��U�wwe��/�����{����T\M��n+���W�&뻋w{��7�� �`�ւPhuWʍ���۫���z�,���(�����<`�2	6�JH���@fg����(�q4��G�ۺ�>�j�ȯԅ)ȓqG'z�� Vۚ>ݥ@fcw`bz������Z�v�vf�����`�gS�@��Ů��6��mҤ4���8*�DnRn+ ��Ձ��Ł���������EL(����vj���mR�3�n�}�
�;����{EӉ!��I$��cw`k�[�4nm*�n�H
�iINC��Է���`���`{=�Wԏ?~���E�.���}�� [�4nm*>�����(ɥ�5�#���@�p����������[�Wkm�ɗ6G����/��x���մG��ڶL��j�g��o�ZX]��r��.���m�I�c��v��4Y��[d��tm6n{��8�,7.��m$m���x爑�j� t��9,Z�D�8����su�;]�@��q�m�5S�&�CoxE�rc] e{V�v��n�ҙ����U�r��r�q4*m�1���\U	�^��>���v"F��WM5n��:Cub�.��AnS��7��Bu#���v�T`�6����?t���_u� [�4���"M�i�9II*�����y@f��`��`�d��yV�m	Jq�����}6�}V�w��{�cu�#�� �nR�+ ����쫫�{w�5�>���Q*Q���NM��]*>�����q@
޹�3C�?\���j"��Ѧ.�\+;^M�[[(q]�sQ���XR2��;�k����6��:���{\�������`n7q`v��)�
��$m�'z�櫺�9�$��]���!��S@~��J�ϱ����+YQq6�S�����,}�
�=�����M�n����)�R����tO>��5��� �ZT�Հt�,�$ۦ�Ӕ���}���׎(޹�3siP��8��uʙ�fK�+m�T��^-]̎2�6�6�(i�#�l���7H����(JS��Ȥ���6(޹�nj�@g�������s�8���/�Ve�_R<��ށ��U��ϳ
�Ju��]��g��Õyߟ}�W�ҽ vß�C�~�<?;�`�ղ���e*.�IԢ2>̪>���}��t���T�fR�
T�8�i9;ѥ��U����X�L*�����@U[�d���`��ƦS����Ŋ����u�SL��Q�@k�9r)7EFTT��Jq�@���X�f�Ҡ3�n� 5�� �M�� Q��nH��@�ͺ�=��{��Fk�Vc� ђ�T�(R�R�*���������q@[�J��f�ڰ/-|%$�(؜�Iށ��U��ͺ�=��T��%�s�UnϽ�����0(��b{�Of(mҠ�seP���������1��iA�m P��q�Q'Fh$E�q;V���΂�k���,�nғ���@�ĨG{j�׮�31��5�\~\��~�u`nnҢ�đM9I�ܕ`{��_u� [nh��U�j�PC
��m''zk�V�ݖ��u`{���@��c���*m�q�@���`k�q`n�w���l�O�RBJ�+� ��Łkw{�@�~�Uu��o�~�l؄�� �ɨ�H�t$�8�)����=�����Q�t=l�0�[@<Fw�l�]o��*a�K:Ý;�Ā�=r�4�n��n��s�7I���ķ&�''f�S ����v�s���K��E�� ;ˮ� ˧�ym�����XZ��	j��6�#�g�m�����n/����v�e����ظ2v��:;���A9�nI�V�g�!�i4$��w\p�]���;К�jv�S:4�vi=�K�����ydG-�xN�nv�
Ġ��,G����B�ݬ~~w|}�&W�R��̦�~�v�q@ۚ76��
��
S��Ȥ���5_�T�}�ޚ^�Tfy������ �ꘘJ�R�� ���V�w�-���@�� ϳ���$��b�I:f�Ҥ������q�Py.q%���T �ͥEӂI��Q������m"�[�.s���C͇qa�e��JE�uՖ4�۲9�pp��"Ƶ�pB����$)�	��w����{tl���+��_u�[nh��K˗������x/܋���8ۊ������}�U/q8qqo.�~��H7����qt_a����U86�7s�nmՂ31����@ۚ#�����4�R	�*�)����k�f��`z�P.76�1������3vf&f�����}��V׮�dB#���~6ݽ������n���K�BA�qy�P��\�Fk��|�n��.�X��_�|�� QR�*�J���r��5븸77��U�(��s]�Q߳
�JuDn1tNeX׮�p��`l=}�z怬�e*.�IT�E#��}���@ž������X�W��?n��f}���Dg���(�W�G�ʈp�F��zl=}�A�nhf�ʠ�9��F�������+x�r.	���n; �}���x�T���؃!�� �Hdk��n�d�l�v7.g�;3�3��u>R�7/<B�򗦦$�	5tX�N+���7q����@fcv������Ѐ�lfP�&6��rU�������j����}�zh@�siR ������3v{=������@ەG9�Y�����{�3�7�$����"r_���[nU �siP#3����\�q
Z%QP:���~�޽�9� G�ؿrWy0D�d�Yٙ�z�R��8�%�����(��Ѓ�������ͽ���au��.�+��6q	;s��lqp[x�5bn�;t����b��@���b���� |۞s�.P��V�ez�[H�rG$������Ĺĸ-�-��Tϱ���1VqoP��Jtӎ���,	���V�$�\Acuh�����[�h���LG{Sښ���G��j�[����@��\� ��hM#u���ے��f���j��t]���w "?n$�2I����9�]x~��`�3�[
"�Y�2�[ݸ��a8��-����($��;�����{�:���4�0�����놸��rt��{=��E&?[���~>����
ù(
78�콵1�3ō���v��5�mh�i�zݻ`�b�{@�TQ ����� �F�j�R�&�l�Uee���ү�����b�hR^�>B�]����‥SR�G=��P�����l��!�\�j��:7`�s��Z�k�U�ٵu@� đ[�y�CkV�Y��Ol2hL峵��l��$�ݶ�qS�.� �)�紋��mmk����]��;z v��3����[@���^lᶋÊ
*�Z,��n\V�w��y�V�V��sihy��ݩu�r��u={Q�1u�ڰ���5��]�J���r*ؘ9Nu������5pK�`�k��r�Rf���S�gn(�����cF�����*8��Ցyul&ie��`�ݢ,�����WUU[U�Ź"��^C�`Ǒ�mY����檊Y;U����j]���W6�y�ag�˸��j�`��sVka�=�M���.$�2��%���4�J���ݸ�KdkhHG'G:ke��􆛬&nK�Lm��^y���Ύ�����Z���D˲ҭUQ�VV5��*��Q�Z@^���,��FC��Q��eZv�T B!��Jd��ؓ���ۆb؉y:6����g�\�%)^Y�^y��v2u��ŷh���=��8e��b�qx�7	RX�+�V�L
��km`[� ���s��T�e�I����36],6�"*Z�/^%k ��G%� ����;\`h���j�^٪WX��m��e[�w�,ɳd��n����n�6z®�.R��)s��X��U�U��mW\nE^%���dv�ʢd�kj!)ڀ.�ҭU\��ۗS,uΛ���	.�FYj��n�"��31t���!�k-���Qg�2��[0[sWW��"]�Z�k��UO(t��l�u�&\����o;�p��W%�6��1�yk�eu�� �J)Ne��e���t�8��qd�}����O:y��,����պk0�(H�!������a�`pz,(���!���'?�:!�� ��Nw�h��/��<������l���v�8T�v�f�F{�����m���=��nS�&:6���ϱ�x�X��M�m�8���]�3���r������#-�e�'=�v�t�$Bc�ی��g��ۉQ��uI�q:�3Y��u��l�\����حѬ'��q'&g	�����������=�<dt�R^1
��]�
����Sl�q�Ry�=��k�ȗ�����~/���Mn���mFcuŬ��N͵���iy���Y�$6"d�\�r��vSB����I������-�n�Ү$��}�݀�z�ԒJTt���(+��*���e*g��؁����d���s{�~���`��g�w�6���R>���k� ��l�+�̥C�!&�5 ܒU I$}�݈���T(-�4\�{.����+�b�D@Ӓ9"�v�P'_h8ەB��T����>������o�6�m8�R&X58$nf�w�����3Nq4�vӻn�fS6c��������݇������Ѓw6� Ff7vq���(+�a���h�T�CwQ���}������Kgc/HOЏ�����{Y�@ۚ#M#5��j17%]��{]
+V���E��U�J� �@�%LA3٫'_i����ͥAG��ok�s3`��$���N;���g����. 75���N��\���?Ȝ@��^���b�� �Y�y�b�=�!��r��άfmvx[[t��(Y��؁<n�3�nՀ�n��\\�������PW�
R�6*q��"���g���=������Bo۴���^��D�M7$�9%��Q��) +m��X�K8q$�z�^~�T~�ٽ��=�g�b�)4���P߷iRfcv�=�4�>�g�ȩ��w�]"[�۫�PQ�cwb=�5�A�nh@�5�{3�pZ����c:���sv+b�k�� ��(�U��.��_��8n�a)8��`��z�@��������*f�f�I���G�w�f=[%���Ѓ~ݥ@��mZ��.qs����I%*P�NK�
�������2��؍������� [���OBbw�+�DL͈��Rfcwb�P(~���"� �������8Q��@)_�SN)�)*�����`u� [nh�v�^�Ը�������T�.l��и�.y7gj㮬Ϝ9Hx6B�%�lp�ӯM]c�k�ni��`7��9�7��Tf7{���c+8��|J	D9,��/�9U<n��޶�w`o�@i����Ʌ2��ڞ���x�*3� {�h��,K2�B#I�2�rU��{]��s@ۚ~ݥ@cA�� J0���w����;���ϳ.���BK��<�^�Ts��ܘ���к�Ș��N��{5ȅԷF�1��Z�f�'!tkn�m`P
݃���+��7Q��z��N$�esՃM�(�搸�:<�@�f�&%�A�ڀ(6MW���Ӯ��7a��fe�V��i����bv����.4�PtP�T1�!1�OnNS[\��V�/���s-��sj41�C�2��mA���
���6�v�yݻ[f��ms�{���w��U=;Q��j��qтM�K��^���%˼@�&���9��DT�I$�F'RD�����3��T}�����7�7<
% �����3ap�U��F�����h�G�6Y�s��<�R�5(�&ړKnm;���ID_d�VҠ>�ӢE
RI$����uՀGs�7q`now����tI?��@��4o\�\\[��r�ϱ�����߷���SI�*rD�]����2�׮�ZqӺe:�:�� ｅ��:ÑT����M��T ϱ����˜�.q(�o�`��JLq�9*���������qs�A2�4~~�w6�.$yf�$"1*R	�;���`��`f{.�}����"�KRI)m)$vf��K�o\�������(�o4�� R��&H7iI:��ŀ}��� w>� �}Vhr�/3i�.7��Њ��!���C��B��u��۰���w��cl=`�v�\�}�~���z�-�%@n�Ҡ>\Y^��%*jI#�I;���`��@n�Ҡ3�n�$��q%��!6'��%*I�������,�eյ�_�^�qr��E?߮�?~nh�64�raL�;ڪ����t����=}���o�`��J#Lm��r9V����@p���-����O�S=��yI�4n�!W�:�b�V��l�ˋ�v��7C@P�D��i��;�5nj� [�4�m*>����d��5�$q�)$wiw6_�H�sn��~�ށ�s]��
R��&H7�I:�t������ ku`c�%jI20r��aTo�7�V� ����s��%ϒ���b�>_&�PJ��RI;�5nk�
�w6X�eՁｻށ��l�8����45+P�ͳ�v�c��j�[�t��ԡ�Nx�<��-��$��Q�NK ���>̺�=��{Ҩ �͖��X�9Hƚ����t��� {�h޹�pif$fQ*&1�I9*����ހn>� �3��x�Ł�e�T%(�&N�{7`qu� [�4��J��K�R�g�������ԕ
H��E$��}V�/��/s{� 1������{�_���A���Bs��Pq@�u[S=�<6@nrD���M�k!.�I��:E�=��p�� �����d��^�N�W[;s�n�6lE��hҽ�3�k�t��8S��0�F�nq��4v��z^���#��Rc���%a�vrv���:4s�N�t\t;�l�0����Etn!HC@��l��V{Xv�)��n7m��t]�c],�?�{���å~�53�\$SԶ��hp�wk��f�#��'$���Ҏڀ������]�՗�A38kt��� {�i$�-���JĒda �RU�ｻ���9\Q��*�>�����*�-X��%D�ӒI$�w����;����ye�����ށ�^-�!R�ȁ�%�p6�߷iP������>�kER1�r;�}�u`{���@73e�wwe��W��5$hPP8m8�E�]��nv��k��{BQ�ʑ6�ln-u�Ǖ��rդK�TLcn6�rU��{w� ��4m��8���Ҡ7��{�&N�� �s�Ks6_�z��TUs�N�����!��*3<��f�����'�!3ɞ�� %�nh�v�8fcw`���,�+5�L���Q���jn���݀=�4�J:d��@cԨ�5	���r'*����{�?r��Uo�`{��X�@{���L�z��GJ:��ٶ��{n���L��.�gƛ�S:�[?>�����=��������{ޙ�m��nҠ31��>���D:"*l�hNK ���9�}�u`{���hs6Y@}�,5PÑ�n��M��Y����7�?�o�އc+3��ϻ�����~���s����ð��:S8rgyFfa�e�`lD�de:���Qq�;�� �5�y��`Iu�P��P�n�4&��+�C[M�`��a� �(`)��"����(��i(J��1!|�P�)��ҽ���`	�<���_��"@���O􅑿�s8�ưc��~�u�a��r�h�Fa�4�ц7��?� ~|
��t�P4�� ��P`P�耽�v���AW�O�(W?֬�����we�g�~����J��m�{�TI#3<���Ȁ���gٗV�� �(��4��r9ހn���%ė����x�*3<����߳��n��gVEWXsr;s,��3�r]��wG�Ն��s�gg3��j�*bff�-�4��J���\�nf�>��E)¢I�4�9'@�nڠ31����E���s���"S�Bj��nK���zbF�ܰ���2Xg��[J�I��'$��$���\���7�٠���H�S� t���?<s_���깞h���B�A)R�ȁ�%�o���ϲa`g��ހnf�ȭ�����MD�rB�����p�G�=s������ V\�)wKu�>��W9�кEa]aȆ�������P����s@ۚ �!f��1ӤA�;2��n�K�� q��@���ϳ.�n�(���% �s� f�� [nhK�$�Ί������hA�������~������x�*3<���\�����4���	J*$��k��:�v��ܪ�fg��|��4m�V��R\�=\����c��$b���ꕹ��t��N���[nv�!�t���6E\unlT��F����zy)��ASj�i=��Og8���A��=s������=����a�;�7&�Y��`  J�����;o6��&�B�p�S�[&�p��ym�N6��(��gE�y�GrHP�+F�84v�$�	o5�X׷cu����`�l�/��}��ۨ���̽$�t:볽)���$h���F��p��n�Kڃ/������h�К�$Q�%X�o��s6Xwvr��7sn�nQZ�R��d���7`�ۚw6�������Ur��[�P�p�R�ȁ�%�}���`n�m*���x� �?M ^�:�)�q������p�6f�X��{���`��`��ʈ#M%�w�*������=}�mʠ7siXUW�8fjq�)��"$IQ	������7V͵���L%Õ���
�l{K���4�)�A��z��v/��3=�_�Π��߻�=���I�%I8ێ1�5ʮ�����x>�&z�
��G��Z�=�ݫ ׮k�7�B�B�MH��rN��]X��k���3se�Wwv{�<�J����Q��P����sAە@s������V-�Q$ƣ��$�@3se���K�{�`k�J���;��}՚�vH��3�Rp]H��$������,un[�f�"N�9wh�vcbF�F�J	J�iFrw��vX�Ҡ31�J�5� �M��
I��)WI]xϮ/� 3w�� |�XsvY�Պ��$(��)H��,�n�^����&��U�zh{:X��-҈�lbR�N�s�76l�hܝ(?r3w���o�A�)���nG$���?f���=���z��,��Lu�!ĚU"L"�i�n�v�u�S���)^|\6E�k.:w]Y�3��y��J* M�5jI:nmՁ���ހf�� �n�"Y��T[��ȧ�*�ϱ���\^�4�74nmU���G�(�_�TI1��m�;���� o��	$�76�kw`}cH�*
�P�����|�z��߾��G�:	EF^���"Nr�����\�
����aȉԊ����Ҡ%�_��X�s@�����ww����;��yu��4UZ�б��6ǋ=�z�v����2,��:y����?rs�$��7%|����z��,��l��
��+�f����iK�(�M�% �sv�\�}�h��T������ꏢ>C]D�
��$�q�X�U �}�ހ{7e��5 �)&�mvn��l��P���=s@��8�l�3ٔ��	��D���s۽�=s@lfk�^�Tx���5Ga�u�P�q��z^5�t��b�2�.�9;2��lW%�2�B����g�7OV��1p�O�zWJ��l�]�n��m�ݰ�`+m���K��u�;rR��9��8V�,l�Efm��:��;�cX�cN�7;7kܻS�0`�.�D8Tq�U^�s7�t���uv�"9R�%�V�O�4���޷h���%D�3��www�9�wճ]9�٧�곬7]�sȀb���l+��A�-cv�l�ԕ=\�+�jQQZ �1�$NI/���Z���׮�����xmD�0%(�qD	�`b�5��eՁ����z�\\� �{�'�RDL�����lz�P���丢��c�V*�4��6E)	�Vʪ�W\�|�޻ �?MlA���L%�nڠ3t���M&ۡHG�@=���3��`{<e���{w�tڎ�D�j�����#[b]�K��]c���q����ҞڟnHr��%�!�DP�D�RI`����n�Ι�w����7;�d&����Q��$��۫�����UzUW*�(#m�� �� ߵ���UИP$�(�`w=�ހ{se�g�e��a`}�QX��*Lm�q��?Us���I(�?M {}�3�(6���*�:U�蔁J� NK �n��)%�q$��2�{��`����G6����2s�3�����lk�Ƌ6D-�����GP5��΋�|o}n��Mgk�ڛV9e����1� x���yb��ȥ"�p�3���Ns�Hz�6M�����`����w����7۲���s�\�ن#�_U�������r��<���Ǵ��B�'(�K �n�f��@nf��z����%���L�����5첀�IqB�8��~��7����snX�by�#�)Q�ө"!�i���'K���Z�]���v�9H���p�MQ��!4�$�B��{7� �͔ ���Ĺ`k�e��Nr`:�rEs� �͖�ݖ��>K�{�ܪ���n�U���7(���=����:Ps���73��^���c���A(�4;q����K=�ޮ��~����t��4����s����W��B��H6�p�3���@Ź��7�ݖ��Y�[r�r�l�T�S��s�7M�Luh�v�單�=E����x�CB��D46�r	�;�1nk�6u����q%�Ļncw`��j$�)Qr�$�?.~��Ӡf�����'v�\��9�?�?z "P��Ҕ�ѹ>l�X�n���k͖�n�(3ي��
�q��,?��w}���~��s@s�s�Ik�L�>��[�J�M��rN�76X��V��Xu�����ߔA��k��H�&Y�5��{߿�LDK�"�]!�RJX����N�߷8��  �(�Cc�%��֖Ɨ����e
4%�#�����	*���J�o�v�ȸB��Ǥ��ӄ�3��J	!�� s0X`���P��(�.% D*⑊�W��DBQ[���G-���`��8�{&�QU�U�����b�ò6Յ��6K�'M�p�h��ۭ`d�cBi:�%

���zf� F�n�U*�^Du5UeH�nzk���WP�s�
ʪ�lJ�7<l���)�E\�K��kj�]�m������f-ntm�p<�n�'�Clݰ	8�m(it�E�	ƺֳ�s����:.���V�f�l�2[]�mNI&�6R�:5�/$G$�4�aN��g`*�ʝ���#˷kd8� �ʲ�[R�+�͂8�
v{nӮ�.-�Ñ�
��[�:[�CIku��w�gn����,�i�yQ�js�*��Xm�Z�5ɰ�ْN�v�S1h�u\�-����T�T-��*��/�9G�����.�s՞g��)�Yʪ���"Yn��m.#4�J�t�I� Hs����2�\Ԫh�v7Yr�fb�V�G��	6p�\m��ۺ�����v�X�9��@^�<^;gK��ˍH�l�{n����h��d�en��2Ҽ�� n���٩�.�'MTf���\GKԥ>�vA��6魺B�:�]=-�@$�w	m�,�[��,-Ay$�Ha;g�k,��ܧ�svڝ�S����:D����g��b�r�յWY�z�]��v紅�QDQ:uvLgnap��s�ׄo.�W��W3��˲[m�\Evm�H��k���L ����ĸ�����nםճRnN8A�ˎ�3UmU����#�˺]q�m�yUh�n"I���Y���e{f�]�k)��cl��n�����RcK؊�F��Stv�J�ҷmjJ\9�y��+�hm\�ސt�����$��b;`e��m���Sf ����YA�I]�\�n:�bau�e���`x\�7UJ�ؔ��q��T�&��;j	1��^a�r���RI6����g�:�ZԺ���N㭛[v�xyKX/]I`��q�IP��j��D�d�+m�[OjR�1����w|i4 `�{� &�(�����
	�@S�'��g�^���9�؋t�/۴�L-�*�)v��2���ѮjB7	�p�5I���$�v�a��Ü9���6X�{��a Դ�ك�U5��������m�Yu�c����1ۣ��$H��P:X��CP� Gvl����Ƙ64n�'T�7lp BG{D�1"�\�	�F�7a�YiL��8�WnWc���vN\v	n���kk���{������h�F���ː��7[m�!-�qge�����a1�N��:���v�������}�3rt�71�K�%�X�s@�����)����@�ɥ����z��,_n�9\�s�Պ��Q1��JR���{��U�ӝ��׵����-�	46�$����8�\������g��w'J$���w`n���DP�D�I%����`{=0��w�@�U��ƒ詒�RR,N�6DѴ8�D+�N��!�tm:�m["L�:D�9\�������R�N��nFP����s�\�F{ݣ臮�l"4��8Y�-̽�r������g���A����. /3HDyt��JjF��w����4�5���0�:���&5���PTH%PR	UV�}�>�Ҁ����I�� .q��P��A"Jlmڸ���4�;���@=�����k�?W=�k֤�(�X{E����'��v�>Gui��[p;-�G]�����Z�V�F�܍�I�Xn~�ހy�c����t7�Y@?1C�#�u(&�SJ����`9��`ct��{�=�QOj"�*(��)����uw����"nT��=$ZcK���]��}���n "P������{=��~�=~�#[��9�r��?~�}s**�D*i�I�iǭ݁����7���Ҁ�s�|��*^�E
v����ӱ8���8���6��`����N�Z��X�\k�ʕT��e�+ {�Vk�X����Y��m:% nq)�g۲���a�ƻ��6_r����"��U
k�ڛ5�(����<�C�?v�~�,�*3�Ӓ6������@����74����s�TP֋6��Cn����s�Գu�}�,�L��w� ڞ��U	*IJ���`s]��nXք�#���!��[O(���7�9M)R4�QJ��7��`}�(�n��o��kd"%�ىmˍ��=�4�����z�7S�*߷gUs�I{5QV�!SNRn6�`c�z��o�ys�r���4��W�`�_����iI$�@�Y��s�fΔۍ݀q%�z�5�J��T�{1=���V��$���v�7���ށ�ٮ�u\�o�z���)'0uΕ`4�y�-�.�l=[���nU���[ ,��P�a�/;<Rm�5�緑�њ�n�ݦ^Q34�v�d���6F�Vku�5k���=hvE���e�ݶ�nG�k���j�M�s�B���:��>��n��������m���mݛ���*S��2��k�d�%<��R�ƚI�.��ew%�}��l<w�5��}b�Z�ˢ�/�+�$���7]Y�Ӕ�lA�훐�܍;�G���TIT�q����_�R���z,�v/�]���Tf#M�i�ڢ�ǽ��-��r�=��u2>ᙴ�M��JA�rN�^�v/�]��n��ǽ���+�I�*B���J�ֵr�=�ŀ�{��#e�Q`<}��5
��T������q`<��z�f�����yW+��OL�#tL]ۦ<���k��q���8�箻v��T���ZҶ,�^4tm�3%w�m��~��27_hk�y�J���P��"�M&�j9'z�n��u�W9UM����`n7q`<��xmD�B
�%�f�X8�X��YS/7����+ ��c���ATq���n>�,[�V�������`t��`�a%)I�$J����۽��wi�O{]��f�Ձ��u8�	�H�Q(�)B��5��9�%�\���'g[D5\�!c/k��7 
RMPJU����������n�}!���zf��h�Jq�E#����r��57qu2=��x<�Xq0MQD�m������V{۽�)�Us����љ���:[j�̆9���������uOn��b��`j�u��L,����V�%*��$Qʓ���[� �����Y@=�w`69�n��gF�K��f꣩�s��\ک�κ]u!��q�cb��:�k�î�)�Nw+3]2���{��2_r�2�㢵�AT��M�v�ٳK�� �nܴY����O�\�s�H>�0M�$J�p�3߿~;�Ս�Z���}� �ᙴ�I���ܾ�\K!����7�>�҂��h\�9�$�.�_Kڧ��Г�vD��N�MR�`��w+q�,���������w��o���,箁�h��c��묧��t�@璸6�Yp��̎�w5}�ӊ�qF�v�}7f�{۽�yc٭Z_f��s0�l*!E*!�����cw`V����=����$����R[H���ܑ�����ij��=��`<��x��d�Ђ��R�n%#�HK����L,��{�9\�<�u�+=��aPU$iSw.>��uq`<��x��Vr���v��J��%��h�JJ��ѹ�������'tr�a@�&�	�������X��.�X6��qX�`���΃c��u���j6]<9-��m��5ǅK���f���E9�	��ֈێ�9��/v�X���Lh�>�˥C�v�'F܆x%�^���C�.�r�
����Q!m��*y%M��!�&��� s�mÎ���}ʽ����׼�˨�ۛ��,#��Xι���gFz���>�ٷF�Ai^��?�W}߯wt'k�i=H9�@y�߮����@8�_W��nҠ3xyf�I(�N���s��w]���r�1�q`<��x|.D�H�L�����k�>�˫?�Wϕ\��?~�@տ�;,�3iaE#Nԏ�9�����{��2_r�:q�7��(�Y���hݭ��^���u�_�������hF?v��ݥ^�3��A��1��v�b٧T�an؜�v{R�Y��Wv�ݶ7LHd���ں�^�l+����VN>V6�,�{� 4��*�a(jTq)����r��s�*�0 d/oh+տ{߷*��>����=�w����H+su�_��	!�w.>�������s�7������G{LQ���$�&�$��9K}��w�j�ߝ����a�=�x��Ff�I$�'N��J����Vrޥ`cḾ���ܩ��nH�J:�J��Q� �lLC�֐{j� �l�y퍻.�9І�����?;�ģq��_f��!c�Vw=���^�v��wx�J*"�n��E�]�`c}��_r�N>V|l�h*!9N�qX�n��b��g�յ����� I	���.��8Q��UM5AAx�̄2K?� �O'��B��#Jj���M�MBQh�i1�4��jZh1��B�"4J�A�N8a�ōc�C�lC�3I*`�FGXU�e�0�8�QID�b��X5T�D�2$�
��� � @��rh�`��V��@�1V&UU�UT�H����#12�%��l�	�:�d�c��D��3(/����A$`d�M�HP�@IX4XX����H�����Ԇ1	L�ᡆ٫�H0#-.��(�@֋�b6X.���@�L5b���t��JP�O?a��ڏb�"�z�>v �G�iA��������k{���=�`wޢ�m"R��rH�U{�9}��s����76N:����W�
��@jRq)�,_f���6����oz,�vD��\�M��iE4t��AY�Ş���L��^��|�t2cn���:;�諧ȒP�黗��=���vƷ�ZJ��~�h�M�T�IM*I�`g�����uߒ5zk��=�b�7J=��Ht��	�ހ绕�ӏ������`<��x|ki*�J9v�T�?o�`f��P߳�����.�_hn�B�B�$�'�7ڞ�ۥ@{��y��|�{ݠk_ٮ�K��CS�"l���#b�te����\�;p�̯Wa�pj�S��c/7@�AQ	�89+��~͟��1n�5}��feՍ.��V-�D8ܑvfn��z�^B��c�hmҠ7���UT��X�U��D��D�q����3wiP�y݁��� -�ޡ5�L$�)�w.>�Y��V}�����k�Wٮ�<W�0�'RSJ�������I���lF?v���ݥ]�V���+	� ��xU���u���iHa�:�v^�i:��N���D&p���,�VQ\{v�[h���Z����I��7
���L	�q�H�5�=��E�6!�R��l:�[eT�o��z�a(���U���J�u4)�鼐v��I�!�M�nZ�XC��ѽW�O�?�h2��nЙn�sSi�h搈0N����ɲ��q�:�o� j�'����펫�k[Z�v��Î����M���{qlp-��̄3�sܺ����(����huI7>�X�����@^�Ҥ�����kD�C�uI��v�n;��>��{�Y5��n��J*"��q���(��A����q����CE���p���{w3]����gR�$���Eb�D@Ӎ���x;ܬ&f#�1�1�2�y���}��"bc����pc�:m�j7n6� �=����5���N��IpX�sH�U*�Y3=;�X��a��w{�9��bH�f:+i�$��黗@����\��,�J�7i���F������>+��"	ԔҤ�,��{��b�]��8�Q���@c�e��Z��EM��
�b��5}����Y�n��3r������Ě�G`l�r��L��w���Vc]cSs���V�;r����s�(�N�J�v�L�R�Ӧ/ǝ�=��t刱��v�`c�e��ݝ�����%�\�}��[F�A$�:n��Ͻ�{���qs�ގ�������rt� >�B��H��ԑ����]�o۲��U-8��Y�U�g�n��28b�P�f"�NHӉ��?s�_��~v��=�������=�譧UM�v�lF����7Vou�h7���}�~��RtF�t�F�-�'�Nݪ�8wOiI]�l����eD��K,K��oDvb�{����h7���lPJ2�hI��Q$��@���hF�}ܬ ƛ���{�c�*N�2����L��T���V4��w����V}��T�Rru�}�K?Oߣ��=�z�ȇ_h6���q�L��y����Hz��_y���U�U�G(�RR���X�n��bͷ`wZ�v����짲F�IJI�NQ���]O���mϢ�,
�����r�9ȑٳ��۾���ԑ���n�Wۮ��{����{䂗�k)ĩ$�8�R�:s�Xֲl���@_r��� ���[O�*IC����+��U���wg���޾�Wh�v���_a� D�)�I8����ށ�ۮ����>��V�X���m�9BL���h���l�b��q��/���r�9YUZW�o��8���i �Q�ڶa;4�,�������Oh��Q�쎑�bfh0�"x�7�씬��J8;x�.nɹ慔7<�k��v|��qe�N��2�uQ)՝�v�F�ru3����*�R�skgU]=�l��ڱyy��#Cg �6zXŷH[�m��v�]�W���u6�d�!G�Sn8s]I�W���񞹺6�g�V�4�no���'�[��l�N��$:�yۙzn*:@�^�LK��;Rq	A�-g�j�v*&�Q�������?b���߾n���HR���BN�o����{�9��`9��`� ��&f���8�����ۿv�ś�����>��W�̢�m" m�jI;�1or��r�1�s`c��x7a�OB�R��I��F/�]��?b�>�n��b��7��jnJuIJt���ێb���p��wG<�������p�uů�Ί�|	RJ7q��ך��=����u�����񔐢��)�I�J;��wz��9����Av\?���������{�bK6�%mSM9��ܬ9ܬ{��{�k聰%Q%r;��������^��b��%��ͤR�TEH^J׀�uŀ�{���r�:s�Xߏ��~��i��Fc�-���C�Y�����;uΌ���H{�v��h\�(��S`'�ݘ�ܬ��N=!��`{�b�DAM��q�;�����H���y��sU�������AK�Q��*T�q��Ձ�ۮ���+%UQ�"xJ��P��^���y��uW������c���H�%M�v���s5݁������{��t�f�D�6�MR��V�{���K7]����g^Oج�{58�
��P�(��1j`	o^�B�����L�F"��N�B�9c���$��))'z/n�W�]��zax�����c�B�
�r�mAH��;���6�`=��x<�X���B�TEH
Gq���4�3���@Ź�����;�`�"�!Ju�(�n����5ߛ��{��R�*���K�5/̢P�r(�9*w�d=}�|�j�ٝ��݁��i�Zs.�%rƚ�rn�8eglԛBf�q��%iTqڍ�1�rvqs��,�J�X9ܬ{L��t{�w)|��َ��|	"�����ܚX�n��b��5}��i��	
&&�S1)Q`<��x6Z}j����a3�m�o1�	&�M9B$�������V=�YS/u����$��ʨ����`j�뾤}�a`g��ށ�ۮ�[�����H@�m�����Q���	��'s`�A��J�zC6�De�cD�%`���M�!�Bt4�ѥ���$�a8�A$*��$��A"8`0�&#�,� BJ�	)a`Ķ�8(=)����!2B@�:�g���Bd�S�e��Q)S��vnG�9��.�<
��֍ngڧ���^�5]T;�^^tj�1�+]��|U���'k���X� CZ�li4N�[@�j�sg���Yx#Cvm������� �m��55�t�5�.cnFP�r�P�u���76SB��V(x	W�ηF��4�ڕ@S���8C�c������<zC����1+.�*���uv��E�\H9@ ��޵�4��K��҇Qۗ-�V'I@��t�Hju7L�!��m�Sֺ�H�-̶6��d 
�V�S5j��Uv���"�d���R��xS�v��
>ʺTeywDp:
����@�j�z���u֠܆��U�~��y�����\�4=k%Lc���4 �|�H�t�0,p�R9yUm��fꪫ9܀�ذ�dP�^�bh�,nGj��u)l�� �K�lT�f^Ck:6�� d9���kz��/r��6�ì�W��Rq�3b@��53]��m�u���]Xy�Kq�%�Q󝗪�z�W�cn,��uA�:kq�;#u/l��l�l��n6j��Z����W��3��P�V�1K�Ի�ޜ-�(��4��N�cr�jWN˫j�*��)i"M@*���O+�P��=uQB���)��v�X:ۄ��ڶ4p��`�a�s�ųW��iP�j;&P��\d�(d����l�#n�rza�;��Vڬ{MΉx})��s����t��� A1O����d�U�s�Y�9���,��I�6�:�Ѫ��R(	!��gNY�ū<�&�܈e��aN��lj�ɚ�e�5�Ԯ�6\�gl�cOen��-��t�.��wK$2�5��2fݔ�*��p�@�7#�Hj�5�������8�[�++ɩ��v�;�۶��n�5JˌG�82f����`Z�X{*�g�ss]JԷ4���VV��y���6��M�����^��]�/,Y;ay�H[$�&u�s��!��<�ī뗜�m��͓�x�B�L���@l�QS!�뮪�����W7�����l���z��v��|U�PO͢)����SJ���@�+��������҈[<���;�z�`���qt��!n���#l�l2eXt:fs	���:T�*аԠL3�۶{���M�SM��,n��k�����-c[Qˤ۰[��s���n�]Y�,:�p�V�n��-aVZ�vE+�nq�v��f^enM�M��;]qn;O.�񽽩��<�&�QyqK�� �=�6O��8J�۶�X�9P��m�ڊ��Ciy����I�s��t�*��ϻ�������o��P�n:��DcD-�v��e8'�����D�*-�/a�ׇHQ�*&{�Ok���P����]�`y{uՁ�{
�RR�FA�X����o��ḿ�e�sti�%܌l�I��b��`j������Y@=�z�f#Hk��f'���;Wۮ��=0����oz9�b��`�f:+i�"������@�����9�s��{�׀8~}�c}�5|n�.�pWnng���L�c�
��ń�uͫ���vų�-*���_�h�'*Jc�Xu���o��o�ۓ������c�ܡG;�1{u��*��s��u�h�'Js5���8�}�;�*��#j(�v埿;����/͟?g���5�H=��QQ����n�c[�(��v�7��7��v+��FJ����oz/n�W�]��{.��5OINJ$bli]F�]'X]q�c��ڕʗ�@�Z�Yl�=-׵FF.F�M���w�b��5{u����Xu��ĲzS*�EI33�_w����%�B��T�������e�V{1�[O�JILM�v��{�U�}�]^ �D�$D�Ĺ����@z7=� �_a� ���z�hcN5`g��{�>^�v��]��za`f��@�m:n@RC��F/n����/���l{,�73��Ȉ�2\��������ۭ%A��g�:�i�x�������dݨ��@X�v:Q��4����>ܝ(�n��61��p)�"T�TOf뽩�1첼�Iq(����`8�zf������R�D�d�U)Q`=��x;ܬ���.'�ٺ�T��7#�9ޅ~�s��}���ޚ���냼�\|G8����ov~�@0�-_�D�Q#�rI�!�s@<s�,����h��9�3��^��Ҽt�%��2��,ۮ�y��v�thSq�:Fv�ݺ*���I)�����}6�}��O�XouX��	�m��)'���o{���������^RG��+?s�$�M�HGfn��]�=����\�\�ǲ�s7�z�`�����I�q�����{L�2=���L�������)w��R��n�ڛ�(�n��m�$���`}O���X�\��M�pM��]+ZB;[Gb�5�Vu���+.�c�����.��X̤t�|��fM>9�2�:�����A�l�[ae����������r����c=Ҷ�[�,��]#<���\-mu6�FM�5�5ճOX8�d�������-Z�=��dF����ܪ�}M�YS��P���u���ܰ�8C7�,����x;)�d8��q�]{��������v& ���c��ѧ����.:"�u�){E���c(l��u���߻�1{u���Z(�=0�=��KxJ)�)�RI7`lc}��sw���@ncw`	r�z�iĩP�Dq9�o۲��z�`=��x<�X��Aо*e*��W^�,��� �+����	D�i�Rn{۽�ǻ�oۤޠ��zt߲�3e7$W]�F(�ۮz��n���E�e�.X�AMm�;��2�AG	6�c�s� b������3rt�71���#\�u���qӎ���l��s�s�\l�VK,�۽��5�R1�j*S�*B��\��6��P���_h��f�}��+��P��q���{w��V��V��X�2b{⠄��.���ّ�h����:P��ٷ�����a˟/g\n�k=˂+;m��ͬT3��v���Wkt'h�f����hݜ��Rr; ߷e�W��,��{�1nk�䃛����N�	�1�����g���݁������q����L��Q�&�`g��ށ�s]���k��*�ޝ��X��X��Kt�i�9)W��|����{L��w�r�f� ���7M�`�l�<��`=��x;ܬ�l]@R��/V�W�7�;K��渦�)7g���h1��f�(a($jS���Js�E;����ɥ�;��s���;;����2�*I�EBT�Q`=��x;ܬ����&:�XW=�����jJ��$�@�3uY3'guX������9ˎQ5
���G��UUR_����=�4�5�~}�z���ĉI��?$�L �� c1*YB$T!	P�!&D�� �$����Id��H��c�pG�{sە����<��8�ܻ�N��y��Ͻ�ށ�ۮ�7��`w�W*��s6��JkrD�j���O,�%-�;�-Ĺ�>N���Q��A%8���ISR�#T�J0��]��߻�1or���`cZ��}O.��IJD�������+ �}V=�M�<��t�`�Oh���N�i��~���θ�9�����V�������&�גW^y�݆����+ �ݖ}�B�*!�M�-�g��ޅF�[;@q�{������B����;�{���/��S*V۴�H^�{+�ƍ�i��gꖣ��+"h0�em�6�f��M"s�ة��jRm�f��e��<��SE���ɺ8�� $��۔ۣn`��v�%�M*��l�w9X�f�eŝ��$�H���6��gm����}�ݻ�n�iu\h�v�����۬��i�;v&�r<e��;b\6�I��AsD��_���}�{�׽{��7�z�.�V�5�oM�vq�:R,
�iP#]��T���<�TR���T�9̠5{�� �nՁ�i�
^���D�(*H�g��� <nh�'M�����I�}��}�:�&�Hn�7s�{L�Xw���{��vwU�fLl�&iL$Ҍ)7�ng��tY���vX~�/n^�����	(���$��@���@~Q����ǲ�s<���O5�][�NH�E@�v�v��:��mc�Z��÷md8����X1�7kz0ݰ����y��@T��߿.q,����l߷�l�K��T�]n>��ɥ�g(��"h!��"jj�.�O����U�����{�U}�}����]�����
�R�Ԧ��{]��_r�:q�1�xɝws-���p�������_n���2�ë<�{��t��CpQ���������T�7up�hs��ӻ��������{N�WF�sgVP��;4nNλF�GSv�yD�ط���s��7qܟ��~��{w�)f��6X��,@�j�j:h��,�۽�|���]Z�e��fZ,��PL�B�	TJJ���r���f~*�H��U_����`��ǃ���'*V�"
k3�,,C�!��b~�`��
Z&Z"
A32��bf�N� &�B&��d��a��ٸy)�R�*��P��dAIM1�L�5B�M*
��e�އ�D��c�UE�ЀjD�Щ1@%!H,��T	��GJ�I���Po� �HK-�EIM)RPĉ�.�Q	HQA�$���*4�B�wȂ/��#ׯi����x=Vac����E-5D��	P]���@P��B!SFQ;��h�*�0�4�#Yk"ƒ���Ѭ;�<�lj�4���B$��s��PO�4�U�ABR����X�f(�L
Gp>�mE�Ca��÷���ڮ�;� CY��y�vb�mAy��vt�7���@�b7�R���N	'��9����4<�P�y݁����ϲ�y)p��8��nN��ɥ��{w�,y��~͖�=�(�R�P(�vr�lF�!;YCs;���u]�}��z�f�Ͷ�Լ*�*�Q��%%)�>�iށ���@����e��X�G�0Gg�v�R����s�ȹ���{L�1�w{����U �+]~cRq��r; x�5q�3�{�wsl=}��gQ��MƆ�7s�f��,�ٻ��ny�ٮT|�I�E4��
���u#���ډ���������>V3�����,�5ҩMI!$u܍eC-��/g��%˵�2�m�g]e�5�.�����Ȳ�?6�Ђ��s@f���\W�?z����N~�6��Rn; �۲��{)P������z�^�A߹�����������'�o��V~����X�m��͖k�e*�DG)(�`w�ݻ��a��P�9�3siP�M�4L	�G�Iށ�sGm �ٲ��{/�W]���y�W���� ��^L_��6ԝs��8
�N3���\V���ݓ975kZۈ��J��{)v������h��ƚ�,�����e��ScC.�ȑE��3O�&����v˨M�c��m*]A�S%Ss;B;v-�gP9��91�kn��;]��f7ls�z��˷�9���h�n��XY���c�E;,��Y�X���\����t������7�7�ͺ���ٳC���.�r:>S��ut�ֶ�&�ㆩ;*M�&k�Wd�.�rs�p�!��xqs��j�L��~ǳ@f�Ҡ/�����z�@=��i�$���w'@�ͺ��/�w��-�v�e�����mD����f��x6Z�`��`k�qjQ��-���M&� m9ށ�w]�{Qs�t�, �gw��H��**RU"UR�`3��^è�3���~�l���%(��m�v��i;3
��Ł��<�kmːLdvz�q�P�T�U�W�Ϯ,��� �+ �۲����T+��"�)�	%X�}���y����������9~g�U�~��m�l1�?�$���������h>nh�6�kw`�)�Zʈ�$"r; �ٲ�x�ڰ>{��b�o�y���&": �ZJ����>��37����+ f��ܪ�줷��"))
�
rW51r]V���V�kՍg�ٴ������cnv�hl�"���߷��� �ۮ�>����$���33S*E@$���o� �nh�6�����D�F�T��q	�n'�o۪\H�{��O��
������z몱n봑��f� 	R$��u�'@���s�a�����>��)�D���{۽��5ؒ7��`{=0�3�j2����Q��#H��q��'a��Gom=9�Ƚ������ڮ7���!�		$�@�x����,�����{��c�Zʔ�6ԑE$v��V=�Xw�ހ�r�݆���ƒc����N��ɥ����{��\kV�����X����i��@���@ng���h�۫��I"��@����~�*��,�>6�%�;�1{u��ʪ_����ܚX�~���H��eHܩ�软ZW��Ŏ CZ����{.��a6�m�ܛP�ƒPC�i��������/䅞��ow������㸂�
���.�}���1�)lA�݀�u���e��{
�TBA��`g��ހ�{�����V=w�~o%ME#��;�1{u���,1y{-{۽�ǫ%��MH�E$v�n��؝(�n�&7��h���MBG�7w�B��ݦ53\ڪU��F�k�[\r�A��/w����^ـ;'Sk�6���ܻ�X#���}�g�~&�9�d��9�+cn%eMu�v�XCf�(�v�)��sɎ�4'�:"c%K�X&4�h�ex x���kt����b���ʾ�Ni�y��c;l����猓�9v&�[�����v�T�`2�V��=�<糣[r�������<A�b)���w�{ݽoZ��Ef�Y6H	�z����h�-Z;u�ێ����{v���?s?��c���$�:�������4�3���@���a��rΤ|0�
Q���~�����{�d��XguXA��Ϻ�v$m3hQ�m�(m�ށ��k�c�ص��7��9=��S)*	�&�R���`{��ow�:�k�=�V�D�%H��m�ө}皕������Xc�=�ԓ��[5��l1���-��=��2k;����K\�lN�=���v��1���|��݁�f����S��Ir�>������"RG�H�� �ɮ��(x8�L���be�{�uʽ��}����AZmk��r m��q>�hF?v���t�7����}��3u���L���J��x�\X�{��>^�v��]�t�ň�M�$J�*,����w'�U��ޥ`{6�������o��婹������=��vݭ��7:v��utj��ێw���m�ϴp�¢m'(m����]����`w�L?W9Π�g���_��q���n8ۍ�`��|�fL�5̀�{��2'{���㣂�%"Ln.�hy�>���O��M � �z}s7����WY���;�e.$]
�E)H�V{߷��2w�E�ӝ���Z�������&II���;�>^�v��]�ߟ�X�n����ն�I!�Q�8AANf��i�[<�=&⁮�M�1Q
�{"ێGq���~v~~�`g��N���]�{�R�m!�%�v�>���M��_�:�X�_/l�h�Z����RD����{uw�|���j���b��Z�;���k%�&�r���q/ܪ�=��������ߟ�X^�S��S�W*�)rk����~"M��%"�*�����ұV��7�����`}��ojA%$��c�D�D�M��.h��ғl����h��0	C��*]z�H�(ӏ���=皬�۽�/n��r�����vٛJ�tD��nE`<�ç��or���+1k�7�ekh�Q7$�I's�jǲ݁���`f-s����ؠ���	$�TҥUVN>VjnU�<�����]�XG��#XTI*q�;��@��5X���}��6�H�6�f�G������?�K�s� W�?�?�F/�f��op� XYThQ��*J��R�ҨĨR*P � Д*R�	*��ЈЀ� �R
҃� �@���ЪR ���(� �@�2�4*	B�P�H���B�Ш4(@"�(�(�(
RҠ:�� P5$�
R�JRC( )JR)!)JR  K*P �@�1DhA�P�8hܨ�  � ����P�U� 7  �(B��* PB9*��)H
(#0� �*P�H�� �@	@���(*�@�
R��#�JP��@ R-�BR�R�J4
(4
�IB(ă����H�@!@�% ���ҊҀ��҂��H3�gu~��  ���)G���_������_�b���D��*�P?�k�o��Aڧ��O����O���A?�O�������?���?� ��x��������D�������������QW��(�E��������r((���=h������������x�!������~���ځ�jo��AE_��Z?��o����?�����������<��=�3� �������B��4*�A (� (�҉0#�#$
L����##��"�(2@���#$��(�Ȍ�#$
��H(҃�%4*% ,JB��B�
���D��"C ��Hʉ J�   ʉ�J����@JI!�
 �HC!H	#!*�C!��@
�H@�H!! ���,
)	�!��� B$��I!$�J�H"�@(#,�� �)
Ȁ�@(0��@2�) �(02�2"��	���,J� ̋�B� ����qd	�@�B�$A�%�  �HBBI	���%aIP�@��!�!�%�!e �%@!YET�  BB�%BP �XBDdP�%Y�e�!da��  �!�aaF�a� �%�eE�!QaPRP�`&@�PHB�eUa	 HFB IB�!� AV�� XBU� Y HQ	F�e�$��P�Q%$A�	FT	e	B@d�aaYFI�b�eda�h@��e�``X$IIF	@�F�BD�TaXJUJ `PJP �@��TI� �`Z���o� "(�(^������y���������O�~E���ݭ���Vu����\������|k��

*������ ��O���ֿ������PQW������"z����@��s�a�wnUx�?����oA�>��T��k����\�������������������'@"�������������_�t�((�������������3]<)��?xa���������g?�����~����0Ǘ��((���K�+^d?���kD�!�������~���^���U���������:Et������ω�������PVI��c
�� ٘�` �����Zs�   !@�     �{     �   ���     R�
����IPTJ�	R�P$R *� AI( P  �  X   �d�
 �I R� �R��Z\Y�9ɾ�X ��r!��b � t��Y;��x�x��5���Ԙ RiM��W��].{ޕ9e+ �N��km�s�;���y}*�  �  
QA� r^�(���J70 "  ����(9� '@; ��AFtL :24 1  � � h����=@ � A�:s�  40tb vt�S� A� � 
  �P�@  �ɽ�O.��q�u�x�t���
W:zr��95֜�t�']' <�t=ź�۽�u�W�R��g�S��ꕞ�G���
��{��>]^�n� �J�g]�{�����}��}<�zׁ��� P (  � �w}��]:�w�ת�m:�����Ϡ}����ũV�t����t�� ��w��e}�gx  W�s�{��|�>�y����{�7��n�z{�׾�� ��-Jnξ�]�wK��M+� }	  @	 I� ϯ�㻭.�s�m>MU������ 'N��t��N�6U�/x�){�6{��\������� �/}�/}��]� ;��n���u�Z]n,�� ���q����9=vg}���  4�Om)R��  EO�CSeJT���C<z�U5L�T �Ob�Q=&�4�dh�%6JR�  ")�����
����?�_�~����T�:v��D�DD(��.��*��
�
��*��ꈪ*�pEQV
�����t�F�����$:2k8�Z͉�!%5�|<��Ù�hjblH%4`�ҁ$Y����.��c1"�D��F+�	GC�(h_��l�V*R�ͤ��1v��Ǆ$.o�44@��o3�5�l��B%k�7��Ӂ���L<��R}#tN8y5��Y�OCłSV�4��<Yg�5�e�6{p �N�7D�24�SDq ư�5�u!4d7����k"�XÜ߇Ck
h�r��R8i!)�7Lу�(Kpד2T�IoE	K�o�)��%���Y����FZh�K��ֳS���#�,�x�x�Z㰅4����͛��� IsA.�L8��3����MIɚ��a&�"j�ZR[�K�
kw���)���3.SF��*Ku375B]h�t:�.ao��p/��<5,�}bk ���R$b�����20�=@B��Yf���#@�N��]F� �B�M1�ZhX�H����:&�)��:HЃM3[e5$WE2aR74��.�i�k�%K�F��+�d����4i`P�5�e,i�6�0�莘P�Ѥ�.�SF�$H��cMj֦�Cn��w��w�y�K�{�����7�����n�s緟o���i0�Z4CF1�!�h4a�.�T��fl!t;6LSLn��6��ŀc��jn���6���dtP�A�����7��Ei5"n�b�=�>����/ov��y���S7Sl-��O6x�XQ�"D�Յe�H)��j
b@��"�X�y�2�RHRD#�D�ul�� h�%R��,�!
�HL�T����XtC �a���1J�HD � ��<!WDL
q�G���!2C
�R�j�FX�4f�n���4Ą��	�4щ���zxa�i!$*A
�����f��k9O)�,��9���$��mYMf��Ä:���
��O���eT�'�WQ䄄*i��|�I
�3��d��R�б�ޭ�1�$ل.�$�ӎߞx�o�xq���	d4F���0*����b�T� �cB%V!$�x���{�Bk	�l�y�)�����L2:���+ �*Ei��i�����$���{�]`F�=|��D���!(DX�H F�!]$�_}I�i��5����<�k����D�z� ��V�A��1�� ��iHU 4�*EH�i�`$ 1H�K�(4 qYR�OC�Ȱ�	�*,
��&�%�	-�!�)���Y�i��t�Z7�|�a��Id���a�V�1\T��U��BYX�D��*�8��"F���+��� $FD"�R$B$B(�"�����*� [�ɜ��Q᧎NR���;�1�j	Ha@�0#�D�M&��,U��!X�XR4 ��(�b`ՈHz)�=f�SI5�B��	.h��g���a�K�M��K�1`����.�!u�ĕ�)�X��)%�j�����B�A
h%��ێ}���޹��=�}�}�m�nϡ��\�����GP���H]�/��_����
i%3y�5�]���5a%�Z	��ټie�ލ��ћ���/������B8:\�7N�K�r���O-�bD��JH]��K�!H�D4B�i��!H]XIi���)�h!�'�HP��)�SDԡ�Ɯ�MRI7��4Ƅ����to��j$a�)����r�|��Ͱ�����V0�3i}nF@�6��7�)=e�<"�f5ӯ&�!���4K5��Aƚ��a�o�|%�����Jk^s!�͑�Ne<��%5x��[����l$���
`�n���HhIuLB4M4�dd�����]c7��.�0�$���M��F4�nF~���k\��Rh˳�5�l!tT�.�HP�Le4ρ��.I_8�4a��0�'#!vRZ"(J�\�*��ǆ�S���ykggj�)Ҿu>��K�]>e�Q��U��P��[�8Wc����%��]���_R쿎O����u.�����v}N��vA\Ns�oT�	�ٗ=�޼c��e��ԩ|�n���:tv�I:�����QyK*�}/��̮�o(T����4�g'������8y��s0�@ķ_i���\C���]xHO<0�
xGZH�9�E 1� H�xÌ*Af��I)�n��݄�>W�|dE�X@�d9,���o�_q�4�f�@W �a(˒�=��<6�p�bP��� H)��k��o���#K��6B�I�d@����	u˘L5u������x� �B@,�+e/�m��)o���g��0�#�����@�*jF�h�G1�Y��l�53�!��)���ѽ�aY��l��h�FmaaN@���.�jcH��)��l�.���Ҟk���{�6�cu�3G.�R��k��"x�<�a�Ixk9�e�Nh�[�6]0�$���$"H2H��RF$��B
ViS�-щ��K��H;Ha�B�5���)M
;$!��SK�JVҚp�$1!Hj@��!H4�XB�fn�-4����HHԔ��X�&�RaR	I�062�o@F�i�"�a]��],R!%�N)����%M1J
$��	���Qѥa��i��!M4!Zi�ˠ��)�70�.��0�R
$�"� ЃX�ӈF����$�E44 @�X����a]nd��	���Wv�
��`�t!�/5���4����a�7J�V�$1�������sM���Sj�f����Y�lH��7��M�y�ىk%5�y�\0��]k�0�<��oo��M�1�۱�cM�<!��o��!nhv�/��������Y�8;|7��BZE�CF��Jj��SA�Ԏ��_5�m5�6�kY�.���Vhf����ɛ�n˫��O7�` %�5���0�2�GRl�v����	B�`�og�.������,���:�<�m�Fj��;qøKټݥ���v��5���)�'1Iti��5�]�!R���F��éS�`X[�0�0��!8B�h���]7W5v@�E.���WY���۲�H@M>��͜˗kN,(�s\ގj���G�@`D#4}�k&�p�0P�^��y�^XB�c�A4�i��7�y�˂��	LW �#�G��$6�H�c�P�$�
��[4pR(A6R����2�LK�HVRy̾oƐ ������Q7�<�L�!h4e���5XA\!� �@��4�ňU`T���$�q�%BHJ�5�E��`Y
h0�4�5��хv�Z���
�V�B��#G_.�I5��p���x1
�*�I��-��!٫uo���[�`L���z��f��,��!�M��"E�a����lo����&�%�ލF��]NL��h!Ii,k�P"GX�*�"膴tFD"�'�V@�a"H	 ���f�I4k�Y@�9	JD�B�Y �� �B
����B���JM�@��������������a����c.�`��1�g4���w͞]l���%�2�l�n�}�g�]�����?_�H    � ��  �`-� � l  K�G��f|�FHz{5շW��֦�.��U �1ّ����2�6`�vum���ٰu��n9���K�\�4���)ඌ[�	2�uh�nzAe쏛������`6���$:,��U�T���T�E!;9�t���D�vͶh��'�-�r��� &�Ԁ�mm���KH�Ѳ݆�ٴ\�l�p�/����86�E��l�%;p :�h���M��X�  &�8T��n<[d�  À   m� �m�m  �  ��!������[@ �    m�L�      �    �����I$8�m p    [@  �� m�m �$���`    m�     � ��n m�@  ��m $��� H   p  6����  ݶ��z� ���m���H    [@ -�.�X�u�� h   �� �|     ��  m���C���	  H���  ���l��   $-%-m�H�i�%�     �    l��Gkm�0�@A�� � $p  k��-�   �kXu�����'��  �� ��m8�����*��F�$h�΋Յ�mm�  ���m��Ia��8*�j 
�m��͵�  l n�L��m[�m�8S�tIm���a�����7n[h��M&��'P  �� 6� m�Y`��[��8-�l� �K� 6���m������  �z�V�h���J  6��L2�d�m�  N��s��6  p6��[f�-����WK��[@�>���7�;e��plsX;&]l�Vu��]8��ysjGXm��I���mU[P�����flv&( $Ht���&�B���k    %%@��P<��9�k���N �u�[hA�l˖{u�)Cb���7\l�t���p}�'o�����۪2-�Z��.��6�P��B�{8��T��l [Ctu�,Gn�P��[`�Sm sm�Z��m���� z� -�Ӧ�gm>�k��n�@`*��qD�ڎ���X[M�޴6�n�
��d�c� ��	�Udˀ $�e�$-�����e��U-�Mu���9Y55�JHue�]�]��]�ڪRej��qr�]���Ҁokm�[EӤ�b�
��l��U=fͶ�l闦�=;ga�.�E�5�����߶�k�R�Um9�5_��}@��evj�2�U�]!�m I: �\lq��T�r�!�`����YD I��Ku����  �]�g-ȼ����ZN� Hl  ���� 	v[��@ 5� 8[[-		i�� ���/����VV��Z���ր  �       �@K����;���&�k�,劶�    h��   ��@ H   � � %�[d�o'GH�G-�M\�� � :<� 7mmÜ���`z�e��`��f�[6�����銳SI�&�w$Hm6��z7eZ����z�^8�[��*�5��F�Nm�)�pH6�zN�'Yf��1gS� �����^�߷��guOP�j]�^]��T��<Hx٪�\e]us�v�h���#�ŴU),l4�X.�j�mm�-[%ss�$��I��[���]/F�� l�if�p�Ԛ��m 6ێ7l�]9���ɹ  [8�vں4�֛i0��g��8֛cm��l��8GN���9m -���l�ZYe�N�:�^N�1������X�ײmwl�$��9  &��A 8�8k��      J��nN��.��k�z�qȰ{;l6���r���+��lur�WU�6��M�k�%5�� �\ϗ/	���F�m�{*�]5��m��@Cm0�8�@u�4&���6�m���}��M�[�`rF�*�j���7_����@@V��f�aY��T����q��5�-ڶD�m�+l�k'P�zY(��jٴ�[4q[ =rkp�9BinY�� �U����kiS��]GgI�����O 3� �P的�Sut��\�CAU��MKkm��U�R��i����{l ��X 㜶�7N��[�]&��bv׳���� *�\��u�������`�`����p�n�M!�J�1Dn�E�h/a�9"�40݉�:��+�q8H�{6�m�[d� ��i�'i�k37V�6�g-�ʅ/[UmT�r�v�t.�q�5�� ��貳+e��1)ުU���;��U��6)g�Y�U'm`B��KB��] �j����^Y6�d�@���I:ml�݁�nݸ l��Ͱ9&�o�>Y�8$�׋T��E�Qmm�	����e�J`  	��i2)y$�l�����      �� ɑ[Y6�2f�d����� ��3U�մ蠶��p Ku��� �m��]lI�6�N����� [A�� 8 �  -�    �-��@9D�vp�m��sr��zy�*�ک����j� U��U*�۰[%�����8l �@�ɭr�[�n׭�9�@6�q�l	4Q:  ��m� p8�$֤�f��UU@l���tV\<��T�)�<��UUU�U#��`)*�����t,�@V�T�[�vj��ۗf�*�)v�eU[m�l [@$��MUp"��6�2�@*vI@�yA��!UUJ�\K>��5���-H���#<��m���m����6^�������-��  �pl�)���e&����4hS\��v��{F��@9K6�%k��Җ�'� ��cvq�܇ I[H۶  	 �t�ns��Tݮ)Bښ͛`��'�a���T�m�R���v��;l$ m��$��*�IjU��k��Xd�hm�5�� 6�k�6ݜn�9� ��J���Ѣ���T3��;e�-�i����A�U�@��   �kz��.��W��R�o�|��� �`���-�  p ��hm��v�h0[I9��v[�� ��g�m      �`Hp^�q�kn��slv��.��&��ì�$H���@ � 6� �lH    շ���Jlpp[%  ��p �fݰ$kM����A&�g 6�&�� 	 m����-�jַ!�.�˛��N��9t�$�ôQ�$[W�h�ڶ  kn��!�� �  	8[&��� �n �V�NH 9,5�p�Ok��0�&NK-UN��� �n�ll��5�` ������o����N��H��}�ʵr��*�8�am�ne�N��Vm�<�Z-���F7IKR�+u�H UUT$t�:�[Pm�f���� �n  -��m� 6�� �"�����[�$�h��m���`  ax�d�m�m���JP m�݅��p H-� �Cm�6�%��     � ���m�� �m��֛n�HĜ �b�	�m�[@m���6^��V�eg�ʪ��P@$�j�s�v�"M�L� ��u�$		�A s������  'Kiņ������� m��8��	��:N ��ځm�l���[FYV�@p�ݻMf�  ����       [A�nU�i� p �$  s� H�  [N� H  �`������� 6� �Cm�m����U-��À�v���Cm���Ŵ�MؖYz�궤 �~��� ]6�% [�[@:I4uqm���{ж�@p�� [V1��l�-HH�j����mu+��ck^�T6�1v2t��*Zf�e�`az��t�5�I�����8)ݖV�5�:�:�R[k�lcj��� ��  �4�\�I	�  -�@-��           l      ��m�     ���$];v�W�6� $    � 8   ��   [@ m�   �  $   �>� h m�6� 8 ���   8A�M����M,�Kkm�l #����6Z�k����Դ�h ��hK*K'[&�   9�s���O�����GD2�cD�	oUK�o�Ny�l�;�l5��訠�@PG�Q"���N�� ���}�oC`�A +��0QC �D��T"�*���D5�6���Dh���`	� q�Ȧ�T)|��v&�O�R8  |�� χ��] ~O��⢟z^!�= �@*|)�x(�� jDU}b�Ă� "�$P���Q"x��lP�|�t�A�@W�G�`� ���< ��U����|�)�P��<T��TĉF+H����0�, ��� D�H+"`.#����Qv<B�T�Pq�|�ϕG|�>@�v��Ea���(��|S኏��@Qp�8(�N
�	#D�T p�
����v���F"f��A8��'�D ���k`@Z�&�H2K[%��/v>�����F�@}�8�5��_��Q�b����TUҏ�� �F z��D�������[�/N����#ӭ�z[�֬"�Z�`m��k�`d�s!�m'l'������	��kc��-��;9BU35*�*�PE�.Wj몕gd�W���B�v�A*��qL����ԫ�P�@R�$u�U�I�m��\�8�;&-�z,]VK�&�5���Ҭ�
�T����l#Z�L����m+�6�(����c_X��֋�bm�	�Z��\����pv�;˯D��7\���@E��.4��mH㜻i������Y�qbv&�J�OO��D�]��ʷ5����n�ls���{Hݸ6��:Kv�F��of��kvȯg9j���h��؉��:��= j�� -�f�7%����T�f]�f\�\h��pV�Su�=/�t���V�n��ݥ�3[g�����2
��تxv2�_B�����Sd�=b�1�`�S;K9Z�x�kqt�"�e��D��t�E�Q2
�F�ی�j�[c�/vG#vU�Tdi-�ڴ;��t*J��s՘�٬�����^mz��t��Q�;s��tYֺ�+Z�˩���T�ۅ�. �9�&�Ub�[���ᵜX�����bL8[I��bβ�n�VA���;M9�3��3�E�q�b���g�����SyGN�N^H���f��1�
��W-���\C���cӖ�(�1���A]5�B��w����v[�6)�kԴ��u�N�[d�M��ۑV�B�U]�E�-'8�*h�m��ȋ&:)3"j&�6�4N��M<��J����]Ҭ�Ѵ"�K�/[ �%XӤ��R�@ګ$W,�a�U�^vYc���ٴ�+�ї����z&��s���'�pg���m�H&`�S@&�쪭GOk��.�����-�I���\cT�RPP���!��G-�: ����g
�n���-��m�`-� -�{8$��YYZ���T���
�\6�Χ�����Ѳ�������r:ID��
(:5"������:���Pv(&�}b����r�vh���֭qd;��:�3��OGQ��P�e^�L�u�"�/Z�VV���q<�8	3v�-N�ɶ�z�����ݤM�ן+�{9;!M`vђ;p<��g�(:�#9ヴvSkg��mh"�k/]r����ڗ��6�;%��]-I���g͜��	�����l�l�NS�\���Klj+� �4��}�{��>�w{��{���ǽ����~�o׎Uvxy�{yˌg�m���7e�����	�gv�yO�Q�������=�j���ݯ�Q�Cg�� �K�����a�����_����*�5g��[�;��U����ㄊSq(����@;�1 ��Lr�T���4L*7Q(�5V.���G d��w�U�ٵ��wJ���71�@tqR�Ih}& 3�)�
%*1D�n&HD�
�ň�\�/Vd�<1�S��v�V췎�5\d��Y��h�*@>�- �Ɉ��X٦����pCRJ�3�u_k�8�����<�+��M�>�$��{�ܓ�ݺ�;��R���s���`b��`t�-�EH�%�=p!R����r�"��ך��\H�{�V�����7]��u�ȓ�����X�*@>�- �Ɉ���V\��nz۱���F��",�M$k�ܜ�����Z��kAsO`��j.X'cw�d��v��Lr�T��c��Tn�Q�j8�]�vu���u`g^�1nm*%J���HMǀyֹ�<���a(�IT
$�DeWy�q��{��ś��$��sR�@�l�P������ʹZI,��_|�X�n��������$�M���pE4�E�������%�6��I.��_|�]ݻI%ޛVi$%"�"Q6��mhx�q7��K�d3���1ض�3cM�RpV�bڊ78Ȝ_|�X�n��������%�۰��Yٺ��$��ҵ1F��L�IN�Iwfj��r���޻I%�=���%�6��I.��D�T�84��K��ai$��u}�Ibͺv�K�3W�$�vV�$R���$�ZI,��_r�}���[�����ל��6P��9�/������(�9�w|��InL�Tn	4��q}�Ibͺv�K�3W�$�wn��Igf���0�_cJ�5�݄sd�{h�W���p��&,���K6B�)��F�l�ڎ�V�\ae;I%ݙ��K��ai$��u}�Ibͺv�Iw6�������������ZI,��_|�X�n�������ʒK+uIB$��iȋI%����KmӴ�]ٚ��$��m�K�D�-iJQ�!��$�\�={��I,�ߏ�I-ɶ�I%����I,+Sn�����$�vf��I/W9ʯm��|�Kroo9m�_~٭�m��!$1� Id���ĄB	,X�`�s��9ʼ�A�nS�QLj"q���z���^��mN�4����l��x��������m�c7˛m؂��ƌ������;%�;K/S&�ۤ_E������-�Iܶ���\&6��/d�W3ͱ&��������w�{�q�[9��v�d�� �5��]�hG;Xβ8���5�9xwl9w�v�-�hI�g���SRn�\���e�6�.���g��=�Mk+i�����e)��]��S��O۔�8]4i���X��Q�k�Ex�^��E�������%�6��I/�f��I.쭾8H�))F	&�-$�vf��I-Y�N�I}�5}�InM�ZI/�3D£��iF	�"��՛t�$��3W�$���E�������%�v�TC��)	�N�Iwfj��ܛh��Yٺ��$�f�;I$��Kb�EIR*�/�I-ɶ�I%����KVmӴ�]ٚ��$�Uz�
��bQ�6�J\T������n��8�<�lk��V�],�P8�"$n��E8�Cr#�[��_|�Z�n��������%�6�i$��Lb�M[�kX�j�^r�~���[|x�:E0O@�G�f�o����-��s�ٻm���j��KJ5����2E%;I%ݙ��Krm��Igf���՛t�$�rV�"R*N)M�"�䗫����i$�'���$�f�;I%ݙ��K�+o�)JJQ�I��I%����K�\�y��$��M���ܛh��]��Qz���sȡr�w�P��v��s�H�����%��
^�xژ��-�	�I�����&��Iwfj��ܛh��Yٺ��$�f�)D9�!R�����]ٚ����r��6׶z�i$�=~>�$�d��I%��["*J�P��q}�InM�ZI,�ޜ����Z  |�����nkvԳ�5}�I*��\n��58�Cr"�Igw~��I-Y4v�K�3W�$���E����1�ER�s�rJ��ՓGi$��5}�InM�ZI,�����%���Eԁ�7�!�r���Nb:�q�%�q��Y�R%�v������HKg��P����5}�InM�ZI,�����%�&��Iw%n��EJE)�@�_|�[�m�K;��}�Ijɣ��]ٚ���\�)��ҽ|p�JRR�M�ZI-�{���ՓGi$��5}�InM�ZI/�7�0��SQi9_|��)���v�K=7��W�s�ٻn
	�`��17��߇9m�-ۥ"�T�$u)	�;I%ݙ��Krm��Igv���ՓGi$�3Z�@����ϖ2��ݜ�n0Ɯ�.٭�Cc���ܜ�v j�v�(�n�c��1��[�m�K;���$���;I%ݙ��IVn��u�Ɗ��K;���{�U�q���xv�K=7��Krm��Iwh�Ţ�)J9�8���%�&��Iwfj��ܛh��Y�߫�I,mh�N������]ٚ��$�&�-$�ww���ՓGi$���tBEJP��_|�[�m�K۞�k�I/-��������%���V�	MH)J�MH��vxjd����牞I�=[�lj\�Ѯ�jx��fdn�i۶*�n����x���:,k	5$7	۶�4G�������[��`����4���}��Iv\Ặ[��{vƗe�L�������d�%ۀ貌X�"΁�c�\;;��@@��ZS�È�,vڞ ���ɘx��ˬݧD��6�v#�;/��48*�R�Nf��E��jj�`:4�������?>��1���s�`�:
^�vய6�JRR�M�u$��߾��I-Y4v�K홫�Krm��I}��1�F�*j M7+�KVM���fj��ܛh��Y�߫�KVm�$q%$�:��$�~u�p����Q2��,���]-��"����7�5X�۫{�K�y��>;�ؙ'"(n\��x�Q
!.ל~�O� ~�j�>̡�+\��17IҔT�nJ�&�:�=g�sN���=�R�t�-fy�;���ŒS�q�XܚXk�V��UUs��|�����N���2D�`s�{���.��*H"$���
"�$�E���8�k��m���D$T���	E`o^j�3�5XܚXk�V��7�)I�Fw���}�Zs� =1�@N�-�f�n��Ӑ�7�4�>׮p��8����
&�NO]YD����M!h�6�2�Zngo$��(41v�ƘF�H�Ʀ����[����2}h	��8�9����zj)��I���7�5X�۫{�KR��X��D�Pl���X���7$��s��<v  	�U�z��+��(Hh��		p9		!�h״R�}�$]��"����*-�bCF,0��HF;����0bF��T����0D��*:�q��@b��D:<ҟ*>�i)H�S�~�^�v������Z(5)�8��W9=�8�=��p��8��}�`�/���ܤH�,���^ɾ_ ��,�m�Т"H�.j�U��VK�'sJV�5�v���7���u��˞x-��KF�
IS��B
P��_�{�`gsn��M?|��{�`wη�p�Jn�n�fj�p��Y�DG�Gϯ� ߫��z�U��f�7H��T�@�nU�;��9h	��8�:lvD)$qԤ'"�>ך���Vw7f�ٳ�4>� �
!�-���rw�	Lj(�>9V��+��V��V˸��'X�8� h�#\�U'[�A��#W쁫u:7k-��.4v�H9�A�r m�`osn�Ǻ���q�p1h�ԧ噙�<����#�- ��p4�IJJJRr+�y���nZ�� 'd���ʓoJ0�2�3v�㖀|�	�%�=1�@w^�Q�)��`�n+:�U��{���^j�7j�;�WZY��n��(9s;��;�N`�s�l)3��X�b��q��۞�{x`H�1���3kX�
��r�m�ܶQ\݃��.@�t�q��vjwNҶurm�s��^u�����M�s�w^$3���m�*�@�.lml�����t�K�G_$.h;Ƌ�8�踫���۳����xҞvo[�]�ݍ[��ܠ�ܗl����F�uH 0��nD#m�r���E۠�BR�(�R�T���f��v�_o��4�ɮ�d��Sq<���jբL�t����ԑtc������`n<�`g^j�7�4	$B�G%mYy�hLr�㖀}�ZvIv��[R�܍���qX�5X׺���Vu� �Y�H�Q�d�����}6	�%�:c����p1j�nH��$p�7�5X���/��=�3�4�7�F�N�H��\ܕNgL�牼���3!��%�/Ni]��6�Y��d�(�7B�*)��y��~�� �;gDD%�C�>�].���JP��V�T��٥���U��y���]n�ԑ�n� i7��v��k�:!D,J��z�Nη���7n��F�!����,Y����'d��}6	�`��w�����Vn� :c����Z�� "��`{��[�Z��R$�BQ����PpωeĽ��,)h��ˇҬ����o�Q��Q���q|��������ՙ����`z�����1�r nE���	|� :c����Z0ǂ�܍9�H�`j�k�;�5XV󔒋P�\B���k�|��)�9���
T�Evu�z�U��٥������:ݧR8(��T$9���s�r�
{���:u�`u�p����7�=n֍�(��	�h��Q��֤8kn�c�����tq�������-�e�f߀���@K�1���r��v�D�R@��!`j�k�:c����Z�� 'M�n�����n��Y����Zv9h�*@K��;�Kb�R�:�+z�U��EH	|� ���������/Z 󹣑9i)ȁ���ͺ�5fk�>ך���Vki��A�)H�D�S��<�Z8���{I8�7Q�[.�q=ܵ �	�H:n6��#��Y����vIh�*@>�D2��(���4���ZvIh�*@F�7[��G#r��!Ȭ��Vw6�� =1�@y͢QF��wFhw���|�o`���-ߪ��}vw޺i$����Mʰ72i`zc����Z��Twf���ۇ>+�6��e\�n66q-���l�tg�I�mn3u�T�����u���۵[z�;b�c��rv��#W.���S����nB�`��㳍$M�L��<�ƶ�[Ocs��R�i�Ż�n��G��;y�;<���N鲸��r�:9�`0�vN�����H�b� Ba���I}����lzn��=Y4�n��լ��O\�����{��~>�iu��s�<���Ll��eun�M���6�*V�f�0��% ��Q'$��Q�t��+z�U��ͺ�72i`uwtN(�!���ӛ�h	�%�8�� =1�@՚9�m�97"�3��V�M,��z�U�ݡ�Ƅ�79�i9���'c��|���+Y)���������`o^j�3��V�M,Y���Y$�JEY���X��"N��p�ZƬ��͊M1Z�s,�MT��G�R��!Ȭ��Vw"�o`���-�6�Em���T�U��o�$@�$�DD�!P�R�P�_����`���\�f��R�(��r��M,�k�>��=��p�ذ�l�W77y��vU���Zv9h�*@ori`|��'r��QP���7������k�0:�8Z��Sf��Zƈp�)x]rZ4h痝x�l��M��[���U@��f��G�e������<�o��9h	��:Q���8�A�{�K�9\�$g��XǾVwf��Hܡ�Q�M�5)�MY�oS���\�p�*P��!]��������:�a#��T�(H��r��T����`��M�QQ8�*��Vwv����o��g�x�>ך��j(��pmJt�iNV�4E���Ҝu������Nn�)�inSu�b�rD�Si9VfM,�M,��;�u`gwn�GQD��RE7 ���	�%�H��/���~�Q�ʒEC����?yX׺��U_�߽���7�����^h�N"�CNEa�U-��+wg���K
�M
:X,����U )��G���s��'�����hNs�jE`fd�����U����g���3�uX���aR8��@�pW9�37�.���&g��;�Z�R%�r�P�U�TXԦȚ��G��=�?:np�7?|��w_�Ҿ�>��R�IBT9����~�W7��ݞ,��W�r�#��G���T�`ɪ���t��l��ES����7���`}���rD�SjH�=\���� �S��?:np:K�}8��AwTH	��D$���^j�?s��\���.������� P�G�
V�)	H��t�0R,B '�ځ%�ddc5��"4"�P�ՌZ��K!)+
1�("�%����k)(�a� !R�6��
)JB��i�
ĤHH$1$a�x0}�Hp�"�!��i!B) ��`�b���<q*X�X�"�	�ca[��!A�!0d�(��"��J'���N��9���!oFz}���+`Chԁ8�R5!�IUIAH�E@�A�F�� ��Z�Z�c�2�p�Ki�FG�I0E�1	�kD+"0`@F1H�"�H���1!^�kR�̄R"�!u4�zzI!����0����f�I�$��Ja��z]g�k��rʹ��<0;���r82D��ٹ���=d��n�IEW[o�;���BU"�]a����]uS���VU������v�U(�ҩ�[W[���0Զ�� H�[-ć�����ݶ΄�ͪ4�,�%uf����]��'DL�uMn�h�:t^�l0�$'RKuJ�v�����%[���4��ec���P(i�5Ƹ]˶�B6�p+p�n�YZ���E؝�n�s�L�ۍZf��{1�=r%�h5���'.��,�pt��n�u6��Wc�pqλ{v�:Yۚ7�}��?�n�Wg�`�ہ��m�@ ��m&�Kk�Tam �*�l�np�55��z2wɠ���I��yܺ�s˱m�E[���b�ti��[m9ݤtl<�]%�K�8�WM��BP�Ѡ�ݭպӱ��Vzr�rZ���(HJ.٨.��ޙt�֛ ��k���m�s��y� �n�v��Í��G�cV�n��ln�x��Ŕ)������zNV)\Z�3z�r�՘8巳���=lj�v���8�Gl���)�μmz�X�q`J�M��ն��eԻY�9vkf��U��dϬIi�Y���Z�1mt!�3�Fi�w\E���M�N�5�RSg�vݘKy����mւG��h�ˁ�>��ɶ;f��u��6�	�Bm@��˜<��ؙ���ugA��F���K�v���`[H1�i-�.XLA��Q�����]��`6p�Z2��k+Wl�% h��c6x���3�&���OJ�kvT��^�Ͷ�k�����L2�waW�]��UUS��Pj-]Q��ɭ���bKv�ISh�����I1�_[y�"�[mR�/R�մ��Gg�+����Q�®Sn�SJ����Ge)�/C�٠5!P�Xu�+ �������m�Z� -�v�vj͛cm�-m	� m�ݤZ9���D����K.�ana��33*t<��1QNUGD��*8�uQ���P�J&:	PTڄT�fq�%���Z�(7E��d5�Ƌ�˴tZW����k��׮[ `���}����l�Y��/G#Kv���N�s�`.�k��gc�O+��1�{c�r��#3��glOnn �4���(fۃ��tk�+ƶ��wC��]� �է�]�n;gm��-�:��f���!���Til�P������K�����wg��ms/\��շ.��-���r�NM�(��]�@�V�t9z����\�Y{�Usv|u�Ӏo�ŀu�BK���V�~��$�B�(nE`gwn��_����%���ͧ"X�%������Kı;�w�iȭ�bX��&�^q&����U�9H�#��R��siȖ%�b{߷ٴ�K�D�Og��iȖ%�bw�߸m9ı,N�L�'f�jj���D̹�ND�,V����nӑ,K���nӑ,K�����ӑ,K�/���6��bX�'�;���k!���-&�.ӑ,K���nӑ,K�~����Kı/���6��bX�'�ϻv��b]�7������]`ps�p�\��m4��ϣs67
�ҋ�Κ�c�Zl�9�ӣ�T�JԚ�Z˴�Kı>����r%�bX��ϻ�ND�,K��ݻND�,K��{v��bX�'���m�&�	I�B��Xm9ı,K�g�ͧ!�@�?*So�<�b}��˴�Kı>�;۴�Kı>����r'�CK��R9_���$tH	��#$����bX�'����ӑ,K���ݧ"X�%���w�ӑ,Kľ����rr��G)�y�	����*!�!|��X�%��s�ݧ"X�%���w�ӑ,Kľ����r%�`~&�{���/���G)�r��������M7%�r%�bX�{�xm9ı,K�~�ͧ"X�%��~�fӑ,K���nӑ,KĿ{�uHwXj�Z��/WN,�����Kز"�NŞ}p֛(�Y�j�s�y�E�����{�[�oq�������6��bX�'�ϻv��bX�'}ϻv��bX�'���ND�,K�L�����Z�uq�˚�m9ı,O;�v�9ı,N��v�9ı,O���6��bX�'�ϵ�m9�:���'t~�k��d5�a��k2�9ı,O�g]�"X�%���w�ӑ,jT�&�}�~�bX�'�ϻv��bX�'�wd�2\�f���V�ͧ"X�%���w�ӑ,K���~�bX�'�ϻv��bX	bw��q	�gIdə�R����A$O>����$�s�{��v%�bX����ӑ,K��߻�iȖ%��{�??���d��ƚH�hNtS�]��dX��xz�'7b�3<�v%�����������%��s5��Kı<�}۴�Kı;�{ͧ"X�%���w�ӑ,K���~�bX�'����YsW2���k3Yv��bX�'}�y��Kı>����r%�bX��/��ӑ,K���nӑ,K��_vk�u�LљXMf�iȖ%�b}����Kı=�_���"X�%��s�ݧ"X�%��{�m9ı,OzL��u��]a�kMk0�r%�bX��/��ӑ,K���nӑ,K���6��bX��<H(������"X�%��_П���5���nf���bX�'�ϻv��bX�����]��,K�����m9ı,O{���iȖ%�b{��;��2�,fKp��������
F�w�\n����ܫmպZ6kp��L�CY��-&�.ӑ,K���ݧ"X�%����ND�,K߲��m9ı,N�>��r%�bX�}ݓ��r�5&�ֲ�9ı,N����r�H�&�X�~����r%�bX��g]�"X�%��s��ND�,K����ɓ3r\4SWXm9ı,O{���iȖ%�bw��nӑ,K���ݧ"X�%����ND�,i�f��D��7��G|��R9J%���ݻND�,K��{v��bX�'{�xm9ı,O{���iȖ"9H�/{�~Q�8ʈ�#��_�p�,N����r%�bX�����Kı=�_���"X�%���ݻND���R9_lž"���q��bt8)6���+$:��<��3>'Z)�a8ݯ\��v�v��x'ϳ��X-ٞN���ٷ^r�S�R�D�<Z�Zz��nǳ�8���y����9�=��%�
3ʹ�v�{�ƺ��8��Jv�z���g)>��j�;m�ƃ�
f9�<�U��ptӨ�,��;��mn�3���
�:hĴ�v�uroW2���V�~����|It~{�������� �[GQ���գy��8-΍��%v�� ��vbb�S���f_S�%�b}���6��bX�'���u��Kı;���a�@"șı?}��]�"X�%���gG���r�s�)%_+㔎R9H�g��;NC�"�Q5���;��9ı,O�g��iȖ%�bw�w�ӑ,KƷ �Q���#jq)�9H�#���s�ݧ"X�%��s��ND�,K���6��bX�'���u��Kħ+n��)9�	P�W���#��U��s��ND�,K���6��bX�'���u��Kı;���iȖ%�by�vN�%�k4LԚ�Z˴�Kı;߻�iȖ%�a��߷{�[O"X�%���w��r%�bX��;۴�K7��������]��cN�eT�uq٬�����SN:��]q[eɋ�;IHGg.��Ȍ�\���O"X�%������"X�%���ݻND�,K��{v��bX�'{�xm9ı,N���3RfI�k4B����ӑ,K��s�ݧ!�)D�K��{v��bX�'{���r%�bX��/��ӑ?�����b_߿K�.[�2k5,�f��9ı,O�g��iȖ%�bw�w�ӑ,K���~�bX�'{�v�9ı,O5ޚ�]d%�[�M3Z̻ND�,�Q?~���"X�%������"X�%���ݻND�,�3Q?}�߮ӑ,K���3��k-�X[�f\�6��bX�'���u��Kı;���iȖ%�bw��nӑ,K��~��"X�%��fwV��)�nk�k\��-X�꣕'��3��Atv��L�Whg��;hHM)x�S�������ow���v�9ı,N����r%�bX�����Kı=�_���"X�%���
5NH6�ȯ���G)�r��w�i�~����b~���6��bX�'߲�����bX�'{�v�9ı,O���ܖf��&���]�"X�%���w�ӑ,K���~�c�A��"y���iȖ%�bw���iȖ%�by����d��\�WZ�iȖ%�b{ܿw[ND�,K��ݻND�,K��{v��bX�j'~���"X�%�����$�ԙ�j�h��r�kiȖ%�by���iȖ%�bw��nӑ,K��߻�iȖ%�b{ܿw[ND�,K���W�C^;V�`�m;c�z4��
��GZ��Fu*А��6z��[���:���Ȗ%�bw��nӑ,K��߻�iȖ%�b{ܿw[D�,K�{�ͧ"X�%���]ˬ���]Bi��e�r%�bX���xm9�,K�����r%�bX�{��m9ı,N����r'� �j%���Κ���a.���0�r%�bX�~����r%�bX�{��m9�lK��{v��bX�'���ND�,K�r^�;f��˭k2��m9ı,O=��6��bX�'}���9ı,O}��6��bX�9S��Aߑ>�o��ӓ��R9H�c���D�� "���W�X�%��s��ND�,K�~��"X�%��r��m9ı,O=��6��bX�'�E�w�����ɖPQy��5���wV��ɻbI:��䜷p��g�'�b��cOj��X�{�{�oq��O���ND�,K�����r%�bX�{��m9ı,N����r%�bX�w;����][����Xm9ı,O{���iȖ%�bw߷ٴ�Kı<�w�iȖ%�bw߻�iȟ���3��W���FR:TڊG|��U�bX����M�"X�%��s��ND�����MD��p�r%�bX�w/kiȖ%�b_;�{�.��K��f\ɴ�K�,O;���r%�bX�����r%�bX�����iȖ%�bw6�_+㔎R9H�u����&�mP��.ӑ,K��w�ӑ,K�=�/��ӑ,K��o�iȖ%�bw��iȖ%�bs��o{�.j����ڹqV�nM�����ң�'���;�;n-�Gf���ͣIf���gmث�9n��n�30N5�����qølv�тa,�3nk��휽[i�9	�鎛ɹ]���r`���H\t�P��͚�z����g�dn)3�p쀆̝�{.�םs�qpO8�U���Ͱ�$t�/�k����ݾ��6FX
�7���;O�ȷ�^�]+��nm�.��۩^-�.|�v�ƞ��-HR�}�ff��E�]`Iu�m;ı,O߲��bX�'}�}�ND�,K��}�D�,K���ND�,K�L�!�0�L��d,�s5��Kı;����r�bX�����*j%�b~���m9ı,O�e��m9ı,O�w�q�L�n�d�I��iȖ%�bw��iȖ%�bw߻�iȖ%�b{ܿw[ND�,K���ͧ"X�%���zC�%��fI�e�M�"X�-��~��"X�%��r��m9ı,N���6��bX%��s��ND�,K���$�&(�4ܫ�|r��G)	�r��m9ı,�o�iȖ%�bw���iȖ%�bw߻�iȖ%�b~ >������[�f$�Z�ќ��^V�ک.�F�����D�u�f呮ܕ��rL5��5��3\O"X�%������r%�bX��>��r%�bX����گ"X�%��r��m9ı,K�{ob��AFTE2H_+㔎R9H�{'������1B;���&��xm9ı,O����ӑ,K����i�bX�'��zk2�fd�I�kY�iȖ%�b{����Kı=�_���"X�T�&�j'�~���Kı?}��v��bX�'�&}��d�rK�	.fND�,K�����r%�bX�{��m9ı,N����r%�b#b{����Kı>�����˭fB̷3[ND�,K�{�ͧ"X�%���;۴�Kı=����r%�bX��/��ӑ,K����SRw0[L���h�\�ѳr�u��-�J�,Ԍ�̲��ގ���Ӣ���[iȖ%�bw��nӑ,K��߻�iȖ%�b{ܿw[� <���%��߷�m9ı,O߰��~�,�2MK5��ND�,K�~�fӑ,K���~�bX�'��}�ND�,K��{v��X�%��s���e�Yu.jK��ɴ�Kı=�_���"X�%���fӑ,`��Y,�{�"�"1bH2�!��U=D^"x�q$/5Đ!b@�Ā��0ĉ��F @���C��$�$aU�񵏉�v�ִҒ$ qT5@��,F#��0_!�0�!$��Y�Ń8B�<EX����D\L@ �T
&+ �A}Tt
+���@�qDM��^��'��~�ND�,K�~�fӑ,K�g��IN�t���_�r��'��}�ND�,K��{v��bX�'���ͧ"X�%��r��m9ı,K�{os5u�e��e��fM�"X�%��s��ND�,K�~�fӑ,K���~�g�������ӑ)�G)����_�B�HnAD�r%:7��^�\�^��gF廱i[���P��sCK32L��5�˴�Kı=����r%�bX��/��ӑ,K����a���5ı?}��]�"X�%�����_�t\��K��ӑ,K���>��r%�bX�{��m9ı,N����r%�bX���xm9ı,O�2�l�52�Z�̷3[ND�,K�{�ͧ"X�%��s��ND��1�MD�����Kı>������Kı>4w�p�L�][�%��d�r%�`؝�;۴�Kı=����r%�bX��/��ӑ,K�D���iȖ%�by��!��B�k$��Z˴�Kı=����r%�bX>�/��ӑ,K����iȖ%�bw��nӑ,Jr���� S>mEJTT&Ҍ�)�Yͥ���f:��7>����t����R�Rn�����Fh��.���ӑ,K���~�bX�'��}�ND�,K��{v��bX�'���ND�,K���m���L�k4h֮\�m9ı,O=��6��bX�'}���9ı,O}��6��bX�'���u��Kı/}����d0�C,532m9ı,N����r%�bX����6��bX�'���u��Kı<����r%�bX����˘Y��e.��f]�"X�~X������Kı>������Kı<����r%�bX��;۴�Kı>�&�z1�M9T	�_+㔎R9H�g���iȖ%�by�wٴ�Kı;�w�iȖ%�b{����r%�bX�|F'��`PT�֠�J(�7�0nP�.:p���%�d	$\=��
�l{n,�[] �1$�n����9
.x֬ې�����<�֍�6`zw��Np�J���l�Ÿ�5,m��m��m��]m<e$ؓ%[���ވ��ݸ�;[������K�ò��A�NÝ�WO��/?�����۶��t�:�ͱ�v{��M�u��h䪇3�S�3�Jo"C�]9�Z� m��k~{��{��:C�S-��0�\�sT���[rf�v�8��I�4�U��Z݄�m[=,�4k��Kı?{���ND�,K��{v��bX�'���ͧ"X�%��r��m9ı,O���3S3WV�Ia��6��bX�'}���9ı,O}�}�ND�,K�����r%�bX�og�
HRB���u���U�6�Yv��bX�'���ͧ"X�%��r��m9ı,O=��6��bX�'}���9ı,O;��̙�sE�Iuu�6��bX�'���u��Kı<����r%�bX��;۴�Kĳ�����_�r��G){�!��'u�Z�s5��Kı<����r%�bX��;۴�Kı=���m9ı,O{���iȖ%�b}�oy�8k-�u�医�z��-�M�du��8)x�>xB�:�V�+H��tnu[�w�{��7���{v��bX�'���ͧ"X�%��r��m9ı,O=��6��bX�'��zk2�fd�K�kY�iȖ%�b{����r�N�dK��{�[ND�,K���fӑ,K���ݧ"X�%��ɟj^���K�ͧ"X�%��r��m9ı,O=��6��bX�'}���9ı,O}���r%�bX�zL흙r��f�f[���"X�@ X�{��n	 ��]�ؒ	"y�bn	"v'���u��Kı>4w��3Yr��̒�.d�r%�bX��;۴�Kı=���iȖ%�b{ܿw[ND�,K�{�ͧ"]�7������ߟ�ӜĠ���3i���n�������K�]�ܹkՠ���q��v�mڲk$��k/Ȗ%�b}�siȖ%�b{ܿw[ND�,K�{�ͧ"X�%��s��ND�,K�w�Զd�˚.jK��fӑ,K���~�bX�'��}�ND�,K��{v��bX�'���m9ı,K�oݶk&�ɬ��F�r�kiȖ%�by�wٴ�Kı;�w�iȖ0t�@���5@���n&D���iȖ%�b}�_���"X�%�{�m�f��̲�9�e�r%�bX��;۴�Kı>����r%�bX��/��ӑ,K����ݧ"X�%����fk0�u��f�ֳ.ӑ,K����iȖ%�b{ܿw[ND�,K��{v��bX�'}��6��bX�&�Fg�t�;w�(�^�n�Ʈ�{eW=$\���{=��Zl�5%n�ۅ�=����V�O"X�%��r��m9ı,O{���r%�bX�����r%�bX�}��m9ı,O�&v�̹f�ֳR�-��ӑ,K����ݧ"X�%��{�ͧ"X�%����f��Ț�bX��������$.T��R�nʪ*n�̹�v��bX�'}��6��bX�'�w}�ND�,K�����r%�bX��;۴�Kı<�vwR4d�5rɫn�m9ı,O���6��bX�'���u��Kı=�w�iȖ%�����D�s��ND�,K��A$�TQi�_+㔎R9H�g��kiȖ%�b{��nӑ,K���ݧ"X�%����fӑ,K���ݟɕ��m�N�P/9��=m���3�u�'Wn*6�=*�9�]r��x�Nݵ\�m9ı,O{���r%�bX��;۴�Kı>����Ț�bX�~����r%�bX��߭������sP�ֲ�9ı,O;���r�c���bw��p�r%�bX�w/kiȖ%�b{��nӑ,K����u35��SXMS55u�v��bX�'�w�6��bX�'�e���r%�bX��;۴�Kı<�w�iȖ%�bw�gڗ��k	�`jkY�ӑ,K���w[ND�,K��{v��bX�'����9ı,O��xm9ı,N�L��sSFkY�Y��kiȖ%�b{��nӑ,K���ݧ"X�%�����"X�%���~�bX�'����"=D���@~�nY�2e�����s����d�\�vTM< ��v�`����;Q�٭fx6����La��ޫ�|sm��N:�q���θ������&B5VL��q�N/E��e�n�+i��ۧ��Ђv����yݬ�p�s���7��M��*	�-��Pq�g�g6�{m�.�4��H=��l�a[�r�[D�K����+�{��?>��C�s�:�.�hH�>ړ�X׹��a�<mm�PZ8�6�p�.z++��4T~{���oq������ݧ"X�%�����"X�%��r��m9ı,O{���r%�bX����%�5M\�R�Yv��bX�'�w�6���Pc���b}�/kiȖ%�b}�?~�ND�,K��{v���R9H�fﾦ�	n�4ܫ�|r�K���~�bX�'����9ı,N����r%�bX�}���r%�bX��߻K��̙�)�Z�s5��Kı=�w�iȖ%�bw��nӑ,K�����ӑ,K���O�n��W�)�r��_��_�i�EU���iȖ%�by��nӑ,K�����"X�%���~�bX�'�g{v��bX�'~�z&�d��+�%F����;��/qp�A�z,Pl[:,Q�o��e.�#G�����oq������Kı=�/��ӑ,K����n���&�X�'�����Kı?|L����XK�kZ�6��bX�'�e���r��4�&�X��o�iȖ%�b{���iȖ%�b{��iȖ%�bw�gl�[��3Z�B̷3[ND�,Kﳽ�ND�,K��{v��bX�'���6��bX�'���u��Kı:h����ɭFd�e�˴�Kı;�w�iȖ%�b{��iȖ%�b{ܿw[ND�,Kﳽ�ND�,Køv�I�Ӛ��Y�u��ND�,K��}�ND�,K�~�����yı,N�?~�ND�,K��{v��bX�'�k�Yܖ�3�F�\�p���ˁ��'C�+��G\-�.�=��;9t����]!%��w�=�%�b{ܿw[ND�,Kﳽ�ND�,K��{v��bX�'���6��NR9H�/b�
�"�EN�QH���ı,O����9ı,N����r%�bX�����r%�bX��/��ӓ��R9H�,�%�q�D�Fq��ı,N����r%�bX�����r%�W�� )�2'߲�����bX�'�����Kı<�zk�sX]\5�f�5�˴�Kı=�wٴ�Kı=�_���"X�%����ݧ"X��������6��bX�'b�Pܪm��|r��G)��[��Kı>�;۴�Kı;�w�iȖ%�b{��iȖ%�bw�۳���&�Y�!����:iSD�=�젶��]&�s5��7a5�K;�f���bX�'�g{v��bX�'}���9ı,O{��m9ı,O{���iȖ%�bt��M���]�Y�3.ӑ,K���ݧ %�b{��iȖ%�b{ܿw[ND�,Kﳽ�ND�,Køv�I��%��I�u��ND�,K��}�ND�,K�����r%�X�'�g{v��bX�'}���9ı,O{�xjܦa35�Ԗ]k�"X�b{ܿw[ND�,K߳��ND�,K��{v��bX�`#�A(S�A�~D��ͧ"X�%�}���5�Y2�f������ӑ,K����nӑ,K�����r%�bX����m9ı,O{���iȖ%�b_�~��K0�L�v�3fevŬ,�Ɩz[��[B�����4D-���
�7L'N�,}��oq�X�'}���9ı,O~��6��bX�'���u�D�Kı=�;۴�Kı<�zk�sYa�԰�BkY�iȖ%�b{�wٴ�Pı,O{���iȖ%�b{�w�iȖ%�bw���9H�#��V�X�8	ʨ�rm9ı,O{���iȖ%�b{�w�iȖ(ؖ'}���9ı,O~��6��bX�'ޓ;gs5�kFkW2��m9ĳ�5�����Kı?}��]�"X�%����fӑ,KTK�����r%�bX�4}�I۬.��ad�̻ND�,K��{v��bX�'�w}�ND�,K�����r%�bX�����r%�bX���4?����@��"�G�@�B+#�b���`!8C*(a4>��xH�Q�20bHFI �B$ @�!�@�1XI#5��Ѣ��2��\CZ�T4<ؐ�&�P�H��H BHA�%> $`  � �P�0�"�"Ϩ��7�@�$a2J��@�?w�of݀��Y�fh�>��T�f7s��&r�N���C��]k\"l�{]�Z�W`�l{�-[m�m�n�lp)2�UJ�*��P ���W��z����Z#m�V�u�m*�p��U ��`H �9�M�� 7���I�E� �m$6�kn *���2���Qc����ˑܵ�n�.6�x����Teg;\�Q�7�.(�Y3��0k�kE۰irV�͸�}����Xwe�J�s�s��5az������\��zѠ��q뱑X����glh�<��74=����.g*����uY96�;s#ˮ������Zݍe��dP�Ŧڀ�m6ԙ�5��=m������͉�����eܛ���&��;9U1�y0�+���)ɫv�n�S=�� [m��H�*�s��ZNz�(���9۶U�:�ɰ<r�6bp�a�*�4�Ӛn��WC��\v��p��m�n���cr�c��x�\vF�q�{v�{R�J��a8��g�Uw����1FÍ�b��v{�K�y_i�9��p@�ݎѳ�6�ݳ�N�
y��ܽ�k�N&uIJ\�/1��l���n4��i᮪U�*�T:Kn}���d���]b.�6F����k�n��m����ɳE�Ӥwg����h�ϖ2,�L�V�M��91��4]Ҵ:5��%h5 1��Q���6%��]U�m�5m�m��#M$I]�mtK׶�[���m5X���WC�ZIـ��^*ڎ�$�$�\�zD����kS�Uu��'�=�7Y؇J��ӵ���:�a�w�-(�f�<�ҭUU+��S@��ç����i�{.�U����Ű�-m���z�A�mn�!$����L�-O ֒U�TLl!D�OU�T��
`C��RB�pۣ��J��֕`(v�T�T�=�� -���`՛6�V]�T� *�ez�]�Z�g���\B�x�K�nfY��љ	�	�!�� v�?"+��L�]��A�^���`r�YDyY���M�X�v,�:�bB��r=7Yn�(0y{��I���e�AY �m{xtS�apBX����^
��K��V{M֔`\�\�n�=���nLt݊m�{\s�r����:z�⎋sgkh����ȼq��ʓݲ�!��F�fژ�fb�yc�r�����Ư[�dN 6�;n��"�b'(:7<]ͻDk��<��  4Zyیv�+EƁ�v��q��aMQOS�Vn:�X+l� i�AuQ�*�2���{����/|}���6ĺ�]��,K��{�ͧ"X�%��r��m9ı,O~���?@E|���%������9ı,O�w�	��30�e�%�Z�iȖ%�b{ܿw[ND�,K�w��iȖ%�bw��nӑ,K���w�ӑ?EuQ,K����L�Y2�f������ӑ,K��w����bX�'}���9ı,O��xm9ı,O{���iȖ%�b_=�̚0��̆j6�kiȖ%���s��ND�,K���ND�,K�����r%�`�����u��KƑ�����(�)�"�0nE|��R9HK���ND�,K�����r%�bX�k�w[ND�,K��{v��bS��W�����D��j����*���.�h�՛I��V'	��
�[��)����ѯ��1�U)�%_+�)�r����{�j�����+76������i���l�s5�'�����C���]�p޾0:�u�BS')O�:j�8��)�+���`w6ig�q,�[�`f�yXV�ՠH�	���V9�@t�s�K@N�-��	(�IITQ��;�f��͞��c����٥���Si5@"�\��^E�fJ�&
���]q;���&��3r��kD�*pp�H�:ME#�;�uX׻8��>�P�^�T�Հ�'뛛���
��7��{��W)#7�Ł�k|���V�v���r�UCr+�~�f�}����А@=cF(�(��Qnk�7�4�7(�M��m7*������N��������� ׯ*�����i����D�v-�vݽ�~��X�N���r��R�$0Q�e�i)넃OB�M3��K��Zi����8n�ە�s-�Ʃ��ߟ�͂� :e��q�@z�T��8�8M�`f��Xֳ]��s]��٥��s�T����J*�RU@�Uk ީ}X��Xt)�޾0ϱ`�nҧ��S��R;��U��}�M�<��nLN{�|AB!������`��$��HTe1���l�=���=.u��� �Iw?����5�-cR*�mtnV�ݠ]�u������ዴ�]��i��u3xn��Q��x>�R�[���Zt� 3�b&��6��R�rU�ի6_���Q2k����)�޾0}|`�S�ݶۃnqRK��U��٥�����`b��KiVkL�ԐR�I"�'M��� :幨q�@z�T���p���BNnM,�Y���z� ~v�b7p�%!B�K���ow~-N<4n)7�m�cgی�;l�c(y��{:�9e�%��;^���������2`ݩ�ã�����"iN;l��v��Q� �;l�m���]Y�t����:nfy��Tta�	J�l1�2ͮ�ޣe`�:Y�6�6UM�f�V��-щt���ܖ�5K�L!Ni�/,*��M-u�L'�7e��:5��`�Y뗻���m�?!;m93Zϕuu˦N+%��9j�:e�(^��M�M�GM��`��:/-��1nk�7�4�|�|���=�ޥNAH�t�jI`b�ן$��;z��;� ���y�EPk���E)8��Hq)��OŁ��ug��]Z��1wu�,�4��J�M�����\���<r��� �ɱ:#iJ�Q�*��՛,W*��=���Ow6���ݢ�Ict�qV�i�i
o���q�=�l:�f�*�����l�6ۂS��X�����,�x���/�����=��)]��E���)��٥���mՁի6X����ʪ��םyz��*p���7��-�@;�1:l�]4����`��,=U�U,�[�`K}�	�`���u�WY��S��R;��U�ꪪ����3}<Xֳ]��ŷ)�q���>7�o����S�ֆ:�1��g�7�8��e� F��N&�#*�`ovi`w6i`wZ�~��s� �~�3�����"����� :e��y%�'M���ߪ���r��l��?�(�*�F�,�����M�	B�UO�ـ~�x��=f�N�jq�)��U\Y��V���@s�R�[���t��۳w%7H$�X׺�s�������5�vq� �*�3B ���$Ԕ7R�l�7��}�}\���ܔ�kv��c^��D��:�.�OD�Nq|o�u`wZ�vq��\������o��QTpJ
0BnU��S���Q2k���;k�pkx��+����~���*p�
F�:ME#�7�����K@s�R�[��w��f�e'"��7���{'���z���3��U*%r���VV�69*
�$W"*�� ��� ��������7�uXn�M�F�6�bD{Z���6ەp��]�l�v;\��VjZ�F�#�T�ܕ`wZ�vq�z�W�A��]X���EN	�L��� 9㖀��Z�EH�nb�������M��W�0��F�j�I"�?k��pkx��gz��`y�`���]��
�&�������5�v.����UR�OyX�릑ࣥ"j�`u:� ��u���󯾜�^,��[D(@������}�p�]	�c@N1,Y��tu,��E�(v
�h�u C�G�C�Zy���e�B��<t�����0�!���ӛ	�tk)�콕Q�K�`0cD6��Y�ӗ7n]m]n7a�)��{uk`�.I�n��]��Y,���M���HcY���eځ9���n�ݴ,=�H�.�4�@�,0HI��6�"�X�A #n�u�;��wv��d���
tQey��6z�.\)7�㴽n+�-�K�y��ѣ���6�QFS��R<��`o^�;��_�_ �5�v��
DJ�C�R�$�?:ns�
"&Gϱ`�_V�s�$���3�IPR$���������Vq��`w�>׺��+6&��r�TnJ�;�f���U����a�qw}����=m8&�2�R;��Z�$��� 9幈S%²�a�q�Pqrk��.��ݛ����k��a�;�2OF�����w��?;|]��Ʃ���}��{<�1 �9�Tu�h�D�NI���۫���ώRJQvk��Հt���?:ns�d{��i�R��`�ܫ5��1nma�D(��Wt��b����U��ɻ��������� =2K@8��B��S_ww���'o��.e�r�ֲ�!3WX�M��J!��?���`��V����`:�t�.4	�#N�n+N�%���8(ut�<I���,5�1�\������ϴ�$�)"EDP܋�g�OŁ�k5�Ǻ���V���4F��R�n�N��J"&Mu�8mwOߤ5��n�=�pM�2%#�;�uX׿]�@� '��T$_A���E	H%R!@��M��#ɴT��"@�T�"��	"��SZ����JX� X[Z¦O��O�J!b���!!�`�H�ĂCX��J�� <�	l�:4)�B�`< TSB>"��A؂�(}dA��U��u%���k�6�f��**#R��I'�!Om�N���Χ]`��8ծ�m#%NqXf�,�%
!���W����������S�;]n���[�;t�������o��8�m��-��m�H�-rñ\���W�����K��6^�����DBK��~,ؽ�T�B4Jt��G`b��`?Ss�k�f�S���"L�w�K�E)P�TTq���+7&�u��`b��`|�Y�H��)���X�I)|�z��`/]`(IZA�>}���ܓ��3캳5.mV�ff��nb�s�K@8��]�����S$jTLq
A�ڔr]u֨��h^'���q�'R��SNf�U��������Gq(�)78Ȕ��y~��`o^�3ri`wZ�vҬ��EDjS%�� �M�r��d|�z��`/[�ܪH�yח��TE8M�`o�x�<�u�DB��u�8mwN�o�#RQ%(�	�X~���,�[�`f�t����|�!N��0�{��V]���N�QH���V�UW=��_������9]��+nxJ���)ݎMz^���R���Ξ��7�����d�cg����]�@۵�3䝰���/*٭ݵ�n�$�q���+HLg�^�]���^u��3�6��܏��u�����-rg����Bem���V���R��Js�[��v:S�ܱm��������zv���� �q��]t�H�Z����uӠv�������ŋ`덵v�jr]m�XZ��3v.�Y�헬��Ŝu
�ћ���?�{��W�~IJT'
*n.��_����l���UW�3^�X^�=$����J@ܹ�?k�`u:� ��s�?Ss��+�W+���ȟ�h�nU*��X��}X��Xݷ�?�|�|�e͢JM�eD�v���)k�y���+��u`wZ�vҬ��EB�R"������BP�＼����g�]���J��Q%N ��mӔ"F�%tԏh��v�臰gvӶ����s���b�����/3m��H�nb�I��A�~�3}�"8�7���`w�_~��-,��;�~Q{�Y�;�~�;��V�[���$�%:ME#�1wu�׺��9��),�����5�v���@'
*���~�� �׋ ��X	(��[�XW�O�8
)T�Ȭ�M,�Y���5g����V���ObT��"g�.��u&�'\0�(t[��:�y�(���tnD�ID8$�QR7��k�6|�`����B��Cy�Ю���$�ܦTJG`b��7�uXܚX���s�\H�*�0�(�!)��~�;�4���U��5X����^�h��E8M�a�rN��0�N������t��릑��a!9�<�`{��������m�(���̂���0:�z�}��u0�ݓ���6���m���2�(����k�}׷!��ۮ�_����@N�-��r��C֢��NT)7��{��ʮRFy��O� �ֹϒ�Jdݮ�WwJ���7"�;��,��U��ʪK5�~�3�I"lC�NU#p�<��8��� �M������Q*$ �� *������>�Mu�(pM�2
E`wj�?s��{'�������5X��W�o�$�R
7%�!qVu	W\U.�/nWBnP��+,�������E* Q�B$R?��?yX{l�<��<�G���:_�V�����Q����&�;�4�;��V/7X�78�]C}jJ����('0��O�����n��l�J�BJ��S��$Vq�z�V�]��%
w�}8���(�Ҋݼݴ��s`��c����U���%��	H�M�8HT���cnN9��9�Wnٺ��]���3�ѣ2��A������6������o\�u��P;Jv�j�<V�ܭ��Ů�8b��h���f��[A<�������Iw<J�m��b\�+���c֗c���}lcfL���smu��ΎÛ^�mw$e^wXo%�͵*C��aܵ�%��` 7�W[ldz�k��}��X3QƤ���k�];+�@Z:�g�u��lv����UC���w{���5=q�-Ya��l�o���Z�9h	�"�3��br�����j�=��p�np���%#Ю���5nq�R+5�{���UU�R]�Ox{�`m*�a�T@���us��B��%�g�N���`ҵ́�y����֭��t�I7��6f9hx�=2K@UT�]���>�t.�ND�sK��!7Yhj�Q�t��uX��0�6;��w�����!�b*#'!�7���`wj�7�uXf�ՀoV�&p��S��$Vq��~�J":(I]��ߧ ��ŀy��p]�C�Rp��NE`ovi`|�T��c���Z�$��ܭ�3v�E"����"!%�Q	V��y`��;�5X}UKV�,�!؇���]�̭s�}
!D}
!D>��|��~,�v����-P��4�	�����ѹ�{rY�n�'epTv(b��Նv� 9M58�)��y�������7n���U���5��Q�A%\��ٝ	(��<��`�>��[����֭��tD���$�`}��VI��^�w0T� �	�!�� 8҃���k��]�>���nI�ͺi)��`�ܫ�<�`wK@N����뒯L�w0��5%���s�|�D%�(���߾<���Vty�����r�j(84SqL].{v��99�u��Ӵr�k�L�;LC�h��JB�8QQ�"�7�4�>�۫�<��r���k�+1��䎥!�EWa�� <�T��c���Zt�_��URF��D��EH�+�����8}�D�޾0>�X媚4�JN2��Xǚ���,��훓���E:(zw��ܓ�G�"$�G��٥��n�X�y���<�`f�t[J�j(�)�#f���s|<|ڍXy�C	�����n�.Fwj*jQR8�4�1!Ⱦ��]X]x� �ֹ�$�K􇺟N�}��K&�F���`9[Y7��3^�Xk�Vٻu��\��Gq�ԘA��l��e^��̟Z�������.�Ɖ
�EF����+��.�o� ��ŀj�k��"��v�p�}NH�RT!��>�۫+�5Y'��߮��^�w$��)^Z/$F�A @H�]#��Ń�0#J�B��LDc�����͞��)�iue)���f�uSj}$Q� bArQ3B��<'����s�7��ඛvm���4�f�o^�n��V6z㡀e�k��z��s:�����c���;���0�Z��^��j�m�
�U73R�P-¦���^ k$��UV� �m��A��֛n���`k�b� Hs-;$��N�(k�m�Ŵ�M���敝���hԪe(
6��k�9���ݍ�L�+>V���MUU�����nz&���&m�ez���Z��9��u-�N6�^��5�1��d�;�iσF��'){t����g�DHFDJ�7nL�Ć�5�����A.��.�k��I��U��޻m�ʭ����ч�mڇ�w9��e�(��8s5�H�(� /h�v_kԊ���)I��ԗ=����޺7:�v���eݸ-Ԟ��f�ˎj/	�Y�.��)�`�9�lJ�q�p��r�:�`�����M���y�*���նs�۷6�`'�g�N6����Y��2W'aW;�eR�P67a\�����:5]�c�qcp�t;(��KgO�(ܸ��C"s�\zH�6rf�Ok=;����k����))���ywB��B)�Ku�y;ut�]��"���-:��WKl� W����e��V�*������Y��
5I�L�;�����筍��̶�Θ�Z�:M��NݶU.���+@�i3]���i����6�Jm��Gm���h�˧��xX�����J��6Z|5T������J�Uv�	�T�8h.���A��%�6��mJBQ;l�i]�Xn���Ut�v�m��[���m9x%7N�ݕGu�+�D����� �'aE�Uej�5&І���͹le#wm�%DU��檃�x5�͝��9&8ٔ��ī�U���C�;>�9rB����2v�Yk#n�J�x�$������w
��EV��T�<��Pm�V�b��l ��5@U++@.�F�(7!���!�b�Ikgs32�%�Y�qW�8�[_7�H  G�S��GIP@]��Nu��sd�����7��l�B��;� ]tW�vt�	=�5����
-�t�hMW&8#e�����M��ڶU,�d�17*a�]�=]�y���2r�N�s�|���Ui�չH�m������%Z�cp��\���q�<A�s��9�#uۣ�vt�[g=N��v�/m6�JY/2�iK��<���o��gnI���v��r�����w{��p�_�ip�i�ላ�q�i�;j*�9���kONt��%ip-؜�e�F��EH����Vq��y�Ԩ�,�}��ܓӦ���k&�:�\�@s�-�Z�EH]�Z�����8��U�tz" �A�$qX��+�EH]�Z�9hSʗ(��ۺm��Ea���Ww����{�`w����P�I*�c��=ϱT�eՓu&�W���u��9㖀��-�6������ā�*��$�6�"Ӕ��v��k;�gY�7(���f����{���� �J'R�'JH�5���`~��}
$�H5��p;�%]Iv6�6����^j��*���7n��y���<�����RFc�S�H���{�����ʐ��<r���3��F܉F��EH�+�5XǛ8�Z��J'ϻ��5r�'Z�:e��wu��zk��9ȩ ���`~��g��⚩q7T�J��U��Rh���g;�]�uz��ᙫu�/K���{����qr$ ���3���`}��V#���*���|�ֺ��#�Sl�.�ݴ����sP��@zc���\H�{�I"E%8�17*��k��=��p�!$��%D�:�6ٻu`}׺����6�S���N�}8��N�[Ł�
>IEu�������$���6����^j�<�T�vs���Z�����۷ 
U7o�]�"�[x�ɨ�TG6��Y�NK�j���D�t�R$���B�/����Hg9�x�=1�@>v]f�NU#��Gse��y���^j�>�۫�RFW��<S��I`c�Ӏ~u�p�gϻ ��׀5+]#b�!�H�>ך��v���{]�8j%���<����wVIy��]��h9 ��9㖀���`m.�l�*qP�Lr�����*�����|�v�rr�]-�劢�,:[�j$dl������K��U����`}��V�{�h����Jt����ֹϦOu>�ϻ�{]�%	)�V{ԜH�$e*m9��=�>�۫=�W9Ij3},׾Vz�iȤ
X�E���h9�@;9�@s�-���`gq
��NU#p�1�x(���}?��S��?kx�J"�"�9�ϡ�h�[�ul�0�m:{ngfjOp\C��g(�GlYۋ����ܻGB�ѦY^�����A�Mf�2��׆�.�8�RKv6�ۇ\o[���ʻ�og�ol;u/��;rYN��5��\!L�[v+	j����Hu�s�q���#�M�R+���,�M��F䋎C���F�ւ�a���e��n���aش�mI��i����x�P�cHʥ��v�E+�hGj�-�pfm�k;4�Z�u�iv,7�����'ր��-�"���e���5ѱD���	V��U��"����<r���.Q��m�集Y����R��j�9h�����H�8�17*��s���Z������̲�Ԕ�%:NI`wj�>ך��v���w6X����/P���IG��]{b�,��/=sӺ��ܽh�K���fLܼ���Z���D��M�"���n�X�����U�޼�r)87B��9*� ����JJ%BQTl����f��y���2�Km��Iʢ�rU���5���9h9 :�c�XF
&� I`wj�>ך��v���w6X��l�q��8���<�T�w��9㖀m�c~/[sm/$��`���Ii��v�]v[#����2As1����N����k3���@yȩ ��@s�-�Z���H�8�17*��՛/ܪHs'ր��@yȩ��,�+r�L�r�7�Xǚ���*�S�r��rs��y�u`b�͖.�Ғ�@�R��̼ݴ�9h9 ���y����ӑILN���q���v��w��9㖀��- ��;��wf���u<ql�u&�ѩX;g��:��U�:BQ{�Q�	P�H�Q��QR9*��՛�x�<��@y���+���S�"�Xc�W������ �ﮬ����r��$�4�dhC�6 ��h�?�����5�Zծ�mE�N1�Ȭ=���S�{�j�v�{�7$���>C����J�GAT��( �3��ݰ>�m�Qr�����`b�͖�s�~��8�o�P��d�? �g�J����e�N��ݳ!�T��9�L�#uqCv*?�{ݾ����М���W�	�}�h<r�r*@;�sP�JRR�R���Q�`}�5X�۫Vl�;�5_�����^��E'ț��7sm�� ���x�<�˰>����Q�ʢ�rU���6X��8�s��	)����\���L�J&� E$�;�5Xc�Vٻu`b�͖UV�JjQӄ	�t�5�xv�����H[+�inۉk,��*'9�{��QnzV�����G8"ݱ�d��՚r��C��ȴ�\�X�v[ԅ��,�:6;��$[/#7����dˤv�=q�����}�n�Y
mtD\a�
Փ���v|=�#뛩�pFc���Tq�vv�� i��<��c��ѵ���WgF��J���õP "���H�����׻���8�em:��[�+a�VY�C&^8�x�ՎP(�kD�� �Ǜ;�#B��)��{�`wsn�]Z��%��u`]K��e�-Iure��h�*@;�sP��@y㖀�3lG�%(��9V.��`}��p�%�JJ��wӀowذަ�*:p)�J��9,����U��f�X��e��7iIJ����c��{k\�(J">��-���.~����V�R�"�S�1:�C���4���[��c3)��&ӉU^��S҉
xn$�:NI��n�X��e��y���j�>�h���*7%X�}�7�� N%�ϐ�S��[��ݜ��� ���Ϣ��W*ry�D(ڜ����{�`}�5Y�r����V�[�`�iF��I��K��Q�D$�{;��7���{]�ǚ��j�!J����7n��sP��@zc��n]�+=�B��N��.Iqp�M��۞�aۉ�u8��P�Po�ww?}����q;8Z��ϵ���9h9 =��&��ĕ'(���q��y���7n�Gse��UčY�R��8�J���� �S��?kx��CP@�QP�n���RB1 H�"$�$-R�H�a$ @���D��YH2�PbD#��X�)D1$A�HB0#d�X�FQM$W@�$H.�R#��L�%�Ѣ�-�F�tQ�CR׍h�� �� �!"J)�]aa�i����@�BR������*H�� F(����X!����@�d��"�Gf�ڿ9�!S�KBe%�����"E�, `Z	 @��T�Ȣof�˥#M0 Fh���!(&���@�]��H�� ��"T�l��!@��h�F5"�#R�P�Q$�Xʁn�
�@� ���JRB�0q0�b}�%]'��Q�8�8}����P�8������srN��U�՛�"��pMSC��`}��V��w�{k\�}>�}8�	�%F��EH���`wj�>ך���,�
;{��Q%ͪ�J�f�URL�Ѻ�����rT�L
��j��s�N��6��%(����|k�+�y���7n�W+� �f�X{OzTt5$�A��hLr�r*@;9�@s�-�c�[D#	ACC�Xf�Ձ��l��T�k�+�{�`}��#�T�����V���s�Y��`f��>ך�8��ߪ��^jM���)�U����8/������ŀl��}�������,�7,j��ƅ�ms��Z"�Ǚ�ay!��;LC�h��k�ƙY��hLr�r*@;9�@sy����БIĜT�9$Vٻu}�drk��5���?:�9�BS#M0��Tt��EI$�Q��`}�5Xk�Vٛu`v��#ZB�(���`|�%�o� �S��?n�X��w���Tl��"�������`~�B�}�~ɯ� ���p(���%�@	T@����n�Z �X�CE>����)������K!\Y�+g<�B�����l�HU����=�ӌ����U���+<ۜv,=)��hN�i6��t�r�С�u��/l>��ۘ➷n؎�3i�:g��l2:�U� ���rd��u�f�<Cn�ScVz9آ��j��_-�rv�T�T jvK9��e�����.��/1��y��Xm�s���̇Z��x94i3=R�����������k���ɪK��;Ej�֯���Wq��.p�	�'g�5��(5����v��PG��X}�]X����y���r������X0�9RJ#+ͤ����9hLr�n*@{�5&���@�����j�>ך��9ʮ%��]X��Kf�D���2�3v���<�T�u|� ;�5XY�)JDB�7$���5��:D&��O�5���?:�8�g��+�v,p�8)�����W-�x��^�N9�%�V\��䅎k.wN��@:�s��@zc���R�S�k)B���I%��y��+��:)%
�(���z�� ��ŀ�]�mf�6R�ܑJ@���j�>��XBJ&G���5���?'I�E�j��49��s�\]�{��},��V��U��f�0�9RJ#&� Ú��Z�����;��(�b�qj�	�cj�k��Yg��n�OWg'f�5;�V)�-��w{�����6j)�"I��|����ͺ�\�+�ᾖ��
D�q��c���k\�(Q'�v, z>��Z�>I$�^��E")H�S��X��Հo��P�Q�""!Uz�\���8���J��ʩQ�*��*�-�ޖw'ր�Z��H�U�&[Y{�Ţʻ�?mk��v��� o��`~�9ʭg���5R'N&�9N&���fٝ���9��7\��޸���R��z]�/D���!�/��{�`}��V�7e��y���k�mN�ڔ��V�����Ͼ��>�<r�olG� FIʰ�,��?URY�|�������4L*'��*����;����p��׋ ��OR ��jTF 9
�\�k���Uw�ۖ˹�H�TN:��0��@s�-�UU�}��g�j�3U���OT�c��DI(�q�).Ά��1�u.�4��Od�T�pCOa����j(�v����Ϳ�|� >$��9ho`�t�Vmnay�[Y��H�&�=�%�9����H�U�&��d�K��`w2ig�����Հ{Oߥ�VWqV�DN8�8���@w8� >$��$�T�\�
JH��IB��sn�-�ޟܮ��=�l�>Qs��B�Ϯfg&�<�����`�ZN.�;m��i�s�U����-i Э͵�n���vݡ�ݺ��׷H�4p���K�et�fz�7���z�����G^���������볹76�n��p��vb����6�L�B���@�w���weT65�ίVG:q�Z�H����]���L���;�r�\jUڳp��:�Rs�����;˝ǽ���񟃤8�;*9�#bY�nS-�������s����j�z��i������8�I0T'+ ?��K�Uܞ��׾^�f����=�TN!�S������u_�RFy���������Ou'R�(��C����-�� ���$� �	��ENTJ��#���sn�Gwe��^��qg��X���D�tܪ�䒬}rjݒZ�9h� ;����x�8���Ӗ3���Ce�U���:�q��N]��4�P�냮�M8�I׭��@{�K@s�-�⯿Uz�[���[Y����n$qXǚ�ꎫ� ��P��S!r�/v��j1!Ȭ�v���ջ,�URY�|�׾VٛcTG���&�X~���� �O�������p�� r�n4�;�5Xǚ��v���ջ,��%Q�\�
�7��-�x^�k�t��'3�Kt��M��� v�������pU*R��41Ⱦ5�n�X��f��3^�wCb�6�Sj�����@s{Z_��@s�-���W9I��DQ6ܪ���X��'��߮�*� ��A9	(�q	,�u�' �kŀMN��6� �`wj�;�5Xf�ՇТ>J"�������}6��Uv�I��@t�-�"� ��<r�����g��B�IE#]I�0���]v^��ݸf;X��4�9�X����qě�ٛ���R u�j�9h��>���8�G(���`�v_�B�5���5���?kx��Q2{i�4� r�r1�`f��;�5Xf�ՀgM�`b�ԜJ��s�r,��:���}ذ|7xDD`��V"c�AL5���]�'~�e�a�f���j��ʹ����M@s�-��+)⭐H��9N�����*�	i��]%�m��n���m��Y՚�X�]�Q�nUJ��V�7e��y���<������w}� ��-G��8ڜ�A�`s�-]�d��>�R |I��9tl��%D ��`wj�>�۫?W9�W)#k=�`f��;X�[D��ٺ]��h7 ]&�<��@tǪ��3lG%H��r�+������p:�8�׋ kT\BG�����(�|Gd#� A
�,c�Z$$�@�V��0�H��F�YZ���*�"A��FNL a��"M(ңY�BP�"P�h4@�J���{��B�{�9��C�Jr#�� ��e�`T�2("����A�� �#"A��A"P��1�@�$�A���T�@�B�u��z��Et0X! ��ffff[s5�Y�ڪ�;��V�\)t��]GM��ڍ��n��D�q�b)I�;Gmt�X�2��K-[[O;l�{l*UTj�WEF�ʃ��[*���IUz����3��5��F�tl崶����6Ŵ !�rf���^۞�,����*�����׀�]�ݪf�:�@��F����ݡ�<�t��۪�r�>Na�ǔ�U�9�	N
�L�2vqԗe�#F0մ���qhɽ>�/W�Ġ�8n���;;]WL%π���[���,I�{`�[tU ����Rm�l؉��6���Er�\L�I�M���1kv�ێڜ���,�bSw�h�ɲ�;rʀ趪� ^�,��d�]�m܁ ��s����lD��UAK*d���7]y�l9槞��������Qs؜SU�\��b۶j�I@�w;Vkn�-��4-�=��y[M=k�3�MN���q]� 5��MY�\Ҁ0d�ra��:��aP��p�n40i�*8�v���[1�:jIy���;n6ӎ��B����D!��֬ɷh�]n�uˬ9(�;������ʶ��Ѣ��\������\#Y�r� �=^V�ym���p��3�N��"a��a����Y�`�*�����d^YM3t��3Z�$j��y9.L]�ly��<cm�29�p�m��i",6�. \�lJ��'bW��
A�j ͞m�$B&[����f: ����������f��cOf�4/ U]��tJ�{�a��7���� mJ���Mˇi������.�mw-�7F��Jr�r�6�R������i�ipKv5&��R��J����\5HU���m��=�vikېN�J�VBS���^Mq�).�UuM����ҫ��v�N6�������@6��9�@+$ko#��,�J�7
\��;v�n��l�Fhm�n�z�Il�󏾴6��5V� ����� ��41�rnoN.��%^��m�N��� +�
����tP�	�U�U@i:*Q�@�>�����߾����e�T�.���gg��d��T�i���W<��O�t뒎�@j��+v�d���څ�������`�sS�@A���/g��Z:t�6)ػ!�l�{4T�[�hn�F{l]�)��M����v{\��ر��[���ɮ#�.����1nL�=�����I��l�St�l�ۋ���#�05�G��.�v�����T�g`�c{p�cߝ�����X�v�I�+�����-ص�x�$ǻl���:{t�]l)Ի��g����|�.���B(�II��c��`w^j�>�۫ ���1w5'R�A�Ȉ9�������M@y㖾�߫�]����Q�N15R��qX�z��3�w��D%:��������Ir[iʩQ�*�3��;�5Xǚ�?s��.��XW�j<����K�Z� �D%]���y�b��������������b����J�^.�������.��@uAL��\�s�Iڸ��Ֆ����Z�EH�I�x�;X�[D��6F$9��n�_ԡ%�|�B���^��N�Z�>�������G%E%&�	�V����9㖀�Z�EH�����Y�R�8'%��Y�|���+�ݺ�1ݖ.��T���8��"�;��<�T�vt���Z�v���wM�.G�գ@�����g���t�K:&�K��u4�vvYW�v2��EH}rj�9~�X9��@IF�֢J6�����][��r��������{�`}��V��X�b�N6�,���Z� �s��jT(�(�PQXB� 
P�վ����=�߾� ���F�Q�RTBV�~�=�~�p�ŀl�n�mk��i9hW.R����Vٻu`~�����f��;�5X����I�ƚwa���[�t�\�{ph]ѣ�[BAC�A����ar���&�|�=�`wj�;�5Xf�Ձ�^h�TrP��*nʫ�g��|�I)�z�N���wvX��'%DR��)G��y� �׋�˓{� s�Հ~�muj�8�JNI��,���5b������"!BJ��d��s�y���nfn�sj��3v�ΓP��@t�-�6�����j�E)�T��6(r����e��Y�)�&���A��fn��cm��4�e���nn�9㖀�Z�EH}#�
��Tl��U%DR�Vu���� ��u�{k\��2jt�y
�J���HU��}ذ�7X|�"!L�����=�73j�q�N
0BnU���s`��Z9 =��l*9(CR�7���٥��y���ݺ�1wu�r���R�ߐ�q
�%-�,���';���U]\v���q��Sw�äg�:��2C{'�$��w��z�;�緮wHn�w�\��F3����fx����z���3�^t&��u���-l'kڶ�wGd��أ�TW���N*_,ڧA�F�C���Ű��h�ͳε�Z�+\ɺ�G=�t`�*lq�^6)Ą]r�  b-W[p�������wwk��o��B]�e��'-�l�p�7n�Ls7oVN��<��ؖAմ�`��QN&8`��V��Ձ�����٥����$r�G��S��`=o&G;�X>�0:�9��7Q�u�%NUJ��V������K��U���u`����*��d��#�Lr�ȩ ��p�J��RTE$9��U���u`b��76i`f�f��8�:C�M5)����Y��w�u����P�u&����Z:@kq���QQ9J�d��Ⱦ��]X���͚Xך��ھ:�IC�����l���J�[�Cwl�?:�8��Ձ�^h�TrP��*n7�����#�R�I�|�y�f�J:�T���U���u`b��76i`|�v��T�%(�!��76*@;�1� :c��9˫ʙ�WP��X+Gb�ct8��mVg������6�%#u�F���n륮�m�n��ـyֹ�~��݋?�)�k�<��U)����=��,��V��Ձ����4ť ؉*"����Z� z�,(�J"�aD@���!d~Pt��V��� ��NZ,��*ꍬ������5� :=����W�PrRQ(�	�V�ݖ��@t{r*@8�*�晗�h�9QBp�ڬ[,i�=Qv�iZ�˛lt^Zt�P�ۂaQ�BiJt�nKsf�G�@G"� �M@;�ͻ�6�r���V^h����T�I��i`|�v��TEIN*hqHX��H����l1�@wQ,�r���r�TnJ��Ur��������`w^jܟ#���X0!�"F!#��!�#� F`E� B1���#�`B#$#$��1 �D!		$c"FIՂ��B�eHI��M '�z/�߶���X�i����G%���Kε� ��X�n�P�%��&9��,-�̳�tf�n��[r�����3t���I�,ˢ�����|}�|�N+�pj�g�ր�EH����lO+u���a)�r+sv��3����٥��y����/�䤢Q�{H����l���'ր�}��3D£��n�*r7%���K��U���u`��`b�h�nD�Q�&�DLr�ȩ >�P͂��#�`UQ=�k34�jۚ�֌����,�jQ���K�6���t	E�g��K����(�b�ޝik��Ɛ��.Uxy�����O������:,��^�z����m�	'8N��q;��%�wgb���A��N�ݬ�u�!Av��l���l��8{h�6�:�=��.��1k���^wS�Yt��9�ͺPŸ͕�IR��ڙ,�[�5m�s&�3���7fCp�4�P�z(�=���^ܶ�.f�����.V����%\�7��ʽN�jݖ��R9Q%8�|r8�ۿ��;�P͂�9h�ɻ��^f�]ff� �j9�@t�-��ߩ �P��i�RrQ���Ł�y-���5 A�(��e�[��.���%	D�[��9�b��w�˕�R���X���N*��)�"��� �����}|`u�p_���~[s���E��M#՘�"���K�w��'O][OA#�Fq+����N�J����6���h��h|�@\ڤ�2�ߥ�S�#rXǚ�j��+�IJ������V��<����w��I�|'�&�p��r+<����R }&�9㖀$�ssM�7kv��ٻ�h9 �j�9h�������I�*�F� ����9h��<�T�P�3L*ݲN�r����z.v����:ݎ	.����7-JQJJJdt�)���DrXǚ���<�T�I��D��˭ͫڰ�ʹLr�r*@��7����N*��`�Ȭ�v�rI�}��� b���8$>�D�)(BVYIHO��	 ��! �!,"��4F�,�E,�V%#"@�d PaH�%b�a�!$�*��R�Bm�YԱ.�_T�=@���6 z���@b�$��!"�G*�m�xC��p�4!l�$�yQ6�P(���@��	)R1�0�Ha �� �B@���hQp"�$��h!)`F����p�	]-`'В6�$����0��$ş!�2'���8�40��B�pO�v1SA�_�|c���!�M
��G �<Q�jxP 4>�|��(���(Z����fUSs�k�� �ޫ�9)(�`�ܫ�W9ķ=�`f���1�@yȩ������̫�ʽ���<r�1�@yȩ �� ú�Dm���H�$bnpJ(�x�=Ϊ6nKQ�nM���rM�M��e0��@zc���R�9�~����V�j='�����>�۫�9�x�=1�_~��u*Y��V�y�Uu������؀�Z����Ձ��x�t�)���	#�;�5X�k������%�")Q*"�N��⦻y�krI���'s&�2kaa��hLr�r*@;�1��m����]tE<���îe���j�����뢀�'Ma.e��v�GF�Xf�<�T�w�b�9hLz��t�8S��!7*����`s�-�Z�EK�9���
�ݣ2�k*�swd����<�T�k������H��N:�"�>כh9 ��Z ��6�j˒�T>9Vٻu`b�k�1wu��^�w$�(h��b��{���<�Sf��:wn��{g�"ұ�Q�����vú^-˴t[������ܜp�>��TN+rh��c]s�d�;Aۚ:���ڭR�nwqۘ���88Ϸm�{n��8���H=d1N����Y6vlXY�Q8�ma1ծ^�Gl`���
�7�nA���M�VYw:Ɲ�ᵻd��C�����n� ��2�ķLgګj�
�"�������{�����u߾�����l�7.�x�h�K��E��غ�<vya�ԋX�K5,d��=[�2f� ?���@;�1�Z���[O��)NF� I������^j�:8� ��\Q3L�L�ͫ7ow��:8���[�b[��@{n���R���X�۫s]������^j�;�����SQ(����w�b�I�Lr�T�����n����N�E����d�,u�kqd���k��W*KW��������77q ���9h�*@;�1������������y�vALU� �T79�y�p5w�v.� ��[�JF2��#�@tqR�9�}& =1�@��du)6�SCNJ�1w5��������u`~�ez��xT�9��7s�K}�Lr�T�I��W���}�o�Vj��B�%��CM����l�n�ę��A���i.A��ml��e�nv�ݽ���Z����5 ����u�)7N"�;��V �M@;�1��?U���~�3ok2%!7*�3������c����NUJ��Tت���{�s�rO{�vnI�^h�T�Rn��JF�1wu�ג�T�I�|�{��W��EYy����:8� ��������?�뗥wM���vn���t�mY�E9���رF�ë��P��ׂ��3�n������5 ��Lr�+uc�IE*�rU�gwe����Lr�T�ꕎ˅��f�^��77P�L@t�-��H�����ҍpl��������`w}�f��>�7%z�B��:�������D�T�:�E`wsn��5 ��Lr��Q�`"���<�˓���,ᨸ�J�m��nz�����0^�/j�ju��\�N����G�ڀw�b�9h�*@{���*I)7J0R7%�������`wsn�;�,]��$
M�E!7��Z� �׋S#����u`���G'�L�ӑ�`wsn�;�,]�vu� ��C��R�J����`���& :c���"���_�=���~o��A<���ٴp�-�Uu+�F����SwK; �i��9{F���涇��[]����zɷg����:�hq�dy�+�J9�,��l۪�F���f�����㇣C������tjc�n�[Bǧ�v�a6=�kc�%]�F��tV�k�խ�54r6*�V�]���3��ܤ��cCjyƉΝN�u�Xg�.�<;Ul b�,��q��]������U���C��j��n�s������*�U�����bTv�Ί�2�f�q&��N6�%��?/��:c���"� �MA�/������0�A�D�G`g��X�۫ ���n���u�)7N��X�۬ �7xtD(�r�� ާӀy�yd�Sq(�	9V�ݖ,�vu���u`}ܚ�
�JI�)��v��Lr�$T�I��\������t�b5�uS[	���u��`8��J��:��+�;Vܴq�p:�8�x�|��DD~�r�� ���JG'�L�ӑ�`wwn�9ʪ��m��Aj��*�P�%��Ұ�^��� ��`[�{JH��CRJ�1wu�ܘ��Z���R��p��3s/hnn �1��I ��`|�4�]F�89H�H���V�x��7XηX����5j�EٻNK�.sMS��_}�2�	9�rΩL�s�[Z:vkp	΂�^zv��������U ���w�b�9h����n��q(�	9V.�n���U��ݺ�>��
�JD`�n;}��$��{�܂�'�=U��W/oݺ�5o���v���S�ȩR{���:H� >�Pܘ��ɴ�rpN$�9Vwv��3���ś����`8���:�qIR$��<V1ER[�6���v�n����C�	ԥ)N"H�R�N45$��7=�`b��`w^j�;��Vki��DE�auu�l�u��%ToVt��ذ�6����k���))��y���"�:���1 �ɈyRa�y�Yt@HU��r������ s�Հl�u�p�(��T8ID���w��5�e�)��`���w]��7]��y�����X[��5�4�(�S��m%q�X���]4"N�ft�2I�^�����%�Q��iF	��1f�;�5X�ۯܮ|�V{��վ�)*q�*Boq��I ���v���M�#�8�H�T�qX�۫w]��7]��y��>�4$��$I�I) ���& :c���"�T��-IFE�0�;n�z�={�����yy�ܓ��*��"����TU�PEQV�*���TU� ����E_� ����AP�B	B!B	U�	B@T$QAP�B �P�EU0�P�U	BAaB$�EB�P��T"��@T BAP��P�P�	E�	E�T$BAP�A�B�)P��B
�P��0(�@T"��U��B�B"�T"00F ��?�*��TU� ���QEZ��*�U�"���AE_��*��EQW��*���"���"�����e5�����D�ݘ �s2}p��   ��   �   �$
T  �   ${�       � �"�(�ª� UT� 

I"J��TU*B�R�P((	#�(QUEN�7� ���
5��(�kő!��s<��`v�;�8�v_�w�<^��)ӝ��t�xz��3Uū���Xz���u
��������sz���{�v�O�U8��9����n�8  |��  >���( SC�J+�O�>��&��{qh,�m���(Y���O�%�H����f� ��f� :\�Af7cu�m`;��W�f�����`��ޏH���k@�
�Р^�]���9����� n�z v��d]�:�: ;X 	�)Af�w:
�;�)e�K� k n��p�v�̠{� tـ,ƀ om���6P ���@�f�   @k ������M�)@����;��{`��>�A�1��)���W���������   Ý���J)�&����y�9{�c��x@-�.�0t��p =�Q���]g!@�`um|��3��s�:��=��k��0΅7vm�  !�7�op΂�\��gc��D���P�o�͸�}��sv�{��   S�O5IJ� hǪ�R@  =��*���  5=��&�U �2 S�j�6*R�  "$)��BDh�4x�����b�����k��;;��;��Ѐ����_�
��S��E_� 
���**�U?��!���.!e�H�Jb���Dk) B0�@�Rh03zu��bD��,x�!w���f�� F5�)��
b��� č�5e���BHhƐ�Hh�"1�4��Ba�H���
�c�4�HC5Is	��a �p�V`c]F�B�k�A�B�H��x�AŀPH�D?��	s`�. 7������%ɭ���˰�p�!sA��$.�4���֢$7�q���@�,�!
�l�\V7ė;B\	s�2���1H�iσ�.iM�/8��6�k�
�
A�D�Ƙi%�G%sD. �2�P�����&����ax�����Mڑ&����5�"HЁ[܌HS)�S�)B,V��Fx��BR����%!�Ƌ$.�P�5 @�F�^@�odx)�	3��i��R"�� �2f�M?��Lɩ��6��i������R�1�c�)B��E����Eq�!����$W�
N:� ���m���i�D!��b��%ms@MF��ə���Щ �����ĺ6�)BR�9����0�*C�Q�(Db���*$� ��@����?v~.���T���7.�&d�x\�0t���Ĕ��B¤aA�#.h����S�$�/�7���!y��^v���M�a4�cw%%���#	�#�xٌk.� �`�+��f�p&�WO4k����9.�.���
s�c)�1# 4D���B�Ini�5�9��9����f���
`��;6�a���M��
Ƹ&�Ռq�0b�,c��\���3[0�0�\�:�����x1�D����?$��L�0���$�&��,�%��N���u�����a Cz)�u�\tf��p�1bI9�5��Й��s|+����D"�~���#��a0bF�N3��2�ӛ����N		p"�!L`@�!d#p%�RY	&FSC�#$dB%T!]��	�:�*�:a.&���# P!A��$�2�r~/9��%4:D���wn����	ro`@/hk�3��ŢH���"��HU0 �`5����A�@��?	ׁCHF��Ej@��i�Õ!k�@B���7��v�Z��4�XS57Y�L/�v_߉M��;k��.d����?�������ơ�r���#�+C �0B4,+<ĊA#Y~9�4�o�)�
5!i������?E����4$�-L&�(�!��`�(���	pѰ�W�C��4%R-�@*�
�R
E(��8<	!L4XNb!!"(@%H-RV5�@*58��8,+��"T�R�Z�*�
1�)�$K�l�u�Đ�IF�B���aP#
+�!\4Ձp{z����e�KSNY}���|bO?FOf�y���=N��[�~�V緥o��N�6��e�в�^Z�Ӥ'�<�WOz��<3�uo4s������t�����i�C�v�M�F!����
S4l�9�2�����w$�B~�F�M0�0eHąb��X���V�[&��H�����o�
�i��k��ap��	-�?f̛���3y��L8˄Hhp>!
1(E��Hjp�CL�i���'�r^F���,�e�9R���E(JF�hCX��`�`�F	������|�!YL!s\�BT�@��%1�e&���s���)!
��.�˘˘Ù>4H��2��eQ���!BV[̟p�m�C�2�Y�,I@i���1�!X3eČ1!�����>H_߈]6ˆ��������~���M���M5x��,���
f��~ M˾0�1��~�ַ��	h%��HRs�~�M�X\"F8p�����aFV$��?}~�j����`B�tDیhF�B�-�ʐ�0!P��1#FcL��F�X�a�),�a���K1�b::0ą1L&f�Uȑ� (�6��HK�D0ѣl.:Sd4a��.���4m��36-t�4fe*B3F��ރq��i�3Y�.aH32�6FR0��c(KsF�0$R�G8�Kȇ�}熓M�7,�S�F���jJҤ+-1�1��5���$���	)�#�dH$"���K)tє!��{	J�P�	��q����ĂB��.�c�:Xܖ˳K�?�d+
�))1���������R4�#'f���ѣL�t���y��?<�{<�ɍ�-���hUĔ7��%Ǐ)�!��~��h��4B�o�.�B��ȜV`?h%�h`m� 	��4��e&+
��~�&o|���ݡB'��.�p������W켚�9�8G ���?�l���c0���o��o��g�GIa��%؁v�v8B�C���W�n��!paP���	Ci�i�nVIK�q�28��	fB�ċSa����!	k�S#��H\���!�#f3�iȑې��@���Y���s"B 4��`2�����9�?4��	�
a2ov��E7��[J�L�%�|�/�� �COߏ�n��H��K�x�A�"!X�HGI"�Jau�\�~���>����a0�	k5�`��$*F�$3VY�@���ɬ��&���Q�$�]�.9!\�6fCLq����Ɏ��&�c��t���'/1�n���Zf��_�����\�!���0a�o�F�"�A��i�H+��cW"P��0��!�4�
$sF����M�`@���3�6ĩ�L�E�ᴉ0�AH�!F7�pp�1$q�8��K�NV�F��P����f�)��Ϙ�2���A�#"B0� F��B�hK��lZa�4�B��
���Ł��@)�$i���B�B�+K�D�9���+
�)�B�:'7���H�;M�v2捛6!(Moz���ٚ!d�Jń	�"ċ
0��Mo��'78�39�5�!���2f�R�%Ǖ�L.0�*D���C^������jv~&��ƞhvhFbP�8M�\�!t$���8:q�!���O���̹�)��]sR��5�h�A

�A��f�[����,�p�#	�6�g�\����'�\[�ʄ)]
��?���%i����K�oD�����}����!�p����L�}�0%W�Ì.�2�t!?�ڿ�$���4�@J�`�04$n]�����,�Bd	�^	������q&����F]��K��$�q�bB%�l���@� ����%�1!
u��iM20�1����g?oe"@bC��SZ���d�X�h$�h� ����%�)(`��}���N$#�H�xm#\t����B���5H�a"�~����;��bMH	��֤n����#C �sH~�!:HW��B$VH��c�d������А���"¸��HD�I̚�����`^��
@�C4�ˌ�
I.�9��9�)#M��0�WN���7��C!	�l���}�� T�	sF�0$�킐?��H�?W[�3HF�-޳a��1�]F2J�"cSF�Q�А�����n���:8q!pѵ~��Y�Iw\K7!%�{#���g���.�� ���Z�0�h�+�k���\�YhKYѡ���!@�V1H�C
b����H�)��4��S|ؓ�޻�kZ   m�q�Iö��)[�t�퇶䳪Y��8M@��6�
v#s-�����È
)`m����`�^�� m��@l-�$p[^6����յm.� [M�  �J��ݶ�m�%�Vm��  -�o  .J�      $    8h�m�6^$�u�m ��X} m�	�-�fl ��඀  $�m ��ͻ6�      o1      �� �  mͷ`     ,-���I�� lH     ��ԁ��m�-����`        ��  	m�l$ Zlඁa&���  ��l ڐ m�����m[@   -��j��m>�   �#m�� K(hp^,����m[v���qm � �`:�m�� ��HH� � �   8pm      m�6�    m� m�  |�� ��l v�6�-��- I9�V�    �`���ڶv۲@n�}M� &3f�zԜ� -6 � 8[��[P[�	 �  � �l  ����@ ��h ��@8 �mm �� �č�-�ж��A��z�ڶ � -����m� %��Xm���m�� 6�Bڶ�m��� m����N� �aQ��jvi`� q暩vzS��RZ�(��VUy�SS=�n�B�)��)����m�V�,p�N� }z�gE�`Hl���$�N�j�A��h       �    &��մI�魸�@	�s�m��  q!$��@,�h�[p �  H  �� 	  �n��  <u�;`�� V���vuR��9F	�t�;,�6�a�h � ձ���-�� �m� :�b@��$�� �ą��Az�u�ֱ�:�8�m&8f�`6�[Cm��(�Wlm�m��  ���\ !#m�[A�lp6�G]�J-����հ �M��M�' m}~���a� ���`�`�A:   &�K��n��:�R�o����-��5N����U@sʪ�[U.�UVҒ�J���u�:�Ϭ�}U��������Y�;$���igLU�c	$�mHW-QeUx 6 ��/R�UW&ĺӻ&��/�Ttm2]oR9n�9T
�L��k�Ki@Y���9j�k�hC�8S�v�b4�U	��J�Wcm]�u
�(�uK��W��)X���,��ۘ����v�-�	��M�$���X @q Y��8�ݴ�\9&�&;ra�ͦڨ:�n�0K�[=T�Pث`(
 M,�Z�yـ��UJ�q����Y�����U���ͷv ��8� m� KUC��	�*�d���늠��-� ]$�@-6 j�a���g6֍�߆�>8:M72�xR��P���N�_��n�H8Yd�H��kjy%��h�nlm�� �^�l�Amm��&�	e�׫ E�C[��[l�6͜.�PhX��j�j7mu���� [@m�5�3��J� ���哨�-�m��6  	4�+�Y��p
���UW�)vs]U,�V�������p9��Wk; �-��2�si6:ھ�v���"N@��ld�� ;n�m�'�U���Umq���U��I6n�l�-� E),UnյK�*�X���gm����٤�n,�UUe���b[-8 [B�m���A/61T�U�F��_@A�uz�n�����U�8А6���yZ�U�Y�X89���@UV��mͶ[@ t�$f�'-ɭ�Ď�m��P!l���$6�� 8��kY 	zV��ж�	     l�]��>��\ ���&�v�m8��-n�o��� �\ �h m�ė��]U�^VUP+�l�3P '$ݶ[@��aj���o�v� .v�Im�eZ��m><}$�Ŷ@� �t����u��H  8ݵ�p以����`#m�zKV�(�������l�a#���gD�e�� v�ZM��l[U�UU�m�U ��A[6��m  m��N����`�UT�u]T��S�$ �[vؑ��D�  m���mm�x6�j�
j����2<Гm��m���n ɷ-U�� ��5,5��=!���m�t�7mU*\�2ˉ״J�Km:;��m�H,�c n�$�$-�V�ئ�80H$��Xk��u͒	 I����ٵ���ѷ6m��:Zn�o	�ղ��H u�d�1 6�Y,� @m�`�Νmp [V� :6�뭓  $Ȑ۱6�� #m��:I�$�l��'*O$�_U}UE�I��Ύ5���s����e�ZRK#m�[@ [A�ٶ�6��'�q!9�k#-�1ͶgLK3��5�Y �
�V��֘Dq�l tٴـ    ����<���]�u�,���6��c�ҭD�>5�,;[dְ��\�w$۶H[E� -���L�	ŵnZ�����Bz�.�v6�1*v�ŶI.��m�D�V�H�	v�n��m�� 8$�V��'%�k[=[Tx������ܻR�Sv��A	�(�*�I8� [@��S�II  $ ַ-�)�jM��]]N_�mR�(�+v���k�Y�e��ة U��� �����6ڀ����s�+�H�� m7Y��0����wo����Im8q��HV�) �@j�� rԫ6���#+�U����l7gn�&�n4�m  s���o�l �:@ H���[��H�۵M����_X��Az��n�� .�Yl+�l�MT�qOdS���5/�4�oj꠷$�㣾�mځ>�� E]$�4;,':��L;mUz�uěl ��2� �P���,�l�rY�d[�9��0�_]d�8�m]*l��q�r�,�0��m�l� [%�I�"��mcqz�ʮ�Jꃐm�l8m��0IV�!OTk6!85T���  h�F�T���Y�-���:	@i��D9�ETlUX��Ƥ����s��jA:-�$�����ZUe����U[*� )��K��&��\�	 �k��m��N�A�m%zl�� �kom�f��m�m�ݠ$ @O+W[z��@W�@��m� �  ������d���lv	3$� �p�`�I6$
<�l�m�� Hm��l{b@%�m���$X�Sh��6 	8еj�n�m�+���4Qa��z�ݶM�t��P�R�ҭ\��0l�m 8a�cZ�mr���L ���2�W��U۪����[@  cX�J ���I��8� -��uP)��8�vz�U��m	�� �e���m�n����I>��/C m8���gL��D�KUup�^�[d�%� p��J ��:�A�-�M��&�����8H n8  �]+`�'@ H�    @�  A�� .ykg����%�m��`�H �8  �Im��Y(��P^K2k�`-�7m��i ӒI�l܎����'gl��ʪ���W� W��V�崐�Kۮ���i�C��k�@�m��n��Ć�8p   ڶs�� �d�%����hh/i�q�n�  ����.�i1m�%nև!m�/Y:��-PR��qclUnS6��R2U	
����7��4P I' �; ��i0 P���5JI�� \�T��VԤt�+)��cbtj��]�zڕ��@smU���\ik��D6uـ+��wX�,F��kC�B�s-ԯ5*�]RN����gS��պ��$��m��mm����f���m�UT�a�����%`�t� p��m��z�� �� VŻ(6�  -�� �%w���6��jR�@����~�]���T/7e���l$p      8�`  -��D�r�@Up��b���UV�ҽ1��@�[!��&�k���*��v9��=]J l8r�����K�F���N�UH�m��m�m��024ul��8$E��v�m&���KwT� U"vj�V��@/'�5��Qm-�#��!q����WK�mR���n
h
�.`�\��H+�و�WL�5�A�r66۬�M�;�@�ݶU�u��m�HWl�+mtYv�mm�f[l\.�  ��	&�)���m���� E� �v�Z $a�v�nݶ�m��Gp�7u�*v�Bj�Ik����
��Fk��U*���@�Dv~AS�a�@ E�
p
Ș*�Ȃ@�UuŔP���D� ��TmM !�j�'P�@8��?=Q��A�>8��x*	D7�: U�`��>!�"Ez(�@�Q�Q�" �E������ Uq@�(�?s��#EU�`�M0I#@��I$ �P4�"b�M�����^�@� h��^�"itA^��kJ���Qb
����S���!�E8�a�x��~G�.�b|v2 �&hQ
��A:)��,W`
 8���
5TSZ���~F�'�L�� ���?��I��II'�c�ڭ�6mD�m��"X��mj���ZU��f�� :i4sm�Ȩ���p<�R\ͳh��[�k�-��9X *��@�l��늸�t��
B]�W��`-��K h�B���4U��UU*����mښ�j��9{v�e����HJA��2�ļ[9f�(&J�w������=V9�G:l�Ҭ`+`٣5. P�m
5*�R���ܦ��^�J$1mX�c:�c��g��S;[��PG2�e�њևa�B6�x�Ӗ�n�]�
�wWIU���P[���N�s��;CO˶�2T0�H���m��@�����2IAW[;l�c
6l �-H���2ջ]�N�[`���v5Yd�f�yì��!��� Z{k,�Qr񓧒�3v\���F��-:��y�\b�
Ng!��#���c��T��LR�n7l����Z���Vǵ�v{
�k"[��&�/����&+���;\�C�2:<��Ѫ�v�r�:G�P���#z�������͢l�J��m4#ec�Y�ʲ�Y��nv��Hcl�1�;�m��Ӵ����#�㫩BK�aBz.6���٪dS!
Y\WUك`qr7j�aj��c@�]��p��y������n�+.)�X�۴���D���R�rq�sO�<Q��<�S]�l:��p g�n���)5!�Z�J;��n4M�ga����m�\Ĭ�ݍrc��Ì�-���mX�c���1�s�n˔�{,&r��΂ѕ;��%N��㜜癉�"fJ(8+Tln�8T`؞�k�Qtq`[x�m�9��3�z���jH�/`k��-�]��*q�M���w�tl����)�(�ݪ`q��!�Wd��F+�k���uA0*�͸!�*4[�j�:J�I�/j�N0�m�enC;P�n�nRq-��
�n���L�M۷[��K�ZE��n�2�e�K$�Պ*��@>e�`,
h_�TC�� ~�8�>�n��f�����LR��#8b P-լ�5�^\r���[Me,��,9� �[�q¦��T ��&3�b�]�œ���k�ʫA��9��_;i۱ծ���r���PJ&�S*J�!�t�c2�%BRg�Vͫ ��B�q�qM�ڪ\��ru������Z�j2��Y8��pa�Egf4�;���ʵ�nv��}������1M��Sf�Y�3&e�\�d��E����l�;T6�ػ@׆&�%�!�%�_���L�V�=�{��<���<�Pl��0��i��;��V&�� �}}UI)ϖ����=�2�c](ISuwj�Wbv��}�K��I��o>� ��')�V���;��`��`��X���} V����v�n��v`�2���`��,���巿M��a�ͬxq�f�0,+%�%�E��6v`�3�!񉙙��vRJ�wX���}�K��+ �H��t��]��P'k ��n��uP"���QA���J9��~�&�}���7�E�{]&!�m����

n��K��+ �r,��E�oS��)X��Wf�+>�:?�X��� ޗ ��4�N��n��wu�o9�O��7�� �I����}�a��M^0r��B�.դ+ӄ+�X4�s�nB�2�f��r,�M�Մ�v+��wS��"�=�2��"�&�t�5h�n��M��7�� ����7�� ާ�`V�)P$Վ��&+��{$��7���<
�
6�W�T��Vdt� ��, �v��+��M�u�o9�NE�oK��L��#�)Ҧ�v�a@���NE�oK��L�yȰ��m7��f������TbDgGb��;����V�=���b <l��ٗ�m�p@�o@ޗd�X�`��X�>��5j����� �&V��Xu9�.�i��7t�+�� �r,��� ޗd�X����M��,j�o@�ɽ���z�t'���7$�AH�Bh���T!�w^�ܓ��}�d-˫5��ݔ���.�2��"�;�Ȱ���}�*j�A�l7E
V���6�Rb�V&�2�94>�߾o�m�]������߂e�4	���yȰ�r,z\0�8� '�We$�n� �:<��� ��d�X���*�SBvհ�]��;�Ȱ�p�6I��r��t�J���n��

wk ��d�`�G�wS�`)ʉV���Z�0�e`����*?���$3޻�}ߵٹ&���C�dD�T-(2��I��5����<
dJ؀��x4G�:�]�	Bk���f�Λ���'c�a9�������PW/�ﭽ��t
Y�3r尉�����Qn�q7^\��4�H�D��R4ViecPL��@�t+N�Nm�4�ξz6v���!vC����l�ܘP�I5i퐳ݕtX����.�D\YGI�����̮GEXb�f����)s&4AK��̳��� �Pvx�U���qի��Z�Mɩ5�Ǵ������	���)�q��L��?�����G"�:u� �&V�k�$�:�ҫWCv��r,�\0�e`�G�Mb���&�mһ)ݬ�L�d�X)����X��9H)&��v�l���6I��r��NE�t镀Gh_�쫤�n� �:<��� ��+ �&V�âT��	�]����0��el�\�Q�F9��0��0�t�r�K��X��<a1E՛��ym��X��X�2��"�=��WMZ̹��k$$3Z��~����C�S��!w�;��ܓ�����>�������@ժ,v酧u�l�+ �r,��� ޓ+ !�1����Hwu���<�t��X���`�e`$��;e�t�M���;Wk �"�>��gǠw�}��o9 T�]��t[ ���2�u�5nא��D���R�g�j�W'�\�@V�z\0�e`�E�wS�`V��-���
�����ߧ'9�%�G�� ���,z\0��� +�]�t�m�`�E�wS�`y]�ʪ�*��+�W�/�L��#y�M	�V]���� �}�L��r,�I�tզ�wn�PS�X���e`�`��XJ�j��ٱl!*EN�g�Oa2aKs�u�l6��;O��du�tt�6���gL
��~��{:��Xu>� �} Cdb;cun��� ��� ��`Ϣ�=��{;�'9'-<�_~�Mh��"���IN|���`�2�RG�Mb���"�t�����:9�L��{�ܟT�B'� "j�xk���N�<T'j��Hln��L������XG"�=����5v+c�V�9���v��CK�m���֥�Y�O�ԗ���v����sc-�f���@�Ȱ�E�l�+ ����Ҧ��a⻷�wS�g���"|�� ��+ �r,�I�tզ6�aAN�`Ϣ�6I��{�E�wS�`����X�����l�+ ��� �"�7�� !�S�ln���`�E�}Q�����`$���J~��v�,C7��7`H[�b�d�#�V	�6P p���6��Z���h(;�3�s�v��yed��y�����Rۏv�ir6��u��q��#Y��ƹF"HQ�ӫ>��lV�uU�k��.���r緘�����..s�5ݓn���m��ղd�'���U�U�j��!��xn![#^g=�� 盶IM�Ê�83E�Y�0�f��5uu5�]*�TY��ڄ�����s�@�K��q�1�3#�XX)pF��AH19hA3t��nxK�*�
��������o9�L�yȰ	�RS^$+���WmU��7�� �&V�tx.�ꭔ犄�U�b���cI-�{^��\���I.}R?} ���< �~��<rF�3�RK��<I%ϪG�%��$��'��@�;<��3�[�[� >�N�9�m�@���/-���{�9m�^�7h��u�Cm�R�eҭ�f�������f�'5�\ 6����.�+��Qi�
���%��$��'��%�\7�����} �ngB��]����o���9�@�@RDR
H1A�Q���vf��:}��%��$�P������V!�׾��)px�K�T��RK��,I%�Og���ݖ�R��X�V o�G�%��Il���Ԓ�s)bI)�;�[�*\E������ $���$���X�K�T��RK�*�������dzu���z��!g6��k��f�@���nF��v�9.^or�9F�^������Ԓ�s)bI.}R?}I/�g�� '����x����3�@7��Y�U6ҎW�?}I.��$��'����sBh"[- o�{��-����7oΧ��`�!YT7J��WbP �� ��
�ct�@�jU:Z ����`D�a� !4?�@n�E	 �Ac�\��� 5b� ~Q���Qh'�~E�%?��Ug=���{�IO��F	%�E=�i[M�wm�U��ԗ�y��y�$�}��׾��)px���n\��~��_|;�����V�Un�X�KgOk�RK�*?����J>��~��]�bI/��y�o}����n�m-��PG6��+fZb
�]i��q$��Qǝ��A�O�S=4��.�(���m����K�ԏ�RK��/��4�}��׾���S�1wmQWt۱�I.}R?}��j|��X�K���k�RK��<���ҟ��_��x�n�i	������߯�#B�'���^����w��@?vn��1�Sc���$�I�{�Ir��$��H��۷��,L�'3Z�eݶ�~�i����m�=��۾C��>{��%��RĒ[ݕ��Kh���1��Pp{1�I\7HѮ�-�f�10��X�Wk11��`��4y�4�-�� ۲G�%�3Il���Ԓ�s)bI/k��a���WMˈ��@?}�<���d���$���X�K�T��RK�wC��;jߊ�]�$���}���Ite,I%ϪG�%�3I(t�$0v��b�{�Ir��$��H��$�L�0I/��}�� wv[MJ�yb�d� ��~��]&`bI-�{^��\���I9���\����)`:�t8�0�^�V����N`��Dw�v�J�n�,F��+b+j�WW"n{,��}g��۩�4u֍#K�r���g-���\��6\m���%[b0\�����6���jF�@X�����=���anQٴa6���p�&۬�s�Ƣ�p4�v��s�Q�mRO�n�XK��̜t9!��kEJ0����m�Rlj�����½�q�f� �58�vERօ�k�h#f�����C��Z���]1��WWo5$��f$��'��%��H�};��&���i�!6�e��t��Ԓ��OIsڑ��It��� O���Kh��Sc3�@>7{����#��%�f$�����Ԓ]�Vx�4�-�� oӽ���{��$�Ξ׾���,Ik���E�i;�t����%�/(Ē[:{^��[�q,�oӽ���];;��6U[��EZ�y�.H�;EӼ,($�Fv�y��1N=)m�bܛL��"-� ��}����x�K�ԏ��^V�IO��F$�_�Hf���ҫ=��w�� �~�����1�KgOk�RIF�QBc.ڿ
��ɼ >ߧ{���C���q休_��{^��Q?�OI{:�K��l����.���� ����} ��� >ߧ{���7u�,�P3�52 �Ξ׾��'"x�K�ԏ�RK��K����>�ߦ��S%�	*�vt6ҜѸ�&���j�i�:���*g�x"�DN6��U[i�n��O�Ē\��~��].⻶����r�|.w��)�����7.��$�r����It��bI)�{^��[��< =���ˊ鍕u��.���k]�v�{�{Ü��TL@C 33���� ݟw{��{IWbg��,I%:Ok�RKy�$���G�%�� ���u�u5��@?}�컶��U}���~�m�wZ����߻�Om����*��p�ȫLQ�@�i�B]6Lͫ��h`�a6�v��i���s���Wv[� ��G�{Ϣ�'I��{���m���:�e*��b�-����N�+ ���E�#�'S�"�]��j�'k �&V�u� ��G�{Ϣ�
��1 ��N�4�n� ���E�#�=��`mT�����*x�:I�V��;0��x��t�X�� �H��m'cb�:N����'F���V��[��l��-�B7fghan�n�Uv�{��2�{�]R<�z���j��o�V��t�X��.��u�9 ���&*V�iYI���u� ��G�{�p�'I���J�m]]���4�`uH���N镁���`%Z��"�;�X�5uv��e`���;�� ��G�w�y�u(�v",l
η
� á�j���6�	[V6U�HҺ�R�Ԣ�`��R�ܜw�˴�v�x;�[��j6�>��mc-�S�nm�t���`A5h�-�]5�K��P��YD� .'tU�:e�.$[�&��c�[��iKO�����g��,gx����ҝ�͆�e)�\������+u�9�[)�d�U*�9��u�:k]i�'$�;��S�I����f�bl7r�HkQq\0���3�?�z���BJ2��	b�`��Y�������w9T� �&V q9� �[,i&����X]R<c�`����*x�:I����wk ��G�l�+ �&V��X�$�0�M7nUv��2�	�e`�E�E�#�%t�*.�t�j�ui�`���;\� ��G�l镀�H��LV՞.�7
uR ��r�l�;�]�Wl��X�)[�W���ډ.Y�<��]R<�\0	�e`�)t�e��L�7�oO�{��Nrp���7<�)�URgI�X�2��p�;i�J�;��*WmU��:t��'I�����K��>R����8�"�j�
�e��:L��\0��xI2���SH�i�bn� �.]R<��X�2��.$�$�]�h��`,a��õ����L�[�x�W>�g����gkN9N�������	��e`���:K��I���]��J���L����#���}��`��x�.*Wi����N����L���aTW�W�Q˪G�t�+ ��Jt�[ch����r��$��6I��r�8%I�v��mՖ��9uH��e`$��=�2�{����C���U�MK3t#�e���ұ�.�>���N��WEn�9�h�v�]�{�V�L�ޓ+ ��#�&ӎR�]�n���	�e`��X]R<{�V WNR�@��wl�wX�&VT� �镀Nr, �2�CI2ՠ��u�E���䟾��7$�����]��0��P�5��5�D��,���"�Bw^��rO�}�$�7nUv��X�}/I��`uH�aO�U�n��/ƚV��RcW���{u����Ys�X[RS�54"h���e��۫�u�Nr,�镀E�#�=�XU�S����Քӵ�{�2�䏔��x��V9ȳ꤈��?�*m]����]���+��t��ꤾ��>��0�j@,;�N�WmU����>�{X����:u����W�<z���T$��m�]2�� ��X�T�gǠ|�}��:t��.����"�LjЈ� �b����B$F!�@�1>�?%���ĉBEIB��7�њ ҀoF��B��0��B�
�BV5`"EP�$`D�!Jߴ �1�B�&,T��"  �H0)	B"AD�1�N�$n��`G�J�Z��)�f���%��21%J�� r5G EJ�*D�,$H¡�r�Hm�n�ka:j\ȋ�%@�$%�h���!I
R"U!H@�`� �T�	B�A++��
b���@���BV0
Z�$xb�p�	�1�D�1��ۯ�XBQ��4�	���&�u�Ȅ�B��(!B'# �"$S��� q�B!��ڙP�~9��J))�aP���^�!Ç98��*�v��M���w��/^;k*��$m�k\�mUM� 볳�m�<��WK���6ܓm�'M�h��[����>>���ە���
�;�����y�QZBzmR��A4%u:6�tEAd�����U�eF8[uhڱ6�-��s�9"�jA)�6X��W�9g�����hv���R�8�=��/��q��R����g��V����XN M�#y4�Y 1�tjگU��g�#=l@d���� ��ԹV5��-Eֽ��G��m��+r��Qm-!&����=���;a�ݗg|��Fn�a�#�h�X���4c^�"j�m��Pq���ه�pv3m�[�ќ[�N�k���b,�����`8S@Gv	疧,��6+��*��Wk�2��3iR%ݞL<���8{{6��T���eB*�К:XCL��Dtа�lԩ��wU�Kl�ĥ���D�m��»�]qq���m�R���䌆���I��渺%7$��0]o���UL�����v�c;E�� �oL�K\WG���ͮZ�� 5�I��`���Ԫ��ڶ�˹�V�n�%��]��6��@���������ӷ�bY������rB[m�#f4�ȹ؅ ���5�72mq�tn�G���c���e�[-��KA�2���!	n�:��f���8�i��)Y��-F�\�Wbܲ6
!br��vk���[I��[9Vpy���'
�73�@Q�nԙ�v�L�\�N�!�<� @�k+���]'I��WC� XȮ�yw��Ḯr]�;`T���0��o!E�ܭUV>~���wl��>��zr��I4f���sa\�]��Uh�}ϐ��1��+�����8�M0ƴ�B��sR�a���py����ܨY,��t��Z�<Cmm/��r��Id� 
ک$ҽ�4N�R�U��i68��cU�Z5*�W�.r�m����=�3;'=���s��A�'O}`�s��[;����{���+�8��D��]L���ֵx��g���c����`R 즗C��,rX��wc�=����1<�qӺΡђ�H�,���#�9�?��a�[�J��|s��ې��P�C���)��]V��j�)i7�k�hm��;X<G\X���9@��k2�Y��+���[Z���ʑ�KiU[t�;���&E�ڌ-�(��6�G&�Fͬ��O�9.��˶�w��ycjx�q��-��ɢ�������[ڱL�������3�ً
򨅷+~����]R<�L���������_}e
��e�A廳 ��G��*���6}���X��� ��ڒL-�Mۻ���]��L�s��U�������?)_�n���mg���*�����z���>�+ �jG���������И��*�꛻XN�`WϫO��X~�t��������Jsm��Wq2�]GU��ݠ3b�V�׋<lv�H깑��Uv;�ӫ-ـE�#�:t��'>� ����,M]��m]]��\2���#}Ӯ[R<�U����J���N�ˤ˻0��,�\0��xN�`'�T+�]�	'n�Ӯ[R<�\0	Ϣ�"�s�P�M�mU[�0��xN�`�E�t��k�s���v��������r]�C=��x�&]�:덓=W[����Y�[t=����E�oI��E�#�=�J�5v�eһt�ӳ ��,zL�-��N��rrZ}g�}.4��Y6[�<�ﲰ��xuo�W�W��\�0���	��6��~ZulWu�rڑ���l}R�p�'SRQV
���xk������$��jG�����[���]�2G��6������ӄհt�P�OV3n�x�#s����v`E�t��jG�t�N%X�W�w��M۵�oI��rڑ���l}$��CI6�����jG�oK���X��X�He0�M7wwO���x��a'��ݻ�~��ٹp"����O}������v�q�,j�c��2�[R<z\0v],-icWAdx�ܶެ��u������Z��̆�v�-�̓g<I�y�`ޓ+ �#�7�� ��, �)	lmS<vU���{���rr��~~0�ϖ�&V9�JB�݈v�]�z\0���7���9mH�	�')ВWi��t�wf��X��X-��.U8�b�_��X$ݻX��X-��.���?z��C,
�dpK(T��n,���Щ�:�*��$3)��Ps�u��5�˒�f����;�iv��JSӹ�\�/@r��I�Nu����aYF
36$ul��oq�ə�yn�G�:�z����͍נjpm�	��'n�aӺ%"��C���)N���s�<�s��������j��.�ힶQL��f�$
����n�L�L�ڦ�l�Tl�����i�C��1�#p{Q��ή��jiS���$Υ&���ЕY�U!`iG0�wZ�W|��p�6>��yUAU��<��:��~��5ʬxkt�.�UUyT��9��:}�V�jG�{]�Եv�v�vR�Wf��X��X-��.U�P�1Ҳ�����&V�jG�oK���X�R�ZWc�-�خ� �#�7�� ��,zL� �%+�Ư�v��m����e9�n�یI��7&'rn7Z��UÄ�Ka��+�]�?y���?G�`�e`��x����Wiۺ�v`E�y�PoI��rڑ�����Ӝ������%
�e!nε�t���ԏ ޗc�K(TH�t/���>��xO�� ��,��O������)�j�ݪ������l}�&V�jM�߹}���X�E3j�kSfɁ+�C)�D��Inv۵�:���:�=C(�n�Uj��6>� ޓ+ �#�7�� ��J*c�e[~1ݬzL��ԏ ޓ+ ��,��/Ī�wN���j�[R<zL�2��+ʤ�>� ��+ �u�]5�T�� �WWo ޓ+ ��,zL����*�}_|���_�`-\���:�w�ށ�e`��x�2�	���L��@ݶ�G*:���m�ul,�t�71q�m�9�s��k:��us�y���g7�y��t[R<zL�c�K(TH�t*�N� �#�:I��l}��{;���}�ײ�����b������l}ӦV�jG�mJ�R۶��۲�ZwX��`:e`��y �2 ��~�E����;O��*c�b��v��2�[R<�N΁��締}���NO��~�U5�i�E.����!5B�)��.CYX�x�����j�+W�����p���=�O���ze`E�t镀{:�.��*wv�v���ӦV��XN�X-�7~������-�X�typ��}���:ea��IE��� �O����SJ�J�7n�ӦV�jG�t镀l} T�2�At�;��[wX�R^ӦV��XN�X�U:�s�����j�r7(c8-��l�_�l`�~�!\p�mē#� ��,��#�C��B,��Q��l�q��Ф��c��[��jU�˸��]h79��\�1��h�ۇT�ps�*玻6ti�{��,�u0�lB�B3
'
ۥ�.e	����pV��(f�����>�ȝ���;f;C�c�|��XQ����)����P�^̧r��.�`
�KYZ9���X\[���lm!s�F/e=Y;����'%��g�m���ڲ����kb������E�t镀�%�R�Զ��m�J�wX��`:e~���]_|�	��+ '))!S+�`+��t镀rڑ�:e`E�rإ��ZN�����`��xN�X��`:e`����J�˷N��Uv��2����:t��9mH����򪯟��l#@F��s�@�7)d:�Fݡ�R�n��ՠ����v�d!��ꭀX�T�.�	���`:e`��xN�X��I%~%wE!�v��2���+�*���<��R^�镀l} T�2�Ah���ۺ�ڒ��2����:t��6�E���;wv�~4����2����:t��ڒ��R�[�i;M�)SN� ��,�L� �/ ��+ %J���LK�3g���ÝL��g���+�.��4�ظܠ7�(�f���:WL[�<��{X�R^ӦW�+����,.�}t�VӴ��"�wX�R^ӦV��XN�X�))�wVݗM�Uz��w��ܓ�s���S�Tz(H)�^�H���$!$�$B�H��q6�#ӴX�?)��P�]�
~Lj�b�A� ��S[�B2A$�F F�� ��R�EZ�^DP�M B$Jh�L	v�$a(I�HqDه"���E�4�%Sh&�>`B��(���
 | |�*�!�� ҆�߹͛�O�}�nI���S�1�MwX��`�2�����&V q9��I_�:�ݻXwL� �/ �I��l}��� ��Q��hivaYG%�%[Y��[\t����0�kn�۱�F���J�����&V��XwL�jtY�t���e�ҫ��=�2����;ze`mIxT�����N�n�TӺ�6>� �镇�U$N���~�e`��T�V�[��XoL� �/ �t��6>� �K�%m;M_�U�wX�R^�镀l}߼����y|��e5&�h� �h^\�G��^���S�]\��9��,n8ej�S�Qm]�ժ����+ ��,��V vԗ�oBԳ�J��;n�.����;ze`mIx��V q9��I_���Cv�`�2�����&V��X]�
��m]'T��`}�S�� ߾�+ ��,��V�:,�R�ۻ���Ww�{$��6>� �����{��1(���*AR�eU	?�T��(��O��k5fy����r�X�Gɍ���|Kkd[W�D!5kl���4�ep�=�O2[���ݍ[0v�j\�p�����'>d�ᬄ0Q!0/\e�z�'F��G	A�>m��sX���1Y톡����.=�9rS#�Û\�:�ppls�ғnG�N��ƹ�7@��B�"�F��è�s� ���T�)Igq,�Z��i2� ���9'$�'^��h-���*L��ݎqv��lq�����P��Kp�nD봦*�X�Wmsv�,�3�~�}��y���ڒ�d�X:9@$�V�[��XwL� �/ ����6>� ��K�%m;M_�U�wX�R^�I��l}��<s�^$v����=�2����5wG��%�е,�R�h�cj����5wG��%���X�].��m��f�yYIr�ۍ��-��u�&	tgŝ1zgZ�V㒼����l����߷@;jK�=�2����
�tE���I�w@<�=���rq�H�����{�,�tx���J���Wh��]��+ ��,�tx�R^�+�
�6۱�b����\,]��ms�3������i1պV�+��r� &ԗ�{$��'>� �y>g�ங4���4�k���p=Cv��sƺr֢�x��9�NZ�����U�v� ��� �I��N}˺<��Jk�]�ڱ���ݓ+ ��,u�X[R<��C�J��ƸR������߷�ޜ���NC��H��b���;�nI�{ݛ�!8s�I_������X��,-��ɕ�N} WHO�[��IـE�#�=ޙX��`�\0I'����&U\锔2����G�.ח L�O� -BktcI��9ņk(X�]�v����{�2�	Ϣ�=޸`mH��]pWi6Չ�6�	Ϣ�;�e`ڒ�����e`�?�-+[��e
�`�2�mIx�L�s�]���wWe
��u�jK�=�e`�E���Uy��<���+ �b��;��-5e��I��H�,{�V M�� ��;���u��wW�[h^6.!� �Q2��JP� W)\�z�^���x��D��X�L� �	x�&VwR���i!;v��e`�K�;���$} T�SĀ�M�mU[wX6��"�$}�L�kd��
��e�Ҳ� �r,G�`:e`�K�=�Re+��j�5c��#��2�l%��2�ڈ��D1��7�y&kږ6B��r"xݶ64.�p=l*�r�ST�l��H��<�$�.ۨ��V.B�m1��R�ȕ��H��f$�9m:z�������:%��۱]� +��܎�G��wն�"�]qЩ7���ۭ�t�PE@��1	�pDA
̰r�4pv8iC�.��sm��&���z6�أV�U��˞m@�vHpu����][S[V�7�;''0������3�"������읋���R�t�\W�M3��,k@Mlj�,Lt�J�P��'�e`�K�;�e`>� �NR�Bm�vU��]�`�K��Ux�'�e`|�� �&V���B��I�M5e��&V#��e`�K�=�R*T˫t�b��G�`:e`�K�;d��"���@+�7~	7n���V v�^�&V��X:�Iv'ʑ�������6�p�k1�]��R��BLnt�q4%WC5���	���K�;d��:>� ��+ ����5�������999�I'(�,gL� 턼jT�J�&ڴ۲��u�tr,gL� �L�d��&4ZJ�v`�e`t%�d��:K��r�Bn���<n�����Ϻ}�z�������΁�s��=eW#t�] k�VJ��3�
�����	;���sz�X`e	�t�i4՗x�2��E�N�+ ;�/ ���R�][�h���XG�`$��9l#�;��E]Þ*���M۵�{$��9l#�� 1�}훒s��]�!߾�m"�;-U���޸`E��y^Rߧ������T[�ӻVV]��p�:>� �t���K�/�C�a�*M��a�v,�V���N0�ܹm�7=�)�uOFn��K~��}�?}�aB[v0.��	�,gL� 턼�\0jG<(E��+lv��2��<� ���������S���lvQeX�� ;a/ �>�<�)�,��e`ΫN�'嶪�'e�����ߦ��w�rO���7%�?@*�@ ,A����%��<T��c��v'f��X��W�}�z;���&ˆ5�S�]9�	�۶�&����t�SK�:�F���s��r:焣˘ݍ��[{�L� 턼l�}�W��	�, ����YFmnF�6g@<���ߤ�䖟y��`�>X�X����E�M;.�RJ˼l�`E��W�UyIw�� ����L��i[M�Tv`(!{�w�rO��lܒ}���ܟȊ%��|`W�?�(E��%c�]�gL� 턼�\0���<򼺪�<�0"�$`D� @�A�!$�!���"�,��*� B5B
�0�.ː�����B��1��F$d��R�FD���-�(�lb�$$��%$��i�F!, �H���A���a#(:"��Ċ�T���A��- ��Q�
���v�m�����#�z�J�cKT�fp9bܕ�%q�X�#�v[�
%Z����-�[A;nu��$8v�mդ���u�n�a�f�l����l���N�g�s���3U$��U82�L�[\�e▕��]©V�-�+�L� �UU�t$2U@e����v�<�9�j�ͦj��K���e��t�]m��6�iBMZ%�mp�j5,�Ud���n��d�/Q��]9`m�H�,`��몫�W;0\+l��u�A� cS��Ш��qɍm��·.=�vu5����-
]��j�Iw�<vrÞ�D��M�J�6�6'D����4g�W�jMv��z���e��(2�n�'.�#s�:H�i0˞��#>�f��68��<ٶ�T f�( nyyN�;r�b+��.�XF��.^��!5l�6����w;�����;q`���d��V�X[��&�T�0KA�4KÝ�.Q,ks`����b���@i�ϴ��MFT.,�e�)�Ikn��{9����n��֌p=m *��=r�<�<���[��.��s����-�V��u���7�@��n{7Tх,ώyb��5�ԵQ�#Y��.���X�t,�e5K��D��- �6����e�,�̝A&5r�%:�-�7@�r�u�������8oml����˻=p���7=M�f�F]��ԋ�^ɶʑ6�$����V�`V(5j�1��`��+V4�ns"�Þ��ʼ�tu���T]CbI�Y wLv�8�4���F抻��'p*���Q�:xu��V7�0���J�*d�R1�U��r��+.�����ֲ���h ����`�� g�ӍO5F�,u��0p�q�ADZ���K�Ɔ�i��h�e4fu6p�ٟU����a��'E�P�M���u�[n�󝚪�ӆ�\`0W7<���Wq�Χ�a��v�Bk%��y�l�aW:ܗj�i9s�2�VW�j�\:��)6�.������'~d��p]�GB��4��jly�z�iM��h5��ۡs׮��8l��!˃�rvۍ֜XŒglYw�����P91�6��ės:4�+�$��N]]b;�D-=Y�w�6�0�Cym�� U���0�D�٠�KH�cQDŴ�RX��dw6�6]�&_؇���l<e�����[;N��#�l�	�n�Z��䱋kq=�RJB�j��t�!�Q���uM��"W]���	�{u9}���E�jųBf4@h�T��*}�Ns����%��j�.� �����p�:>��<���Pw��~�i�P�"�eX��xl�`E�N镀���yUU�$t��e��J�N�|�� ��+ ;a/ �.U�9�_��V�nݬ����}�` �.y^R�\�`t���R.�v"�� v�^6\0���'t��9K������]aqn��Tc�%��1v�����i;�y����������	�;,,+�Y�mE��>}<�bX�'}���9ı,Ow���Kı/~�����bX�'݇�K�m�vͰ2���9)�NJr{����>?�GHhJ�%�bg��ND�,K����ӑ,K���ߦӑ,KĿ��L���۩Iu���Kı>�}�iȖ%�b^���m9�,K�{~�ND�,K��}v��bX�'���h�̹sP��WZѴ�Kı/~�����bX�'~��6��bX�'}���9İlO��p�r%�bX���w=&�.k!��sSZ�r%�bX�����r%�bX�����Kı>�}�iȖ%�b^���m9ı,K����.j@Il�v��'�L�s��GL�3؉��О�ܽN��\щV�@ɝ-3|���,K��}v��bX�'��m9ı,K߽=���?DȖ%���o�m9ı,O�=��%�5�]f\�j�9ı,O���m9�9"X������r%�bX��ӑ,K���]�"X�%�O���,ц]k%l�h�r%�bX��z{[ND�,K�k޻ND��"�`�UjEj,P,BBE���;�w�iȖ%�b{���ӑ,K����8Y)n��֌m���ӑ,K�����ӑ,K���]�"X�%����6��bX�%�ޞ�ӑ,K�����.��3.�f�a&����Kı;�w�iȖ%�b{���"X�%�{�����Kı=�w��Kı/���Md�\�2õ��Ӯ�VY �4�r�=z��v�F�f�nP��*�9�0��y���*X�'��m9ı,K߽=��"X�%�﻿M�"X�%��k��ND�%9)�������k�U���9(�%�{�����Kı=�w��Kı;�w�iȖ%�b{���ӑ?�A2�D�>���j�u�P�sSZ�r%�bX�����ӑ,K���]�"X�
C"dO����ӑ,Kľ����ӑ,K��	l���a��SZ��r%�bX�����Kı?{���Kı/~�����bXO�{U�? lS|��}���Kı?����4�Lѩ����j�9ı,O��m9ı,K߽=��"X�%�߻�M�"X�%��k��ND�,K�@����Ku���MkD��챭�g�,�n��]XV�%��^��t�kb1�
ͨ�$�y?^B���/��?���Kı;�w��Kı;�w�iȖ%�b~�}�iȖ%�b|}�,��Fk3Wn����Kı;�w��?��DȖ'�����K�C"dO����iȖ%�b_w�k|��%9)�NO>�ݟW3m[��SiȖ%�bw��ӑ,K�����ӑ,Bı/~�����bX�'~��6��bX�%����-t]�JK�]�"X�%�����"X�%�{����"X�%�߻�M�"X�#b}�w��O㒜��'���J��^-Vm9ı,K߽�m9ı,N���m9ı,O����9ı,O��m9ı,H/���9��2�&���ѽ���Dd ���m �6�u���WB$p6m�`ke-��dI�P$u����5!,	�N6u�ޔS��-�j�`X����9�d��#������l0ؼ�S�&i,c��c0���դ�3c	��T�hX�ͱ��1d�^��`�i��d6��Pۖ�֫\݉{Hd��Ĕ�HK��Ncyc���e�w~{۾�?��I��d*
e�T&k�eѢb,$v�\pܛ�{��R,�,L��4nٳS+�'�����/'~ﹴ�Kı>����Kı?{��ND�,K��{[ND�,K��>�����FU����%9)����]�!�(�"dK�����Kı/�����"X�%���m9lK����6K�h�u�sY���Kı=�}�iȖ%�b^��kiȖ4X�'�ﴛ�H�����I�9�N����%l��n	 �藿{��r%�bX����ӑ,K����ӑ,K�����"X�%���|p�R���fBۭkiȖ%�b{���ND�,KW�w~�ND�,K�w�6��bX�%������bX�'�þ�Nɿ 2��k�G��.�ݨYI�[�r�&ET�e�V�P��=r��n�o�ߛ�o%����M�"X�%���ND�,K��{[�"���dK�����6��bX�%�����-t]]ZMf�ӑ,K�����!Qc"X�%������bX�'~׽v��bX�'���6��
ؖ%������]e˭9]j�Z6��bX�%������bX�'~׽v��bX�'���6��bX�'��m9ı,O�點�,�e��j\ֵ��K� �k޻ND�,K�w~�ND�,K�w�6��bX�%������bX�'ǵ=�[m�]SZ&�35v��bX�'���6��bX� �}���ӑ,KĽ���ӑ,K�����ӑ,K��Ӿߚ`a<�h�e�J%�v�uѢ'Gd,q_��w=�Gvh�j���yB��0�[�N'�%�bw���6��bX�%������bX�'~׽v"�"X�%����ND�,K�wǚY�5.h��Ѵ�Kı/~����Kı;����Kı>���iȖ%�b}���ӑ?��,AC"dK���ג��fUؚ�{��rS���������ND�,K�{~�ND��)�2'��m9ı,K�w��r%�bY�������m�vZ@V����%'8����M�"X�%����ND�,K������bX�'~׽v��bX�%��g���.�.�&f�ӑ,K�����"X�%�-�}�m9ı,N��z�9ı,O���m9�S������ς�SG���Ƶ�����(=J]��e�k��7�m���e�+Wn$n����sZ6��bX�%�}�m9ı,N��z�9ı,O���l@�Kı>�}�iȖ%�b}��\�B�fi�5�5�m9ı,N��z�9���WQ5�����M�"X�%���p�r%�bX�������,Jry>O�%3[2
l����%����M�"X�%����ND�,K������bX�'~׽v��bX��zo�B���r���9)�I�X�{���Kı/{�kiȖ%�bw�{�iȖ%�U�+dO���m9ı,J{��iufjfh��Ѵ�Kı/{�kiȖ%�`��^��r%�bX�{���r%�bX�{�����9)�NJry7���˶sU��kg��x#��܅F%�Ƹ'���(m�N�7�=+�Tf��fU��
����/!y�ߵ�]�"X�%����M�"X�%�����Kı/{�kiȖ%�g'�C�ϫ�m����y?�JrS������ӑ,K�����"X�%�{�{[ND�,K�{~�ND�@�"X�ǯ��&CR]�JK��ND�,K�����Kı/{�kiȖ%�bw�o�iȖ%�b}�{�i��rS���x�|�Z;;2��,K,K����r%�bX�����r%�bX�{^��r%�`�2'����r%�bX�����셚��%�B˭k[ND�,K�{~�ND�,K�F#���]��%�bw���6��bX�%�}�m9ı,O�U��������U!�JJ�	[hRt����7A;H��.�<�%�H�Oh5�=�@:!�ۗ�4����Nm
�cl���Ӈ�{
�틡��=�� ��3���g�ᎂɓ-�Y��
�R�s`�Wpl�]ն#���n|e
� r��8�;�{yy�XJ�Iu�D�3�c�yJ��e���Cn���n�6�i��q��H[�duL��{ۑ��V��6u�6ȼv.a��G�k���|r"�ٕ�|�{L����ȓ6������^B�>�����r%�bX�{���Kı/{�kb<�bX�'~��6��bX�r_��7ܡXF:�ʷ���%9)������!��$r&D�/�����"X�%���o�m9ı,O��z�9lKħ���K���Au�6��bX�%�}�m9ı,N���m9ı,O��z�9ı,Ow����NJrS�����4�q�v&�^�D�,K�{~�ND�,K�k޻ND�,K��m9İFĽｭ���%9)������˳�Z@�u9ı,O��z�9ı,Ow���Kı/{�kiȖ%�b{�o�|��%9)�NO<��٦��(�c�GL�`�5���l�� �:3lM�̶b���\�'8J�8R!ZQ,.oy?�JrS���w���Kı/{�kiȖ%�b{�o�iȖ%�b}�o�iȖ%�b}���
Z�˹R9gy?�JrS�������rSQE 0Eș���ߦӑ,K���{�iȖ%�b{���""�L�bw�۷?��k3Rd˩eֵ��"X�%�����M�"X�%����]�"X"ؖ'��m9ı,K����r%�bX��=��B�LՆ��]\��r%�bX�{^��r%�bX��}�iȖ%�b^���ӑ,K�X(�����ND�,e9/��|o�(V�pe[�O㒜��b{���"X�%�� ��{��[O�,K������ӑ,K�����ӓ����%��g�)p�!��)���ux��ʸ�����F���[���'q�M�������m��sV��f�Fӑ,KĽｭ�"X�%�ｿM�"X�%����]�"X�%����6��bX�'����&�f�Z��ֶ��bX�'���6��X�%����]�"X�%����6��bX�%�}�m9ı,O�v}v��7*;��rS��������ӑ,K��{�ND������
����:|�Q�(lS�<@h)��C�H�HB9H ��S܄�d,fp� ��0�"#_��9��Є�L@��hp !@Z�POȿ� <��mD
� Wj��<�pC�$MD����ӑ,K���ߦӑ,K���oі�����fjm9İA��m9ı,K����r%�bX�����r%�bX�{���r%�bX�}�Oh�[���k5�iȖ%�b^���ӑ,K��@������~�bX�'���6��bX�'��p�r%�bX��>�*�j�V�F���ei�zݧ��D����<���/��b�^9�Į�	[�ֵ��Kı=����Kı>����Kı=����9ı,K����r%�bX��;��B�LՆ�P�W56��bX�'�׽v��bX�'��p�r%�bX������Kı=���iȈ�bX�%��fy�]ѭY.kZ�ND�,K��m9ı,K����r%�bX��w��Kı>����Kı)�zy��sV�i�Y�iȖ%�
%�}�m9ı,O{���r%�bX����K���
.X��}�iȖ%�b~;�^4��L�kS��kiȖ%�b{�ߦӑ,K����]�"X�%��w�6��bX�%���m9�JrS���s���K��q5\�.¦�����:1�W7�̜&�&31�c}��'�7gm՛gg0��w���NJrS�������Kı=���ӑ,Kľ����"X�%��w~�ND�,K��ߣ,4[��j�.j�9ı,N����Bı,K�{��r%�bX��w��Kı=�{�iȖ%�NO|~>aJ�^TL����%9)�D�����"X�%��w~�ND�[���]�"X�%��w�6��bS���x�o�%t�a��e{��rS��� �����r%�bX������r%�bX��}�iȖ%�*X������Kı?|{sڅ���f�,�jm9ı,O{^��r%�bX(�{���ı,O����m9ı,N����r%�bX�����Y3Z&�!�86,gh6�c\*l�{g��rJ�@�QƮ���m=NF��H��\�*����w<6'u�uԽ�\ҶI��+j��BU9�b���N��c �nc���6�\����e#�D�PL��6r���bd�ħK`�β�x9�/Y۵41�ȭ����+(j)t��\�6qd\mO��̈�f��[gr���Ɉ���H�*]��4g�X�!BdIR�X�]p�v�k.y� mfjj�&���O$�)���a�+{��rS��������ӑ,K��w�ͧ"X�%��w~���&D�,O�k���9ı,J{��4�.j�3As4m9ı,Og}��r%�bX��w��Kı=�{�iȖ%�bw���""�"dK����,��Fk3F3.��ND�,K�����r%�bX����Kĳ�����O�,K���f���%9)�����ZͲ��-���bX 6'��z�9ı,O{���Kı/��kiȖ%�b{�ߦӑ,K������!ul�5v��bX�'��p�r%�bXD�����m?D�,K�����ND�,K���6��bX�%�|_Mk-՚�Z�5�:����[��U���;#��[��b�01av��cI�XR�f��G,�'��NJp�/��kiȖ%�b{�o�iȖ%�b{�ߦӑ,K��{�ND�,e9<�=�LJ�Q��+�O㒜�K�{~�NB!�]ʣ�U`Tı,O{���r%�bX���iȖ%�b_{��ӑ,K������JdӬ�%��M�"X�%��{~�ND�,K��m9�,K������bX�'���6��bX�%��fy��&���.f�6��bX�'��p�r%�bX������Kı=����K��;�o�iȖ%�bS�zy��s5�֦�34m9ı,K�{��r%�bXG�����O�,K������"X�%����ND�,Jr{��}�ë����MR�嗯3�"Z�6�X�^�&��2si5��hׅ���tc�Y�m9ı,N���m9ı,N����Kı>�}�h�"X�%�{�{[ND�,K��=n���ֳZԄ���ND�,K���m9ı,O��p�r%�bX������Kı;�����,K�5�RKL-�CZ���ND�,K�w�6��bX�%��m9��C"dOw[��r%�bX����iȖ%�b}��=�Y���]8�W5�iȖ%�ؗ�����Kı;����Kı;�{�ӑ,K��;����ӑ,K��u?��1+�� 6l�y?�JrS�������r%�bX����iȖ%�b}���ӑ,KĽｭ�"X�%��>���n@L�a48�ͻ�0�*�p�Gh�08#?�z�n�h9��vu���x�s5v��X�%�����ND�,K��m9ı,K����r%�bX��^��r%�bX�޽���3Y�ffh�r%�bX��}�iȶ%�b^���ӑ,K�����ӑ,K�����"�Ur�D�)��.�.jk&6fh�r%�bX�����ӑ,K�����ӑ,ı>���iȖ%�b{���"X�%���ޜ))n��f�f]k6��bX�'�׽v��bX�'���m9ı,O��p�r%�`A�E�ʀ;P һ�=�߿�i�rS������?׳��Y�\�.oxr%�bX���ͧ"X�%�����ӑ,K��{�ͧ"X�%�ߵ�]���%9)�~���F�p!�����Ô������5g:��6�CJ�ۓ�)k�u�SR5��"X�%����ND�,K��{6��bX�'~׽v��C�L�bX�����ӑ,K��u�o�Q�:��[�w���%9)����ӑ,K�����ӑ,K���m9ı,O��p�r$+`�'��L��.[���A;�{�bH$��{�&��'�}���ӑ,K���]�"X�%���M�&��̚u������r%�bX���ͧ"X�%����ND�,K�׽v��bX�X��^��r%�bX��w3<�\&��˖涜�bX�'��m9ı,N����r%�bX��^��r%�bX���ͧ"X�%��^ק���扭e�2��toj�s��ci�L�0S$q�為�:�9Խge �i��)W>�!�ns�ֱ@���(us���Tٺ��=�7Y�����8v݉/mۘF�vy�mq��ۓ�^���s�n`x�Oa�v�MY�ɱs����ga�ϥ��\d����z��i6�v����\\D\���Jڃ6�V6a��T%�3[E�����K	��.�A��[p< �Zw9c�B�逖S�"�[�����s��ݝitۚ���h�}ı,O���6��bX�'~׽v��bX�'}�p�r%�bX�{���Kı?{Ӆ%-њ�ь�֦ӑ,K�����ӑ,K���]�"X�%����ND�,K�{~�NE,K��ǯgڵ�evm�s{��rS�����羻ND�,K�w�6��c� ,2&D���6��bX�'�����Kı=�^�l)�]d��$���r%�g�1D\���~6��bX�'�����Kı;����Kı>�w��9)�NJry��
;d�7e���ı,N���m9ı,O}�z�9ı,O���m9ı,Ow���Kı?��G���F��R��4[���gX�3יj*���[�x�3�:,W��{ޓ��4@nG'y?��%9?�����r%�bX�{���r%�bX��}�iȖ%�bw�ߦӑ,K���~����$3rw���%9)��w~�NB"+P,K��{�ND�,K���6��bX�'���6��bX�%����6K�ӭf\�kWiȖ%�b{���"X�%��w~�ND�,K�{~�ND�,K���6��bX�%>���]6��34m9ĳ�H�&D����6��bX�'�u��v��bX�'}�p�r%�`x�/{�ND�,K��zp���3Z��]jm9ı,O}�z�9ı,?�A�����ߍ��%�b}���ND�,K���6��bX�'���s9M�(\��C�g�ݹ�;nmҚ��Fh��v��k�X)|t=$\-'l:�ND�,K��m9ı,O��m9ı,N���m9ı,N����9ı,Ox׼[
a5���$�֍�"X�%�����"(�%�bw�o�iȖ%�bw�w�iȖ%�b}���ӑ,K���zg��Y���C[�Ѵ�Kı;����Kı;����K�?Ǫ�-`��B
ț������ӑ,K�����m99)�NJry�~�^WK�0����'�%�bw�w�iȖ%�b}���iȖ%�b~�}�iȖ%�bw�o�i��NJrS��ޝ�f��
E᝛�O�,K���ߦӑ,K��X�����m?D�,K�����r%�bX��]��r%�bX��wӚ��e�̗]�9:ۖ5 �lF͑���i�:���c��
�.�8p<-4�lu�[�'�����/��m9ı,N���m9ı,N����AND�,K��}v��bX�%>���]6�D̶f\Ѵ�Kı=���iȖ%�bw�w�iȖ%�b{��ӑ,K�����ӑ?�Eʙ���NJ[�5�ь�֦ӑ,K��u���Kı=�w�iȖ(�bX���p�r%�bX��w�O㒜��'�ϯgڵ�evm�sv��bX�'����9ı,O��m9ı,O{���r%�`EB*!bw�w�iȖ%�b{���V�L�K�a5��ND�,K���ND�,K���6��bX�'~�}v��bX�'���m9ı,O�=�9=f��� ;WF��|��:n�X�,-p-�d�a��*	�k%f�Ҷ�Ϡk��~oqı=���iȖ%�bw�w�iȖ%�b{�ߦ�Q�Kı?{���9)�NJry�~�^WK� 7-��ND�,K�'��]��%�b{�iȖ%�b~�}�iȖ%�b{�ߦӑBı,O��ߌնۓZ��nk3WiȖ%�b{�ߦӑ,K�����ӑ,K����M�"X�%�ߵ�]�"X�%�}��Y.L�љ���r%�g� @ȟ{���Kı?�����Kı;����K����6��bX�%���.�u�.d��4m9ı,O{���r%�bX��]��r%�bX��}�iȖ%�b~�}�iȖ%�bpډ�=�#�$(`���� DcT�!�Kyp,2���PH��`�?1??$2F4��#$g
�1�9�8! *0YZ�b!�`A6]��[��޵�jMRܽ%rӑ����ڹ*m�$��5��tm1�6�pn���t�:Ym�s��l�����omn�6Z�Kh�Y�a6��DµQ���*�������`k<EJ�*�UJ�l�v�v k(몪\�Jس����X*50 ˔yV��m��R�,��v����up���z���ݎ=u:��]@�Uj����6�I[�;&S��`j�n_0A�vS��Wc����]����ZB�J���ў2���N��.��Q����ݙ�;8|�A[66��6������ �ubٮN�2�]�'	Z�ʃ��h��.M��U��CC��a9��h��pF�V$�ݴ�Lc��,d�PW<�[��N�qOd�;�-��k�����s�<P��L�wX5AV�nn����.���8���\��6	��\4�%1�@)�ER�K��� k��j���14ph��.iN4���d�����Gk��v��r�p�v��t0FS;=�Zp�Q֛&gv�b e�v1���v�p y�:���P�7%e�Y�y�H��C�l����M��u�q@��9�Zw�)v�ԍ*��Π�8&�e&��3Yc�Qn���k�9XJǰg�[\h�QK��\�vw$a8�p�.�ۛ��pݜ�h�䭪C�����9����M�B9@�S����P6^6p�s:�v 	�R6�õ�ؔ
�6.��f#&�7����jUX�:��ʎT�eMk�Uy!���n�t��g�FPM�1�=�Y綎+�I��F*_*8�<��v��47N@��Ch��Q�[L��F!���GV�U��X�Am;<�H��!69t��$9 �U�UK[G6�8Ü�c1��
���e��l헓���u�U�-bz�D�<f�Ŭv������`�u�uԧOcێϱ8������"����2���m�eY��9��4�WL�ܥ�9�]aF�`]CK�yM�� ٙ����-b�z%���O��DWʚx,DD�T]�8���'��&�je�ho6�X�1&63�e
A��t�]��C�uɊZ�'g�2���n϶D� �ٵf[3m��f�%��*g��l[7ld��n�8{.�,ؙs`����Rj���T=�øm��4PrdT�mb53+Me�.��K��b�n��ˮ]�*u@��/]e +v�,����	8[RZ�B�|�b�����M�
RY�R:�'X�;.����{ץ��՟6ϋk����6gs�!�V2�mp&�\Z9���,Y�2���\���}���NJrQ;����Kı=���ӑ,K������TD�,K���6��c)�NO����F���X7���%ı;���ӑ,K�����ӑ,K�﻿M�"X�%�ߵ�]� ,�����'���eⶀ��D�,K���ND�,K���6��bX�'~�}v��bX�'}�p�?�JrS���xϷ��l�M�ܳ���bY� @Ȟ��?�ӑ,K��u���Kı;���ӑ,K������iȖ%�b^�=�[�.h�[5sZ����Kı;����Kı;���ӑ,K�����"X�%��w~�ND�,K�}�\պ�{TyM�F��� %Z!���,f�i��L��5�f�
\�,��'97��ɐ �k^3SiȖ%�bw���"X�%�����"X�%��w~��T	�&D�,Ow���ND�,K����%�i���5�Ѵ�Kı?{���* �D�,N����r%�bX�����r%�bX��}�iȠ��bX�Ӿ�4�m�HfK�3Fӑ,K�﻿M�"X�%����ӑ,K���ND�,K����"X�%����?�+��nS���%9)�NO<~��9ı,N����Kı>����K�T�;���iȖ%�c�xY�awCn���v�}>��7d��:u� �r,��y����X��fĲ��g���k�x.�����p���og�h�Oo?�NsY��X\ⶀ�����ݝ�\0�"�瞠�O���_?�j�v���n��p�7\� ��+ ݓ+?W�I)_|���N��+N�;0��]�>��ٹ�5a��$����+�<o\�X��`�\e�$��v��X�X�.����+��S�?~X�~g�R~+
��6��2�z\0�"�7��iW��pS]ZFM���B�b0�Ӝ�d�;$e�1�62r魘q1
���we
�n��7u�>��u�X�\0vL�kd2�*V�v�Qwf��X�\0�2�z\3䏾�W�awCn���v���0�2���x�ϯ� �|��.RHM�,��� ݓ+ ��� �r,+�<���W��e`��[n�������K��.�L�vL� �D+�Ɲ�wuJ�]ӝ;l�J�78��X(�J<� 1�����͊���N��+N�ݘ�`�2��2�z\0g`*LwV_��ݘ�L���;��V����;e�>�*��ăg�������UcM����e`��a�y��%;���:O��%��I���cI�`��`��ot��6t��6�C)�lwn��v`��}�Uy�I�����+ ��� ��y��53�XdXݮ��,�D�3c[���Nq�l�Du��`Ji��]	k5���l�e�⬑��Y��V��]�lU�-f	v��稙T�٥�n7�1K8Ir(���7ezvے7�'��h�`.K�S �J�9���
dܼ]ưp���{�pۗ�v�7a�݌� ܖܩ�W����hW�ʼ������hw%3��N9[�r�{p�q�.#v\4�\��(z0���.Deɸ
��<�߲��2�z\0�2��.RHM�*�]�`:e`��`��ot���ξ��m;w�~[WwXϯ� �{�V��V���7J�E�i�۳ �{�V��V�K���JU��U�Wj�N���7�e`:e`��`��z�ONP�G]m�w73�kSb�f�ۗ��;N��\=>.y͡��e`�[
؍�ٞ[N�X�.l�`�p���,.�njMS%��s��p� E��X�\0�2����@�]7wwN�wk ݓ+ ���&V�9�J�Xա�j�?����ݓ+ ��� �镀t�r�TS��wH-ـ{�e`�`�2��N�{��}J�6�W)���Ǝ5�Rl%=e��z��[\�]j7�W�6��m]Wng��)��n�yȰޙX�L�ݓ+ ���7J�E�iի��n���7�� �e� �r,�-)VR�V)�j΁��_N����ӧa�9�r���Xt�XڥKI:B�e�5v`�X��`�2��p��)`��N���1;�z\0ޙX�`�X �K�����X[|��Hg�g��Ѡ���.�6��hT�ր��	��efʳH*�}��?y����2��p�;�W�6�;O��� ��,���lﾺ�'}���y�I9%���_a	n�3(U����e`��nˆ��X��P�tں�j�ۻ����yT����`~����vnO�_�*|Q�� dTF "+��w�rN���/t��]����7\� ��vL��\0@\��.��e� �C�k#�O�nLWn�!��m�4������2mQ��I/z�ؒ���3������z��e`��n� CeKI]!]Ycmݘ�Xl�`�E�l�+�rI�Z�}�a��]T5����~��uȰ��nɕ�{[Ҳ�
������-ـn��\0�2�>��%�߻��=��?	�n�+�*�69�&V�.�`�M/zQ��Qc��gZ���c�xr�P�RyS#ndN	@%8�ݜ�2��٦]RTf[hR���hT�3�1;�1q�u�=�����z�l-�[; ��q��],�C ��-a���^���G=n��S%ӗ��q��:���4NsOgaY8�p�Rhy��Z����'��[e��U�B�q��v�[%���b��H����>��t����{ۜ�NQ�ٺ�457<i�ڍF[ �^���N��s�c����kWi�f���(\��<�ﲰ�p�7e���W��z��|�_}E[t5w@�[�wXt�`��lr,vL�-�)*Ct�ʺ-]���7e� ��,?�y���<��������)P�J���WH�-ـl}�&V�.�`6T���.�CY�Z�ܓ���f�ʂ����s�h?ߖ��X�%e���Vt��#�Aρ1�]b��ī4�8�0�וXh۲�L�WI�l�bcwXl�`�E�l}�&V��+)P��e��?���~����GAH����O�����\3��^y�GJ���ƭ&ۻ��v��}��nɕ��^RS�������$��*��.����򪪗w�{X�� �r,gL� ����Е���[�wXl�`�E�l镀nɕ����e;�Wb-Q��z�Xsx-!1�שZ�]��ʋ]ut�/n�E���'Ǵ�6�D����7�^���V�&V�.�FB�*���]"�Wk ��+ ݓ+ �w{��Ӝ��><�|��������>��ٹ'�w]��lN�XA�����F�����H21D�@>N�Z�JH$�*�F�E�E`J@b�)A�Q �H�� ~ڱ�!�@ �
*a�S� g6�\�)))��Q@�	X�Y&�-	X�����X1`����C��`U�T�VUa@�A�X ���)F P�IX~�l�7�$�@� �1��� oLj��$��b0c �M�6#Xး�`a!0�$	(� � � ��,�,"ԁU� Y�L"HB0�HD �HD�����XA�V8�-5-Z,��d�,"0�`]��Z2�C &a2��r)%SLh.���!h�1bBR�%aB,W5����&.�i����B��ePI�Ąa���yRV\bBD��EЎ��zCЊDW�� �Q����o�*�7ڰ��`Eҝ�+�7~[��;�� �}�Ȱ>�*�o}���mt���
��Wn��n�u�X�"�=�2��p�?yU�/�?�i�Ƽ�B玬��vl�ppcQ�S�H®7m�=���i�]Q�̉�n�+�f����@�d��;���<��W�Z�G��~����T4�;c.���ݓ+ �u�XΙXZICi��RUn��`��n�������X��e`t��i�Q�j�N��NrK珿^��O��vL���F�*$*���]"�N���V������k�'}��{���I6�l�ݱ���N�I5�X^�p��$n߸~�����Cûmۋ�#��~+�*�M�z��e`��n�� ��+ :G)�$:c�*ؘ���.��UU6H���	���ݓ+?U$mt���
��n��n��ϖ�L�ݓ+ �r,z�ڶ�n��~v�?UU.�ｬ{ﲰ�"�7_E�N�JT4�Z��� wu�{�e`� �u�^I>�;�'���7$΋>#D� dA�����w5����m����$m��]Z���%��P���iq@��q�f���oN]� � ���n�=am�f���x��t�r
<�Vd�&��9\�4j5�W&r�![G<S�٠��7��v��;cvR�S��!
\�iY����:��;�5��;d�A˶|��]F63SZ7�X�����-ό�݈pܳW!'$���%��R�X,+F�F3���z����Ӭ,�=u����\ݛN���
�ۻ�s��n��L��Uz��ﲰ�W�	*�wh*�خ���X�2��2��p�:5PH,��"؝�d�X�X}UT��_����`T�R/�ue[i;�vL��\0�"�6I��#����XҦ���.�Uw_�/@��+ ݓ+ �S�;�����Hy�6���7&%����0Y��Ei.}s��I��k�3�,,
�t�
��~�����e`�e`��l�Wj�i�f�q�3WrO��vn�D|�l��{u�I��`�E�N�JT4�Z��t����&V�.+�+ʤ���,���-$���	�Uv��`~���'��w?�X�2��2���RH�v]j�f��X�2��2��p�	[��`;�j��e�-��u�ʸal)��6��3��8Rlٖ}'':�[0%e�wt�bv���e`�e`������A���`*�?�@�h�H��z����߹���r��>~:�o�X��g�*��"�/�t!����Y��rN��znI��w�sBA��K����;���6��e*ګ���[��yK���`�,vL��Ȱ�.ն�v���'k ��,��U���נN|��"�?y���������b[=�Xyk��f���.�٥�9Eoc�<�vrF�n����(U��y��v`�E�n���XZICi�I�4���;e�?y^RGs��w�|��2���RHiӶUեv7f��X��a��K�ﲰ	�_��KQ�B����B��`}�y������I���}���܀�R5X=�ADz��o{��ܓ����)��Mywwn��&V�ˆ��X�鼶��	޲����&�V̠$u�'7H����X�,CfV-̀��u�U뱞p�bJ�wX�.�`���7d��;�J�*I�wwO�N���X���vL��r,z�ڶ�N�i�	��5oG�{�ea���ķ��,�ϖ9ʔ�i:�i�t�wo �d��=�"�7_E�jޏ �I(M��ՠ*ջ��=�"�7_E�jޏ �{ݛ�i<����Pp;���2�њ��s��8,�hx4�k=�d.R��Z�%��6���k�^}r��6:x8w;<�VjX;r��i������@tǇy�+�Y�cu�q�LQ�̠��ȷ��a�71g�z6�0�`3'���l[]fN�*��u�z6&�r��e΅Œ&^d�n����Y`�k]&;��!)������ۃr�T.:��Au���_v΍��-ݵ��Vtc\�D�#y!���a�C�
��q��]���Y�Ɩ���͙���N�WE��ݜ�9�`��}>~����X�.�Z��![WHvSVݬy�X�&V�K���,䈫��xR����]�wk �d��=�p�7_E�o>� ;�%]l�vX�cwX�.����`�X�)Y�I?.��P'k �}��,ݓ+ ��� 4�*�T�ڻ-�������V����]����,�r�ns���9�u�]�ն��+���y�X�&V�9��,s�)����Cwk �d��J��ŀn�� �}�P�cI�T��j�yȰ��`Ϣ�=�2�k��CN�e]��v���`Ϣ�=�2�yȰd�.�J��h�V5m��7�E�{�e`�`���=\���4�U��2n���=W.����љ��H�V���3� ̐er����%ՑZ������o�nŀn��k��+ bI���)$��y�`{��X��`�X�)Y㤓���v���`ϥ�Ҕ `�H�!`Px��[��ٹ'�����?}�۳V�Ӷ���;X�\0vL�ޗ��I|����>�}>嘺.��L��=�2�z\0��`�p�	(��Հn�M,U՚:�F:nuv�6:c��I]f�Us��s��ڻ
�8�]`��`���7��{�e`uH�:�j��We�0��`�p�=�2�z\0d�兪M�E:��n���ݓ+ ��� �}lq�C.���v`�X��Y$��>�ܑ ���TJ)�{�L ߾m�HI?e]$��yȰ��`�p�=�2�PC����M]A�݇j�pW�X		[PA�si2�Q��EŠ �[ty��芡��߷�ށ��ݓ+ ��� ބYV���vմP'k ��|����X��� �}�Y<Ubt�v!�ـ{�e`�`���7��T�!1�vګT�]��9��,{��&VT�T�t�tZ�-ـn�� �}�ɕ�{��m*�|<�*�
����� � ~���$0�q �����T��*)��]VV��
o�^���A)0c@i +�1B%�A�+2+,D��X��% HRP�H�) ��J$FV�!)	HB��!ģ�)�B 1H��l)eHH��� R��hJ�X0m
�!RV��R0qjԅT�X�� A�@�%�`B��`�!V1��RYKg��6�Eb@���(D	�a��9<�}��dP�$�3@�جB�i����m<�Y.HH6��5���嬧(����sk���;��<�4�i�ze�V��E!Ŕ
��7���k���G���TJ��@]j��K��Uj�yꪍLJu��Cae�i�����bI�t�e��\��U˷7lU*d�N��1���uZl$�s���v�1��*���8�ln�X�����DP2�,[l�U�y��Lq�N���>����"0<Z�I6�6D��\�k�CVlmF�,mJ�W8!-s[H��"�\G�q�"�L�{V��7N�<���s���T6�N�'6U;Y.d��N]]���1�Y9��ȅ�m�F�ɡW�p�ڛ9���I]�(�1�'z�-u��ݶ���,�nqj٭�pA�@���u�v��ڍv1���(`	9�0lh�Q=U�U��[�l��@&;2D��-smr/"ݔk�ƃv�����8�j�@w�m�{��'3���� Z�R]�i+;2�L���:^����*�r9��cPI�GEq��OE�u�L�vd93���wb��������0}���h�Ke�+���Cm`�t�L��K �,n�Q5���a�%ļ*֠b�t�f�y`Ԕ�HĎ��!-���9����۷�ӂr,�|n,��l�ѩ�,M���K5�#hA5�"ʌ���~���wÞ�� ����:	r�s���H�=[=�:�e	υUY6�kE�쥂ug*7s	n������K��Z�mV`�gvPd-l��	x���h7c@s	Wn��� ˲ٴ�j��Z��9+�N4Q���t�q+c�A� 6��p:�UH;Q�q�42Z�Sm��L�N-Z���[�+��l ��1�l{j�F���� ݧ;rC��\�6ҷ��v=��<�ڪ�m�Q���e@5ե`�:U��,���D�+9���n�7c���%��uHc\su�G&�	��B���k�s��$�_��Up@O*��"*�T��WȊU_�E��Y���Sf�EU'c(G8�����4�*�'dM 앸��޹x*ݴ�9�n�&cZ�Q��pQ����7B��O;n1�c��tDgf�:㙧ֺ���F$S\\a"�7+l�)S!l���I1��ݶ�-���b��u��2���vYt 1��޽��+J��8�Tb�3-�B�G��MR+�.��H�v^Y��#=�F�L:�.��Ns�O<��s���S7`�#c7&+���ڗk`l���F�&��A��Z`M]���|�vL�z\0��`V�)
�5ue;.�`�X��`���7�� $�9�B~
��I��`��n�����t|����=��*M�j�ݘ���"�=�2��p�7�U�m���m	��7�� ����;��������X���N��q�
j9�M��.���(+�9�f��Z��Kz��pP�N�u����Cn��&V��X�`�E�T�$�n�l�um]���Y��"TL�>���I���n䟿w�7�g�W�	Ri��V��]�����7�� ݓ+ �r,ޔ\��I�hacVݬyȰ�2��"�7\� ��9H(V	���eݬvL�z\0�"�7�� ޒ���i�)U˙��g3/>NZ���"�:�õ۷\�:���� @���aJn��3�o���m��v,yȰ�2�{�3�J�eڻ���f��X�`�e`��l�YV���vմP'k �r,ݝٹ��*�R�(�S/�޷7$�}�Y<Ubt�v!���{�e`��`���7�E�T�$���l�b�wX�.UU}^T�/@��� �d��$��j�ؙl�@��m�i��X���ݺ����g�ku�v.ˬ۫�.b�ˮ���9:���o@�����=�2�z\0	(r�M��Ҷ7k �}}U��RF��e`>��u�XU��TP����x�k �d��=�p�7_E�o>� 7��B~%~]$��>�<�����;��`Ϣ�AQ9��ٹ'��M�R�L�ֲJv`���7�E�{�e`��`_gۥ׼`)��f3Lݳ��h�e�$`ճ��6�w��;�\hym@ˮAU�j�`Ϣ�=�2�z\0�}�Y<Ubt퍫Hn�`�X�.�>� �} MRP��e�����`��`��,>��K��<{ﲰ�S�T����Zwn�v�E�j��ɕ�o>� ���-R���l�Sv�WH�vL�y�X�>� ^x��.��]Z,V�w��࣠�;��.]Ĳ�D�R��L�։�(�H�=/�]��tp;'^�u�
��R�����y�A�,e����e%.��Q����'>IM��s�k��r��C�\�<e�;s��W�S�ݶ�=F��.[�K�U��u�pb�
4G]��/-�v�D����jƃ\$���7��*n�m[h�k�R�6L9ʲ�K�˓���{ww-�%l���'[sjd��q�窰x��,��ǎn8Y��W2��	Y�e�+5���wj��?~��7�E�n��WH�z1J'�we$�����,v�E�z�G�{�e`�Fg�J�c�v;X�>� �t� �d��7�E�v��m��۶�
n����ɕ�o9�O��69S�V'Nخ�ݼݓ+ �r,v�E�j��.�b��E&QwE�7.�nS���VݞuC�p���8�uas�ـ�'J��V�� �r,v�E�j��ɕ�t}NJ��wh*Ӵ�`��,ʪ�����z�G�ot��7�E�IMH�[W㫴[)�X��x�&V��,v�E�E]�E
�v��˻X�&V��,v�E�{�E����!?�J�����`��,�r,ݓ+ ��gJ�3��=t���^M�*�`�5����Qr�H8�����]�\�@���鼋 ��� �d��7�E�ʯ6C��i6�wwwh���`�,ݓ+ �}�O��=�T�E���wLv�vL�y�Xo�����<�}��X�RP+Iһ��b�wX���}�9�ɕ�t}NP�Mӻ�i�v��}�9�ɕ�~�y���y.��VZ�5���;�����q����/;�a�M��Y����R70JV�����n��9�ɕ�o>� ݧ�`WIb��tջT�eݬݓ+ �}�O��=�"���h��]�HcwX���}�9�ɕ�{��]*N�-�ev�'��|k���~�{�rN~�vnD�9 A��,d"0��D�Q�`�1� �X0X��F)I!���a!���$|���z�}}��ݶ�V����{�E�{:e`Ϣ�;i�X�I�I���O�D�5f�Z�-�׆�'Uv3��x�������E�����լ/\ma�UwHv�~�e`Ϣ�;i�X��X5I@�N��+�� �}�O��=]#�=�e`S�H����
��;Xu>� �t� �I��o>� �Mt)[�~;*�ݬ��<�&V��,��E�E]%���V��+�v�d�X���}��~��巳�I'$��5rb�2�,l�J��J���L�l7&�=K;8%64m��e4BpԺ�QL��i+�V�x7�n{��Ɋ�]�k����#;�d���N3]�v6-r�#<�gsmm7S��@
�!���R�����r�� Y����X�?]��N������ѳ�K���S#�|�5���l���,��jZ�e�oM�8�W`��9�Ӝ�Od�=a���B�p�ǟZ�#=�봏\ȗ�MNm�X��ف�w��a�ˊ�-ܵ�����{���<��`��z�~���|���Si�զP+��wS���`�2�y�X�J��4خ��E7k ��E�{$��=��`��,��JAm5e��[�XUU-�ｬc�,��E������}�����@ͺ9�Q)�`���}�>� �I��]-�YZl�7\��5�H�qcNun�фv�.���h��"��36ЛL��i����X�y`�]X�y`�c�ԃ��6gY�ym���ONIɼ��=�e`Ϣ�;��XU��@	�+N���`�2�y�Xu>� ��E�ъP	?�X�u�{Ϣ�;��X��,�&V�#Y�Ҧ�nզP'k ��`��d�X��, �AP��ݍ���Ye*�a�k��]���%׃2�q�:�Nh�m��AM�۶�AM��=��`��X��,z�E�{�H-���]�wk ����=��`��,�} zI(����h�5wX��,z�E�^QB) ����+q���p�=X�a��~#�&�.���N��"V���� A���%@��������Ѕ�~\MZ�M�6;P�*�H)	��X�1 $XE�$Y�)I YK(R��1� Rp5��ddH���H�� 	0 �8&HV$E�$�~����~%! ���#��#mI�0l	�k6��6-X�i`�B1� �~ �F+u�0pP>����ki�ס4�	�'ƠM���~�i �.���P�H��-��:H�W�E�1��d# �
��T1
5��C𢿕t���|�mGB+�f����ze`���t��PZv����<��Ү|��|�zL��}6��E���~;)�)�X��,ޓ+ ��E�oS�\�.��բ�� �nI�*C�30)��R�0`�����s6VB4�� e��v�d�X��Xu>� �} wG�~+iU��wX��,��E�{Ϣ�=�eg�W�����g�J�M�m��;X��� ��E�{$��=�"�=�eZV�۴�AM��7�E�{$��=��`O��	D�($
BJ�/9{9'�~�w�/@��#� �8YA�k �I��{Ϣ�;��X��, ���K�[nk��B1Z���eb70frė��f�6yc�gq��룙�j�f��5��� ��E�wS�y�X�L�.���t��PZ���wS�y�X�L��}}^$}���,��+�iS�)�X�>X�L��}�O��"��R N�U��I���=�e`���}�>� ;���	?���i���}�O��=��`N}��ܓ�p��A���=35i�m�s��luے^P!�wm����օ�<�N�b^SA`�!��B˹tKq��;���fH |9Z9�6s��'/T�c���ۇ��öD7-����˹�:�cf��-�ƤW:i�i�k���ۂeۣ���أ��!ęP�@�-	�۩#��O:�Q��؍��ntb㶹]��2��y�XI�:�x�n�s�3Aa�kQ��998t;���[ub�F�8)ù<���K����74l�]cTmfhm��Xjf�R[�>�M��^���,ޓ+ ��� �N��i[m+�v�AI��7�E�{�e`�`��,d��Qce�e� �v�d�X��Xu>� �} MRP&���i��wu�{�E�wS���`�2��S��ӻ�iڻXu>� �}�+ ��� *h.�[Al1��gi�ik�ea�܄ܽ8�9x=�o��3����<\��r��ۣ�,�&V�>� ��`WG)I%��kT�35w$�{ݛ�'��y^myUUV��`S�`���8� '�m*�n� ��E�oS�y�X�&V��y�ҡ�j�P'k ާ�`��zL��}�x�W�i[m'c��
Nנls�{�e`���}Ҥ1YB����3�n�S��:
Y��bD�i���x�uۓ�M�\2�.�Z�A�z�����?�r,z�E�o>� &�(I�ݴ����`�`��,y�X�&Vy@tr��n�ݪN���7��Y$��w�r
#���H�C����{+ ���,�U�^%j��*n�X�`��X�`��,*�� v�n�Rc�X�&V��X�>� �r,zL*��5v+iӻ�-M�jsی��Hi�����C�;r׶���[+m��h?iU��wX�`��,yȰzL��Ѽ��P�5j�x
�`��,yȰd�X��kzVRJ�i;�PRv�yȰzL�y�X�>� ���EJ�_�˷L-�X�&V��X�>� ���>�T94�s�o]�נy~���]�]���X�>� �r,ޓ+ �{��Ϫ�M��s�@�K�,�fQ���u��p4,�Hh�r���l-fIo5�[ӵv��9��7�� ����7�� ��i�׉Z�;J��n���X�&V��X�>� ��9H]�����ޓ+ �r,>��N|��_� wG��-�lM7u�o9�O��7�� �I��{:7�]*&�]/]���E�oK��I��~�w��߹9$���K�e�ٮ�[�X��&�t��ʍ-�Rv%e����w1Ӂq2&�9��j�4�)w���X�ei]��`nb�Ļ�q��� ��Z�pD�$�&˥�0M2�����O<u�y�.���Q���uěeb#	l�N����`��d02���#e�;�n{Au��F�ܺvb��!v��h�ѣ��$���}�\���%Wo=���~E�`qQ�,��Ԗ�մ� \�՜\��V�u�)vm9Μ��
��gn��.�[3���krgR�������{$��7�� ��`����V�j��N��&V��Xu>� ޗ ���M'N�E�wu�o9�O��7�� �I��{��^5N����]���E�oK��+ �r,gX��+WI�t��v��p�=�e`�E�wS�zAc��n���@�nmL�ew��7&�<59�x��pq���}��f8�1efٔ��G�
��~��0�"�7��_�<��>�� ���\eѩ���ѹ'ﳽ����Q�!�$�A�A"0")(b�jA?�q�����s�`N��0zL��Ѽ��P�5j� +��oS��p�=�2��"�=�递��n��

N��.�&V��X�>� ާ�@Z�U�n�]�X�&V��X�>� �r,�<��ß6Ѯ�[�,���r�d$�J@W��T�&+���8�ۊ�`Pn�A�t�M]נt|��}��X�&V�k�!x�]ݺWb�X�>� �r,ޓ+ �r,�X���
��v�7tݬyȰzL�.���<��O�����(wY�]�;���"��R Wj˺���`�2��"�;��X�`tqZ O�]��m��yȰ�}��X�N΁��'����1��j4J����2e4���jf�nq���nӏs�o\ra��P+��wS��"�=�e`�E�{]��m�ݫ���yȰd�X�`��,z�T��c�L.ݬ�&V��Xu>� �r, ���M'N�n��wu�������{�rN����I���n��'����＝ߵ��[f�W@j�o@��`�E�{$��7�� =���i���d�;
�R����)k,�K�����B:[*�9պ����r�CSعm`��{�e`�E���AҜ�`l��@	ګ�t	�v`��X�`��,z\0�8� '�We$�N� �r,ާ�`��{�2�gF�˥M	�V]�ާ�`��{�2���`[&!�m�ݻ���ޗ�U^l��)�N~3��rO��**���**�� 
����QWE_�@� TU�� TU��?�P@T#P�QD`@T �T B
@T",B �EB+P���T ���P���T"
�0(�T",B+P��T"DT"0��B	P��E��P�0��T" @T"��T"(DX�B DT �$B "@T (� �P�@T  ���BE��@T"*@T ��` ��B"Q 0�P�AaP�B0DX�B+E�$B
�DX*B*E���T * 	P� �`� �
�P��A`�(�Q#P�
DX��E�*B*DX� @T"��Q
�E��b��� TU�� ������ ��PE^����
���**�� �������
��� TU��**���d�Mef�Ѭ)�f�A@��̟\��|�( * AP�P
�� �h�	KF�ڵ�v���� ��� (J@(�R�%U*�% �$��X�HB�   !$P�M�*@� يEB��@   �� � G�/t������7ͫ�\���@���(+�l���ͫ�����sۥ. :8u[�����Ë��=����7�;t�ԍ��W6������R�.��B�����ک\  �>�� ��A����>�j�l�ngfҽn��R�� �+{�J��*̓�s�t� }�As4Ww:� c�}����t >�ڔ����>��5x}�;������P� �� �P�@m� ��� O����L����˶�۠��=�S�s��s�fj�;8�@r�۾����x�{:�o6��p�ܪ���l���U,�������h���Ҧ����;�z�کp��� h��H	q >}W���.<�t(��t�;�����馛��PRݹ����P7,��, nR��}�z)J^w:P   �h��t�J�;�(4�c�
n�:)K�ҝwp(���AJ{�:i��Х70: �ΚP  � ���  
( �y���[������Jn`����^ۘ�o�7bҖa���X<������w���a�  ˘ۼΓ}�@z�;�;����`��Lt3o;�q��`�}a��  ���&j��A�F�"x�T�&����&M2��R��"�  ��U��U= @���$�@ 4 DHSeJ�� h�O�?߿������c�?��|�;;�w��9��
�*�5���*���EPU?�*���`UQW�UEX�
��O�IO��B�����HBf���a&�˭�)�jX\e0��Mַ���i�3{wO��[3a��(o��sYp��/?��J'>ĝ����ӄ�HH�W2��|�'=X��&�����:>�䐆�~g���5�B�@Jf��Xg!�B���\=��#�2L�f�NNnC��fbJ��He�g3$H�,�w�w�f�˧T`Sv&7t��[p��֡]�sRXl���]noi�C�	.��q"B�`K�P�H�di�!LI�� ��K��H�"B�@	H�`8�ґ��`P�W�B) Fc a�!@�7BRV!FXA0���Rɨ\`��-Ha1�D�a ��)%�`H�
�*�h�%��HČk�LKLH/�"&0�)*���ộJ� A"H���[���y�jD�F��� �!J(P!`4��E`W#���`����M~�ۓY�i� ~�� �ŤlP��\LN I!� @�@���`jm��$HF�)�A��4�XaBa�08B�,/!��g�*��b�tC���nć.����!x��z�亽~�F\�m�}�/�%6��9~Ɍ)$1`��m!��ā��.Y�d��ºϾ�)�MԔ�qѠ�*Rale0�"kZђ���B0!(n\&����n��qO�E��H�'�]|�~�"B�HXYHR B�H�4�%%0��`�ee�#�%27
d�ȳ)��۲B�E���R�I�ۙf��0�A5�MBr��#���-	BQ� ���RX���JA�
���B �(a�0ٹd�	sC$i
I��SCx`��#B1` � �HR`�&fC \+L�$X�4�)�&�h����$�NԖ�R*#�\"�ywg��.�3�{��5=x�!9��RH�5&�ٚ�i�!FI4��h��oߩ-	�3 P�0�'�&�]L�$%r%@�A�Đ����^�8����rF�!�j`C46���v�.�z�M!�!�!&�$h�o��F���a�7������,1��t7t7UH0O&R� r`�d�o����'�P�g��.�s��'����).՘��|,�����/V��C��R3.�sD]��.���k|!
`ʢbn\�{Q�E��X9D!��T��Ӿ���!��s��F�PѸ2)fq�0��pi�ڌ!w����N�E�?f	���G��c	�!�
C	�uJ����}B�E�<JdB�"<���Ra#���IV\p"��%"�!HB��$��"a�p���u�YYs�hѲޖ�w�C�����MK�0�XT���(Wl��q�a4�h��Lu(�bA��!f!��C	�B1 ��6D�57�(q���'�]@Q���B�<iJ!<	q�))IK
�"�2���X����D^�J"�*�i"5�O$�Lh`A�
`B���a�	�@��)5�q��04;#�"B$S5&�+
�0��0!LɁ�&��`?"�b�ZO��B514�hp�ġ��*������*hx�hB��!R��H�`������p?����4l�T a �/[k�پ)SSr�y�I�{�ɪM�9��C���?�`B\q7�Ih���ia�Sx�2�憖��,6S\ɽ�adH ��`B�B5R	�A�C���	!��s0��@�%���-��h�ѩB4��V�і�-�@��Ӡ���֝��@� T�7���X��[�jB�)H44 V�G���G|H�q��$qXP��!d�\4�H�"��"`�*!��x�� C]���{}����TJ2"5b��	��C��&	�!!(����$I3eX̐ �A
F��M���f�2��GkNo��JS!�Q"ԒBB�o_pː!�������K�@�x����1�岌�熓�Hp,��˲1�Q1���I,hCP(qH%!M��X��t?�&�ČIT'*��\���8�0p�����.ٔ&d(D��"F��a�٦����m���p!E��,2�2! ���10c��c@nH^$t��Ƴq�t��Թ�c䟰%�M��vhp�$)������4l��09�/̦WH)�cK��I�R^(p�Û�����?'�O�	��Bj��S֮;�MjE1:�^]�;��NT�P��Ź�!�V��g'�2�"U��I�BLY	���!�b�K��i0��&��W+��<֜�-Ȅ�$8��ۂ۶��`���ٰ�@rW�3�e%�6�[��b<��r�K$7<�ܔ|��
]��.���k[�a�Q�h6E��b\"S	>�����%�.FÄ�?h&�����a�n��sb�(� ���[�[��;�s�k) �)������Ԧ,�L�Iu/79��4�s�F���!� At�R�!V$eZ�q���t;�u�e!h��M~��8l��C
���4�;j��F�H0�[J�\�,�'��p0������v�R
�v�#%����yGkog �y��K	��H��ݏj-U"U�eQQ˄���#�e�����N/�������l�: �\(��ċRF%�~��$kx.sKpӚل;�-!�/9�f��*j̉1F�Z3U�h��8�k��
�ap���K�f���d�0dnh�46n�K���]����fo�5� ��J`CX�%�l�x�3��?3��|CL$F1+�aU�>����n���B@��.`J�$�(IB
Ro'ۺ��]i:&}�~�\%��M�4Ěi,4��^K%��ya�i)���!p��%��`��C�eK�ȯ���f�߿�x�fn�aE�v~�92��7�aX�#b�4 @�3*)r��Ǟx������ Z!`���Q���d
f�i��$ ����-��\akl̆F[�^c2��\ւ0ͤɕ��ki�y��&kK�+Zl��⺄�����s�9&��A�!��������Y�
?sۜj�Yw�D?//�z�����x��1������0.H\4`�ƬX2��c�5�9L M�$.V�!��J80Y4�(0t��y{�q�n�M{P��15����ĉ��	LX�1fN%��W'���HM;���DLr%w<C�]JpbL0�e��� ��㟂��ɟ��!��N2�.~�.�&���;8�%�ܟsFЏ�D�)�
��=P�Bر��^�a��\1�_y��ana�6%6����f	X~������r�w���F�a�$0ff$i�*J@��)c,
�0����Q��)1��6
G��Ŋ�š �4 �Z�!
`ĢB� R1�H�Ė`¤R�,b�P�		$j�,.E�0�F,&H@�	0% d �Z�h�a7`@4�6��)F�&��"��]	%�C��i�!P�LHa�B� �~�<1�\.@��bFN&��%��eѣ
E��/ �L0����0�NkA���W�ƚ��%Zh؃h&ӊ�2�%�&�e�maJ1�(�Tx��&SN(�`~ ��Q��"���,bPH�c�0��L4L 4H5H�`�Ce��hDt�(F�L϶�S$t�!��BS����6��1c.ė5�$�I��C�W��k{B�M#�́%����]@��4L�k`FBi`��\��9xp�d�r�%�i�({��[i���I(���`�w!*�� �Đ)Ԧ��oL��q4���d�H��0?E��v$��?;M��a�!@�o�3�ٮl�k9�7p�,�
H�I�!LaL
�8A��3Z�B#F%0��bK�)�bD�bF%q�܄�:쑒Ff�!�ː$$ Hń��B�t��b�ܹ#�e�2}Ӻ{����o��    6�  m �h    �` -�$ �`     m� m�5��>�M�g)l�1�v�W��]eu��2au�$����9����� l��:� �nZ� 6�     -���m�  �  Zl�    �-�� �Z �  �p#�ӟ�H  �@ Mgk��h ��i&��	S(U*�UT�R�"AJڶ 6�����Hp [F�	  m�m6��pm�m� ���	TsO*�@UT^e��(�9�$ɺ�Iu����L6ܒ͎��% ��Ŋ~�>5�j�
중όT݀�QP��kh-��$H�a�!�l  ږ�k���6}��>6� ��&$��m�t��H9�m���6�Nk�Đ��ڐ�9m��  m�� 6�q� ���`  �e�G���2�P���j�;WK6��t���]�kn��U�v"z*-h�j�L  v�8.��cL�[u������ȵWJW�OD�� <؍�#�H�h;i�.H]�P��Um��S��^:v���#T�WdZ{8�m��Y:���(:ܖ��N3"�iu�+v�/K]�5;U�!�;����Q����CeM����.7M�$�V׮H�8	�t��c�� ۤ�m������΂N�-�h6N^_+Um��6���tK�]�ē��^c^�ҭ�[��Ň	�7 �,�j�� @]7�W,� �Su���0W-m pUPkJ,q�JԴ巎	 Ŷmq^�[�R�Թ`T   h��ghA$˶�ā�6�v�;[OBF��@���.�x,�n��7KsE
��[9�N��Q�FX� *�1S��x` �5ܚۉs�in� �; ����3���T	(���������lKn�Wl$ xl �;q�u�:[($IZ�nl:@p�m��ز]��A���[Uu�T���/Z�0� ��gk�@�Wej��G��Ӂ��m�q$� ���u��r�3�\�R�Àu�xqm]�^��� $�ڥ�닳*��6�8�W���j@�V8(��ӝ�ki�U���[H���
��J�7MOcg�ӋNN�Zn��Hj����Ӳn�gk�D���d����tU��]�����T����R{��#�� 5,YG��lp���v��R: �ZmmCv7/k����.�@q!ݶ��u�[),�#EӖN�2 �x����2�UR�4�*9�*����U���A It�w�}��ΓW,7FW�P���HLdP�l�P   ��l�l�;g�p����m�.ګj���eP��M�ª�W���^�z�$�	�u�Nɭ8,bA׭ m�m$��i�J�p�n���*��x����ݵĵ	�iI�Uڪ�@m��%h-�"@[xp_[$�^�e���-�:�Dr�P!Z��*�.�� �P^m@�`   �����8#��PH���ȶK���nė��ֲ�� $>��	    n� ���-�N�t��ն���   Y����-�%sg����f�5E^���K�(m�[@���X��msE ��m�I��蜑p������Z�ۙUZ�T���i�c�#U=�w;��޷����k�����z��$�v�� l�n̗t�k�����v
�[t�v�E �[���\N&��
U����%��q  8Zm  W����S6�*����^[��{ uX���ځmp!mr%�m��-:��p.isi6�6�h��Hُ����Ř2�mpHU���ly.�r�����*Ղv҃�mPUs�Ӱc��2�C9����8SQ����Ume�r�d&�D�8-�JQ��x��x�]B*�;c��S�g%J�U� $(�]�n�ðE�87m&�RP)�a:]]J���]j\5�7NYf� �jۜ�WyX�'�t��[s[3v�5]Z��1�"s]x&��
�}DP��#ۭ�KҶ�l�˲l��vhw.�*��
��m25]+<k`"ݸN����J�u]Ī��ƪ�e�5$i �ɶsmz-�k�$�\dV�)��ԫ<� Ck5i8���s���P@����<o��󧃆(
���cWM��㽜��y�"�muU\��Bv��PC�ɰKUr� �n   UY��:��a�4�����\ -�K�
�^����I�m[p8]6A�.�f����	o]����8��X5�E�  �H,�N��m�ჶ�i��lත��� pM�ֱ�Ā�n֍� �>�i;	F�\b�mu�p���\��+`�$$6 ��Kh  �a���hf��W�2[Cm�]�m�!"�	I� ˍ*��l�+m�5��gn��n����V�p-��@����[V඀���6ݜ8���8�6�[H[��8[B�;m�бv�iŷ��ܶ�  m�l  @ �Ԁ��h	$��m��m�    ����j��l    6�`	 vݰ ����K.��h)��a�!��`���n�a.��Z�ж�XE]��iu��p   Bڐ�   ]4�n�"@ '5��ym<�[���5UV��������m� �m�m��$��H�f˛l�c�� �w�� h*�iV�V�W��:��l���%��[Z�8N�Cl� @��  �}��[��nձ,��@ �^�y�Ãm�m $  p6�Xbޮ�hlN @ p[~�}��~$�h��:��Ӱ�4Y0�D�6������%����Ci>�}��,�-�$a��� Ե!mm=4k�B�rԫA�t�vZ��U���V��hY� X�UUT^���G=�+�U]T���v�6i� ���\Lm��8���$ m�  ��<�*�P<�C�]�����m5[[*� �  �8���[M���n� �^)m��H����n��� (y���wV�R���qm m�H��Z[z�X�`�Ͱ   ��m�}a�-�ۮ;Z�Wl�c���z�z�� se��6��M��I*�vY@���T�c  �/  �� 9��}� �        @8I'6]v�@Pl@�PV�5UV��l�6�0�e�@�j�r�����y�v� �k�$�m��ڶ� u���m ��l�5�]J�+UO+TO*[S'3m��0[d����n�i,���ͶH
��������¬���㝱V�H�d&��K�/6�
�
���ծ�᱋(�T�R��UP 3kf�[Ɠ8�v��]�ղP-� �m$�m#m�[@ ��p�i���.��7k�V��*ҭrƣ6�P �mN�֛-�%��*�qv��MO+V�Z�Z�`��is\���\���6��n� sj���y�, � 7mm�\ @	6ؐ�6��&֛` ��n���n  ��m���+fܴ�  �۶��YS"��Tm h-��%���օ� -�$��6�  M�� �M��m��$$ m� I&@������u�8 �m���Zƴ$[\ �lm�m�    6�@$�[@hu�M ��m�H�Y�xI��  ���Hn˦�l�Kz���� p� 6�ڔ�����b�y�[Pn���ܺ.�X
�l���U�U���V��Xض�` d�ݻd���m� ��Z�od���)�l�Z[��mi�] � kmڕۖƪ��ڤ� ���/H��䎫f���;s�m,�j�Ui:ؘ
������U�)Xb�y8�`.����aZ�K�")��d�m��2�����[�L�@����m)P� �[R� �\p ��&�   l�sk�\��  H  l�A�kX�U��w��ΊVV��^��@   �  �M�s}�� �V��d͝�薪�UB@h�m�@ $�u� 5� n4]�@���m����@ ���`]�&��m�������lm�` #� �@ 	���c� [V�$8Hl�H�5Q�;5U]����T۶� 6���c�-��s���:t�^� ��Ui$�ioSm���i)h-+i ��&��7i�fd2Z5-m��biV��+e�,\U�[j��.ì,�0�@sm�y�\D�.� I,�;]�NYF��%�m�,�����  ?m��$�l �������c�А �[p巀��  ��l6��`� v�@��h��     � -��� �$ -� .�-�-� 6� p���� ���� G� �$6Z p �  Zkd����;` p$�m7��{��{�����������b����@����?�*�@W*�(1���D�B:F% ��DCH���]�iAڪ 
�<�<x| ���H�P �?P�|"� �S�"�A�����"F�.��O�0J(0��P��|�T~@�����P�O���C�@4���F$@d@�����R1��B$�#�`�!#���0��`
�����(��b/�'���� �"� b��P�
?�@:����t�V @��m 4~:`:@mN�AC��TN�|��"��+A �\@����� �X�QPЏ��������v1��J�"��TU����"ăf-���ВEh�H�$�	�Uv�:�rm�gZ�`r�愒9wM�g�<�P�-Ɋ�
1�)5H�vv۴�m�"�p%��s΍�iD�Q\=P�nH�g���etuN���ҽ�h�/3d�C���k�J�btv���yq�9�Q�ܫ�z6�l�f��sqI��mK�����s��Ҕ�U/On�Q�;Ƌ���cA�OL��Y�9˱Mp�����8x@b�s��vxûv�Y@#���rZ�&��jz^7Gg%v��\�8��{k9Zf�N��ld��j� �YU "Z�^^�[2[�&��øb�jn�^�4��J����	85ӷ6Z
�JY�Г4נ	8��vvٜ�IX�RV�F��]�ܑO':�A��)�Sc2���J��C�*��s�.�wa�s�<!�rc=t����Iϖ�=�vۚ�ۜ׌�8L��&�Jc�;����L��h��sێ]8:��{ml;e�9n-����3UI�{gx�9�k�d�lp�m�^�R��Y���c+6{�WvX ���lv�;cX�0��n�'=��O6��i�3���GF���eS��izu��b��<�U<X�y`�l(��δF̻,.��v0e�T�Yx��5K�r�=���c�]�y�۶�;�+�ۤ%y�"�=��P@;�Aڌ� 5GR��,�����&2�K����ke�i���!�%��Y�� 2Y�Ж
҅���3<�ogTq����ۯoVM�g���I斡�m-�{s�<olh�-�E
�#	���I�L���I�;#< v,�����+Ю��۷ �ge�!���b8j��ో�l��PPccV�����yݳ�n�]��l�O<r�K�-�������f�˰�5W�U^�Y�:86�:m�A<f���AZ��s�bLpet��iZ�K+���	��5���&�w�8�[;-`�fݒI�iΡa�h��Zs�1����D���N��ʭ�r��jJ:�P�Zѭ֪ ?��?��PX@$ "��6"�P\CO�N|*�BO�j�3&ML�C[a�A[I�)tv�(`o	�ș���6�c��b�7���h�auk������n�+Ҷ0�8"cd�v�֓g�]���]��p�Onࣳ
X�1�Է.�lb �F�lJ+�K��K@�'[XC���Q�K���a:�n�M5�u�[s����E� unGC<��1ZE^��`6ј� q��)��������w���E��=��wg'&wa|��.a�pgn�DN;s�i���R{%��?v��<�(����f$�a�N����G󣕊H�$��=���ߖfbl���=��|�o\0)��m"�M*Н;0k�k�`޸`�.w["ݺ�o�v�k�o\0w��,.�)M��S�e&�`޸`�.��x��X�tJ�F��:�i1eu����Z�&�<f`�,5�%��+):؊���N��[��'�{��`�����`��`A����R(B�@<���q,�$�D��UO�蠜��w� �}���r�$Jj؆�1;����,��,��� =�/ ��t��_�E�N���}���ޗ�{_E�w5���;�n�����ޗ�{_E�y��^��C�HG��+�jU Eq�9���Ց�`�BЉn]u�m�'̸n�[�7HZ���c� =�/ ��� ���@󜯯@�9a�BK���9n�澋 ��� �u�����	K��T��6@�NJ�=��y�Wצ�X�DH
�d�� �`�3X�<���9;נq��>���hWCWv`� {z^�}���s��o�J��P�נ{����,yȰwZ� 7������e��k�tgVc9(��'����y5��3��vy�Yp-j���fZje_m��n���"�=�j, ޒ�	�7N	�Z.�wv��"�=�j, ޒ�k��Ƣ�;��`�+v�wZ� 7����,yȰ-��[T�t5I]&ڵ��^�}��n�ڟ����EAj�
��ĳ7�]z�>���BK)�����X�`� oIx6��Yr���`����6F�����6�g�mՈ]��9:�.��,���K��ܛ��o9��Q`�K�=���9ԥ4ʷi ��۵�{��X�%���`�G�t}���l�����X�%���`�G�{��XP�J����&'ww�n�� ��<����/ ��ԺJ����e��k�=|�f��ĳ��_��wﮒs�}۹'#B�+ Q��H4��*e�$`�"�!4B�9�i>Կn�[�[�l�"X�ɠd:�u�sj�bM��,@��UB	j���z�-�	���їv�nNVyw^p7*�[U� ��nZd�v��W3�t&�8%�Z\�K�wF81V@��,���ef�����Iq�q4k4�2���Q��E�pv8y3{<u�c;3��v�N.Ѻ�R�m��ӯ���{��q�j�=a�@z�t���m�,��J�[/e�ή�#<9+/U��U���4���jnV��ݸ���)_X�;M�&K�vݿ�-|�zK�=���5t� ��R�k��+��V�zK�=���5t� �u��	%�&��v4��n� ��� ��<�֢��^s`���)ղ�v�]#�<���d��{_E�j7�Ji����n���G�$���,������~��ɴȭu�]�؝�[���z4/oI[��6d�m�s{P�`/L���ӵe� �%���`�G�yw�C�������&&�� ���w��B!��8�-����8�ó@=�{t;jm�u��m`�G�yw�Η�{_E�{���C�R���K48vh��n�}�dx��[_��%I_��w�:^�_�o\�x�� {���{�|}R8�!U#�,e�U�+z'm�ů;.H�f-�����f�>ٻg��М�r;������`�G��%�Η�u�}�	LQX'%z��ߖb�߫�A�^ w���=���<��R������e��8v���n�,�*�⢇ʳY�k�rO���nI���Y�մ������|�f�糝z]#�w���SLe�����}H��ļ.��{���a��h��I����q�A1���6���*�ú�x##�/WF�-d��`t� =�K�"��}�z�:�aje��%��8v�}#�=���"�}U����]�X�h/�l��>S��}H��ļIl��m��L�����ok���z����'>�w[�ρh���۳@�� �����(�����< �q/ 7�^�}����-Q0T;WV"Q��� yΝ���,��\X�޳�+CSX[�e�F�Ʊ�	FZ9�P=�K�{_E�ywG�z5]MtN�l�B)],�9���X�g�s�j��ywD��II������w�n�� �� ���<���=|�]��X���Q�k�<~�@���< ��xtVȨ�C.��uj����K�<�G��/ ռ��9��rIإnUr�b��e�3�7 �ҔuB�5v��@�Q�n���z�<�i[�L�ru��N�q�eC�N�P�6݋1�ݮ6�Bz+�[��M[���k)찀m�L�s�mR��4!�U}ٮz�)��F˥�!c//%�%Hv�8��`�Vn�}v���}�B��3��j=��M��`N]ܶ ��m�^T���cK�M����%�t�mr��>�Nq��=���ݾ���l��s���(N(+�3�쓽�6��k��[��k���uv��$_�� ��|�w�����l��I��2�wt�(����K�5wG�ޗ�yt� ���S�6���������`������-S� {��t3�!�V֚n�Yk�7��]#�oK�7�E�z5]J�N�l�B+l�@���ff?y߯�ts�ޗ�t�F;���*���.�����Ý�[��Y�SB�F����p��bm��wLLn�� {z^��, ��x�H�]K���
�zֵ�'����@(�H��?~od�T��w����QQn�]Ֆ�һ���^��<V��y9נx�����U2������5l� �} n�x�l#)4�+��'o ղ<y�X�%�|�f��$�3��k�]�������-q�\�9��O����.jz�5��f\T鉫�0�Sn߀��� 7d�ˤx����
Pʻ�J��;�x����S�����Ϣ�=�&�'l�ʙ�Y�x�����{4���<�"p3ƿ���3AM*� �&:t�:цhe�ce�jb��Z��ha�D��Z�1�(�T�0����ok��]�����Q � Ml<��T8�	�j T ��x���U���*�Z�k�<���"�Q	�v�ݼ�dx���[#�<�G�lq�t�]&����+���j� ղ<ˤx���UW�������n[���^Kd�a��xx��'Y�W�w�5�%��>݋S�*FӂnutM?�����<V��]��[�U��¢�T٠x����,l���M�O���Y�G�[�I�j�(������z<uȰ-�����:bj�-�۷�jޏ �r-�9w��)�(~QЀL��7 ��BR�e�T+�n���G�uk�[#�<���պ�]H��m+��D�ͧ�P��@�6�U���� ��?��O�7�#�M�.c�]���������<Wtx���H(�n�mZlln���dx���[��]$�<��]�����Gm�@�����.��[#�;���bV�uj���5oG�yt� �����@����k��UT��;٠yt� ����U~�8D��]�M6�kb�X��ͣv���ڎ��3s��r���ջ`@{5Wkt�on�:1h�����Gɫd����8{n�%��y�s���޺�<�љ�K%î�c)(s��nMϓ�h�����WQ�=�l1���g���<�%d�*r:k�ẗ́Hh�MEU��#n��I�딡�j�;crp���l�b˹�]]���s�e�[��w�>��+[Km%��x����0�vsJ�LR��%�mejA̵��R�Wq��*,�?���5wG�ou� �����S�&����M�x���޸`]#�<�G���Q�2ݪ)]���ou� ����<Wtx�UԪ�����:C�0.��]#�5wG�jޏ �AD��;b-����<�G�j� ս��<� �eЩF��^��#9�8*w�fA��v�wB�[:z*��u�MV#��be�U�[���[��]#��_��W}��$��_0u9)b�Ge�@����1%���{4-����ϩ#WE�Yn�Aut@��T��yl��W���)>x.��v�D�&��bT]v�[#�5wG�j���<���LM]1���v�]���G�yt� ����g���m�U�<"*�bW�7t��k�N<;L&�02�˒�D�9(2�\�)]���j���<���\�f��c\MtNYT�Lr����`�G�j� ޓ+ �A��j�VHIm�����=|�f���X�{��\�Ii{�ՠq�����m\v]	�+���j� ޓ+ ����xs�����v[��j���7���>�߫�k�|�)�� ��D�S���N�p�+]4�l�W2�,�	5(e�2F |ʛm9�Ʒ���R���Α��$�����B��I-}���%�f =�0\�8	Yi����ω$��G�$�9q�I%��?y$���Mq6+5��m�� o�����^�Iy��I!t��$���B�)��QJ�ݿy$�ˍbI/>���$.��������@?�}i;`�L�t�I%��?y$��;ĒZ����K���x ��ڷL�.��0�
ํf僛�~�>p�2;�ݍ�c#jgE�h��j��fخ�hln���I���$�����|o�o w������Џ2�T����I-}���%��OIy��H)������t)�3V,×{����$��G�$��Gx�K_t~��}�ȦxV+.ٻ���{����Ik��I.]px�K��FRb���@��y$��;ĒZ����O�����~Nw��lX�:!{�[ecE��]��]3�ff�q"�9�f���Z�+a��Q�(Q�x�>�ϓ����
c����C��$��W<���v�\
�p�Z�����`�<د;��s�iru��"�Pr���4���TaA����t�+���t���:�1۷����M�R��%"gv��/6�.��rRbtݥ�XHBLΐ-'^�ef��Y�l2� ����'4䓓>i��a���PM��{�M�u�n1����v�؜�F�n��N�g��Aݧr�~���?y$�u��I/>���$-��$�'���j��+�����7�Ϥ~�Idw�$��G�$���H��f۠����{���w��?�6�����J|��X�J9Q	�[i�����$�iϾw�$�����K��K�?m�������7��,�*�ĒZ����K��,I%��?y$��7���o�]t1�r0
f�"�^[G87V.�v�Ƨnֈ�kmtm��k�?s��q��CdX�]�����O w����
}���'���o} �~�yg�]4Mk5.��>�s�8�8  ����K�/������{��[o�ֻn�����6"ಲ�;�@)�{�%��?y�ܗ�RĒZ��?y$�u�Gq2�k+��+������@>>{w�$��G�$�[%�$�U��Q�1]�R�wo�I.]px�KϤ~�I-r[� ��}����xe�WX���u�NN�h���iz"��o8�l�Xz���!��[�3n(�w����{�����I-}���%ˮIG ��m���6Wy��������9Ͱ}����@;�m������N�N�#ʭ6eG��}�w��}������~�����y�{��~�> }+��M��f-ݿy$����I/>���$-��$����������]��0ˌ����?y$��;ĒZ����K��$���|vlivՎVj))B/���Z���a6t��,]4��gq{�O4ˍ��o�I!l��$�������'�$����} �|�w\L����6�| =����%��OIy�G�$��Gx�IW�|P�Qm�e�]�������B��I/>�����	�f�ͷ@�w��﻽����| 9�}��-� �:H��@"�@�4�R ��0 .	XDЪgo;������ӷں�6��w��S��π����K�\$����I%�4�������/Gf]68��(.����ѝ�Ea�C�j�cv�v�ܢXL4Uπ�﻽����$�����W�֒}�I%>��w⚙K��9w��||�� >���$-��$�����Z�c.ۺe+2훼 =�w��@)����_t~�Ir�Ē^p8k�q�b(����$-��$�����\���$���w{���S�k�k+��9� ���I.O�x�KϺ?y$��;Ē[>u�2%dR��,�-�XB�-Yk"# � ��*��@� FbF I��� ��#D�a�u�"�R�ee�$HŁ%�4@a�.0�0�)��#�)� �q�ј`GV���Z��a�d��D� �k�8�H��rBi�$]�J�$���*�65%`�RQ��e)�#P�H�%A! ��X��.�����l%e���� H��A�9�M�Ɩ�
P��(D��G`��HBI B1�H@�@
�,Xa�#����e�1	JB��`�B00H�E�Һ7ld��$���0\��Jā!H����[B��B q��K���Ip%��RT`�b�� #_��D����(�%B$�V0�[���22�W�F"1� 1�,�*F��w���I������Ͷ Hm���l�;fM�Z��^	 �˳f�W-Ux];�P3�3ZҚ[��Y�@���0[w16ɲ�v��n��8]��j��Y�@	i��[hԶ�0]GX��rv+�3�Nv�゗�n�it�ٸ.�Riv�E�����aD͈��5D�er�gh�s���E������;8�r���r�
ݵ��k��wb���j���m�"Fy��Ψ�%��v@�<]b�M7X�R����8
š4ٜ�QA�DA��]C��G%e��e����@���mG�5n9:�r���[���e��uX�۾@�������qi���t9m6�쉡���;(�ɶ�e �-f�f�aHQ��n���hq�I��]! �օ�E��48�6!NF<��m������(u;u���q͞�Ռ螧M۫"sD�ˡ�n �1	V\�L(-�,	1q�+��]�oU��ӭ�7R[�v%��L��r�:N�y��X�ո��]��f���򅲥Pu�=���j�l�HQr�zA��5>�cX3I\�;��m�8��W�6�:mR��Z[g@U����9��fm�pT�t�jE贊cx^6Ef��d�-���kbV�bp�b���w�F�`X55+���P���F����4ތaڌ®�QJ$�A��6��wg��7.n������а�'h�6a��E6��6 ��l��[�\�sv�u�	��C�Y�����;[v4�@�i���"M�M���:����=�%���ug��=��PƦ�W$�E3Ӹ��^88`�Kn; ����"d���
�X�`���胳�	�l��S�����-�^��(�45J�m!�T��;Sj�}��1]��dעʣZ�UKۻbn1�CjN ���fkRmNJu�&�8F���L�C>R�Sŀ@��ug힤�;0]t�v�Q��]ڪ�Qt��Nl���J��D���8[��׈����.L̷Ra�X�@j��"8�z���#��'���ְɭSVU�@uF�ۖ�:�F0:Rۄ��B���B�-U��\�c�����L��k�����T���q�w�%��R%mY���!��yl���l��{p�r>��F�g�u��\�㎊�l�3��̘���g��Jϓ���=PV�v���/볂5��6c�q��:q�ɒ(4��H��|�f�h��Å��M�ƙbەI1p� 0C ����;\�4�]7)�s�����󹝍=Й˹'^8��yZ��0���q��|�v�w@���I/����Ē^}���$-�s�����} �1��
E�.(Y\��~Ns��?�bŒF>����o���=��w�� ����u�6��_��B��I/>�����m���<I%������}�w+�ahs����I.ND�$��t~�I�w�$�e{wJ�kVa˽���x z����H[#�IϺ?ӥ4cM���s9q$<��7C@��u�'v\$ݛ�*�Tݮ��K��-���e�-��}׀�^���.�9ST�v�L�����^U~�Y��]��K�@���Y�6w��)+�����5I��7ze`]���K�9u��v�����7d��<����/ �>� ����$���	���<����/ �� ݓ+{�ЧyOK�U�sU����W���,�.w&�v�}%�:�L���J�*��o 7d���,vL�˺< ��i7M݉+���=Ϣ�7guh>s�@<����%�cgx��>`�%l,Q�k�9���@��z�ĳ�3����Nu�w�z���,D*ݘ�\�< ����=Ϣ�����&|X���$ϩ\�E@��9(I{�!�9t��]��΅R
�Ֆ��ݚ82kE{[^悗�	`�����JMu&[X@��Ĭڛ��uH"�I-�{��j��������}x�TpV��,��=}�f���=}��@=��]�r�ߒ��__A��7j��]��5I���/�~Kd�����:�����I[�9,�C��>��O�w^��~����:&�*A����7�w�f�}ߢ�"�Ӕ�e������'ޯ��� =�^�<��7kΈڹD�a�1��lŖb6���0X�Ԗ0bR�_^ũ�Ϻ{?g�cj��y[�<I�V�< �IW�wK��;ߝ_Y%`9
��Z���o�H6}����0�X�So��[����t��{z�ot��<��4s�7��uH"�I-�<������V� v�x]�Q)�Uݠ�+�0�2�-���%��^�X����K%	,!%��W�s��D/�t�3Y��%ӷg�g=Y�(0]me����v���]��uG��Vu�=�f׏R�p=k�˺N|/;+�k�tff��l��[���W�7�v� �Lk'/[3>]tn�	���X�v{��rv6V�v`x1�\��۶���*��F��- z�8���yE`+��>u�7}&���:C�$�����٦w����{����<o�L�.-��Yvb�6,r��Q���ͷ#��t�/ݯ�o�t��u�\V֜c�U�}���9���yz3^0�{�� ���������drYf {������_�$oK��:O��-����]�v6��)G-�@��^��镀yoG��/ �q*�tt�wf��+ �ޏ =�^�놁��J�d�����U�x��f�{����zL��t��էw#��d��ǵn�{.�9�˩E�l��[]R�H9�$Tq�5$�	0��@=�{t=��&V���IJL��t�E�r[�y�/Mՙ���$9��Z����y���1f6���j���XO���<����/ ��� �����N��m
��`[���K�<�s�C�1��Š_?���Q[i�v��%���`�2�-鼶�{���)63,n��l���S�[�.lk�l�)�ٔ*P���Tl]�ض{;����=���7�e`[���K�;i��AJ�ttӻ��ot�Ͽ~�H������k����J��T�*�<~�@9�{tՋ3s�{9נw���ӭI3���
�]� ݒ�k��2�>�������s�������1
In�糝z�L��z< �Ix�Ќ�Pmt�gY{��s�p�Uѭ;˺�5s��ܖ�uօee��V����ՀyoG��/ ��� �T)�N�ʶ�;��<���t��{_E�ot��t�U݂v����o =�^�}��+ �ޏ &��V�Yb�����,vL��z<'D�T?�Q3>����>���ܥM�� ��wv��X��x�;۠y��^��ff%���(��F�I.�5��M�3�n�V�'nb��с�Vo:qPD��5��CSj�{m�>�����x��X�X�"���*�������/ ��� ݓ+ �ޏ �뤥&~��H��M����,vwV�$�M��ߦ�s�}ts�ga��@�wk ݓ+ �ޏ 7d���,�.��uvU�'n� �ޏ@=�����u�����5f,�1b1NO諒��S V፸�]�ei�i'�>s���nrm&l��u��kn�gh��&6��z#���=�$������{gv1'j�ݫpY?T��O-�ڔ1w3v�i��k�R��v宻GR <j`��f����-t-�r-ÇA��a�-Jxx���t�:6�͉�mѹV!N^r��r7^�����n��e���	�:��)��i���C�=�~՞Z���F�3��go��[ﾕ��E�r��6���X��ncF��VS"�l�|:}x��X�X��x::�U*��۠y��^��y�Z�z< ���Fܤ�Wm wM;�XΙX��x�%���`RQ[wBLM�HWu�yoG��^�}��V����D]5��v��%���`�2�-�������K=�uC�TL�V)KK%+TC��çɮvNR���X�մ�̋u� �z��ޫ�qt��߀�s�nɕ�yoG��^ Ww!F�v�W@���7d�ί��̙�R�q�~��}t=���<}|
��n�U�'n� �ޏ 7d���,vL� �AJ�t7j�ݻx��k��2�-��ӑE�ʤnP����g:�{���<����/ ��2Yt��͐����K3h� "Xm��ha����g.-#�B�h�d�9-4y���<~�@<�{~I,Y�y��_|O�r�H�e�m�`[���K�=�p�7�ՠx�u�"}h�<*l�y�����f�:��I�P�H��`	����c�A4��`B P!�M��&�N���$&��"F)a��A$HB0��BCZ�8�H� �i��łA�cФĄ��ZHH2D�v�!`A�";�8��'� ��~�U�	�"8~G����Qv"	U� �
	��D�����/�~_�Cm�޾ٹ'׽�nI��%)3�v�Qt�����{�V�< �Ix]܅~v� �	]ـn���<�G��/ ��嫍���ls��=:���m���Wgh^����\Z*�;5��Ÿ�4�`[#�l��{z�n���tDZ�CwmZ�o =�^����V� zs�R�l���Չ���޸`:e`[��l��v��"���b�i�� ��+ �ޏ ;d��~z�!�S�-��E	�ƛ��<����/ ��� ��+�o�c�4��Q�y���Gy]��ɒz^Ԫ%�/����KS�h��-�9^#���v���l��{z�l镀yoG�{yS}N�cT��{��@����z< ����
0���:wf��V� v�x����Ӎ���d�h}����4����=�p�7d��uEJU�6ջV�����/ ���|x��V�䀘PB)D*T���Q*! 5�D?쳙�eN'Yиx�	��V���fƺo<�S���#����*���Tjׄ�����=>ٹ�N'�u��Ѻ��i�2r���Ӣ��v����nM�����-N�x;j]�[��
��Ҧ|[�l�����S'��v�۲e�Sa���t�%ӧsZ�;��mб���̇'g������!��Ϛ9��3�F�
�K�%?���������+��n�8��!�y疌e��nܼ�v����-��e�Dv�0���52���~���Cw�V� {d��[j$�۶�m]4�ـn���<���l��{z��N[]�	��Ӻ�<���l��{z�n���<�6�!��]�x��o\0ޙX��x�Z��M[E�wx���L��z< ��x-��D]ۻ��zH�{��z��%��n�2�M�˭�\��8��R��7Q�� �m4}�u`[���K�=�p�<�rJ:TR��	eZ��vn��%���,�P�w�^����7ze`:��*�Sm[�իv��%����7ze`[#�{آ�7A;A�9m�O��(�2����3�׀v�l"�V��t7wk �镀yl� ����=�q6X� }Ƭ!]��(���e�9����T�g\#hTݛ��Lxv���^�m�'u�yl� ����,{�V pC��nRK�t
��]#�7_E�ot��<�G�wu�JlC-���nK4}���=�;�MıfE�$!$bY�KJ�_;�@=�;ts�c}F;v�N����7�e`[#�t��n�� ���J�Wh_��ۺ�<�G��/ �}��+ ��?/���ԕ�Aɺ��;��t��)�%�Yӣ�����E4r�q�m��ٛ�$��x��ޙX���dt�~-�+�j������`�2�-���K�;b��CC����n���<�G��/ ��� 7�Iv���	�cI�`[���K�=���ԌK3��uh�C��:GSxT���K�=���7�e`[��ա;���0������,o$�d����6J�k�D���{FvВb��t�v��wx��X�L��z< �Ix]�I��ݠ�N�`�2�-���%���`\�	A��h��.��� {����,{�V C��>�샖VU#�h��n��':��X�tx�:u?
�
����x��X�L�˺<�dx��:B$R�w�%�]k	�r\֤%�U΍�'mk�0T��4�9��[u	+�W�mҜޓm�1��5s]��&bw3�L�h�d}�c�"u-Ȯ����!\B[�'N�_M"Χ9�m��<�Q��M�[C.��q�][P�U;.���+��E֛r-�����Q�{(lL�p�Ě�t�wQ����ͤ�쁥1ug�/+��F�H�C�ǣhݯ<�Km+��y/$�$_<����Z�J@u0Yu����%��mٲ���Ÿ�B6��(��	��&��l����zO��.��-����`�).�'aCj��wX�ty�U_��#W}��69��7ze`P ��-%t�An��<��,w�V���օ)�5J�]4���{�E�n���<���l���B�E2ݪ]wk �镀ywG��/ �>� +kPJD���ݶ��1���[�%�1�c�	ì�ۚ��ӈ��~�|c}�Y+���(��BYW�z�ߦ�y엀{�E�n���uD�I���*��4�{۸�g���I��s�@��wV���;4��Mu1ܖVGG-�@�>� �镀ywG��/ ݊�JM��h����n���<���l��{�E����T��T6��'u�ywG�V����69��7ze`��bb�X�UN��r��΋ #�@\ƽ�k�g���ۄ6r�tk�k���<�G�{�E�ot��<���;��)I��heV�v�w\0�X�tx��{�U(�[�@+�Wt�=�;�@��%��f,_Fs���=�oƁ���l袎*��eZ�� {������R�>�`���_U�m7n��v��%��`����vh�Ms����e�,W+Cs�Sm��e�sv�v�f2�T$=l�t��}6&�2���G-��=�oƁ�9�Z��x�H��ƉJ�]�J��wf��+>��]>x��� ��� 7�Ie۫��5lbwX��x���޸`�2�(EI˪�п@�?g�}4y��s��f%�e�E�H������nIϾ�>�*�*��f�缽4���}���|�RG���P6��\���vq���y�۲�Y]�Ӷ�]�O:t�%���K*�P�V���9�wV���t~��A�/� ��RG�:nA:ڴ���ٟ��!����s�_Ɓ�w���:&��v9,��K,��^��Wꪤ���WO� w���m�H�%tr[t?f$�O�w~4�ߵh?y١�33o�w�w��3�:�*jJ�%�������w������9��FOL�j$&���!+mCH%��H�b	�������a[!(ƅ� �#�^r]��8�,� '��`L! �1�BH�#	$H]	pa���PG ��p� �|l!0�(��H���)Q,~Cj�D����!�!��4�bD�`��F�"b~LMBRU �	� �D�H@9$�8��`�"B0L��N:F�_� ���Qz�B1��B���������/��m�����9��+jU;\�NnJ�N^ѷ9qI0�:]%�u�%^�cp��[J2/T{v���ԁ�+5@%1a����=8�8����Q2=��3��<�p�*�T6=WQ��Κ�ٜT>�ͧ��\�h�{k�DHv=�����>$��5��ͬ3�NJ2vԻq� �lv"�xNyͶ�i�:N{%��c8`�ض�&�� ^ށ��yvt�h�+YbX�F�Mr�n����ӭ�i�vgXT�&�m5�+�\m�.���RcF���.c2��ɧu�l�f�p��]G!.�Ҭ�{�y�v�v��(F��v��w\)Y�h�<-B��vRGyR2�Q�9Ŗ�mI�T�sY�[eCa�[�TFa��9M��k��mD���S��Q��²�q����5b3��;3#ڙ�j7;�:̕5�D��Yl�R�.i!�f�R���mqM����8 nŭ�n�'͵�vg.oV�]�,�;|��גP�}UA�	w ���g��N"g[h�'���y�j�L����B(���`X%����m��H#�m=�N�RY�N,���6Iu�m�A9܏mȴ�%a-�B�t�S �);P��78CmAdel�ڜs͈Z��r[�m;q��p 67;���>�b@e��()�Ω5B�5G;F�v[����`�۝����-�u\��ͅ!j��I�t�-�$  u�b��.�9ȸ�Rg���T�Ӧ˷���:SNc' �s��B�siR˥Y�R���̀�=�v3�i"Tr���K38�vە�U��U[�PA���{C�(�[Tnc!Pn���d�+�<^��'v�m2nH���j��N43X1�`4U�f6�;��`ݤʗg���*UGۘn]�eUڕ�gںyؘɧXp��j�E�kmQe�Z�����V�sͱA%�mc4������ְV\��ڕv�����]R�H.X������yX�;'L�R��9]lq����x`*��*�â W@4�q*�!,�/�}*`�	N�FZ����wCJ����kX���Џ��A�1��)c��)��u�܋�N�+�ey!��)����\���ۋZY�˘��z�=]��S�\����3�;�ڛ����p&S�y$�U��6�j������gm0��ͷg�֕){�v���Rty�*�m���D7$G���v�3��؁밤��.�x�:0ucWm�P�kN�ɞ�q�O9�#v���lЅ� � �����E)�ARoӜ���<�â�j��wP�|�ӥ���}_�,^0�;�����N}r�A�P;f��:<��,��V�}_�~���%�_!��.�E؄���|��X��x���wP�PʺwJ�h���bğ{߼Z���h>��C����;������E-��t+�h[���� ��� �+ =���ݱl���ʱ#th�����Mb�nU ���3f��7d/�{���ێ��r���<w�I2�-���k�luF�%tr[t}���Inb�?~��V`�ﲰS��H��ƉBr:[$��9��V�����}�����@�;~4����VV;	$� ���tx��)��Հj���>�G ��@��;4=��s����vh��BuF�H����yp�����pCU#���ZU9�����3m�ܺ��Th�,�<�/M��uh>s���xï��4��l�UJ�@���:t��<���9N� �u� ������ؙJ�wu�yoG�r����	�yBE�E&�Y����^������:'�NV6[M۷�$�����X��x��K%t�lV�M�����L��z< �%�!i�m%7L�Yk���Kq\0F�а�1Y5��K���F�f5��G�R])��-�vL�u�X�K�=��]JKv�h���i�`����^�r-��uo�K=4�֐RG�M�^�wﾺ�����ff$�~��Z9;��7z�(���WL������r,{��ܓ����rb�椪8��f���t�z���R��P9k�=�{��n�� 7����X���~���~|��׶��Kb<�[n�:���ik�8g��)�EkT�QiS8ŭ�h�T�����0zK�=�E�oI���R�'+$,�v��;ۿ,I$�)G���	���V�� ��F*J�
حX����r,zL�>�IwK���}x�ƉE&�J�[���X�L�w��yl��|��R��m�.���wX�U� �<��Y$���f�^�b��"HBt��U�����K�O��.�[9���0:-۔��Ӟ�e����m��f�;N1w&�J޹݆f��v��u	r�Yx�F���z�j�x��es�g�i�v�;7��s�.n��Lcsˮ���`�K5c�r���n��Ȍ�	��&�5�	��,����f��csqҹ��n;5gbw��K׶�y����+yV)6ӫn��>�>���{r��؍S<Vy�v�����m㮸��k����9%��+NYT��Sv����4=���=�{����9�|�s�7�pR:��S$�@��޽��16s�ՠs���@��{7��������2J�@�@��+ ��"�~��R+��X��pMI
H�|�1?}�z_~�h�"�6I���R�I�-�E�e� ����~�޿�^���w���o�z�`o/��	l�G�W���V�	�r'Ql���OX�a�0J�.N�q:9m�������ՠ{�)��bř���`|���h�Oџ�����b$��d�Y����H��"�"��r,�����N���gd��\lfym��� ��<uȰ�e`\EN[�$�T݅z,ı>����9���@�&V�,� ���R��t����{e� ��~����}���ϖ t�����_��\-S;3j�J-)X]���w�3��8�g�U�l9�۫I�>qu�:�[M��uh��u�;�߱,K����z����H�cEZ�޲, ���l�`$����U����bJ@�}�g�)N+��߿~�����=I�$ffbP�w��s���{ȻF�w�ҒKf�ؖ?y��`���7zȰRG�M��%���KQ$��9��V��%�wO��q��� ���%6cm��m�jvz���ݻ���a�[���D�#s�Lx睵K%b��c�ʴ}�:�y٠y�oO�/w��V��������&�%l��yN�?��~H���0	��w��ߒı~K�~������J�����l�X�Y l�x;��� �C��[t>Ē}��x�s��h��n���%�Գ��������䩈��@�ޫ�@��˾�_�7����2�	�����WiWi�&ꋞ9�X�P���K-v{vv2kn}�\�gY��`��ҥ�6��)3|������l��vɕ�������U�`�󯘕+��ؚ�7wx���2��W����;7�Y���,JC�Y�	��r���m�>�ߵh��u��$߯��4�}��.3���.�㒭ؒ��wO����~��������>�x�_��}m��70��
�y٠}�~ıNw���w�ڴ}�:��\��~b�t��e�Ijj�q�t�K��=�ڞ���<�
C<�	��u���8�j+4�=mY�d0�6*r��T�k������3ɮ��3�Mf�C[`64b��fIaع�y��㈱��Er�gۄ.�Vh{#�OqێF��Z�뤝�3q��%��d��m��p;ll��=�e�ٶ�������k���3�q^�c��!�k�f�zBB��l6�+�D�N<��Mۡ4�Vv:�����.ѭ�%",$N�"T�,��}��9�;�@��S��,�z���@>��BI�v�Q����տ�f$�9���z���@<����b�l������(K.��g� � {d���V C��Sj�;��l�L��yN� =�^��y�Z,Y���= ����6��-��wo ����+ ��"�<����y�'4���,I"w�]̎ysi��y�:�33�fpK3WO�s�;�`�'%Q5eC����~ՠ{��v��r,V���;��N�ѹ'����U�(�g��� �s�l镟���9||��v蜂*n�M��|�=����f$����V��:�Ɓ�8TuG	
�h�X�z��u���ՠy�)ס�Ŀ,I%>������~�8(9pP9+�=�L������za����,��, ��[�^�v�B��J�:R���M/Cje9���)(�8���5;�f���I,Yn��E 얟�Wu�t���w9�}�wV�t��:�,%���֥4rw�>�UU_�7��`>�+ ��\0j�@u��c��W�y��^��;�Zw2�f����8�����gLU>���/�](� � � �P�(D��4ʚ��&)�� 1'6�$TM�0D?A `���
��x��b�Sb�@�oy�MnnI�g:���#:�RUSVT9ez%�~��}�� ޕ�`��`�:ղ�:�,$���x�M��/ٙU���?��������2�ЗMS�["�V�۵��ڱ�oJ�C
�+��<���6R���3a��*�6������ذk��2���U_��zU�`к�1��C������,d�X��^�9;׿,Ř���~�8(9pt	�X}��X���w9�r=��q�v����V��c�:��'~�z�I���n��ϔ@���@��X�IF�-jS@糽z�Ȱ�2�ޫ��U���J���Nul\mQ�v�⺹U�����غ�m�8:{�	�+DV���,6=6u�,�nց��,w�V��p�5I�{dgSjKP�u[^��w���ı��U�`���{_E�r�R+-��nVBJ�=�4_{٧٘��y;��;߾ՠz���YU�W���SC�/��{7$��w�rO��vnO�F����`"��1ӺiP���,�Y��{߼^�:�Ɓ�gz�����⥚���b��:r����p^=N��1�p^;v���j�J|.�y/Ont]�������k���\S�i�9B���Wl������]��4�Sl[r�]����꛷7U���Kų*�\�&�7V����UۏgTUlv��Ł�1դܨ"njI�Dg-�P:N�s;d2�4TL�:����!suM0 �R��KDҹ��W�L��xMbA��b'�
@���U<�wnbv��g�N��n�y�Dr[gw�ffn݆��. �2J����@�ʸ`�E�n���!M���_��u�nʸ`�E�n���տ�fb���$�߈~d�Ym�֝�?��n���+ ݕp�	�ӰT%�����|�3��:}��n�\0G�`:ch����j:�-�@��噋9�>~��|�k�`��t�R.�Ҵծ�D��R�n�X[mw0)�[m[]�p�A�k�˃�r�U�{�)נy�ν��XoL��B��ڥl(�J٫�';�v�
�S_g�w$��~ՠ{�)נs�*����6�Sn׀{\� �镇߿UUU%�,�`���E��������'v��X�)נy�޽�,I'�/�=��u
"�Bcal�@��S�@���^���O�z=�uh��t��K[�M��Y���ei0s��x�I��:��(c1��tٽ����d�6�ݻYv�k�o�|�k�`�����Ē^0�;O��w��򨰄����7k ����+ ��`��{�KM���l��E-cq�9mz��w�ᇪ�~���E�{\� ��z�eD�8ʠ�Zf,O��ߍ~s�{\��~��S�ެW���Wt�J�Qt��f�:<��XoL��x�M��K��a>�"#��ZI^��)��,:��ƞn'n�sr	b�K� &���y�Z�8B+H0�6�~���ߞ��yܬw��z>� ������+
N�`�2���Iү� ߟ�,��׿�bX�8����DWQ1�YV��*�0G"�=�E�wt��
�D6�ݻYv�ـz9�r,���7'W~$  ?�S���n�H}�����.�X�4ݬ��X���W��|�)#�$�����Wl�����N	�s�B��k<��-�om=�-�G�H�demIk",����uh��u�>���Y�0����?�t��#�%t�wX�Y�$x�Ȱ������&B0DM�_�}4r�7w��޳�n�]JLc�E�;�+��{\� �镀n��`}U���ﾚϯ��2��'-z9���=����<}�f�糽zňY���?�-{{���a�n1nbm��u\E�̌un��ML���9��mŮ�'��f�7#�����7&�Gj�uh�@'��۷�7�z���=�֝����&�v��-q��;�npi� ې˃7�F
�
�.q�G.�Y��Җ�7�lt]pFҧ@Z:�祖�/S��7j�܆�Nm�n�H-����f��ѫ�	�R6T�5���9����O3O]�\��䷕㛤.x�rݩ�Nq�ל��՚��J(D�9��[�Wj�
[���ϖ�$x�Ȱ�X�"Wn݀��L��yI�s�@�9�Z��{�bI�����QY	m�:���O�z9����%�7�v�=���M��#+�ISd�[V�~��RO�Xt��yI�r,�ФV[��I�]4����E�yI�r,��V�k�m:��t�.��5c��N���N8Ti潝%=ڷ`����ND|���YXT���~���=�E�wt��7zȰޫ��Ȫu�*c�h{;׼ı/�̐���Xt��yIu5)~b��aIݬ��V��E�yI�r-�c��"�i%�h~K1%�/߿~r}��`�����r,��V C�3�8�P-p�@�����f~Ifg;��?@��j�=����?.}��`zȚ�DՊ��[�Q[�Ÿ��(��/	�l7�@��j��\�F���|��`�2�޲,�H��1�Z�ISd�[^��s���$�&�s��`���n��h�[��:M+��4nI��MvnI�߻��
��� ���H�)�AG�'�37�����?s�ڴ9:>�h�n���+�f�$x�`�2��Ww��!�;���������X�3?$�%��~�z{�_Ɓ��{4��~ӥnZ�6��m�p=ػd��{ й�f(TY䥮9�ۮ����+mذ�v��X쫆�$~���^A�O�z9`|(���YV��V����E�wt���߫�U$�5�;Il�Jh���h�;ק��������@�>W�@=���SuBKD;M�o �r,��V�*�+�R@��P����nI����Y�e���vP�ݬ��V��p�I/ ��޽��uŶ'�`�W-n49�،��l˕3�Z���Zq9q��3�m�m�b�Һi;�w�� =$�����Ib�w��V�����]�u��5l���^�r,��V��E�Vbēgy�W̎���n۠s����+ ݖE��/ ���%�h�t���I>�x�s�����n��ŉf?y~���}��!mU9���wX�Y zt���XoL7$C����Ab4P�%@������	��P8�#�4�J����`�B@��$~q�5�tC���L��
�QاT��v)R�B ���G�TXAX�HHH@�� s)���B�$�s��e�!$���v{OG��Z�b�۰ ��,��:^'�\b�˃j٪���Ӱ�U+��V�S(��[@{d��㭭��촣P曇��`���kY�"����yLwm.4��`�n��R�p��4�I�ѳ�l��k[���8�g OM�[���ݵ��Z�4)J�����Wk3��P����!M�L�.4ls��\�I��=j��g�,������Ĺ�@�5�W$���Ζ��%.E�t̜k+Xe\m�);G�������iqn^XI��ɺ��z맪�xP�v컗��E�=��A8Ut%ڀ�l��Š�V"�ܯR�h�V��٨� �hҝ0@�f�Uܬ:S)�T�-Ϋe��N#��Юa���)C��M��ypTj�)���n�f
�\�dE@��uXȜ[�J����\���]�I07k��v��j�gɉ%쮊6�n���4�a��hϷ\�v�ʄ�sn��[&��Y��NŴC�y׀�Fj�v���łc�x�\L&.��6�+D�q�]���UN5/�ݶҖ���5�d��Ce@�:U��4���`:HX�٨��in�Fcan���
�yei�(�QvS SZ��j�����C+rQcvh���\nu��]��搷h�I��X��6�9E$A(��tӝ��tҜ�=����['d�mll�c�k�sk��V������+X�6� z4�ŭ�h�2�V����nx�vk����Nͯ	t�=R��$�u�4!�w\�=��jx�[']��v�ܻ0���Y�L��㰻*�I����a��8ؔ���g�"�M�kdd�]�ChMMkp(dT�bN79",����t���n;Fvn	�t��@*��\��&ֱ�eCge���`�U�s�a����W��W�ӱ�7,��i-��S���YV�mu�h�IЃ�Z���� �����1Z�H�r΍��k��M�)�6Zi:�%E;e���6 s�A�#�hj	�fs3Z��Z֍h��|"���1C��:'�S�F ����	��%�nY��Z�K�������j����tj��%�im[Zy�^�r�3�Κ����βW\Wn�	��Z.7�^'��<�;Id��L�u�n�g�Y���ҕ���q�C�4H���k`�y4��u��Q�O�.휆Ns��ʪ�8=��I�uC4r�x���uld�uv���W�(�=���"�Z�r��*j��wE����o�oAl	pT>��N��Hsm�u4�1s�3-Y��i�X�u���2^÷n��#=�v��S���Z�p��y���gz�{���f%����i���k����u��-�=�E�v���7zȰ)#ϫ�W���}߶FV�#p��r����j�7zȰ)#�=�E�r�9®��ҁ�U��bY���=���M�g{w'�{���䟽�ڹ��]Y	�+e��H�k�`�2�޲,-�^�!�6�hiK�c�A��u(�`;B�-�Ė5���)��J�k�s��䏚3���+tR�Bv����wt��7zοىfx��ﾺϯ������N�`�2�?U~H��"��/ ����X�&�S��>iYN(��V��K>X�%��"�;�e`N�6�ݫ�`�L���^�r,����,K9�>z���_}۰V��Թ�ֶ��bX�'��]�"X�%����6��bX�'�ws�iȖ%�b_�ﵴ�Kı?�_���a���w:�+�Y�����F^]+��-�A�ͬ�j7��'&_<تi�5�en��Kı=�p�r%�bX�}��]�"X�%�{��ÒD�,K�������L��]�C��[-�@��L�ND�,Kﻹ��Kı/�w��r%�bX��׽v��bX�'~�m9ı,O����\�a���4[���ND�,K��}��"X�%���{�iȖ8��(@��,bH����H�) �Q,Ow���Kı>����ND�&bf.�0�ʛ�q�n����X�'��]�"X�%�߻�ND�,Kﻹ��K��X��I��~���131~�?���v�	H\֮ӑ,K�����"X�%������r%�bX����m9ı,O�k޻ND�,K�>�x��:��U9�-�^2��B^�����[&�@��4��5�MK2�װ֕�T�-�n/L��X�}�~�ND�,K�����"X�%���{�iȖ%�bw���"X���M}�ƾ��k�)JJn/LKĿ��kiȖ%�b~�^��r%�bX��}�iȖ%�b}���m9 �y�^C���~�(�p#M����ı,O�k޻ND�,K��m9��D�Dȝ���ӑ,KĿ~���131s��䌵�I ��֮ӑ,K��{�ND�,Kﻹ��Kı?g���r%�`~P8�Q3���iȖ%�b~Β�zkY��..���6��bX�'�ws�iȖ%�b~�{ٴ�Kı?}�z�9ı,N����Kı;�=�)���k�\n�+��d��Y�2B-)pV�30.�9�^F��ۇ/7�t�����Ȗ%�b~�{ٴ�Kı?}�z�9ı,N����Kı>����W�&bf&b�;��	�v �c�jr%�bX��׽v��bX�'{�p�r%�bX�}�~�ND�,K�{�ͧ" �TȖ'�z����[�RI����]�"X�%��{��ӑ,K�����r%��ș����m9ı,O�����Kı>3��=B�a��kY�iȖ%�b}�M�m9ı,O��{6��bX�'��]�"X�%�߻�ND�,K�흞�r�-(JZԦ����L��^ϻ��^	bX�� G�����?D�,K����"X�%���7��Kı0�	`,T�
�E�~��|͝2�k��<px�&�:v� �[r�Mm�<�˩�Z�m�hK[s�����̥ͅm{,�d�;KYkr�H"Qa�kiU|T��<�m�k�lv��t�6��x2�����T��m�����ծ7�6{xk#�I��9��؛��Yj����K1�N�s�&���T��2�]������l�fN�!ݯ<�Km+������I��m��)]�4�-�luu��'/c1��H�v�*�ˀx-�ݲ��~��K������r%�bX�����Kı>�f�6��bX�'��}�ND�������{�T�iV�eO9=��%�bw���ӑ,K������r%�bX����m9ı,O�k޻NE1G����V?�Ų�):�r�Ñ,K�ｻ�v��bX�'����ND�,K����ӑ,K��{������������~vyR�-`�'�Ȗ%�b~�{ٴ�Kı?}�z�9ı,N����Kı>�w}w�&bf&b�;��	�� u1ۛND�,K����ӑ,K�����"X�%������r%�bX������������?};w�Mr�����F�X�x�m���Oe�jSi�m<�Ҝ�q�wTu7QK�J	�^����L��]�}�iȖ%�b}�w=v��bX�'��}�ND�,K����ӑ,K��N3�救VE [*�^��������Ӑׄ؀c���b}��iȖ%�b~�^��r%�bX�����Fbf&bk�:�
�JZ�^��Kı?g���r%�bX���}v��bX�'~�m9ı,O�ws�iȖ%�b_z��$�i�Ԛ����ͧ"X�%���w�iȖ%�bw���ӑ,K���w=v��bX�'��}�OL��L��>��G	u��+�9ı,N��p�r%�bX����ӑ,K����iȖ%�b~�]��/L��L�����8��������lַ/Z3��"܆�!�P5e�1/��
��+V�d# ꄕn/L��L��;���Kı?g���r%�bX���}v��bX�'~�m9ı,O����g��`�f����/!y����fӑ,K������Kı;�}�iȖ%�b~���6��bX�'y��%M���ٸ�1313��]�"X�%�߻�ND��p�2%��vo�iȖ%�b}�wټ^����������
K $�iȖ%�bw���ND�,K��7��Kı?g���r%�bX���}v��bX�'�}gI��0�p�&���r%�bX���M�"X�%��=�fӑ,K������Kı;�}ͳ��^B����^��h�\eX����v'g�>��_)(�v:�'<����r�6oksvB�Ue�P%-jS�^��������߳iȖ%�b~�]��r%�bX����ӑ,K���w=v��bX�%������b)I%�qxbf&bf/y{��r�	"w���pI��u=v��H����n'�A�dK���̧�[�G���k�^���������ND�,K�o�iȖ%�b~�wٴ�Kı?}�z�9ı,O�ս�˭j�&Mdə��"X�
$Pȝ�M�"X�%��{�6��bX�'��]�"X�TN��A	W��AH�H+��I(
@F��D�׸m9y�^B�~g����V����99ı,O���6��bX�'��]�"X�%�߻�ND�,K�o�j���L��_�Is�ϿF�D����m��z��M��mOp�8��T�.7.�em���P��bŎn��J��;f����LK�����9ı,N��p�r%�bX�}�~�ND�,K�{�ͧ"X���_N���RX �)-{��1X�'~�m9ı,O��M�"X�%��=�fӑ,K������ı,O��Γ���Yp�&��6��bX�'�tߦӑ,K����iȖ%�b~�^��r%�bX�������L��M}�tʱ�T	KZ��\�bX�'��}�ND�,K����ӑ,K�����"X� !b}�M��^�������_?��!,E)&f�iȖ%�b~�^��r%�bX�����Kı>���6��bX�'��~���131{:3�!TN+3���Ԍ%<=��m�N.vu�F;aB�aƻ�X6����b�c��g�ݱ�Ͷ�Fɇ�bݱ[%�|�Gۊ�%��d㭹�*�x�]Oe�f��<�yI�r���'k�5�u�V-`�m�6�h��*�6�X�%�g?���$�k	��P)n��
��v)Kl!F���]���M�\�C��i��֟!��Ƹ@W=Z������ y{<�Ml�6�0�8�3gыc/\��J�:��^�ݴF�gҩ��G$����+��&bf&b��~�n.D�,K��7��Kı?g��� ��bX�'��]�"X�%���c��[m���$�qxbf&bf/y�~�ND�,K�{�ͧ"X�%���{�iȖ%�bw���ӑ,K���_?��* 8:��Sqxbf&bf/���6��bX�'��]�"X��B #�2'���ND�,K������L��]�t���7`v���Kı?}�z�9ı,N��p�r%�bX�w�~�ND�,K�{�ͧ�&bf&b�w�?�B��C�����bX�'~�m9ı,?�"��zs�m?D�,K����m9ı,O�k޻ND�,K�t�fkXZ�G.�Y���8�>&��G�L�F�To=��Z]�v�)	�k��o%�֮g���B����{7��Kı?g��m9ı,O�k޻ND�,K��ND�,��M}�t�n��	JRSqxbf+���wٴ�7��� ���U�
�'�'u�z�9ı,O�w�6��bX�'��ߦӑ?�C*d��O��?�R9j)I,�qxbf'������ND�,K�{�ND��@dL��zo�m9ı,O���ͧ�&bf&b��l��Y!+,�p�K�U�?w���Kı>�w}v��bX�'�｛ND�,K���縼1313{X������6��bX�'���ӑ,K�����iȖ%�b~�^��r%�bX�w�x��&bf&b����#�a(�V,�Ň&���7mn[N�g��Ez:)u�>Н��Ns���٫�Q���r{y�T�?g}��r%�bX��׽v��bX�'��m9ı,O���]�"X���]�t����da`�,�^��ı?}�z�9ı,O��p�r%�bX�w���ND�,K�w�ͧ" �L��_N�G�RXt���ᅉbX���p�r%�bX�w���ND��C�I���ojZA�VB%R�X�  �Dj��RP�I�0�JP�0X*�(0�

"�V�B�	�b�% c�a �)���e�% `N;��m�D�$"
H���HB�#1eRb�Q!T"��P�*iB��e]���ʑR$`$X�RЊ�� �H�I"Da	hQ*�Ģg�ֵ/f���bD3L���i�I71�*K�$y���aBRP�m�!s�qd�r����)0�000�%epi�����°�*�Ƥ�
��I��9�c��-��l 2�J�$�Dc$[�$%,�"g��E��h�@*J��(�,-C��YF�b�� @�Ā#�"D�B�0�! ��s�1	U�R��Oف�Œ�Aa4�@���A~~]�|
@h��x��?D�M��}�ND�,K����ӑ,K���ل�uu�q�&��6��bX�'��ߦӑ,K����iȖ%�b~�^��r%�`������"X�%�Ovå��[	R���^��������7�'ı?}�z�9ı,O��m9ı,O�ٿM�"X�%���{���~���-�	���u�{f�M�v��a(�5/�ź��ۨQ�l�(�n�fd�ı,O�����Kı?w���Kı>�f�6�E�"X�+��M�ቘ����w���1�܄,��5�]�"X�%�����"X�%��{7��Kı?g}��r%�bX��׽v��bX�'{�/�sS3Y�&�˙�iȖ%�b}���m9ı,O��{6��b�bX��׽v��bX�'{�p�r%�bX��޷���5��ܗE�L��r%�g�������iȖ%�b}�]�"X�%�{��[ND�, 3"}��zm9ı,�����&�í��3�������O�k޻ND�,K������bX�'��ߦӑ,K�����iȖ!y��})����f��]�ng�s�8|I���Ld�a�w#vШ��lh��]O$mΝRIu!s5v��bX�%�{�m9ı,O��ߦӑ,K����iȖ%�b~�]��r%�bX��wn�յ����m�^�������ߍ�����bX����m9ı,O�k��ND�,K���[ND�,K��ã��H�������L��^ϻ��9ı,O�k��ND�,K���[ND�,K�{7��Kı/�O{K�le�)�����^B�rp���=��r%�bX��w��r%�bX��ٿM�"X�%��=�fӑ,K��߼��Q����)��r{y�^B����ӑ,K��������~�bX�'�����r%�bX���}v��bX�'�y 40�Q�@HP*@$$���5�u���� U�i'�ų���sc�콬�-Ґx7m0G�z�ʚ�ÎY��Z���v��d�W�^ۂ�$A�u�qcWC̝6�.�lj|��]��Jr��c�Hts�r��P뭰�:�� v���Ҷ��%[�Ý6�nG�3�8�3N�z���Yt�Qƍ�F^�����<G�Z5MD���r\� 0�nB
������ϧ�<t1�K��&��9A�ݎ�d�u��.َ���&���ӶKcg�9Cr�:�U-��b���L��]����ND�,K�{�ͧ"X�%���w�`"X�%�{�}��"X�%��w�&`���]��'�����/'�{�ͧ"X�%����ӑ,KĽ���ӑ,K��ӻ��r%�bX����ChfeŬ�.���^B���뾻ND�,K���[ND�E�,N�;�M�"X�%��=�fӑ,K��{�_�u�I.�.f�ӑ,KĽ�}��"X�%�ߧw��Kı?g���r%�bX�����9ĳ1w�� |ev�87m���11,N�;�M�"X�%���=�fӑ,K���w�iȖ%�b^���ӑ-�/!y?v���[�ど-q��n��^�c��M>6n��D1�e͵[��`�2Y��&�e��jk56��bX�'����ND�,K�u�]�"X�%�{��[�?DȖ%���o�m9ı,K��O��$t$v!H���ቘ�������qr�$�*�Q02&�X�;�kiȖ%�b{����r%�bX����m9ı,O}��_YMd�2k5d��j�9ı,K����r%�bX��w~�ND��B"}���ٴ�Kı>���v��bX�'�՞�L��јf[�5��kiȖ%��bw���m9ı,O��{6��bX�'�뾻ND�,K������bX�b�����X�XA�a%7�&bf'�{�ͧ"X�%����ӑ,KĽ�}��"X�%�ߧw��K�/'ݕ���Ħ�u�8�ቴ��l��w6��lmJ��cb&���<�䏙�P�F����'�����/'�^�<��Kı;���iȖ%�bw���l?��&D�,O����6��bX�'�x��W&�T�]H\�]�"X�%���~�NC�DH�L�b{����ND�,K����ͧ"X�%����ӑ?��̆(bf/�~q��+�q�m�ӑ,K��g��6��bX�'����ND��E�4��dMD�����r%�bX����6��bX�%=��S��Ӫ2QR�n/L��L����M�"X�%����ӑ,K���ߦӑ,K��ӻ��r%�bX�ާ�@�	�H���ቘ������ӑ,K�{�}�iȖ%�bw���m9ı,O���6��bX�b��X��}���A���BT�X[.�e�;=�s�G৘��k1���,���]�&�VK�֯�Kı=�p�r%�bX��w~�ND�,K�{�ͧ"X�%����ӑ,K���K}�e$�E#v;M�ቘ����û�r�ș��=���ND�,K�k��iȖ%�b}���iȟ˕2)���_���L��A�a%7�&bbX�g���iȖ%�b~���Kı>����r%�bX��w~�ND�-�/'~{-�.*��`s�������*D�����r%�bX���6��bX�'~�ߦӑ,K<��A� � ,](Qn'����ND�,K��|W5sXI.�.f�ӑ,K�����iȖ%�a�1�g��6��X�%��w��6��bX�'�뾻ND�,K�-�?U��u����
�ٵ�!�e�r�i�tVSm����SS4��,X��5�W.Z֦��Kı=���M�"X�%��>��iȖ%�b~���Kı>����r%�bX���vK뢗FY����SiȖ%�b~Ͻ��r%�bX�����9ı,O���6��bX�'~�ߦӑ,Kľ�=�&��&�5�2�iȖ%�b~���Kı>����r%�� `.DȞ����ӑ,K��;���ND�,K�k�����!+-�qxbf&bf.s���r%�bX��w~�ND�,K�}�fӑ,K��>���v��bX�+���YK(�L�����13�N��iȖ%�b?��{6��bX�'�뾻ND�,K﻿M�"X�%���"?��qz~Գ�����kXMV�ʜ̤�����~���.�H�˷W���͵�8�i�NvKfG�.�$1ӒB���'�nv8Z�S̯)����}��i�;�t�&3�;
tv-�{v��ʼ�m,,�Cp�Vb���;����0sC쏝�G��ᇷ:V�n6�{-��3���$�gf���7I�;�	:���l���j�vz�ű�5:M)���%(Zww�e��K=\/F�v�z���˒�O1=��d�M��n8��4�cV�^z��Z� 값��񉘙���?}����,K����ӑ,K�����iȖ%�b{���m9ı,N���ÎZ�*��f���1C1{�ߞӑı;���iȖ%�bw���m9ı,O���6��bX�'��2��j氒]H\�]�"X�%���~�ND�,K�N��iȖ%�b~�wٴ�Kı?w]��r%�bX���?�[(�	-�����L��]���m9ı,O���6��bX�'�뾻ND�,���ߦӑ,KĿq�󩲫i`�e7�&bf&b���iȖ%�b~���Kı;�w��Kı;���6��bX�0���~�����4YY���l��N�����>Ms�@cK����g���t��gh��I���ֳiȖ%�b~���Kı>����r%�bX��w~�ND�,K�}�fӑ,K����fOY.�[�Y�%�kWiȖ%�b}�w��"@k�2%�ߧ}ͧ"X�%��w�ͧ"X�%����ӑ,K��um��R�܊��i��1313xw�6��bX�'���ͧ"X��b~���Kı>�w��Kı>�O��6c�_9=���/��Y5��_��ٴ�Kı>���v��bX�'{��m9İ?��ݞ����K�f/�~G�䖅��Q�,�^����O��}v��bX�'���6��bX�'~��6��bX�'�｛ND�,B����?B鰸Ʉ�2�f�]�X��d(��F;&xx�WMF;��:�$�>Lyd\iu!s5v��bX�'���6��bX�'��{�ND�,K�w�͇�`�'��&��	��r��ִS&fK�֦ĐI�};��OD�,O��{6��bX�'�k��ND�,K��~���&bf&b}�:�T����)u��Kı?g}��r%�bX�}���9ǈ�� �0X(@B*Dz�F����@�"r&���m9ı,N�۾�ND�,K����P��m���131s�w�iȖ%�b}���iȖ%�b~�w}v��bXʁ ȟk��ٴ�Jbf&b���H~a\m�e`��/V%�b}���iȖ%�b~�w}v��bX�'�｛ND�,K���ӑ��/!y;�����7�e��"����vl��O���v�n��N��]xK��*_@�:�L˚�fkSiȖ%�b~�w}v��bX�'�｛ND�,K���ӑ,K���ߦӑ,K���<{W5a�[r�E�e��r%�bX����m9 lK������Kı>�}�iȖ%�b~�w}v��bX�'~�I��-#
�rY��1313�����bX�'��m9ı,O���ӑ,K����iȖ%�b{;�/�d�ֱ�ԅ���r%�b!b~�}�iȖ%�b~�w}v��bX�'��}�ND�,� 5�j	���w���Kı?g�����h�K�n�4m9ı,O��ߦӑ,K����iȖ%�b~�]��r%�bX���p�r%�bX����L��j]i֣Jk\&�v'np]�+��]p�x,q\V(oks{d�1(ᙩ��ks|������'��}�ND�,K���ӑ,K�������X�~��,K�zo�m8bf&bf.�ߚ��E�(X���Ȗ%�b~�]��r%�bX���p�r%�bX��ٿM�"X�%��;�f���/!y������-K��%�T�9ı,O��m9ı,O��ߦӑ,,K�w�ͧ"X�%���w��'�����/'~h~������K��iȖ%�b~�f�6��bX�'��}�ND�,K���ӑ,K�����ӑ,K���<{W5f���K��&jm9ı,O���6��bX�'��]�"X�%�����"X�%������r%�bX�t��@�R�%aI`@���%"V�(Д����`D�)�4`)�EšbFF��Z��I$�GS Ŷ�+ F� K�qH�C��
A`$�)ii$"�-[TP����P�B� �b�X��!A#`T��F @#� �� �ѡ�B
U�H�# �F%�	FH16�Q6`I	a��*80C����$�v��h�"��a#F!$!1�����B5BZ�V�$�3T��cRB! �D1 A"F)� �@"�D��!CJ��, E���)Eb��?���mŶA����
MuΚ�!)�Cͫ�j���;l�n�U+��9�\q��2�n��ωg��e� ��	[�qL�y¸r����zx�=�SU)��j��,�궴��Nv���T�Gm���!f%��hܑ�6�	�C���ݷ�7:p�w�r��!q�Fݍ��z;��Qv�n;)�YZ���z:�ۢ���]"��GU�q�l��)Iֶ1g��#�Q�R%aX��M6�Ǳ�!��ӻ��m�v�Z�ώ&���H�k�*�eia� H4IV����A@�0�N��wc�VWF�h���M��)�x�Q-��\eP�[t4��� j���H�k6��5U��,�[`ݨ��v�:���ф�]4���4��[��P�:qæ�$b��,�M��:���l�b��n3���L�:6�&��vd�H�K;vy¹~�����&�Mƌ�ss@�raݫu��]R��m�λmz��XN7�}�p��Gl<5U��!np�=��Dm�v��l�u�+���m�ܜ�㞙|�)�G)�.-<�D��i9�q��֦XF���{z5sl�xJ)c8��PNۊ�R�j�VV��ӷ�8��xN�bUZ��L��$��e��Tـڝ���t]��� ���'P
˷<��r6"����-��R�	����ݏK�R�R��"��$��W>�Ti��4�l�X����m��C���O4q\�5�R�og\�O*�b�[tMy.{s��T:�9��s��B���V^��77"��	dC6:U�������9v��Ĵr8mO�]� �{A8�b��te�k#m5lApD�j�SNN�l��nD�z�����ҳe��`r��=�ƅY^v4z�{aqKUhԪ=�5�|�iQ�J+狚��%��2@-Ob���S4��6�F�,\e�h��K�3�ܯ��{Ko[7o9`������H$dY�K۱ �n[�nKT���*ʭ��5j�;Y����3�$���s���9�1`(uU�E]�����G�� �U�%��ֳ5�h�fl���V��e�ջpu���.&�u��H��ŷ��4��cs�K�;;��Zx�^��n���XH�T���Ѽᶇ�g��Qn�'O[���.{7��H*rݞ��˷I��ԩ�XI$ &Nr�X�hK��¶^�;{H�۞^����I�q��m���ժ�In���	F��SMf�1%β����gC����;c�Gks%V�94j�w����||�=��Y+h/�5��շI����.���
d���,����/~��8g�|��epZ�w���!y�D��]�"X�%�����"X�%������r%�bX����m9ı,Ogze�L���4�����ND�,K���6��bX�'��o�iȖ%�b~��ٴ�Kı?}���9P������w���pVS`vg���B��b~�f�6��bX�'�｛ND���C"dO��]�"X�%��{�����L��O�>�?�U-n�)��ND�,K�w�ͧ"X�%���w�iȖ%�b}���iȖ%��'��o�iȖ%�b}��2�I�k!5&e�ֵ�ND�,K���ӑ,K��R=���6��X�%���7�6��bX�'�｛ND�,K���p�0��B��)k�q6fϫq��/���tn�y��=e/,b�>�]��G���{��%��{�M�"X�%������r%�bX����m9ı,O�k��ND/!y�޴;�GW]v3���r{xX�%������r"�A2&D�>��ٴ�Kı?}���9ı,O���6����TȖ'}���jdҥ�:�������L��\���n/�,K���ӑ,K�����iȖ%�b~�f�6��bX�'�k����caTnK7�&bf,X�^���Ȗ%�b}�w��Kı?w�~�ND�,K����ӑ,K��N�A�i�NJ��&bf&b�{�ND�,K�{7��Kı?w]��r%�bX���}v��bX�'�|voܪ��.����:]�f�#����U�|g�٪�Xk:$�oۈL��ӑ,K�����m9ı,O��}v��bX�'��]���2%�b}�p�r%�bX���ԗ�d�pђ]MMe��r%�bX����m9ı,O�k��ND�,K�{�ND�,K�{���Kı>�z�'��Vd��2�kZͧ"X�%���w�iȖ%�b}���ӑ,~�!`�DhH���w���Kı>�wپOo!y�^~�����GZa�i�=.��V�Z�`]#�=���;��;i`�nX2J�9���ؖ/d���7��`�2���D�h��M�0��6�M�֤ؖ���M�d�씝`��;v��D��R��T����Jh>w�@��� �镀{��`���m:���U���g:��1����Z��=��vhg8�`�J�t����+ �u��.��k�.愺c�	��%Z,�~���z���i'?gݻ�b r}�xnI9��I{0�t�2�j����}�镠y�Wנs�m��ojVZ�qEd,���b�
�hɻvvu��3!�w�B�9�봽1��d��-����=���=�2�wZ� ��5����m[�	���7�e`���<��,���:X�#l����r�����i�YIo9��:O���R1��Bn�Ҷ;0.����`�2�wZ� �}DCi���M6�`��`�2�9���;٠<1bB�x���X�B^�D�ٶ�i�/!��I�M���~����N�.K�L���Ŵ��c����f�˔���n��v\�i=������ۙӠ�GcK��«Än�8�u��d��)S�!��7	�N`����p<��V �\�v�g`�u�z�GcE; ���!��^L��l2�μEL䎽rt2@�5�9�V�L��{li\�r�ܷ~�������v9�qV�R��Ӣ�b����l�+���s�5v^�f�k�!�Re,e��+�i�NJ�w�j�=�j,ˤx��X�愡HV�`էu�{��X�H�k��X5r�AЮ�,��`]#�=���7�e`��EC%5J�hm7wo ��� �镀{��Z�O�߾�ܟI��S��X9mx�L��֢�<�� ��� �ꋾ�2�v�67-xz�ll%�u�{��]�����A����wc�9@�L`�3wX����$x��XoL�y:�B�8�NBS@����1%�eU~�lZ�,��V���n��!���e*�i'o ��� �镀{��^���{4��(��)]N�rW�wt��=�j,�H�k�]�	B���2�Ҷ�wZ� �<��u��;�@���Xڪ���U�+�z���vr���sf��q�:&^'v.b��b�]Z&YmZ�<�� ��� �镀{��X)5R��tҴ6�wo ��� �镀{��X���	�6��+�ڷh���v���=�Mvn~��+D
)���qx���4�9נ{���e�hv�Ӻ�=�\0)����`��Z���V5U	��Jh>�@��� �镀{��`�:�*We�$�똪s���+���dV0�Σlc-�c+Rc�v�Q�Or?m���ޙX��txGu%)2��)R�Cv�ޙX��dx����U�Yj���V�N.�����`�2���P�@���B���-s���� ߾��ɋF)� �H��  �1#b@�,b�
�g��|Z��j5�uF�$r[f���,{�V����<�G�}_�W�K�w�'<�r��h�7b,���ۙ�.���q�ŚSۢ��u̇nm�BV��I����'�X�ˤx��撑�Ʈ��;b��=8�`�"�7_E�ot��5C�X˲��t��c� �9��,{�V�֢�;_P�uv��WM6�`���7�e`�j,�~[/��$���ʷi
�c��ot��=:�X�ȴ}���8����,�:2M���aIet^���֩,7�VC/G6ՖE�r�]/.	�~��}�� �}�Q0����9u�a��w9]�����t���X�j�}-�>9zԝ�Rwc �qs;�.�c%�ǛKx�X�`��حs�Ц��ζ�"���:�歴�
q��4)n�����m��P�=I,n	�^�.ڮܭ����F[tb�Ր��s�k�����YM���9�s�NrG��Y�V���]f���	j�9襕W��W
���[0���J�!|��Z:%
I�Y*�}�=�N�����7�e`m.�EJƭ�[V�s�`���7�e`�j,T���ҺM�Ci�ݬu�X�L�ӭE�{�� �-��WM���Kk���,|�~�h���z�����bK�/~z{})!T�5,%Z�Z� �9��,{�Vu4&rs�̩a{\��i�i��թ`�aHƖi^fǱ�W��n�ۦm]gTp��¶׀�"�3�y`�u`gm�XN����"\@���u��IbM$���镀l�`]#�"7�)I�l� �1�X�L�Ӯ5�yt� ��� ;x*���t�v�����=�E�{_E�ot���]Dj�e��+,�m`�"�=���7�j�<�/c�9����-lr�n�P����٪�\�[]����\�l1��Bdx���ŵ2�Ce���v�`��`�X�\k �>� �-��+������=�2�N����,��,���v7t���lCwX�Lf�}�~�R+��bA�4zD�X�$X�j�����"�! �bA�"B�$�
���_�$�	B��[`EhJ@�D����r��G���	�~	ebV+"�	x!T2dHDĆ�p�c�D�0#��⿐�� �HB@�$R�*h�@#0 ⑌Zŉ��[��;��C�*�(A$D�l�.�	'M&i^O������B'��5��R�B��q>`H�\].�HB�Dp�BMb��녴�
!m\�� s��H�aq�D� ��J�[H���O�A�&B1�)ѧ�`�$���&����H�`P`ѡ#X�� �BI�O�x�J��>@?
��+R(������Ax �DS�T7~��n���ٹ'�ӫ��r"�%���Ic���=yϖ�镀M�2�	:夆�-Z�UГ��n�� �t��&�`�ν 醙�2IY
�C)hY\<����"g���Z��,���nN��3��p\;��.�M��=�2�	����X����T?5WV:n�Wn� ���{�E�n�� �t�ϿW���R���MZi���ӳ ��� �}�镀M�p�5H�������Vӻv���`�X�W	�R�����$B	�E�k���˹'��#�\�8�!%��s�ՠy�WՀ{�E�n�� ����T2��l�����՞ǳΟK4�H�8��6����E�ۈ�Bm��]�����<����,u�X��V���;��c�m�X��Y�Gs�,d�+ ��Qgɳ�~�jH�+�T7+�9�ߞ��t��=:�X��XGu%)2�����v�wL�ӭE�{�E�n�u�9�k�F��R(ݲ����Nu��9נy�wV��I,31`�K�$��9y�9'{���=r�;&�ݚBNql���L�Y��ԱgQ�n���Ɖf�k�k���[e��`.j�0�(��45��!k)�)#@X�M�]6ae�0
"��~�y���͖��n��gquc[d\�1���f��f�N9s����w�]Yݯgv�v3�c	�эq�4��)l��$V6���i�v�i����莦��v.�k��e��+ez3����ž����֨ҚҜuλ���������T���xˋ��n<��i�ؕZ.ؘ;,��@>��|���`���� �Y��	����W�n�� �t��=8�`��`e�α��&�!%��s�ՠy���ŋ���=����􏯲�֚�M&�N&V�}��,��+ 6)R�-���0�V˺�=Ϣ�7_E�{�e`�L���)M�Cl����r�1�B�GKl�,-�D*Z��#V`���2�&�C��ԑI[xT7+�=�s�@��zq2�s���JRe[�&�d��ܓ�}����+E���#Ԓś��2�^��Nu��;נ��DƭR(ݶ���}z����7\� �u� �H4"������e�k �9��X�\0�j, �D���h�����7\� ����E�{�� $�&�uԲ�.��-�i��q)�:{3�8{IM�i������[$eccw���W�{�^�ε�r,uȰᨣ��2�/����gZ� �9��X�MZ��}V8��ہS�:�9;נ{��^��`�bX%�I�^���}z�n!4�.�E@����X�\0�j,ˤxGu%)2�J�c��7��l�Q`]#�7\�-���}7Z#�L�5ֺ��Ԭ�6:�랱�˔l�����,�ݮn�6���y�"���6u��s�`�E�ou� �H4"���l�[V�s�`�E�ot��6qp�	H��V���wn���X��V����}5���"�*����k �tՠ{����':�f,�f,IO]�^��H��(�UC%�$�@�/M�N� �}�镀l|�N����W�3�x�n\N�vW\��p�3ںə��&�	��p���q����!)�y�νu�X��V��� ���&�E�H��I��7_E�{�e`�\0.����JRe���E���=�2�N.}U��Z����|����K��ҰM��wX�˺<u�z��uh}�H7����-T�������,��+ ���o�����i֫��f�:볦��UƮև��� :��\�Fܭϗ:@֭ٺ�5�u�p!�ӗ���պ�!Z��{-�i�`�x�.Ӻr�6n��Ov�vS<��e�Z8��5���(u� �76.z孃C���{ ���pj9�g'k�(��n�M=����f`8v�s%kr6��Ÿ���nJ�9v��N{b�݈�V���j��8�IH�ej[���,�9=�9'g$��$���/��zȺ^;ˮbȜ���܃�`�3p9�� Bol[������!�����N���>�`�X���,k��!RE�Uv1��X��X���,u�Xh�Q�J�Vd�e��w��y�ν?fb�T�s�,c�,�r�m4�Ҥ4]&�f�}��,��,Ӌ�'[%&�V[h��J�`���=Ϣ�=8�`��`m
�)]�M%����	���Ѷ��&nݱ������͉�]	��y�&�p������Nu�N.�Ⱦ� �s��$|�뻥Z.d�Y�]�9ߦ�7�h��iB�PhP�B ���%��H D��	P,Phү�We�`���7�E�H�	���lE�Yc� ����,y�X� �D�I۴&��wv���`Ϣ�=8�`�"�&��"%h�e�7wk �}��� �9��,vEI�-���֕�ۚ��Rl3٭��k�Q'Y�D��X�3[�!�X�vRֆ)h�k�<��@�x����`S���+��4��lv`�"�7_E�o>� ���I��I��]��.���u�X�������� �����&�7$���n��'v�ht[ݬy�X쫆�r,uȰ��R���諤؋wk ݕp�=�E�n����@���X�
��I
�UvK��ᒒvT�N��N]A��ƻE��cqWwn鎓Uv`�"�7\� �}�*�E�)5ui�v�۵�n�}UU�#c�,�꿌��,����V�����`��`����X�`�QGe�WC�N�Ӷ��X��>[�{�ߞ�ﳽz1f	f?99נx���B7J�u)f�}��X��X쫆�Y���8�`���>��Lf�UH�LѴQ�X&,+�im�Z8+�;hu�,���vJ�`�E�{�E�nʸ}����A�ϖ�_Seݶ��7k ���*�{_E�n� v�*���wE]&��ݘ쫆�}��X��M�����ն�"q�M�g:��"�=�p�7e\0\D�I۶�(:Kmz�����3�wϏ@��zjI�g���*����*����
�*��
�*�UQW��UE_�EU�U�TT��U`��DX*�DX
�T ,Q(Ab�a�+E��Q(E��E`*DX��E��A`��`�E��DX�E��DX"�b Eb�AbT"�E�� Q"�, �E����Q*�E�E�1B�`DXP�DDX0BE��b��E�AP�$*B(1DX��*(D$ 1B0PB�TU��TU��UQW����Ux�������*��*������������*��UQW�*�����
�2�Ȅ����@���9�>�e|     �� 

 ( �h�� 
   �   ��  �%*Q*�

REI*�JTJ��EAR
@�H 
Q@(�U�Q( Q   @P(   
��`��iAc)��bk���xv{�@|�,}���׻�]>�u��瓯K��sҹ=��5� ����O��Jp ;:S�ҝ޷<���dҘ =gA���r}P�`��p<         }� :��֞O����È1:� 7v�i�Y׭<}�5��t�  �湟^��ݼ �^�K�)��� �}�+{��Kŝ�w��Zw��_x S>�..�mɝ3����YE� z(��@   
U� i���qw#st�����5W��@���ؑ���wXu}�uA��9L����\5w�����-Pc� �ޭ\�]S����t^ۖ��� �-źUrk�+�����|�ꗀ< �  P P�P ���g0ʲ�϶�O][�q�{����[���9:�&u�Ž�� ݔ�oF�ɻ� ڼ�J��w�_> ��)c����˅��k���{�m�  ����5���m�n7+�  � �   $��A�_S��Z��g<S�X,���� �M4� �LM�6X((� 4� l((�`�  Af4F��c� `4۸ ��M4���( �J0 �h s�� ��:14��4  4��T�*��5 h�T��OU?=U)P  Ǫ�)5=@�1241تT�(� T��%6�JUM4�&C�
l�Jj�4C)�T�����?����*����dV�m�����f����
*�Y�T@QWAT��U�� (���@QV*���ޞ�����Ձ@�4��N�����BC7���5�ؤG�BH����T�5��' A���Đ��X�	�0�!+�͍RH[h㭄�!0��BF�I�$u����������B1�@�	7�R��K��@�ҔX4hdB!)�F5����4�v��8�%u�G�8~��F�����k$w��-2MI(kD��F�鹣D�!�A A�$O�O� }#�2h8��$�l����>�S�r�!]�z�7�+7�#�P1���T�8���x���0>H�� 0!��L!��c���:��w��q%0�2j�Mn��f�E!��!V[�&�%�B�Bf]L�R.��E��&�H��IaI��јB�G�D����Z!%/0!��N���'��r@���?@���A0uA�h�$H�Na���`30%�5
��%&j$,�P#���`�����ˣl�Zn��X[�s�����!T� B��0C�p������jh8FD�����XU���y!�����e$$$��#$ިJP1�D�a2�b@�DcB\	p �0P����!�R��"I?b�cBIm%l%@��U!RB���>�Fv)7#�2@�c.��1��l�d[����1^X��fL�&�[�
Q�4�X���`P�D�1�X�SD(B�1b�ЛLY&�$�H!L02u6��࿝���3F����.S����	�ɬ�"q��m%ɠ��]γY�:�������@���!J��f~�5��L�5���ٓ?i�B��#LaF$X�q�GN2#�P�0�%5���.�6��ޗI*B�����Ca�a��
igؒ$�(�E�_��RCC|��&�.�o���MM�D��~G��X�ک/��$�*������a4��Ѡb]k|� ���$�O��	%�2��ct6�"��C��GbB#D���ӳ�!LC��9�%0ѱ��H1��b�aL���S~]q�%aq��u���5O�TU�2��lϋ�Лe�p�CG[aYM~�p��cX�5���k
�a���L��In�L�9�����0.]2�B��M57!$��L�k�gw�B���I���pu�8�`@��K�h67�BXS�+��|�o�[�[�\�ư"B�j� �����A4�O����]ǉ�9�?}�#�XB��1��ZZb�K�h������M�o�/4b�"Ӱ�D�,R7��.W[���ƵÉL��$ �"�n��V[��of��"��
a����Ì	���x	��B�Jf�X]Ĥ	�+5���
n�yϡ΄V�/8߾�bT�O�M�.ki~$f�����j�\���@������!I�z�}{��q���e����B�	!� O���j��@ B+"����Ԫ~d���2g�?L���Q}�L�WT"�h�HⰦ� �>�0���Y1ͼg�~���\�2�"0��hٹϏ�%Lt�5�~����|%�h#,E�?`~�S��!8�����3.���+�E5-('bS.-]K�a��D�)�L6k⥙���r�O80��.�1��op&���f� W3Z�7d�CN$)g'��il�.�H%	p�o�&�� �!��ŁLѫ�Gf�!&h�i!���
cI
B�"\&�����!"IMJo��r!!XR\3|�\��)3{�	��
��
1Zb@�0��+�0��[#�IBE��0���8CS!SL�d��V,&a�0ַB\Ѷ�"CU�aM��M�Y6�z�F�j�ё�5�&;H3F�\���L��p�H��$S�����&�O�;�)b�wӰ1�X�0�:�ĉ$��Y����8�����l������!ܡ�՟��yI�PL�%3���#3�����D HP�ֿBK���s��5��։MFӼ	���6�H2��_�ƞ�(���)��1��t�D~�ōq!L�XE��i)Hw>��?Bԅ\��ILbL��Y��6J�"3��Y3/3�	BC7�������V�ᵔ��x�h����4D�3f���K�0��e!R\a��0!LI5%�4�&D��q��_c/=��ݚ�۷v��862���HƤ�(F��������ee�%�%1���u�ˑ!��+��pѭ75��~����&}>���K����jw��\�K�S\����d�.kp�sF,'S3!���IVH��!&�&���!��\J��jա+��#ߒ���L���^ѳP��~>_��f���f� ��,I���M}M�8���q��M��rk���dMR[Y��S>G� ��_�_���Z���߾^�p(߀�3E]�	O�2j\�k�������J�:�#�A� ~#X0 �ؐ
����� HָiU��R5*c1���"Ƅ:q�a���#����wIo���3Y��pCC�o{!sDvj�?j�4#��|����&��?}�O�S2�o��t�c�6~>@��B����"mނ\M&���?a�#s[�&������of�sF�����ю�W������l��^R1�e�Z�#%���9��s� ����H\XB��C���]h�FZ�#��A2�7���b�\?HNO�q'B���O�?s�n핱#[���f��������9�L?:��[�W	��,qȑ&$��2d���F�4Ln*��Y�Q��˴$QHE�YA��Hm#,�,3"Ip%�f�7T�&����u�ǉ ��衫�{7sdh���c@1!I��+���"R0�hڐ#���XC�A+�	V���I	�i�8�4�	��@"%� T I�� �x_�Y���j$JOى)_�0�F�bB,5M	
�MϾ��.kg���7��`�r\�[/5������\t˚��(�R���?�hC����0���+U�!��.����H�頗��Xl#B��\�Ë�����&
4g?`r��i��?������s��L�f���q�\t��@�:C�w�/�8?��D�p��~���_�l���1�lv���SAB��H]k|������N'�?k#$�!Mk7�'3����s��SD)��B4fjg�^s��2]���!��< CW|�D)ѳ\�CA5���XЋ脅ģ�b�~�7��B�X�XZ`B��K4�©�5,5�2~�n�q-P4&!�����}�z���C��2u�Z����{�?�Ĕ`��\�:����	L28����V�N��Ĕ�1�:$4n�&&�ĄX�� ��$�3��)Z�_�seѳ�㤐 �cP�cB1K��䶑)I5���1�kt�FĬ��!�#%���R�g+�y?/� AH�T�Y����{�D����|��D�K�_�+R~��ܶT5�-�D����� �#Zf���p��~Kc�he3K+�iH"�O�Έ�5�RB P RS��ߍ�Aro(Hh
��� ��B�!����h@�+ 2d�ތ���D�ó�%$������JI�Ȥ �#�&�I
��͒��?^�.B���M_��f��l8�Z`F�Mi��p�P1t�)�B�? ~FD�(d���rMH����㤐�0v� hH�&B�j�@�$*$�2�1"AH0!"J@��p�����F¤hS5�P� E�IL���!q ��^nbF��qI 1'�p$���a�l
D���̬0m��df��)�#F��cB1�a��f��i�!)�.i�aM��M��3F��	�P�D�l��L4�c�p!p�ѷy��4�$����A,��he$�%t�	��e����:�����ыV*BK�|O����	��O�h0 T��D�c
c�4������C��ܘcm3�� @�SN��!\�s�o���fC$l�#n�p���H"G���	�`Kr���R�ۜ���'I��_���� m��m��   [E���'�kksm%��I)m��zFb^n�GN�6q�hܷ  	mv�A�鬟}���Ol�tjn�
Z��� RRKn���f[@m&Ğ���m�� 6��mm�P	l	-��    -���h�i H �il�� 9 E�K�|�_�� [[l  -� $    �n�[d��-���C��@Zt���8z�-�m�`x� $ �f�@嵶� -�     ��@8 m� ��m� $ $m��mm���nr@m���	0�����m����N p�ޣ�E�"Cm�lxjU�Z�N4����檨 �6�`Hm� �@	  ��;um  ��.�-���m��+K��[��B9B|��U�Pr�dV�)�"�rh�M�%m�礶C}�_���m��ƀ��&ͭ���@o;<:�Xr��\ m�j[��]Í�d��շv �P8#m���m�C����d2�PUU��U+��m�$�/Z ݮ���׵�]{F�  &�i@�I]cH�i���[YI/]��쪽-H(G5UE�rd�4�[�m���^�N�m�[P9� (��{d2�U6��®̫tv��5 OC���\�n��Nn�F�
���y��U�UV2p�K	[\:
�kX�@U�=��N�)Y�m����`)��!���.�td���l�$q��V��Ćyw���S乬���C�Xc�����v��O�#nbR��/f���`	�� �	�@�R��H-�m�Cvͱ��Ϋ���:�'L��&��A��&� 6� m��(	�ͯMr����h��6�1$���-���۶���i�IoS��ܒM  �t� "D��d+u�m�O���ɸ�M�I����ڶ�Y@  Z-�\�����t�4��Cf�  [I8��m �m���`gZ�� v�t����L	tZ;GV�-���R�P� w����� ⪕ݚ�o���]�:� �W��rIm6�@@�79-p�$F�լ$� �k���h$:�e�9�f5� :]$ݍ�9Y7^94��pH���K=Ri�̷ON���m�c�4�\Li��i��y�������c��.Y-ʶ���&�WR򀪮�mKUԫQ����U�AVC��lH�'I ���L��kJ�峬6 �����n�H�3-W�Ն[�]��D����s,�*뺪 ճ;��r�5*֧�U*�ŕ�^���2����A�՗���.�Ӧ���t��R�7���K�M�g����
�ڋ�%�Pj���$m���F��#'.�����m� ����WOm���b��n�R^N��}8m��  OL��k"Aʹ�4��[�[)AUc�������e蛜�mO*U�.�-[R$k;um�lm�D�$�SsK�t�8:��i1�!s'��sC��9-0�\:�Y�
Z�T��F8�sT9wktk ��l��d9٬g2��`M�j�������>`�m[���7l,��Um^�Åӑ%����T lje�iUZ��[vH�S8<2F�IgVw2_|�'�W[�@����
����V�`knW�Ü	 �l.=���2m�m[.Z��8�j�꫶UCL�[=�Ut�g  [M�7K�2��J�R�W[JK�q:���G��kda!�n�#^�;n��m�I6 �Y�[�[�� ��v��Z�[��W��`�t�TR��H�y  �(7'�����[n�J��
N�gM�lnԫ6;���v��t��m�dmTUK��U�AYm�U�e�ʵR��.���Fs+��*�khq�l	M72I6��~��L=�qUW�n����P���Hl�$� -�h*�$:Z�뀕��j�k�˶M���6K�����-5T�ۦ3� ꪺ�
@3*>���� m�rV6�[�Ē%�k, ���&��I�Է��ν*�֬g#�6ܵcM�qfkh�4n��� :@7l�^� F5,UUPlJ�H�2�a.�j��nl���J��RT�c���- /#���j�j�6%����*��`4�5� M��5��Z/i�I�l��8m�m/[��N�VJ��p-B�*�Z���u�;\��P UJ��T�J�Vį���!��� ��p�А�m�t�4�$6�@p�j�N���Ā  �8-.���m�h�-��l 5�� ��S5UxV�v�m�ڲ�T�cYVv�-i- *��-���`�X�\m�m�bM��6�  �������^`�m�궸
��_��r��m� H mms����M��m[a���$��m�pX�-T�-��l �����X[dŶ��a��[j��siU� �vj��pn��m*���q$����f �v� ��`��  !�4Ͱ���-�m���tؐ�Ӓ[M��I$�Z��� ۶@�a� d�qm@m��i T�<�f�b�U���vo6��l�kV��E�i+m���3��(Im �z�M�[%   z�m8�v"D�]��� 8  p�l,1��H ���@ֳe�H$�i7 �����;m����@h � 6ٶÀX����� �pr�ֵ�]z\ �>���Z�U���i[��������o��:@$[]�k�l����m&�-��A�8t���<�+�!X
�g�����J�l  	 m���(� [d�Z� �m�m $ ,\���:�J � 6�n��(>�[��@  8m'n�UUBh .@6��5R�V�m���f� ]VMm��H8��ED�r@ H�$� $�ȇuۤ�m��ԁ�vmnN�H  N��Ui�U]�`-Ssn�[L93m+U�n��a�YVu�������1�OKd�%�XbНU�m�l�-�7$����q�W!5�IZy�*� ��ej��,���A�U�@��G*�&q�%
R��
G��e��Ħ����P��jk�C�%ƃa�;mp�9�]�-�N��vԫ�v�ب�m�t��(�9�T��Y��Ս�*���;p2�N0�M��U��&\�V��[�m�	   u��mH  9t�I$,�    �u���`�Y@6�	5��!��7�Ի�m�  �n�A���@ k5�nm�ͱ�Ŵp g�m� ��p�;����NӖ�@jL$$-�$�m���s���\� �M&\U+�<�vE]��	�Tc��V�������-�d> [dm�!v˦���2Hm4��U�@\��[[l ��k H�E��ÆG�6��	&]p��`�۫(m[
�U�j�j�:� ��m��4�f�ͧL[@'	��H� �Xc��& �I�I����m$���2r�^� �ioZ�l�:&�pl�� �`6���@�;Vm٪������ݶ���]�[@��WT��B�
R^�^ �z�;m��iڱvm&�m�m�6�ˀ-۔�r@�Ym`F[T�[ڀ�x�Tx��,��2F�m�Z	|�]�1�FWE��y[U)�-J�UP�n�m���u`>p�: ��bV���:M��ջ��Kf���mI	K\����[u���z    mm�X\� U�8���ջ6�m;Em�Nے]����\��@ /�[l�| H p-��E� �.���:91uTjj�s#�ٳ�l%�9%��i6�n�L� ��8�e� �t3�����O<B�`�!� ��6�:�K�T�9�<KS�⧲茓�]Ӷ����p8�\�L�3v�m�x��f�T�b��UWT���z�S���-�k��|�[݁ٯ  ��5�ֵ�i6�t��6�8�
W�I�*���UUG5�m�umU �mx  m���c��߾��v�e(5��h �	e��b��	 @	 :��}km��� =6�6ݖ� $6�6�fݵ��� m�HsV��q �� �� �`   �-�[,� �� �'n� ��Im 	 �� �  m�� �Բ��^P%@j��Z����� �ZN٭��i��� 6C Z���`8 ��Y�I6�l�p �X��M�      m� �m���m�H [@P�g [[l�6X�l��` lۖ�����UC���UK�)X��k��rکw3��NZLM��RZgc���c!�B����wH�.�Gj��]P�̠)oXi�i�I� sm&m6��` �  U0� ��ѭA� ��	 � U6��)����ۧ/����h�F����Q��'� �`���.�J
�@]���� �D Qb�S���@*:B�(�P�#�N��B uS���B�����ߕNO�a�M�N(TڨT��"' �^�!�b�VD0> 6 ��D���EH�V@`�AF��B"D�~�~\RiT 
����8���F(i�jc"�$b!�� @��""� ��#"$b��F#"��a.��� ���: �U1�|� i��T4i@�k �D(��� ފ����C� �`�`@N�<�§�����X��_���A���(uS���W�� 6( 1L �/�����	Gbi��UЁ�����#0"�l���l��;@sY���V���m�a�0�KHR��F�Ή���si��X�Y�aRZ��y甛[Cv�!ɯVmRbN.�j�%<�Vxx���[��# v�M���"i�5obꮌ�i.�����n^�9�@�[���cyn�۲�����ѥ��$<���9:�&�&�4*��X�U�mM��9����ۣK��6�H6Kc�6*�ls��pr�&��]��l�e�t��lt�Eԛ������GI�˴I�c3u���<AC1�\Ix#P����]��m�,�e�UD�H*�%��;9�'A���q-qlV޶�i��yA���e3"u.k��N��	.���;p����M�涶�l��Ԇ���s����"N�z캇m�g�6����#l1p���W,��@oz7J��j�m%��C�v.6le!��7v����ش���;�[�]!d뛞�\������N�3����=g�F��ڞҮ��y0m�!j9M�Zk��*��e4�O��Q`���ƅI!�ەm�f�-��uaBv�C��8$�v]a�ڞ簰IǞ�`7X��^�͕y]�7T�)��\��c[�Z��XN��^�(�ɹZ�
�,,8�Y
�Im+��e�C���r��3]vx';�{o;N��S�WnY]u�tdsts����q��v}p�IKX�`*�ke%���Ǌ�m�)��@L�������ڭ���y��eC����E�c�z���gD���G�[9�A�:-�tc g;��$����79jpq��Z�Qv��^�t��&��Tn�.[��a����u��Ϟu�h퍳eb�mn�b̪��m�[hz��1ȖM�c�̧Z2ks�b2�֪�ٛ�i��7j���)T#c�XH��ɳ�6��NP*5*��ڔ�L铔3���@nZ��8��-��OY4c�Uyn$��e��<f6Z���$ԦJc�j�W����(�( @A� ��*���� o0�>�֋u3Y��Y�q�t��+��%��]{.������V�Y����؎��1U�=Q6�㤒��m�'V�K�x#���m�[s�p<F�!�:�ɩ�ƙ�E�!��+�+��!��&<�Vľ��m�]� �&��5��4<f��n261�*{6-p�[Q�����l0�Ac���4�c�l�"q�:�\�f�m���.3Z&f�T�Ё��n�<���ヸ7&����w<���y3�vrc��q˄�[��Zk�2dI`�}��&� �&���&��	��ϲ��PT���,K�ﹴ�Kı>f�\�R�d���h���%�bs��nӐ�ș��w=�7ı,N���ӑ,K���ݕ7ı,N}����H���������oq�����;ݸ�%�b}���iȖ%�b~��ʛ�bX�';��v��bX�%����L35�.����dMı,K��w�ND�,K�ovT�Kı9�}۴�Kı>ϻ����%�b^v}�j�FKsV٬ֶ��bX�'��쩸�%�bs���iȖ%�b}�gr��X�%���ͧ"X�%����&�ɕ�2Oe.�8�m8�.��G[c���v�c�����ݱ�sl/W&�]��=�o%�bs���iȖ%�b}�gr��X�%���ͧ"X�%����*n!��������z�T������X�%��}�ʛ�*+�)"��!�A���Mı3����Kı>��eMı,K�׵�/�&Re&R��Yw	$������f���X�%����iȖ%�b~��ʛ�bX�';��v��bX�'���t���L��^���ݦ��r��k4m9ı,Oݽ�Sq,K��u�nӑ,K��>��Mı,K��w�ӑ,K��޹�h��u-�K��֊��bX�';��v��bX�'��w*n%�bX�~��6��bX�'����aI��I���oV�(�[q1�]��d+rizxs���t�z�sȗ�f\�C0��D�HъE�c�w�{��7�����w*n%�bX�~��6��bX�'��쩸�%�bs���iȖ%�bw?��*0؝�I��{��7������iȖ%�b~��ʛ�bX�';��v��bX�'��w*n%�bX��������%Ȳ��)2�)}�ݕ7ı,Nw_v�9� �@H�"!�DdF�L5"w;�ʛ�bX�'������)2�)=�V��$�G�ִT�Kı9�}۴�Kı>ϻ����%�b}����r%�bX�k�N��I��K�{K�.�%�ێ+����r%�bX�g�ܩ��%�b}����r%�bX��{���X�%����ݧ"X�%��n��)�j�f��(j��nig�k�Vw]
�� �%U���ٍ B���r]-MY��;����d�>��xm9ı,Oݽ�Sq,K��u�nӑ,K��>�&�X�Re/i�z]�PC�`�%Ŕ��I�b~��ʛ�bX�';��v��bX��נw��h�����&8%�rJ�}s��u����Py� ���i�r!H�x��@��^��빡?w��ܚ�#1 ��tT"iR�IA��x?����rF;��)~�@;y� w�P�sp���o8>��j4��!��[qV;X�J�M���%G&�-7s!-I���KU�# K�`����k�5���U���nh�������(�#���}V�W����s@��M��cy�F�QLN7�W����s@��M����\[$jD&�Ȧ28�{� ����� ��L���C�`ӎ��7�M0�IR��s�?o^�{q`*�,�H@�@*����"!p�*��DH�L1_~~a� �TZ6�n�kA��l�n�%x�Kg;r:En:mgi��;s%mQ��gk"%�wKp˲��=��Ȟ:�N�+��f6�u&�9�v5�9�wn# ]�E�9C��͝n�z��}
���h���ڄN�ֵ���vd+p�2!�������e<��*rt"�f�D
- �l�r�a�cv7q���j�q�nrm̋����R��6�=����.�<3�9:q�l��r�jܙ�Mk4�&�ۻ6���ģ[�f&���CN	F(�p�/����*�W�wu��/�S@����ND)�N\x�����$ٻ�� �l� ��j�:��ǋ#�bpQ��@�빠^빠}]�@�ֽ ��dCjH��B�f�{���v��Z�{:�3�$E$�4��h�ݼ����7��X%�쮻.�hi���5�"M�=<ζ�^ݶ��q�b��Nzs�%�4M/KD�E�,6߷߿d��P�� ����j�{�r1��D��r�{ۋ���T�M*��R��T������߱`}{� �����To@�ą��^빠}Z��\�ws*��2�y���\�$XUT����~޼����7�n�}cU��n4)oqh{��9*�������X�׀{}���&�:�ծ�$����!î��lJ�,v�
%����nBc�:uvlN�g���� w�P�-��r }N}�2�wc�,~��Ϊ�J�l�����_�@�빠��#1�"CQ5��s����;}�ܢ�U� �s�7U���_u��;�.őIi�#/=��7����Py� ���׮-qG"��zw]�����v��uz�Ԓ�dr'{f�K�v��~�}>{�$��<HY��0�@��9�6��D��$&�π�����Ÿ{�@;�� ��ϙ~�=g�Q��}]�@��^���s@��M�R������	.���9q�����e@�$�prԬ��ap.X��x�����`��X��܀@q+ �5/��l�u�
Lj	Ȓ�$���4��h{��;��hz�du��c��N款�G1��Mv��y��vw�nչ8�nk�a��Bc� j"9&hWj�*�W�wu��/��hݗb�q�1�"�r\x�����UU6n�b�;�ش��h�qk�9�I��dq��ʀ:��\[�7��{�M��9�HQ9�����b�@���������5�a0���L�>��n �s��e@YP�=��Wb�u���aݶs<l��dQܽ	=���c��:#t����o�[y%Ҕ7=:C���my旉���^cj��lnm���j3�@�q�c��m�<�.z�O�x$hȔ�ܚ����9�S7l����:ԣ�J�p<1������4|}����ܘ���a����8�H�rOnKvSk�����۱�Tݹ�Lm�l�cHV�[�MjK����J �L�R�W\uX��W�lmW��:�uA�-��t<[GF컋�VIK6���H���6߭�� ��TՕ �ϭ��-J�Y�8(̉Ǡwu��/���>�Z]����"�(��%�I���� ��^�*������ذ�u��m�L��ɚ�b�@��zw]����˱BE#���G����:���w{��m�<�U��+i���c� A�y�7�L�L��x�.m��R�kؠ;�9'�����c�28���hu���Z�z,�iO���Nf�y�n���H��V,R<CP}b�@�u�@�빠}o����a1G�@��Uhzנwu��/>�@���<�GH6��-�[��e@�n��[prԬ��Uډ��r^�{q`�����oG� ����J�'�k�˫,��M�G�5�tI-@��v�5�$�t�#��h��ל���䈎7��4�)&|���}�*�
�k�;��h�u��nBLMDK���=y�6s�u��ذ���weء	"��d�-�Z����7?H�F)I!T��Ci��9��@2��pg�d�q��tA�`�J�kHM.S#��4H�1#4JJ�b� B�BF0v�G7VH�!!$��IR��� -U��%�4��D��P8*	�8
C������� �����؃� � � � ����؃� � � � �����]a�M]kFf���f�A�����lA�lll}���b �`�`�`�����؃� � � � �>��b �`�`�`��wt��.�fi�˚�ѱ�A�A���w����k�v�{ۋ ��T���C���Ѹ���䠆��I���I2��M�E�]R,�����Ơy0�����w���p�r�̨��:߭.��ń����@�ֽ�g��$[nh�8�?{cל���+MEv�jKn�~�@�* �y y�� oW ��"#��l�%�I���>�/n䝿��ܘp>�9�)�5�U��mB����䓿����3Z����ㆁ�X��;+�y� �5�6�6�͌���������
4]1"Z�^4t���̍I�2E��ֽ���{�4��V��������$L�=��P�� �ϭ�z� ^��f
,r�N)3@�}V��X��*�W�wu��>��Sx6Ʉ�R-�}m��r�̨���o֗D�$�M
(�
����w4��>�Z��̽S'��������;-=LMn�=rN,-<�癎svG�����	l�ڔ�=Pzۜ�:�=�ݻQ�u���o7/m�C;�f��A�WCvܝ2l�m��x�vۆqг��|�D˾n�/F8۝p3����=ѳ���2axnewN�Jt��=]*��K
��Hn�wm��jם���s��`�-�v4g)eP��]K���q	���w�.�6�eftg�9�=���py����ջ`��6YZ���5�ۨ���2)�[nh�)�}�*�
�����"$��P)&h����[p���ws* ;\���rbj"H�}�*�
����w4��;�.�H�Q���@oy�w2�����[py��H�2)&I#�@�빠_t���X��*�W�}GqcC�2b�l�\���]A�^ۨYnՎNnθ/�[*�[�����Ȍj6Hc�8�π��~4��V���m�RU_�n�b�;�S�%�n�D���b�W�ffbE^���Jh�EE��$�M
(�
����{qaʒo��������{Lx�90YFE#�;��h�)�}�*�
���ו�E�LQ��Oz�w���[p�r�̨w��;��B�=�`�v�@���[���l�Dӯ/^�\땸����F�ך��#O���>������P�� ��!#�(��dj-�Z���>�Z�\Z�FɎ[�\�����7ޚa��U$�ʕ$�T�RI/���=x�۷�n�5���F�Rf�{�4��Z^��������&r8hv�^�UI.�w_�=�ذ����F(\&D��"2܀' d�����px��E����ܦj\NJe�r1c�F�6�%ߏ\�\�os* �y y��իLx�L5�H�w]��Jhu�Z^��ו�dY&H�X���^�M�aV�W�zw]� �ΰ��8��Dq�@��U�U�^���sC��)�wv]��ƱH�)"�/��@�빠^�M�U�}�����nb�������۬j��[�3�;Q���sM`Q��X丘���ɍLq8���>�Z��z,���Dc#n)3@��H�}m��n�̨��%{��S���b�@�}V���s@��M�QaJ`��Qh�7 ��T��@>��n�Z��F)0�F�E�wu��/�U�}�*���h?�/%�1=�J6d��W`뤫�u]t�R�#������5��u�dDN����[qb�SjV��m����ks��ۭ�'k\gmd��nn̖�c�r!�B�B̩��p\�f�v�ɺ;X)�ۋ��ks�v���y=��8���:�Sӄ�m��uE���vG�z�kvs�=I]HΎz؅��37>zGŷq����+l�flx�]d���6�m��7�w������ |d����ˮHn%���Ku���`D��+M��!�������$2L���I3�}��Z�b�@�}V���s@���'�G0j"5=p��ۀ7����Ps��wv]�E�8�&&F��*�W�wu��/�U�}�*�^���<�	ōLd���w4��hu���uz�\C���"6�4��>�Z^��ꋊ�jHG��f�tu��;;��6�3�6ᇊ����#8q�d�kqM���Ol�\\M6�m���G��گuzw]���4��E�q
`����]]]�;}��Ȝ!���_>T�te@7�� �ϭ���_��R`����G�wu��/�SO��^����˯�^VDL��2F��$���@>��n ��?|���}�~j�d�rH�DG$��U�U�@�빠_u��U�����&.��\Dt��{�&kx�v�����]m��k�^sט�)�I$��q�L�E�U�@�빠_u��>�Z�\Z�G��B�r�{ۋ:������� �z>x^��x��Hbd�"6�4�����6�UN�Rm������/_��4cL&(�4��V�W�����}�s@��TY�S�B�-�Z��b�@����iDc�2a�D�#f1F��;5���\��7k�sI:�UVs����U���(�k"q��w4�w4��V�W�� ��(��$i,RL�/��hu���Z�ծ���#s�#�f��X��*�W�wu��/��h��Z��I�'&$�Z_{o ������*ʡy*B���E�Dc+�"& PHD`� �0 �Q����/�Z���G�8�pdq��ʀ<��y�� o� mn�ƳMgb�]2.�������}s١c��V�뜇s�V�N���p�r9���A�b����݋ ��^�۷���K���X�����8��	�6���U�Uֽ���z���Qdn8�#�M
(�
�נwu��/u��>�Z[*Q&�G1(��@�빠^빠}�*�
���ו�LNb"���I3@��s@��Uhzנwuٹ&�tN}$"K�4�Y��R�G�
Ե�!%F�b$R]�d�a�ٙI�J%���΄�� 0� $	"�$Hq�6$`�bA� ğ�0F ��l� @����"@�Z�$)oc�b�`@HX��m�l#�$��apj�0
�(H�5�\/ "2�ChF�(Z%HV��� �s`���
�JƤhR�XL��-��dA�BXѕ�FRR+R�#��n�,bE�c�P��l���H 6Gd�P�)8	@���4[ �0�+%*U"�h���iJ~@B��p8f�V�����6	U�h����J0�+
�� ?;H͏eDJI��,�]����N������
Č̠��ݺ޵3.kY�WC%7.�P(U^��������ȭ@r��Z�̐T��N�&�9Cc����t��<�F�6k�m��w@Z1`�W�a��BD�t��<�����9rhQ�[s�m�M�btWF�[�.Ɍ6�md�6ͪ��\z�9�g���;�V�d9���w����ѫxx�Q� �����dK�ԇ=�p 0�+7n[[���������[,s#Tv �Np�TOkufda���Aخ�v�8�=5�6�C�3t�qV�`<9��cv�����M�l̳��OG��<Y���o��x���Y=:�m��5	ӪkX:��TrivT60F)�rr2�ƻ2�mjݠ����h ţ>���gjWd�8��uo=gh!�;v��uD����Nq�Rva!Gmʜ�t��BۓڇY��q����T��p�8��v��Ld�N��]����;v1�xh���;u�ԫn��ݬ9�ۚ��a%ya.�Ef ^l�X�t���UR�<��/��M�Ҷ���]��Ès�&�[;e%p����'l�r�ʶV�*��5]q��� ��+e�g��m��ѯ�>�������v˷N'���Z�꺸\�y ����\z��!w>%g���D��,�Z��#�?��m���kΓl$��d^���@���m��Վk�v�q�j��N���'{f��ؽi�1���S�0낮�VTZ�]Vh;RvČ��8�ͫw]�эX���6�5�n���u�\AA�z3��[�ъ��kc�J�)�Ld�e9z�ǝ�ۃMW�t �O�l�_o�xۂ�{u�8.	N���G�,5=���pn� �C��X8�����G�	3�7!ѽ��n@oy�4 AJ-��s��B�ٛ����M�\dr�\4��M�n�h��@���2�L�52���t����I���P�[2���UuF猢�d5��8��cWN�ήqX���ݲ���W��n�-vd�{������"jh ����A� )�\��'��mf!9d�F���&���.��=Rg��e��l�nm��O]���a�M����۲<MGChV��7a��y9.�,8�{lۆuzzB��ô���'ز�t��D��B���8����Kڶ��3�Z8ūr�ͭ<cK�{j�[�v�� ;��]�7E��5�u��}X�bt�z{a�ڷ3\F.ݵD��Qxh\vx0��w�ܦ=5+{Bt,�%nu�^��zi�7/\,��=�E{�[�f���:鉥���:j��~�G�z�\�\�ws* �2��3/#�8�8�&H��*��ٙ���m���~����X��=z�Y�8�Y$�����7��Xu7��|�~��@��Tc�dN0�����]��>������P_���ʼ�	���f��X��*��@�빠^��K�©���"	!��I'�ň8�ȼ���aS��v��k�㮋g']�mIc���8�Т��$���}�IwK�ԒW���|�^��Ԓ^�jQ&�G1(�L��-���ٽ�tf�o~�xs���v<Om��u��ʪ�ݱ�����1G#Ib�#RI~�����%�n-I%}-_|�]��5$��.���#s�#�g�$��Ÿ�$���}�IwK�ԗ��o����|�K����RF� �ę"��$���}�IwK�ԒW���|�^��Ԑ���~(���t�Ź�����%Sv˰C�F1�]k����,ZrI��i�$�I�$�t��I%{����%�n-I%_�|�V�#L��	G�ԒW���|�^��ԒU����%�.��
����>��2�.Y�kG9m~ޏ��{n�����T�&���rf3I^��}�I{�ֲ28�B�QLZ�J�Z��$���jI+�g�$�����I%�v�<jdq
9���|�^}Iw���K�Ÿ�$�~���$�38ߋ>s���ܾ���ɷ�6���5v`˸��m�]{6�".�<Y��3P���*7�����}�I{�[�RIW��K�]F����Փ$�!��$���%�n-I%_���I.�u�J�����$�e���$k��$S����_�$�t��I%}o���%�n-I%��|�oLn<$|�]��5$���g�$��Ų���r@�DH$˟}��-���YQ6㑠q��5$���g�$��Ÿ�$�}���IwK�ԒWӂ��8<^�A�Kk�s��={q�b,��
�荧�v�H�?��o���Ξ����������ԒU�W��%�.�RI_[�}�I{�Z,��(��IBbԒU�W����Uwovv3m���/ߛo��bx�o�nk���G������%�.�RIz��>�$�l7����_�$���D�9��%�H�I%{����%�a��$�~���IwK�Ԓ_X���I$�j"9&}�I{�[�RIW�_�$�t��I%{���-�O�&�q�K�#sY�L�[����p��9,c\u�T톪���x���m�Z��v�ش�\]n��m*�pse��Z0n�k���b���r�uK�o)n�s�-�B��k72�ϬӥUѫ+��`ڙ��uf��f+kh��^��u`�<:��n�6�.�mp�x&� ��6%�[����clgs�[ƶ�m��¼��N�6ܝ������w�����>�����S�ng���o���u���c�96�'kdR�XZ��"	q�LI�)��$�;���I.�u�K�����IW�[o���x�oۼ��.�\E�f���k9�m��wvo¨fe�{���T�_�n-I%�ֿ�I+\YY1G�I�#RIz��>�$��-ũ$�����%�.�RI__��2<m8�&)$�7��]Z�I%�ֿ�I.�w�����}�Iw]z,��1514(�5$�?Z��$���Z�K�߳�K�uj5$�����NNl�桷Fz��#�S��z���rK�z��U�)Zku�����7)7�$�s��RIz��}�I{��F���ֿ�I$��D�c����X���$������RUwo�n<f6��n��ͷ�^�~����C�����3���������Z�I%�ֿ�I.�w�����}�I��M&�#1H���F����_�&߽{��m����~���UW����1�߷#�x�IŒ4�����wqjI/^�g�$����jI.~���I,����tt���;���V�KGex��]C7g��[�O"�#Y�|��sE��5�u���߯��K���jI.~���I{��Z�J��_����&��g�$��ը��*��oo����m�o�<m���/ߛo}��Y"ÎjbhQDjI.~���I{��.�TB�o������wwf���v��#�J9���|�^�w�����_�6�۸���J�W{=��6�|oH�,s�9ILZ�Kׯ���%�uj5$�?Z��$���Z�K��ϱ��ƈ�{)]1v�ɮ��n��r��&q�E��벗��ã����Td�Uw���>>�׫��[�k̨}K���&Lb�	���/Z��ڴ^����s@�uF�����dq��� �YP�P�\�+�<ۖ��#�%ǁ�T����`�� ���x�T��U��J��{�k�?}�����i#�9��չ�yzנ{��x��ŀu*��5��M�HG`���'\C����淶��xͬ��nyRv�
=���T���KYLE�ͷ����~��v�׮��nh�W��MI#�ڍǠw��@�빠{�[�yڴ*u�?����I���s �ۯ���_s�7����o�`Y$�!��$��z�nh�j�;�ՠz���*촍&&1H��d����� יPT� �ʪ�����{�����y���$��8��>('�N�]Aj̣��4�8�3����[�����Ŷ+��n�f3��ç�|\�d����X��Hs�nyۗG.ް+���R���nW�k�~m�D4얻�;)�oZ4�n����D��9����N��J����6V�C¬n���"���&�c�[��9-�$�z��f�ą��R��@�I�X�uF��ݍ�cGt��0Q�ͻn��&sѱ���O.�Зn���D�%c�4��lGV��g��?��2��*ۋp�<�$����I��[��z�*��p�[�:�J�ޫ3=�fW����@5RTw��� �\X��x5#nAGr���Oޝ� �_s�>�w$����X�N�-LN@m����zyڴz���kŀ|�ݼ���UW���0�5{X�.-�nݡ���R�5�<���Y��-��I�H������X���;�~��=֭��ֽ��Z�9ܟ�H�CQK�֍�?}�ݛ�R��E,�t�@�;V��[��U�lLL&Fb���<g�����[�k̨�]������L����;��@�YP�e@6�r�{*�]߮��	�-޷s@�R�h^���ՠTub�dx�cS!�d�eݝ��m�I	�q�<U� �p�kek�n�z�c"	����j��=�j�;���RT���v,w��0��r7r�l�_���p�[�n���ܨ[+�c�"jcj7��v�޽ٹQ]`BD �vTڕĊFD1�A����$�[Fp.`�SC�0`������ ! ����#(G�� ��IF�A�q$
.�2��ĕ�u*&0R	h_�*��`F�Q# ���R�A�#�*5P�"�H� � �T?��U(�8�E�U>@�E�P �#��p |�nhVנyS��xHdr4�/{� �YP�P�\�v�� ���O�$r!��䙠{�[���zyڴz�����;�4��H2d�\�C�g�e�טἝ����۳�:뗨.�n�$#D��RbL�L�<�k�;�׀}��.��=����̑���q�W�3��v��ue@7��@6�^��ǊģN7���E�{��h�r�z� �Ÿ�$�����W0�q��=m74/Z��h�����uYspq	���J4/.@;qn����* �_��YBd�L�v�@j�g�n�k�k���VD��VA�u�f����]�.Y�c���*���z� �N}��$�%�H�z����s@���@�;V��)���$��BrL�5RToW �� �YP���M#1I�8�L�<�k�;��@����=n]���6N�&Fܹx�{� ��w~_��r�X����*� ���V�j����P��QH�n#�E�DQq���x��m�s[�G;:ku]l����E�Q��]�k��ܤ[����n3Ϯ:��%r��v�٣��R��՜v�؀��:�kn�6ps�/9��۷<�GmҼg&�o/ �d�k�%����D8Wc/�#��]��\����	���6��E�u9|��l4��x�n3�99�9��D��U��84��Z�#GR�I��L5�NӵN�������ѻQc=m�l�cs�˫t]:�8n�Od^-2��4~��%@5i� ���v-�i7�Ȇ�L��8�h�]��ֽ�ڴz�����`��8	�4#ިޮ@;�n����ʀr�Lp#����MF��;��@����=Ի���ZʝdC	�Lh����7VTyP�[�wb��ʩ�c��$FG0Q�ġY��X苴�tl��8;g�I5cg�]9��ò5���{� �FTw�ط �Y�{-Sf91&BL�=�j�qE�H�U7���w$��{f䟺�s@���1�E�#r8��m�5�TyP�[�s�ʺ|z�Ŏ0rH�;[� �R�h]��>�w�S���a1L�H�h�e@:�r݋py� �:���ѵ[�u���8ێ�[;,��D�l5�\M�f�&�E�����G6�,���Lj�:�r݋py� �FTo����$$sQ���j�=z�h�]���zʝdC"�$�0�-�~��ٹ'�;�sn����%If7����~׀~f���rEp�D)$��K��r��@�v�׮�^�Zi�1�c�d$���zv-�5�TyP����fR�P�f�gpes��NG �s�(o��v(��eГ�Mur��q-O�o���׀}��X��qw���x��Mt"X�ɀ��E�z���=Ի�/Z��j�/�S��m��29#��o#*׫��[�k̨st��Q5&�4"L�9zנw;V��ۋ�XR��V����<����"��I�Q���j�=z�h�]���z�`*��N"fI�� k	Ǎq�䬶'���n�w�=Mi���׷[0�E^���	"�=z�h�]���zs�h"���I!j!I&h�]�^�@;�n�2�Թyw��S�ę	3@��^���Z�]��K��{��q���b�&F�q�ط יP�e@:�r�{*�D�FL�-׮����9{���>�;۹&# � ���~q���.x��q��	����6�ں{�� q����v�\�Zk�Y;s�s[5�����`Jr���g49ڸ.#���v�pm��v��������|t�3��ey�Rs��[\�-b��#�-��Mek�k<�<{6B�Bl����ݸ]�2`��Y�>���\��-t���%n{��s�A�{' ��ls�;l��E��F7T=2Ra��!����@ɣF�74\4�Kr�َ�g�ګ�W�R�:N5��*F��TJ���"���o"i�2!I$��w�~��9zנw;V���s@�.��4ܘEi�"�<�ݼ���M����v�,�K��yu�H�$Ȥ���zv-�5�TyP�\�}��޼��	�$�@�빠{�w4^���ՠ|�s�$#S���7�� ���v-�5�T���`�yf��7E�q�ű�u������P�V�U5=���e1s��u��z� �Ÿ�ʀo#*�͘�n�8ԅۗ/ ��u��IUm*_3�2��ʀu����U�Xz�d�1
9$Z�]��K��r��@�v���7�0���LP�L�=�e@6��v-�;�T��a^��w"#�팑`?n��R[�����ۚ��s@��A7ZK�9 ۣ=@�������g%�9_\n�3b�F�kX����9�$��c��J7�Z�~Z����K��yu�@�S��r$Ȥi�I��qg$���ذ=�޽ל�6q��X�rF[��H�w.� �W!u_>W����[�w,� �ݶ��c�eț�ԋ�R~��v���n����I?w.�����W-�y26ԏ@�v����o��g�u�~��<��@�QLˍ���`ԄnN�u��q�a�mwE9	��4�u�N� t�Wc�\�?o{�s���[��'�$���� ��n��mzs�hݔ�CBSa2\$� ��n,�R���%vk����������n��V]2��oB$�绷�{׺�ꪦ�{�`�; o���[�"�7�w/�*Ovw<{�lܓ�ݝٹ6�`bA��	RV��UK�I*M��^����ˎ]�$��$� ��q`�R��ߗ�<��=�ڴwQ����b�b��&K7	��(�0�f9VQ��;����)pN�"<@�18�hjbD�4u.��mzz�_RU_�n�b���m7#�e�Dݐ�`=ݼ�_�T������xw��, �R��qsY�8�F��zu���Ň*J�&�o0>����n�Lr��R�I��~X��������T�'�;����14%0&D)�4�j��������>��ٹ'W�$ҏ�1�H,$c
�tGv��|�~"Hl[!�"��,�� �F D)��|8!���f�42�\���Fd�Ni_�D�a��	�$!#"Prq$c��XFƭ!BH��D�D�J��6�A�5531� D� ��R��9��@��`Ȓ$bly�L"�&1�CC�X~b<E"8�+D�$!4<`�#����$�A��� ��D��,��0	�"@���ј 4@D6�:��@t1`��$��t#w���əu�,�2�N�5�;��<h��>8�;.�ק+P
�`��^�(��g'I['4�2C��δ�.;V���<@pR�i�8	jL`���'<\%뫲nմ��kv.�A��-�I؊I6���F�8��\���:z%�W��vM.[��sF�X׍]c�wX���l�%�M���;L��Y"���d�J��wWh��[V�$�$��<����m�Nӛ��=��[�%�������X�9$���i�agIe^����ݫ���9i�v�Z|*'p�U���[c�ywkm���:�Y�C5x���m���u�r�ļu.�k�NAgTV�7n^;.�v�D�n��0�3�Ѝ'E!�$D�۰����Z����v֣��N0.�Ŗ��k6�,��m�*��
R��D%�����w���`B��v�����O�{Vy�yy@t��s�W��(�8Ý��;��y��[��3g��e�p��!��4��ln�O�l���8��T�����XI�n89ܺ��m\<�7���a��K�wV�{a׹6���O[ʴ���L�9r�gVݶ�"��'V�\��]���]��-qiU��E݂㳱]*շUmM(�<@q�&�u�d+v.; q�3T]\��<�tJD@]6���+1�w[WQ�u��;h�^���hH��H;n�W[fX�@&,<l�ٍ�'�Lӝlt��uZV]{n��&s,񭶒�(-��P�����(��������sq�����P���SEh	���a�N��*	����<�����:�m��i�8,@�=pv�.yT6��c�c$َ�uaڒ���ns�92j��mA�Jl�!����Uݒ5L��G#�-��k3H�\��]�]Û������Ag���Dn�2`Zɹ�fw;u�r���Hzۭ�9ɴ�iؒm&`mz%��Q�0��mNѰZ���xU6:�3�6�ݡu2[�N6^i�n�wa%�v�3�ik��m����r;$pv���������6��@-T�І�@ 6�~�r���ML�3-�b-��8ً<]lz��Mt��u�^X��0�Y�2Be�:NP�PGx���sʹ�Mɶ�W��/�60,�搞��e�zN�v�Ag�܍F��]	$�HWe�.�+���z���%�pWT�RY�:�zt���ęj��8�豷N;I;x��ҥ��s�#ٞN�݄m��rh]�j��Y�G90ٞӴ�;lE�',rpY6u/k�m���b�l\�[�*y���5�������~;�P�com2OW_�@�v����ʩU~`{x����-ے7.�m��d���* o#�ڹ?|���gύ�q�jK��D���ذ�K4�٠w;V�}Kd�7��l�,T��x�� =�� ��u�r��{�, �]�ۖ���M�	 j��wb��e@7�� �j~���~���dw0�
:S֎ܝ[�3ۭ��Ҡ'\7=M��\�z����|��C���2V_�����.ܲ��ʀ��mz&6��(�h��m���b�����;�� >��{׺���$�����V��dE�#�,��b�[f���Zu��uYt����&�I��l�;��@�sC���?}���Y�m85�IG���p� �FT\[�}�����m[�^�X.�܏n���k�U�S��s�Y+�'K%��ș$�qF�H�E�w[� ��n,�٧�U/�;��������14䑡��L�=Ի����;��@�s@/e�%!�"LI��`n�0z�^�*�B�H�Im�Ēv�E%Y����x�X�MQ�c����+�\0?������xw��,�K��z�M�]I���Ʀ1����w,��2��Hv-�������L�t��nc���\��nF�Sۑ+�E9O��l��n�ܯP��k�W�_��o#*��wb��eh�e�$x�'1���f��e4z�^�n��>���?��$�9�Z�v��p-�C ݾ�{۸�ꪤ�~�;�����푗p��D����,�i���f��R�HN]��N���䓟O��9��#�$I3@�R�h�S@�v���ŀu*T��Vrwm��)#����\��m�s�r��Þ;�v�s��!֏�.�ZJ��" �x��O�w;V��n����>�H�19��cR�{׺���$��;���`���,�e4lT9�̑�8�h���>������8�7o������S�E$��K��z�M���9'���`���B��7q]ڰ�J�j� ط �YP�P|��/�Fj��ۚ�ur���I�W4a�s�)�uE��&u��k�מ�7)���l;n��ҹ�h���l�وzcKx�P�g�u�q���Ѯ�<ڗt���K�͚ueӜ���u�!6�N�nǱùy��ޑ��C���JQ�ט(N4g��+�B�&�GJ۔�x��G%ݴ�5G�ku�/j4�-��u�s�m��xk��P�q�X�4on͎;��w{߽���}ь�)��tA��p����6�$�'�(ش�L�F�p���7X�nȕѢ�!�z���n��>�����U_Xo���0�]�jH5D����,�J��=������u��%M��w�1����S$��u�~��>���uS~{����X���۵ae�bv�r���}��`�������>��� ��]"�� �y#I�3@�v��b�{{����ŀ~�w ~��\rB�̂�-H/�}���[i�ns�]Vq��WN�]�g#up<S�4�A'!"rH�����>�����_䒤��UW����������m�Z�	"�>��{U+��o�X�u�}�Ŝ�RM��ڜ
Ki'2G�j4��~4�h��h�ss@���A�8%��HR�*T�ӹ��ذ�ڱ`n�0���.[jH5D����,����o/���`��^��%�YZ֮��hzq�zz{Yg�%��ztݧBIX+�l8�2&�$�7S�$I3@�뛘۳L�^��J���w� v��mA�2�N7�4[)�w��@��ŀ}�Ջ?�U$��UI]��O�VI�j8��� ���{��X:�WUT�7��74[)�[�^&nc�r��rUI��~X�yb�?n�0?�{��������#-����Ȱ�ڱ`�U}ݜ~}}� �������ݐNm�tn���n�ͭr��s')l�ӗ�9���#�n÷v��um̻5��3�`�f���׀{��\�~a��X�~�]v]��$���`��^$�l��ŀ{��,����I*J���ٯ����$����D����� �}��v���Z�-��Dț���X�?v����������m%J�*��v��hݖ�S H��y3@���U9߿g���Py�Pޯ�����9:-���s�Ld�ݒ۱�����:85m�dHI�j�h��Vm��?�o ��q`o�b�I~a��~�k�ɓ71�8ܑ���ho�b�>��x�۷�ԕ$���������iL#��_���nh�է�I&������X�b�vIr�Z�娰?�U?t�x�w^�n������?v���{ֺ"컍�Icd��?�o 䪿�*����|�w�ŀ}�����UIyE����7e�jKjX�T�=a�������z.�0���n�ψ�Վ��;����j[l9��9U�SG=sř�Lv m/)lT�t�/����^�t���8���'z�[��:͒v\ۍI >Z���1m��ɺ��X�s��hvwk��-��u��v��rZ��ئ��q�x�z�eμnm+�:�v<X��&D;.�s�{=�3��}���b�〣>��;��lt�����*�ώ�q�][�T�u֧��^Ĕ�\��뎊����b�>�jŀ}����*_�k�u��wH����;��$� �}�R��g�����׀{۸���*l;Wu���!�hN7�4��~Z/Z��w4^���}�.�FB(��M�������,���XT���w<���Zd���"����n���74Wj�9zנ�.Q�)�<��7-�y�nz�8jG�l&}�ր ��[,Mu8"�X��ʪ�^)���)v�"�p��o�)Pqn׫�� V��eg�&����3Xhܓ�s���E� ,DR�UU�J��~�w���V,�*M���tE��M���q���x����M���,�}� ��^�RLi���E#�;���=z����^�%I$�_M��� ����"��2(��l�,���X�T�{�s��w^�n���֍2G��$��������u;d��u���Z�D��sJ��X"��L[��w���j$�E�8�L���~Z/Z��w4^���}�.�FL$�L������R�����X�yb�>��z�u�H<Ī	�=����~�s��C
X�4,�S4!���J��k�cVŇ�@��H�cHPI�e2���S�"H �`����\D�|4P��h��M�1q�F+"�#�K��8'�P��� Ȉ�Eڀ>EUK�Tc�ߞ�����k.�����\XJ����_���y��zu���(Tc���<c�&hm���/�UT�M�������X��Y����bdo9�8`�d�8��k���\�b�n�N��\�x�p��h�M���Jspq��q�n��{q`o�b�I/�>��x���jH��,�&����e@5�@>�� �����Wʪ�q�%6E(�q6I��X��{V��ֽ���^�Z"o" F�r�E�ʩRO�� ����=�n, S�R
i�(k��?�~����]d���dmȴ^���w4^�� ����ꤷ��r.�qI.0�7`�@h�iN�����G]����ql�s����~w�Iy�츭���rK�����X�\��>�ՠr��@���4�DIn9q`o�b�T�$�����߿=�����Tc��7�ɘ�{� ��v��*ow���X�~�W�v��wc��%ǁ���I������X��X�?�%T�ӹ�{ϥ�%��"j9/ ��q`�*��������������%��V��#�n�cVg�]��n�;�1��� ru�k{u�\�v�ecE>��&ܳ����t�S��'c��샃�7:�	ط.�'=68�q��@ܹݢ�lp��s�Dsq����]E�ҡs�b�9�t�m
m�u����f��k�/�"�muR�!s��ڮc�Kg;�8zGp�F3�[�F����и0;u�raM�i=���d�n�q�����pf%�h���l��� ����W\`��������l����L�������ڴ^���w4
�-�$�LQ�?fW��Ÿ^�@;�� �IS�UIW�T����xչ-�v�DR�H`��2�̨�J�}_$y�x\��A�$��^*����~X����>�S@��^�}�*ID�H\� �wLX$��������xw]� �C��N5�Bb���cY��Z����,v^^ͧ=oiy�ve�Qvѹ�r(�hbP��}l���ֽ����i��U��֓$��#I�Hh_��o�����7��{�7$�߿��ڴ.�Ǒ��F2bȤx��ŀ}��,:�*M����~� ��d�i����H�f��i��}^��<�ݼ��'���`�wFKvD���L��}]�@�W߿?�����=m74qT��B8Hб�8�8�����z�[X���ζƅz3q��
)��]1��6��dmȴ^���w4[M��*U���}� ���v]�$��d��PT� ������>|�g{T9�7�28�E�{��X��Z}����sv�����T�,q�˹n�r�X�$������<�����T��y~X?u��n�p�����\����_�k���R�\[�u%I{ۈ��ڱ����F�M����q�z�mq�VagL����T%z.&rS���w������܅�4I�ww�,���X綽��Z�:����!�&ho�bΪ������7���{ۋ?�*T�v��d�n\�C�v��>}�x��ׇ�S{�ذv�ŀ}�i��$m���di���h�w4^�����/���C�߽�ܓ߽�d�dDw, IrH�{ۋ ��v��������;�ՠ^"N��(�5�˜z��uƝ1�k���1�1����.m\h��QD��׮nh+k�;���I/����ŀw?�cW�$w%�W�T��[�ws*�5*}�]J��|��nƋ���w �_s�=� ��ٹ�~VנyuV<R1� Ț$� �����ڱ`���*�{���y~W����!�&h�ss ��v�}{� ����
����B(�n�?�������V���E��s���s���/\3���#�.-)G*�ՈvD�ɸu�wr<�nn�u�ϰb�Y�G;�<G�ܝf�*p�1Qtn{���#���4�@p�4�����dU�ZF�؃�;d�ۍ�c�Lv#� �&
x�·g]mq&۳�X�#g�K�ժ����I��r�����[v��ֲ/*��(��c�Q��;��'��w{�ҟnw�+q��kT��idyޞՆ�5�9&0�T8+�lQ�z��c~�w{�����ܓ./=�V�߳��v���e@5RV��u54��(㘦F܋@�;V��n��>������I%M��:�E�r��$� ��ŀ}��,?�UIS~��x����yCYm��r��K���ꤒW����� ����x��׀w[��wUu$O$�r6�(L�5Ÿn-�;�TU%@7�'���qrr���"�KKa���-k<�L�1U�K�*v��o�{���矐�的���������;�TU%@5Ÿ��ȉڐdń�h��m���K�URWf����{��x��'�c��p$��z�nh�ՠw��@�s@�nX��r
(�'&`*�����*�����v����=��X��s@������(㘦F܋@�;� �I$��I$�����|����V�z�,.8��I����?�}��]��Ϟ�ۉ-���$��գ9�.J��[�[8��#�~��=z����Z/Z���T�K&5N��=z����UUSg�����׀{۸�{^��p�F�(�f���Zyڴx���Z  AO�����Ѐ��U*J������ŀw��ŀk�ڽ�����CDqh�j�;���=z����Z��ȉ16�1dR=��,�RUU�T�Uo�/��o��<�����N6`2B,��3$ȞG;s��Z��[��vn<�v�+��[uv�����ˑ`o�b�>��x�۷ԩR��-��s@��?G��&D�8�3@�u�^�@;�TU%O�WϕWf���s#�I��ۑhw��@�sO��T�7��1`��x��j�ʻ�,=��{� �YPT� ��w���0P(yT]}�f�������SCQ8G3@����=]�@��^��n���Lk�0�"PP�ç`�!<���9��N"�vcm^�Ѣ7#g�ڴKlt�P�6�(L�=]�@��^��w%IR_�{��X=�W�ڹarU��\�W �*�����u*�T�<��H���"j9/ ���TU%@5Ÿ^�@>�|��3�I 6\��$����� �_s�<�ݼ�UJ���w�k�:Z��q���Ǫ�-�:�rܲ���6A �n	�|P��"X�`F��s�+����XWjH��0�sB@h�����$*,� �X,T0�m��+X$ � 1 �m!�h���*pB.�(Dj&�14�)���<b)"G����!�ǂ$FR�D(TU���N�Hrg�əu�]h�ZԺ�N�;V��ݳ.L����O'	���V�X������.Ҩ�WN,$p��&m5*�KpuRd�+��9�Eѧc�.8�4r8��e ��N�s��Dj�'E�zz��Os4��2v+r�;F�ܑ��݊ίZ�}v2F�i�`z6\��뭞c�`xޫm�fn$��p��t�n; 4#\�����wBK�5s���t��i�n݂�NF�U���q�u�s��uv������4u�3�
n�
�'m�w2�a��gp�6��3>��gy^��Ѝ�hr�'��TXx�O�0����ґhl�/E����S`��2�k�3�B�sM���v	&���:���=�a�9Ȁge(B�Yys@;�8��.�g�`D��U�㵍,�+G.�����Qbdc$��50IBcT<r!��\ov��nq��P���c]]�݀M�v���}Zvرq��v��Eulgj�Ц�:����7<�x�;�+[q5ư��oc*cHp�!R��`5�sDͳ��gi%vMQ%jJMz��]���'=
۪�+m��U�m��<�.�9�NH��q�9��r�!/[nϐ^��G�t�L�l$1ӗM՝�J�@��6lp�sV���+�QEQ�=��B���N�`v3�!;�]��sN�4�lW1����2b�W�	��܎ֺ��2;���uڜ�5�1h5�����t�c���l��Tm�eM	n��prj��gd
'H�.F����2�[t���Nn[���ݞ�5u\��c�,�7>�셌]��ն�lqb���lV`r �q�97/]C�٪hRٶL�k�úk:7^'o[�d^�D���v�8��+��ֈ��T�l�k��g�0�MO"������웛�� ��j(�[�bޡ�	����6�m�%�#�g]m���GZ�VU�t$�q(֘�&U�R]r��c=h�=h{�P]Q��%u����'<�;xMs����R\���Ueh	5��q�Y(�����=����l8��QV�W�� � Q�(�?T���gߓ�M �u��R�E��K�Y:ⷧ��uts���Hr6�-��xd��ag��M�ug�v!jq;���ۇ-D�s�v����&u��ݬ��;+�<��e���$����c[V�`��c:�6��n��{p�r�n�� �r;�����s�8ؼv�rl�qڰ.�u����j�q iŲZ۞�x|�Y���1�C8��ͳ���{��=(�9��9:,�ˁ��/a:�db^��ey����g�H8�Gs&9��ڑpu�@�n��>��UR�I~a��wl�-���7$zu����������ΥJ�$��j�5c��[��=��~��� ��z� �YP{v�'R�\vG.�n`*���ӹ���x����U*����~X=��K`���Z^����h�74Wj�=�a]�b��)�Җ��F�^����;n'�1nջJ�^+��NU$�H�ǒ2�ww,�&����݋ �n����O�UT����xϟt�v��.@l���1eR��U&Ͻ�L��v����?�U%I�^����"`�P��u�?^���w4֛���q'2c��894n���q`��*��?l�x���ӟ�Ȇ7$z�������^��5��x��=\]8�jT�[rW.�u��}h۔��5�0st���u���q���$�/���q��K������%��\�7��� �\�WW�D�HR#@��^�W�z��X�f���RM���_X�q �v�x?w^�n���eU$KR�AT�]�&���]�rO�{��.�ȉ�DBbȤzu���5�绷����%�J����^����Jo?����^���y[^�W�zu��{�Kq�<n8���(,�ώ7Cv㦤�m㵭g���fL��u����������}5Ƞ)�|~�-�Z��w4�T���jq�d�
Lm{� oW �* ����-��.����cN7"8�q�����z�[���M������x��(���'�h�T�Wj�9zסsU�*��;��Xv��M8�q29vӼ��\[�u���e@5|��???�8��p���uV�6�/����]`H��tm��#u�[�ɪBm�Yt�%٬X�#�@�;V���s@����}]�@�t�&�I��LXI���s��ɞ���_s�=��䪩���zJv��$�m�������^J�*o}}� ��ŀ��WC�B��;�K �����*�� w���@�()1�"�;�ՠ~�����������`m�URK%J�IT �@;�t�t�fMf\�,̴�3���qs���۳���ۉ����yP�����͸�h�X�e���y�ɠmD�i��N�ԋ����]v3�\����&~l�����6;b��mIٝ����8������q�D��y�����%��db�s��ts�-s�s�\[k=[E�qy��N�9���]V��v�3��N��nɑev�ny.Cl��vr]��a�ڹ6�1%�moN���K����<����Ju�7����8Fr�zh����?~J�j���� �Ÿ�^*�
diE�s4[u��h�j�;���;���D0s&�Ľ� �����*�y �O+J	H&&���;�ՠw[��z��@�v���ȇ1��1a�z��*�spqnۋp��7�!�5���ɫ7o6��伺L���'K�f^�\�K-:�J9��\g��V }�k��\[�v���e@��])#��\� �ou�%^T�������Z�w4W�h{��ێ$I�ڑh�j�;���=_U�z�V�oEq�Hd���nI�ܲ����-�;qn �W���1L�(�p�f��Қ����j�;���-�'	��L$?�y���a�u]���Q=ok�nz�3��E�k�[�0"lb���h�j�;���=_U�U�<�m(% ���Ǡw�u��l��b�=׼���o �oM��!�E	�	"�=��h���ss3�SJO����z�� ?i�"e�r����z��@��^��v��n�^��S$�h�ՠw��@�s@�}V��O�
�����R[bۤ���۲�`įz3q�܎�&n(�m�!�4�Zyڴ�w4W�h�ՠ[�\x9���v�I�n�ϗ�+���{�����O�T��M������qKn8�=P��\\[�v���e@;��&��(���U*���������{���w$���f��
Db� *�1���t�*�V6��LM
C@�;V�ܲ�����>|�]̣?a�R�F͈ඹG��}wk�.^o7Tv;\i��E�����{����s(�qڣ��~��%@5�n��p�[�Q}��I��#�I93@�}V��v���Z��Ŝ�%M�j�WM��8������ �Ÿ�ʀk����q4ۘBdq���h�w4����UU?ogv���r��K���"�=��h���=�S@�;V�g�n
�A�fAF�F��Jy3�n{m�۪�[5u F�����n�'4c.�vu�.���-q��MX��u�M3�lȑ���7vS6�;��C�s�l�8���<��g�4Q��kN8[*�0 '�e[8v���0Y��8g�j��n��v�V�.���!���n$89^�m��G8`�`�i��q���&�Ѕ6���(�;m[A{��w�8k[7L��r��Z�rݭL�.�-��<n&7�<�uur����h�;����x��L�^��IU%����s@���n(��p24&��h�S@�Ÿ�*�sp��/,�w�;��0}{� �wqa�T��%T�������?�绷"����ݑ4I.�2��7 �|��[�V�E-�r��mܑ`m�^�T�K�$�.�����v����>�n,���b����ֺ�3��$�;�!,OM�mۃ�8]��"�h�y��՟8������?�v��^e@5�n�����=AwH��r�}{�IJT�Q$��� ����b�Pߧ��훁��y�n�*J�;�>V���]���G�{��`m�^T�z��x����l�X7r9�*T��y�p���v��^e@;��Q�Ȍ�	��Z/Z��h�w4W�h���x1̋�Ē��`�v����@��U\����8��o��{ڜO5���S"cj7�^�-׮������z��ɏ���&]���2��7 ���n-�ԒM��ϤRے5$��rE�{�y�'��{���`E�H�"@��Z��R�X F" @���W�D�
$J�Mf��	Bą��%m`�	��!HRe��a�	��2`B:\%7��H`@�IR�!bVVY��q�G���i��(�Uq���"�Sm�! Ѷ�U��"@�#�!H�!��X�h� ��H�,`���!J�HBq�cR�D�,��t��F�h B$`��H4"�1a!Q�B�Rb0�V�1�$fc���A�kh��
�࿖�X%XՊT#@ ���Ype �_�� � GQ,B��$UE�@WH��]��:�S�Ch h������
�OȨo��}�ܓ��Z?䢙��qȴ^����^�����T��o<ݼ̶����&F��@��^�{�����_۷�*I?w���$!jԂnn�������փ��r�����x�n�ݘ�+!r֊.x9�226�$^����s@�}V�W۷�UK�I/�;o�������B��Dqɚ��
�k�;�ՠ^빠�e���b�M5"�*��@�׺��I7۽� �^��<��fۻۊ]��.��RT��N�v�b�>��hO��_�z/Z�ǍDD�9�G�o�q`�T��g?��}��x��׀�V�C�Y2�!����ύeա��M�;q���Nl��4]]5P��������sp�rۋp�T �-�D���qȴ
�׿��1#}}� ��ŀ}��x���-7r�%��5zyڴ��h���*뷀n�m����]���G�ʩ>�� ����|� �Ÿ=�謫p ��`m�^����{��������ٹ$��) ��@ �(�@Tŀ��t�J�18��E&��"V�
ᗘ��Dní��>� �e�k<�s���]pW.d5�x�����}�-ՠNãwnh'm]O6Ԏ��(֕�f���s�����ƹ�5���
v{=�t�p�A;�cRv���R��M�t�q�L��<�݌��m1�[���ڍ�oc�g�.�O2P������"���k�+=v��3Vᬙ�W���7t�)�!PX�f�8�	�c�R��]��N��HyW�q.��g�bc�\gqD����?�=��}����W���x�볮ݎ	L��j7��v������
�נyu�<x�DMc�a$Z븰���T�|�����< ���HH�s$�mɚ��
�נw��@��s@=KG��I8�8�Z��o �U�����ذ��� ׻f�p��'%�^���9�(ژ�*O]%l��ە�v:��ѳ!Y��ynͤ�� �Ÿ�ʀk���\�/M��pQG������b�TUR� " �� ����=��Z^P�x�DqȰ�l� �������J���y��ذ�ֶ7W,N1ܹp��UUI����wc��s*�_$���̼DL��j7��>�@��s@��S@�ֽ��,��$��Bd��Jv���8OO]Y����aݫ��K�ٮN�}��wg��<X8f9�E�����}�)�W���RJ��z�� }��HA�$���"�>���䪕&�~�}}� �}����J�a�;����e�r�x�w^�u��R�J���Wo}������r���I6���=��Z�ʀk���W �p�3�zȣ�wr�x��ŀrI$��y�_�� �׺��T���;�-E��۩�;ckh�Ϟ�Тtk].u��x��g�"x�����,1�"�#�<�?��r��@�;V���s@;��	�`��Q
;r<�����URI�}}� �ob�>���*��[LY2&6�q��m�5�T\��z� ���e]�%��$x�U_�*���������	>���ܟ��	DP�"�� @ �����܁��d��I�'$���Z��2�����_s�>�n,�{q����g��מ8�T�Y�2l8�6��'[tq���N]q��q�������獊���f���}��@;qn�2����zڙ����H��@�;V���s@��M��z�+&@�"n9���q`o��*�_�*����������z��U�<JaLRI&h�)�u���W �* w7O�U��2��� ��v�UI%�����}�rO��]��iq��"UT�I��~��~��ݲ��l[���\"��s����95���RvC��ř�Cvb0޺�!�c�����z�g��O��i2�d0D [c�K��[C������ss��0���2v�o��}�	�?Q��qƞ�lw)���6嶱^�)�6wm������N�[	lU�D0S{u�]<섭�ƻ��q��c��ۍ%TMsvzq���3���q�a��]vzi�%v2�hkm:8NG;��֛`/1�.��RH⵸�R�L�%��%�ͷ��� �*�y o9 ���eY��8�\B�K�=��,�%J�g�g�_�@��^�}N�6�9��LII&h�7 �y�^�@;VT z�����8�8�Z����h븰9%T��y�n�Ywr(�R����n-�;VT\��o9 �����nng�f��s�HsO.�g�з�z�ٌۧ��s����7}a�g�v�-r���wb�>�M0��o��%�����ۢ�!Zn"0��rE�}��y�+�ϙ�Z�����jʀ���ɴ[��v�x�}��y��xu%M^��s@���Z]͕�o&9������J�'����7�ذ��� ���.��x��2H�@�[��z��@�^��ֽ��H�i,"!t��v�ݼ�5YM'{`m��:�I�\�;��2��8��{�~�ԧn��]��_��@���@��_��[2 ^θ�r5�0NI�ܠ��-�n����:��>�|�샑G��r�����䟿w�7:	�H�� �"A@�D`�TE�X	�j��/*����禘��m���e���	��&�h����Jh^��*K��+����p���`��'%�ި��m�����* iB�II�<C�S!�@�C����9ug�^\�f���BC��2�zf�#�\��[���W �� יP{� ���ZA����@�;V�����v�,ݳ�����>{�b��(�y#�@��s@��M�Z���x�M�.�r�Iqۑ`uU'��� ׽׀{��x�*��T��T���U�U�U��>X�V��\���C�~� ���n-�5�T^�@6��������KElZ�n��v����:M���vp����+���\��t��7M��S�/ �׺��w��i�UI~a�{�������x���qH�u���Jh]k�;�ՠ[�J4�Jc�"r9"�>�M0��o��&������nhuYa�51N8h|� �Ÿ�ʀk�H|�c����	ƙ�@�;V��s@��ٹ'��{��A��4!/��O�QMpe �
-+ �XT*����F�Ь!
�R�0B"Kj�Vτ�)�#���֌L�]p���HEi���J�#(B�+)!iHД%-����J!	X�"�eaXV YB�B�RVR1�HA#	B��(6��8���l1 "@
�-P�X��"H%!R����X)R*0%#��W� `�bD�T"8�	�4*S��D"�!,�a%
QK*R�`��?�����	�B�Wd2�ڞ[8�m���v;^�pQ-m*�f�VS0l��*�ڰt��0�V�X���O�S���N��k����1*��p���SYv�7hg�����C�{]���8%�w7h�y�#[5�p�Dn�٭�َ8��m����i�q�.=��=�kX�0P	�
�n)���:���^�Zݭ�
�f�-��3��9�L���qs�*l䜸G��q�6����{v���//F�v��ݫ��T�ې��.���"��q�ܝ�}O�q\m��9R�6{�8{p�m����i|K�[��X�qgi����Ĝ˭�ηTΝv&e͌�@\{i��n�S�7��]Ӊ1�I�r����}8}���r�N7���R���FtZ�r�������8�v�Ņ����Ì��M����ڧM��'N�9����Ѻ�0󭳬�v��gݑ�H#k[��m÷i��;!��7l{i�:��x�`W����!�wn�2<lg�#f�T�� ���@�r�.Ѧiy )Μf�9s��ӷr�f훪�ŀ�@1�i���+��v5���r��Z�lHNmʱ+�'��[��*򀻌N4i+�EK�؞Q̰i6���@���:�E[.���Z��nb��]�[YI�lwCN�$M5�F$ݶÅ�������lCq�.i",?W�e~hڸNї\�6�{��Cl��t�=r�@Ξ�[�3�6�����Ui�.
 �,��%7B����g1;;)�-N�;4]�L����]a'��/��:ՠ�c��U��oe:ڜ음t�#�m7,rrmf�j�]lq�(s\;s4p�����,�k+ɢ�C��&ť[�ֹ�#�m�óU\<CA��y���wg��6�"��m�B��Q�m��j�%pq�N0��� �MW��L�>��=T�hT����mV�8b�Ͷ-�5��V��0�,��!�MٺJ�r���b�x��l��cv�nN9d"fܴ�V{c�*��"ǝ��֍f�kY�  :U�E�E��!��ut�� O߷$ч�\3RXd�2������V9�tX��HpQ٬�g��LCm�q\>X����o�dfz��]Ϗ\��Q�J��Bn�W)d�v����ѻ-���s����1۶��:����g����s�4��.�D㢰�c�ml���,���ծ�0���sn��6� k!ь�s��gN�M͌7p=+���A͍��D�����a�m��n��_��w�O�;�պ�:{].C''mwj��-�a��#ek�[�����w���}2b#��y#������z����ֽ��Z�-���L�G0H�T^�@6�rۋp�?Wϟ*�$�_���7�<�C@�~zz�^�U7��ŀ{�q�~�t˴BHI�8��;�ՠ{���=z�h*J�S��u��:�E�Dd�K��G�}�n,�$�ݽ�~�׀{��x�~~�ᆵ�tĜ��Q�m�b�9�g�{gF��I�B�h�s���l��s\{מ�@5�T������ʀ����iۉ�w$X����U���(xD� A�&{7�w$����7$��n,����{ֺX�E$�vK�x�?~��ʀk�H�.@6��W�fIl�Q�D��?�$�~��� �l� ��^��v� ����
d���D����m���W �*�)��~����%s9:��јnr�z�����5o3R�m�3�y���K����ː�\�o,��_*��w�߈���kDRd��$qǠr��@�[��z����ֽޕ���]�$��n��>�M0�/���$�	QJ�I5BH�JO9�x������Y钳Y3E0��ִm9ı����ӑ,K��;�fӑ,K��}�fӑ,K�����"X�%�{�5Ќt� ��ۑ�/�&Re&R��{6��bX��1�����O�,K�￿�m9ı,O����9ı,�.���糛���,��.ܭ��!�urĴd�etl�2'������}8�K�˓Y�ͧ"X�%����ͧ"X�%����ND�,K�k��ND�,K��{6��bX�'��{4k!�ճXj�CW5�ND�,K�w�6���ș�����6��bX�'���ٴ�Kı;�{ٴ�Kı/����-)n�!��YK�I��I��ۜbr%�bX���ٴ�K�,N���m9ı,O��p�r%�bX��;�kY���	sY�M�"X� �Ȟ׿��iȖ%�b{;���ND�,K���6��bXW`D_"9�Ko~�)~)2�)2����8H���̚ˬ�m9ı,N���m9ı,S���6��bX�'���6��bX������_�L��L��ܛ�r\��=XĜ�(<��S�r.�Y���[��ջ=�V\+XWi�\걑��}����=�{�O��p�r%�bX�{���r%�bX�w^��r%�bX�Ͻ��r%�bX��f�J�����WZѴ�Kı>�w��Kı>���Kı;�{ٴ�Kı>��iȅ�b2������8�n��)~)2�)X�w^��r%�bX�Ͻ��r%���"dN����ӑ,K�����6���L��]{�Ĳ�E$�v9q�/�%�bw>��iȖ%�b}�{�ӑ,K���ߦӑ,K�����ӑL��L����R�.+R�pw/)~ı,O��p�r%�bX����6��bX�'��޻ND�,K����ND�,KB�y|L0�I���Û\v1D�9�S�竴����Le�1�V횳r����6�-�#�����toe&;b�6{s�;���bG�+�n��~ݝ�=u�g�nv�/�l�W"���كG!��ݔ8�z�DY;&ݸ��*���ǲ��n�+�c [O<�ϛ�E�!�۰�j�.ͲY]ۧ�6�C�h����
��֯m���R���,�Ei�:��[%��1����{�������˻g=[���#Ճ=�M��Z+������y����1��8{f̐hqKwq6�ȽKJL��L���g��Kı?w^��r%�bX�Ͻ��r%�bX�w���Kı/�{��R\v9hw.C)~)2�)2��;�'"X�%����ͧ"X�%��{�ND�,K�w�6��bX�'�{���d���jc�w�{��7��������9ı,O��p�r%�bX�{���Kı?w^��r%�bX��}�v�q8�p�vI/)~)2�)2��{��r%�bX�{���Kı?w^��r%�bX�Ͻ��r%�bX��f�J�����W5�iȖ%�b}���ӑ,K���{�iȖ%�bw�{�iȖ%�b}���ӑ,K����?KËF���zӕL)e���Wk]�z1ղ-�&+Dsmlz���5w�Ȗ%�b~���Kı;����Kı>�}�iȖ%�b}����~)2�)2�_���X(�A�n�.=�"X�%�ߵ�]�!E6�r&�X����iȖ%�bw���"X�%�����ӑ,KĽｬ3	�4aL֤&�WiȖ%�b}���ӑ,K�����"X�%�����ӑ,K�����ӑ,Kľ���֦�R��ۚѴ�Kı>�}�iȖ%�b~���Kı;����Kı>�}�iȖ%�b_t��4�5&�\.kY�iȖ%�b~���Kı;����Kı>��iȖ%�b}���ӑ,K����g�K��e'3����۝ۇ�b�Иwsm�������غ3�V���O%t�M��{��ŉbX��^��r%�bX�w���Kı>�}�iȖ%�b~���Kı=���p�4]Y���fj�WiȖ%�b}���ӑ,K�����"X�%�����ӑ,K�����ӑ,K����z䮲fh�E֮��iȖ%�b}�{�ӑ,K�����ӑ,`�P?�bq���`E��]��Ȝ��k���9ı,O}��ND�,K��=�4J�YK�.\�h�r%�bX�w^��r%�bX����Kı>��iȖ%�b}�{�ӑ,K��w�鬖.F�[�ˏ)~)2�)2���yK�,K�����"X�%����ND�,K��޻ND�,K�ކ��X�o��n�.�'�3��z�$��Ga�v]viЗVd�I�M<���7i��܉bX�'���m9ı,O��p�r%�bX�w^��r%�bX����Re&Re'�㤅��wm�R�Kı>���iȖ%�b}�{�iȖ%�bw���ӑ,K�����"X�%�}�ޘܹ�5f\.j�Fӑ,K�����ӑ,K��u�]�"X�%��}�ND�,K�{�6���{��7�������VR��i��܉bX�'{�z�9ı,O��p�r%�bX�{���K��>A?V0�@� @$ �� ��I�c!$��a�)��bĈ�,`B�$���5�{�iȖ%�b~��̸K�WF�Mff��v��bX�'���m9ı,O��p�r%�bX�w^��r%�bX����K�2��*�T�o���"�H���"\w�ݎc/>$�r��,=��sv`ŷ\ܚi�����Ͼ��|9�!ܰi�rE��Re&Re.��ߖR�Kı>���Kı;�{�iȖ%�b}�{�ӑ,K��}OrM���.��s5�iȖ%�b}�{�iȖ%�bw���ӑ,K�����"X�%����ND�,K���շ#������)2�)n��Ȗ%�b}�{�ӑ,K�����"X�%��u�]�"X�%�{��T�%ˢ�kZ���]�"X�%��}�ND�,K�{�6��bX�'�׽v��bX�'{�z�9ı,K�=$-�A��m�"�_�L��L�������bX�'�׽v��bX�'s�{6��bX�'���m9ı,J�:�b����ܶoZ�˭\@�H�6
�8�$�bۧ,p;�ksq�M;���j״ux#Y�򔛣	�g)g�)�p��㫴:�M�p&C�nwc<�<�^E��g� ����u������l��<�C��L�Gq��w+�ͳ�9�Xw�3ɠ�.Gj�w��m�au3u����v#�-1��O�q��s���83�Q��J���V!��ݛ���7��:;�s_�����sS5��̛Olt��-�2m����h�۵�K�v����mO0����l�ӹ.,��&Re&R�����9ı,N��siȖ%�b}�{�ӑ,K�����"X�%���zs1�֬˫�љ��j�9ı,N��siȖ%�b}�{�ӑ,K�����"X�%��u�]�"X�%��wܙ��r��2k35�kiȖ%�b}�{�ӑ,K�����"X�%��u�]�"X�%�߽�m9ı,O{�����&f�J\�ִm9ĳ���;����ӑ,K������ӑ,K����6��bX�2'�����r%�bX���?�M��[�Rf�kZ6��bX�'�׽v��bX�/~����Kı;�{�ӑ,K�����"X�%�����ߦ��߽����s7Wm�Z��r��Ah���ƹ��Ӫ��7m��׆�����*@�-�t���
�����	�~�q=ı>�{ٴ�Kı/}�j����f���5��Kı;�{�Ӑ�
�Lr&�X�{���Kı;�{ٴ�K�e-�w^R�R�Re&R}�:Im���D��Z6��bX�'��m9ı,O��z�9ı,N���m9ı,N����Kı=�=���jj̸\ֳFӑ,K�����ӑ,K��}�fӑ,K��{�ND�,FR�o~YK�I��I��������㙣35���r%�bX�Ͻ��r%�bX{�p�r%�bX�{���Kı?{^��r%�bX���{YL3SXc�Ժa�;��淰�s���v�4/n^�jc\C�_��%e�rK]H�����x�,O{��6��bX�'��m9ı,O�׽v��bX�'s�{6��bX�'�����c%�0�5�Ѵ�Kı>�}�iȖ%�b~����Kı;�{ٴ�Kı;���Ӑ��I���,��q˷n�rE���K���{�iȖ%�bw>��iȖ4(�H�!�:1��-)Kx�@b��0H$!Ye,
�fӌ�"��	�0�W�C\���@�����T��6.��c�+|�K�~�{�!��������`p��_�H�|B�d�r8�����$H���!H�  ���* Q� D�!)%�� �q�X�!�		�H �FcJD	%��i��^E�ZB!�:�U��Ӯ3$��*��C$�J�!B1�A�b�C[�H�c�@ ������.����ZR�!$����$��7���%XIH�B�lZU�H�+X�Q 4�T�@���ȱ1!�A� ����Sc�"���,�)�b��ê�T� 4��Q0O�!�O���B
@��h�|�&�M(�P|v'�9��ӑ,K���}�iȖ%�bo�_[�	N�nK,r��_�L���*���=��fӑ,K�����iȖ%�b}���ӑ,K���{�iȖ%�b^�ަ�&fh��5����fӑ,K��{�ND�,K��p�r%�bX���z�9ı,N���m9��I���ͳ��#$d�(�������lt�c�5��O.����-ٙ1l�uR挚�˚Ѵ�Kı>�}�iȖ%�b~����Kı;�{ٴ�Kı;���ӑ,K��t�d�ԙp��f��"X�%�����ӑ,K��}�fӑ,K��{�ND�,K���ND� �2%��������艹Zc�w�{��7���g}��ND�,K��m9ı,O��m9ı,O�׽v��bX�'v���;�#�"�n�%�/�&Re&Q���6��bX�'��m9ı,O�׽v��bX���+� X��)RB0�D��Ng��fӑ,K���ۧ�ɬd�ѣ
j捧"X�%�����"X�%������ӑ,K��}�fӑ,K��{�ND7���{��~���E)��u���k���3���n��i�m��Ѕ����q��͵���fK�.�kZ6��bX�'�k޻ND�,K����ND�,K��m9ı,O��p�r%�bX���_e�	e�Gq]�.<����L��[~�(%�bw���"X�%����ND�,K���]�"TȖ%�����wqHE.1Gr��)2�)w���iȖ%�b}���ӑ,K���{�iȖ%�bw>��iȖ%�b^�$�ː�H�Ȳ��)2�){���"X�%�����ӑ,K��}�fӑ,KK��m9ı,OgN��eֲ�$��浚6��bX�'�k޻ND�,K����ND�,K��m9ı,O���m9ı,O�O�D�@�Ξ���]X;���.cɝi�t�rσ�m.���.8à1�r�k<J��^8�����4��xѴFi��Ĺ7�v����0&so��P�5Ύ�Wց�ət��鮑3Ϋ,C��Sg+cH痃wLm�%L��r��*�cgX[�������`n��6��]�;g�׶��p�6 G�.n4�t��ۙ	P�R�����y�� rg[�����r���-�]�,����q�5�b������g��֯\�3�3���t65:"nV���~�q�����?���;ND�,K��m9ı,O���m9ı,O�׽v��bX�'���e֤�e֍k.Mf�iȖ%�bw���"��bX����m9ı,O�׽v��bX�'s��6��bX�'����&��2�Ѣ�sFӑ,K�����iȖ%�b~����K�HdL��￳iȖ%�b{����K�L���!���pw.K�I��K���]�"X�%����ͧ"X�%����6��bXb~�w��K7������?Q-9��{���d�,N���m9ı,N����Kı?{���r%�bX���z�9�L��^��/��V� �jD��i����87ݱy+�ӵ�-#.q�%ʷs�8�ͭ��5���5u��r%�bX��}�iȖ%�b~�w��Kı?{^��r%�bX�ϻ��r%�bX�����l�j�h�]kFӑ,K�����i�tZ$���_y8���%������Kı=���iȖ%�bw���"X�%����k5sY&���ֵ6��bX�'�k޻ND�,K��}�ND�,K��m9ı,O��m9ı,O����]j�]]f��ֳWiȖ%�bw>�iȖ%�bw���"X�%�����"X�%�����ӑ,K������Ԛ̺ѭeɬ�m9ı,N����Kı?{���Kı?{^��r%�JL�����_�L��L���6�2�r���x�&�wu���ۄċ�y�.���!k�2 �.y��t��]u�#w�����d�>�w��Kı?{^��r%�bX�Ͻ��r%�bX��}�iȖ%��K����Z�c�qܸe/�&Rq,O�׽v��bX�'s��6��bX�'~�m9ı,O���6��b]�7���ߧ�%�R��Bc�w�{��,N���m9ı,N��p�r%� �TZj&�w}ߦӑ,K�����_�L��L��{��lwWj8᫚ͧ"X�%�߻�ND�,K�w~�ND�,K���]�"X�%���u�/�&Re&R}��%�w!H���h�r%�bX�{���r%�bX�����9ı,N���m9ı,V�{��_�L��L��,��;�$�N(ꮭ�9$m���vH'�����dռ�ήkR 3�<�q��.��������D��w�iȖ%�bw>��iȖ%�bw���ӑ,K���ߦӑ,K�w������L�3�X�����{��;�{ٴ�Kı;���ӑ,K���ߦӑ,K���{�iȖ%�ow����ǳPC]Hꟽ���7��,N����Kı>�w��Kı>����Kı;�{ٴ�Kı;����&����F���6��bX�'���6��bX�'�׽v��bX�'s�{6��bX�pb&�Ȣ��=�{�iȖ%�bwކ�&�umշV]\�jm9ı,O��z�9ı,?�#�w��6��X�%��p�r%�bX�{���r%�bX�{G}���R��h�`�Ɔي��R�"�3�i�.��˸��m"Z�*�&6��bX�'s�{6��bX�'{�p�r%�bX�{���r%�bX�{^��r%�bX������.kRf����fӑ,K��}�ND�,K�w~�ND�,K�k޻ND�,K������oq����~�{����*��Fӑ,K���ߦӑ,K�����ӑ,�!�2'���ٴ�Kı]��ߖR�Re&Re.�[�2.�q�ֳSiȖ%�b}�{�iȖ%�bw>��iȖ%�bw���"X���[�߿�����L��]��ߣ�#qˬ�L�fj�9ı,N���m9ı,N��p�r%�bX�{���r%�bX�����9ı,O�$�������һX����ԛOv�;����"��e���ܖ�� ���>:7F�}��g����Mۭ�:`g�÷�n'�n��8h��͎�ˌ�wn.m
�q�q�LJҠl�p��G9��i\�Ж�t���}|�*��9Ǖ�2s���;k��%��m;�^{�E:��c��:ĹE3i��cG��Ya.�ܯ-�,ie�]Iuu�@��!�Dw��O�+5k\�cc�ܙv����}�ݮ��@_�Y���+v�b�vg�'�Pi�duY�v%�bX�w��6��bX�'���6��bX�'�k���D��dK�]{��yK�I��I����k������-fh�r%�bX�{���r%�bX�����9ı,N���m9ı,N��p�r%�bX���Vk��u���SiȖ%�b~����Kı;�wٴ�K�XdL�����ӑ,K������ND�,K����\�ԙ�˙�ɒ�5v��bX�'s��6��bX�'~�m9ı,O���6��bX�'�k��ND�,K��z���j��WV���r%�bX�����Kı>�w��Kı?{]��r%�bX�Ͻ��r%�bX��-�������K����&�����l���vrN���#�9r9�Y������*��]�����K���ߦӑ,K���w�iȖ%�bw>��a���"X�'���O�&Re&Rܻ�[��XGr\2�"X�%����Ӑ���H0O��)"�PJ,
�
���n%��׽�ND�,K�}�ND�,K�w~�ND�,K��ܗSY���f��Y35����Kı;�{ٴ�Kı;�}�iȖ%�b}���iȖ%�b~����Kı=����f��f�Z5��5�fӑ,K�����"X�%����M�"X�%����ӑ,K��}�fӑ,K��wOfԓ3F�.�h�r%�bX�{���r%�bX���z�9ı,N���m9ı,N����Kı=�vOLnM=�����ʣ�n9X Z�R	�ے4��h��˅/GU��ݪjҮ���{�K���{�iȖ%�bw>��iȖ%�bw���"X�%����ND7���{�����D�	��c�w�x�,K��}�ND�,K��m9ı,O��m9ı,O�׽v��e&Re-��j�䌻Q�(伥�Kı;���ӑ,K�����ӑ,tE�W�+��9[׽v��bX�'��}�ND�,K��������um�[eִm9ı,O��m9ı,O�׽v��bX�'s��6��bX�'{�p�r%�bX���R�ܰ��rH���)2�)}ӹ��bX�'s��6��bX�'{�p�r%�bX���p�r%�bX����Z�V,��|�������'5Ϭs�s��Y�xM�um`zr��7��j�a&r�x�Kı;�wٴ�Kı;���ӑ,K�����ӑ,K���{�j�Re&Re.���Z.H�.E%�K��Ȗ%�bw���!��r&D�>����"X�%������ӑ,K��}�fӑ,K��wOfԓ3F�.�h�r%�bX���p�r%�bX���z�9�� !�2'���ͧ"X�%��{��ӑ,K��ާ�I�Xe�ˬ�W5�ND�,�PVD����iȖ%�b{;���r%�bX��}�iȖ%�QZ�� ̉}�p�r<oq��������H�������Kı;�wٴ�Kı;���ND�,K���ND�,K���]�"�I��K��gI#HYm\��e�c&�^8����f�j�p^�[���n�Ɇ���ə�Ip�Ն���ND�,K�ﹴ�Kı?{���Kı?{^��	?DȖ%��￳iȖ%�b_������lђ�ն]k[ND�,K���ND�,K���]�"X�%����ͧ"X�%�����r%�bX���R��e�"�_�L��L��N甹ı,N���m9ı,N���ӑ,K�����ӑ,K��}�j᩵J�r�{���oq���~?����w"X�%�����r%�bX���p�r%�bX���z�9ı,O{�/3R�Y�5�ѭdɬ�m9ı,N���ӑ,K������~6$�H�i7�O�ﻛA$O�U��U���
*�@QW�QE_��D�?� �EQ`��"ň*",�� �@�H��H� B �@ 
�X�� 
�@"
�`
�U�,@�H�� 
�R" �� (��`@QW�E_"��U�
*��U��@QW��E_��U�H����@QW���e5���Pd2]� �s2}p��P C�   �(
J
 �       m� ���     �
�D�B���%J@PIUT��H$(
 (P��T���IE
\  �E(    (
1��O>������QNmB�`��U7X���R�ťIX��U����T��%T�� �f        h (  @`���B�Z�Sҩ�R���R�� څFZ��Yj�S;r�*媕@  �(   �� �J�gn���jUU�u
���GN w���Ż[qu�{� �J�s���v��q�a���{� ����a�g��{x��@9�L����p;���8�z/ �T    @0hP�������g���3N��}��}������!��4�1��9�0 �띯��y�w��<�ֽ��ݠ���z����9o��w�y�.>�{�Y�Ҭm_f�oV������}���    �f�y��9�z�;����n�l(� ����2�t27^;ye� �)Y=�9�d�  7���{6�t�� >�xo��w����c֜���O^�� ��\ZQ���=�������h� J�(     {�
w�yN�ܔǳ�N/K����U �Gsh�˧���/y�������sn��x  ^�M;g ;�� xt���`�42��:w }�>�3��W3]�����)� 4�)S�JR���O�5T�� �<z�R�P���Ob�Tm�  !�T�Д�R���!�����5%$D 4x�������������h����BS�p��F{n;=����AEEz�r��ڈ

������TVEAS�������A����0����?��>���/��E��N�5��0##Na�2H�5����w�Y#A��\�6���1�XU�K0��ӭ�k
��f�Y��>�����S�7�����nap���FbXa�4a��==I��f^��u�,��9�>�e�qA�7��}��_5� Br��[����,�ρ)D�a	�%q�&�4LY��Lm����,8���HIL �.�<c0l5����[��X��&��Up�k&-�|b�����Y�,�h�F;�ncFØ!���޼���tc*5,[�������}�y�y��Ip�L�=H�$c�v��g[~�o.q����s=�A��`MČ p�i�9���F�d�1�l�#G��c�.�i�F�^������$�5��3��8sz4��I��Q�7�Vh��Yd�&8'��8�����N:v�8�M�)�@b� ��1��ȋ4��5��TA8����pח���l8���b�~�>��;J���9%��ดMU�w�.����'��!��c DA!���T�K8�I�N͏(�ı#Ѿ0AѦ�4�j4l�s#	p����ooT���=�1{���n����Y��F:6q��[�$a����ѳ�e}j�o�6�'<4���5���$�x1��kLkF��ݬL�61����������p48���a��mx��	/ ��'#A��Z�90@��>�8��6�h6�4n1��p�3_y���0PRQ�����٭�N�1L^�ky��qtmq1$�D2SD%��F��0��F	�V��# �Ha�����K0�2�I��BP���P&�������u��<��b� J�,��b�:'`�Q�l>OG������_쫾h�Xca��8N��H��m�,�I��3N�Z�|M%����{�y�p���#A��Pf��Df��^k�2F����ϼ!� 	xi<�C�t$�Ϗ5�%����l����u)œѵ�#�v�a8Nh�IL	<
H�H�2�l�4�O��d�F��#��0|ַ�|�{�cs�c�a��_sy�O��h��4�3[���#��f�6k\7�o�y�l�=���s[���K5�7�X�|�͞;2���19��nލF�.�00�t�Ȫ�����6j����M�#��Nl��\��y����|$��c��Y��q _V���-\��s��&��;������[mn޶��6�X>|<�ѱ�y�l�tFj1��|��Č���a)��1�z�c�c� �A�LB�K7�sF����x�k|
0��~Y��&l���>}�3^x��sA�螺xǆ��<�3\�`H���vS�Ŝ;x�����^�n"`"���{��lXYQ:��F!\�����ع����g3z�|y��|��z�A�#4�$f��fč�p8�zi�<��`j����|(]�6kMf�,�i��|h��g<n6�a2#~m�F݌��[њ4ٖ���������{����o���z���ǅ�ޭf6Y�2Z�5�(�0��BhM"[	m\��_������l�-�Ǒ�0��s�1��$����	����h'�c~0��4�!���81�~Af�D��X�$�j�C��	�;�>r��Ω����߯o#Bf���3ύ���8bQ�.Ec\1���y����S�9�T�d�߅���7k�8����,�=���k�|�ig�߾���<�~�=��^X�$K�s?���E��������s��s�Ƽ�҆�4m��=��4l �6i�3kes�$sfp#a�C�<�-e���y�~��64�{�!%��4h�F�,�3��³[�0�*�I��� d�M��&20$�t٭&a��Ѳ��h���3[��c��L�
C ����|x���&1��o>(�Y�n�гD2Io��4;0ѳ=��N;&��O��V�F�kAh��h�4��`Fi��Y��]��F�&��l�0�`Bb�$3�G	��eڐl��cA���Q�g�F�s�V�Br�4��uLw�?�N$h,�h�4Xkn��ih�0Dfj���Xr\�pN&a�>c�AI��n1�n��N1�a��h#caF���4��5��H#6��[ܚ��Ѡ�H"$�$��1� �4:#D�,�&f��1��
LX�̴n8�АiX޲��4�I�'(!�t�:��^�����aĜB\1�@@�9���b�DsX!z�Zހ°��7�[9�'=0}8�3K�30$�m&���٢0�p�20Ѿ$%%b:�=,�!��p�|���14��Y���I����6m#�L�'o�Y�[����`hjI�c�´�[����(�#2,3L��I�u#����i�`��$!&�ѳg�$��e�o �����F8d�:��6�E���h7�HIR�8A��J&+#!3�y,O�Α�b�[�0�#$�j"�If��fm7��;�4y�h>�C�Lc�Fs\(��-��� �0ٰ��J`!a���s|#�e�9�9�߼�xy���SZs/�����5�n�b'F�15�ha��|q�&b0�Z6[ׁ�r�TsE���H#a�I ��嚷���7L�C)�ǆ�M3���X|C!+����8a`�!��H��H'�
pt\��oe��	I$a=������(����ܒ��#0a�NBB_0��Î'��I��88�/�R�4�h4��$DI+$�6�"ѶHdpڛT�A�,3�i����Յ��P�±�X,���(�N�+���xl�o|9k�����f�l�8��\#���[��f��6�G��"t�52i=��(�0c�a�7�z�!���p��26<�3ˇ�7�г�1�ޙ�e40�$�FsH����0ַ�<瞶k6F.�34�-��99\C��q��s{�PB��9���4�oXpqt㑭a0_�s5��e�l4Fj{�7ﾇ�||���I1=@�\M!�@c��a��8�Bt08��S�x�z32��xK�o�f������`Xm6��20�������5��H	� ��ci0�9Í��a�t��j7��3M��s��i[��D�����F4a��1��������M�H��O96��1�4O����3^�oіsq���
	�{êj�}�y����N��V:(����ǀ���H1�o���Ho7�[?�$�Hư}� �p���4����;�,�C8r�Vq�����zmv��S �FhŒĜu������0C�>>��Y㎷>��sq���-�7����0p~<g5�����׾����\t.��ai'LH�S��Y�w�;M8h�i�3[>�[�� � � ����{��Ԃg����Z>o:Y���f�,v@�go����s[��<�m�/T|�Ă`��3,2�#� ��0 �� 0�&$�3$�Ĥ�i 0Q��Y10&E�����A�������z/������O_O3K���x���8$���$�I����N���<@�}}�XZ��>��&� �N'���I���LQ��J$�hM$��0	�C��\���0���d0I0d�Ґb��Ht�Hl\_P��c�o p��ӻ��m��   ���H lp  �H���l�n�[;]��[G �� � 0kh�,�M�n�8m��m��
���K�����NP��e뗭K.�l-��2[E� ۔�:^�8u�f���pSF��B޹�n���H�$�u�[	��u�K�h���P�`�M�6ZC���� ��u�� ��R�lŴ�UVҭ�U&EP6���a�� qm���@m�N ��p  �  -�h  ��h[@    -���m��m��M�m�[M�   ~�	 �[ͷl������#���` n�[n  ��{m�zP �R��ަ�	A  -�  Ԁ  ��  [m�6���`�   m��m�0 8;�� [@�   8H   mm ����  4�`  �ɀ8۶H �[I`$� -��m�� O��}������s�$HI��ic;��o���l�[�A#m�m�         q"C� ���m� �I� � �` l����`�  	  G ��a��p���j@ �`  ��bΖ���� � [I6�`5�� �n [D� HYˤͷ �nmn� H8    �6ٶ�m� 6�qm�� -�  @ m 6� h    ��m��j�r۶����z���m�`8 ݓ�0v�@���m   p>� (��� 	ą�v����'It�kdm[C]1t�:@ �͖� 8 lҴ��m�R%����C�sid��(� I�m�[�V-�u��b�a ^�(k�� @^y��y�&��Rʸ)�m! �smm�H�٥�	  �`-�Im�[Rppl�m�ĝR�r��/���&�۳��O��m�-��	8pH����-�ۛm��p8��c�]v���9���*�їL  �I�oV�l	"�"@
���iT��n��Ѱ -���\��9 [@H:\������ ��մ�Kh��$$ 8l�g���k6��j��\�iz� Hm H�d��v���Ȟ]�  ���<-�j�4�9�m���8����  ��i5�7/Y� �m�t�  !K��-���v�M�M+ ��vm�� m���履]��*�^ �l[z�Wrp@R��K��_�9�HN�%�$��J�2"1�6,���;f2N�e�7�v@큁�B�Q�:J4(l���*�v.�V��@evB�m��n�++��U�m�c�ڠ:��@�v�� ښ��m6����j�U�*�㝞��i	��mYA���U����F1���V!�gg"l�B"�-UU�X��Qˢڭڮ��c�!-��u\ul�i:N���mr�\&�v� �I4��`nۤ�6㬾�mI�ҭ��N)/-����j�6j�ɞ%�ڪ��\ mN��ݰ�Q� *�c���6){K.HH��9�v��Kz�����M��N����Q��Q҃�#��-[uN������@w�[k�b���[Um� �� ��\��UY-���1.v��m��`  �ZI[�3�trIe-�ą�/S` H�#���KD�I��۶-��hH6�෨\�t6�$k�L��p� 9&����t�5�5��,��ZlZl  	 $ۣ$�U��U�B�m�����t�7MR�3a��U ҳ�'(�g'�����:�{v� -���$ۖ����ٶ�g&����հ ���N8�d��N6��� $jV��8��A�m�: �`8( �2h�M��'$�J�N�� �6��pm����M���������ǰ��s�G�!��6�ڳm"@Ҷ�dH�z������}����j��E�[����	1 ���۶ʁt���Kn�N��;lՒ�n�r]�Lq����� *�P�������ʭ@U�Kn�j�iy�V��
���q�]@v]�b4�H΃���;K�6 9Í�$Y&E�5�m��&D�8,N��4�� >^�_���k� �j��\�F"�����ˇ�u�naV��Vl�M�<�US�u��km��-� 6�^��vw�����]@�Pq�d��h-�$����n��� H5��V�IS��I��,X�ezL͠ ��m-��Ѯ���j� M�i���e�II  {�-�$�\��o -� H @8����6[wmm� N��:��m��sBmw'@-���p .���d�۲��N�*�પ�"��\�ÖӤz�[@_��M�]$�C�����t�  �m�  m��   �.� �%.  �"���   �>�   ���j��p����� c6�u��Ś��ާ$ l p�m,�H5+ M��v�E��Ő���9��im '@�3T�i4�gY-��v�*��I��'glƴ�2�����
�8�H=[�I04�`H�k2�6�[ׁ��lx� iqeP]<D��������Im��A7$f����[\������hǵ7h�1%���Δ��N-�G%��v�-W�����]\���ݗ�^[t�`�U/(�U*�}��}�iPٷ"Z�	)��t�!��X�N�(�m����N]�m�F)W>D�ً��x�K͹@( #u61*�ٶ���ͧE+*S�68��]���^��[��C���xn6�fn��wB�������:��a����	x�uN�����[zM�iZ�R�'�� N�N۶�f�dlۤ�;n�'i��v���  #C�N�E��v�z�m� 4�n�h�)M��m �e��ZI�S`&Q�]F�O*�UUt�9vZU����i��,�[@� m���$Ml�X�[����6���6H �� ��[M�r����}F�Im�l�WJ�̷S��U�d��y�U��۶�����QI�:�e��8mi$�d����r�'��̜K�l 	6���m�m��d�f�C[@ mPWQ�"��F5B��m�մ�f�@  m���"M�~/��m�l�ޡn�H�  	8�۝�Z4�I  ��m�b@��@[/k@ 	Ѳ� �k��l   �
�v��*�ҭC���
m&�X�� ���� 6S`כ[@$$  u�h�$2�Jٴ�J����K5tzt���m�u��q 6� �ωӯ�m�lۮ�\���p �ͰM��� �.�A���]�۰$��%��۰p�`ge��n�P�
B��a�j��j��v�.�� �[C��$����_Sm�����ڶ   � i  ���K�[�RJ�TQ�$�m�66�J�l� !{m f�����-���Q�����f�K��m�cm� |    m�       ��n�p$ � [%t�YE�Rl,�mM��!���		gIR�i��[��h,4� 5/7+J�ԫUJ�@[ڸѭ�@H��$   � $gF���6�'D#�B��U@�UP]�Q�e^�cֶ��� -���
��
�Z�e�*�Ԇ�(d@檮��[Y�l�l-�$ �Y-�� ��F�   �u�6�9,�*��-UH횞I�Yݻv� �sm�	�Ų��T�J�v�m� 9! �Q��巀�lEj݃j�
���]�	��O(r�������U�=23M�-�m hֳl��$�v�Kۋu�6R�	2�%I˵�9ۢZ�p��L�Y)�k,MWE��熡�P���@ͫ`�� m��ln�!  �-��-[�U.� �*�*ء�m��   	-ēY/f�� l��k�� �>r#�`��K�a���	ݖ��	 �(��7f�'YI6�� �l�%���㭒��nM� ��1%�$�pH�F��ݶ� \�l5:w"��UNZ&;lmuT�F��:�Z^T�C�;J���F�t�l/bKl�����&�UUҽm�*�^D���V��kXh��A'��p� ���*E7e�vݱ�m��%;fCZ^��x(����mi@�@ 4Y��n���a�[x��`���h�[S�gK����{&� �AT�d(*��.�v%�J� @ -��m� ��m�    8 �  �!�H ��$�UmR�*�HM�W*ʙ�	 @ j��      8mm�� �[pd�	�R�*��T��ή�V�{ݼ���{���EAS��!��U���<G����*˵W�P4�]*@��ǂp��M`���Tآ:�P4
���؁��� O �ϐ�B
���iW�`����T�xuE�t u|��S�a`VU�%�``����M���*z*a�@F"b�U]*�
�
D�>��� Ц�U�Q�P��=U}F T��m��`(	Z`%`�JU�fR$$�dQ�$����R�a�b�|EQN�ҩ��EWk�|
ȃ
���`#�W�⨾���] �ABD��R` � P:����'�(|	�FH.*����+��T<=�@_�`�tm p��N( �UN����2J!"Bl� /��QQ]���(z�ޟ�����k��q!Q(�t�-�1�[V�3�Qu���Č��u��I[=�nnxx6�j�ބᬣմ�0�����c�M=3��)-v�UX�k�n]�w4�j���j���V�R�)�m�Y��Aր۶"Ɲ}�q%Ӷ�N(��	��)�^���@M+�[`6��@���pt����%�N�9M��^�9�,g���!���Ѷ���D��Ais��Bq�in�Ϸ��v�S��[�����Z�7��ئ)70p�nn�����c�Rw&�l1��(2KK�ٳ��ycb��h�^���N
,Z���D�n���&5t�r�b�v��l Qi��f�S�+��@98:}:�-�ש]�E��po:�F<e�m��:��I�r\[��:n����s��Ɨ�62kQ�tƬ����K��{:|��ɵ���U<�f�-�F��&��5�']��������r�[��bdk;22�Vؗ9��۰q��`�\csW. �U�.���$Okjy���H�;�Ȕ=я<o]n.�j�*۵U�� �.�Qm�E�mfYx{Z��ۮ���S;�թϸ�ˎ�V��e��y�$[U�3F$^�৐�d����7�{G#�ۺ�Q�M�I�dAD��1!Ʒj�iֳL��B���3n���=9�x�5�'e�C��h�"�py3׳� \�.�_< �C�-�mU�a�u�eɓ9%�*�"@�m�ݻkff��m���0Is�oS�]%���
/�p���/lr*�m��U��p�T�E@ H 6��n�f�Y�v��#*d�Κ4���N�j֧݅k��/g�$x��<[��r��ֲ�m��'[����b��W[���9��N�\�k���Dj{.�ӗk�j2e!^3�3I�m����	��{S	%�˯,EK�����-ӣ�[�Ź����3��CrX�f8[۲�]]�1s�mUg=�[eڬ�����V��̜3-*�����ʸ�2�H�"��M*�z��������oՆ,`SU����3��s4��3�*�����©�����ݭ���p쓄��ͦ��+�T�T��nY2]s��)���pm���A�pga�������њ�6{B�uh;3�P����dL�'�Jn�b� �1��et�B�%':H��6�9��ۤ2UtW���a^.��)]����Uuv��v.���N��y�{���=����ș1 l0���L���c�`w�ʎU˰�����p'Ɔ%��}���|��� 7��ov��,X��zo� �vȼ����R�9,� ��ן�bI�����=�|��׀]���s���\�����0^Հo^Հ�{�Tq�898�H��`�� ޽� -�0�`�q������`����f }v��j�;_�IX�v�y�3ŕ5�^�ZZd�;]C��k;�n���lA6q���8	��(ڑ��� ���j�5wk�/j�a�_#Ӆ��o[�*����6=T!VTXA� ��E$A_@ >J�UU>t��`yl��$ٌ�,�1
N9!��j�5wk�v� ���b���&� ��G��^ [�`�l�-{V{��^O�g8�n?�=��]� ��X��x���Z�ƚG�a8��z��;���3H뗬d�Q��7���v$S������ >�fkڰ]��ݳ /u"�i�&�8��)&kڰ]��ݳ >�f��D�@��am%��u�ݜ ���FfJ��0��j��y�U�u�s�|�o���\Q�#�v� ���j�5wk�;v�C(�"�L ���׵`]��
�׀�����\�DD��ع�[�eJ�v�wr��ٱ�p��7g$�b��H)&kڰ��xWk��l�6�q��k�	(�q`�ڰ
��u�J=�v<��;�}�┥'w�=��qR�K�,�3f/?o�1)J=�v<��;�}�┥'��س�b�ovDݲ'j���9��J=�v<��;�}�┥'��wC�J�M"$�#)*������: (x����\R�@�����N8�r�m�g��w_w8�)I�����R��w��R��^��JR��������yo4cru��꧗nT�n�ԏ*�`'Z6.�w8����t�r��l�v�Z���1/��by)Jw;�u�)JO/��%)N�w_3f Y������,��d�Ŝ��;���┥�w�JR�w_w8�)I�����R��ﻜ�Toz7�0�v���R�>}��y)J}�}�┥'��wC�JR�w|R������GV\h�v՜3f-�w_1)JOo���߾���)C�۵g��~6�V���m�,���������y)@~P'?w���JR������)ߵ���(S��#%pJ��!!&l�R�&`���0	LA����{�۷I�QY�$��X����̝�;�������i7�;+t]��lm�]���B8�z�;�����29��:/Wg7C<[-Z�n4+�Q��g���7��2l��ͦ�8�6�gk=+Ͳ��m�vh��8�O[���<c���õI�h5vu����L�;p���Q�u�]m��)��w79VrN�+;����Z֛n an(\�Z���s1�kk�J�A�l�c�!��q����mu���u�:�s�T�Z��>3f#��~�ĥ(|����R��u���)=��Ŝ3f/���"v؜�&7-�b�(|����?�I���_�g�)>���JR�}�w�)J�쮺�T��X�ᘃ1ogu�1b^�}�%)K���┥�w�JFb�ݺ9(�]��U��f �A��ﻡ�)w�w|R�����c�J�[�����1��������zJR�}�w�)J>�v<��;���qJR��ﻡ�)wܞ���l���8��N�\�B<�M2��*֤��`�m��v!b3�S�{v*���>}��y)Jw�}�┥'��wC�JR����)I�ߵZ�l-f�n�f���)ߵ�s�`����TuA]���R��w�%)K��w�)J>�v<��;߳wM�Y����ff���y�)JOo����{��JR�ϻݏ%)N����R���~�5;���T�Z��?���`�?߽��JR������)�����)=;݋8f �G�{���b�R��ݷ����w�JP�Y��}��R����hy)J]����)=��5��8�d�.��M���:��A�nF����V֧DAM��-�c���f��A�%)N�_w8�)I�����R��߻�)JP��{��)�o�k[����+��e���3b��v,ཋ����~���JR������)����3f Y߻	��-Y,�g�߻�)JP��{���	�U>tnS]���R������y*��{���V�X�;l��1b�}��y)Jw����)JOo�������b����$ф-�h���c�JS����)JR{}�t<��.���R�>}��y)J}ڮ���@�F��fy4����x�Z���
�J�I�u·]N�mpj�>��e)=���JR�{�w�)J>�vg���;���3b��6���^
S[�j�oC�)w���┥�w�JR�w]�qJR��ﻡ�� �f/��ԉ�b����ܷ��3'�����)�u���)=���Jb;����3,ߵ�T��E\u�-Y�1�!b�]��b��n�,�)}߻�)Bp{B��	!��z*��s��ǒ���w}�Z�Y���m$���3b��v,ᘃ1����(|����R������)K{�_��	������b6����;�0�O�U1x���x�u�DZX�p�2�s�6����zJR����┥�w�JR�w]�qJR��ﻡ�)�~�5��"�m��f �@����g��	���~��R����hy)J�����1i�`I�Dv�4Z;h�R����s�R���}�%)K��y��1���՜3f-�wYl,rZ��-��1b_�Ŝ3f#���R�>}��y)J}�w��)JŻ�m�Ix+T����3�{�┥�w�JR���┥'�{�g���գ�l���(�u���qpb;�?\o��Iy�Շ�ql�N�qƸ5�{v2�ŷT��n�a����a5]�X�tP���2�s�́��y��mm�6�7v��qT�S��7^	�C��Զ�G�;������� �\n�Ӛ���v�KcNs��lem��cjn ��	ݡ�e۹�Muv�;F�:�pU��Zm^�c��{isY�wwv��(��'7W���ǆ�Y�y�����vXGvlG=�'+�nl͉]��=7�NڒKI�8Z*����A��f�����3��┥'��wC�JR�{��JPo�٪7*�Q�-Y�1bݝ�qJR��ﻡ�)w����)?��Vp�A����trev��l���┥'��wC�JR�{��Jń�������3�=����1t���F��K%�,ᘃ1����3
;��y)Jw��s�R��_}������7WB�k��f �D>w���R��������8�)I۽���)w����)K�k2��;��h� :՝��4ܺ�G5�6Ƹf�<��N��l�ΰ�-��N���{��v�����)JR}}�t<��.�������݋8f �]�n��X�4������)>���G��P�E	6�Cr�{�w�)JO.�b��3��|�A����[�~v^
�,prş�b�{���b������R��u���)>���JR��{�b,p�U5A�y��1/㻰y)Jw��s�R���}�%)Kwv�1b���j�ʥdE����JS��{�R������y)J]�{�)JRy}��y)J�������H.����f�'�M\�&m9�gr8���k4mTL=�6�U��P�������R�����)w����)I��{��)���)JP��_j�ef���,��p�A����ė�fb_]��C�JS��~��R������y)���2)S�k��f �A������R��u����|�g��Q�����<��"$#�Cf��{��)h#��080��{6*�`��I3�A�e�ع,�dV�+�3t>Xl��hbا�����1�Be5> �|6��4'�,#��&A�LE�0�̳@F�b;eM��u�4) |��*BpC����C�b�� ࢑��O�@pU4,��;�>���JR��}��JR���j�]�-f�j�ټ��<��;�w��)JO~��JR�{��R��_w�JR�����"�t�{ݷ��绀�v��ے��>�p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg�߿o��(J��J��(L���(J!(J��30J��(Os��h��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B~��߳��(J��J��(L���(J!(J��30J��(W�ř������VVU`�"�;
����4��$WU�] ć;l�9d&m3��l����og�P�%	B{�%	BP�$BP�%	Bf`�%	BP�	BP�%	�������(J��"��(J3�(J��J��(L���(J����8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP��o����(J��"��(J3�(J��J��(L���(J���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'���ս����������P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'��ߴpJ��(O3��e�J��J��(Mf	BP�%	�%	BP������<��(J!(J��30J��(H��(J���(J��;���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&~�����J��(H��(J���Z�(J��"��(J3�(J��?��_Ƴ5�[�E�[޷����%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bo��<�J��(H��(J���(J��"��(J3�(J����ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	��~��<��(J!(J��30J��(H��(J���(J��=�����P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	���~�Zw��k5��Z޳[�y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�{���(J��0J��(H��(J���(J��"��(J?~��~x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B{���G�(J��0J��(H��(J���(J��Cz@�Yq�@� |<��(J��?y��	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	{�ܿfVj7�{3z��[��%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�&~�����J��(J��(J3�(J��(J��30JBU	W�����h~����A�A�߾��@�@�{}�c~�b�r.K��%_7۲Vw�F��	��۳3�%��幘����mf������(J��(J��(L���(J��(J���(J��=����	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B~��߳��(J��(J��30J��(J��(J3�(J�����	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bg�߿o��(J��(J��30J��(J��(J3�b�/=��<�#-�Wl��BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B~��߳��(J��(J��30J��(J��(J3�(J�����	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bg�߿o��(J��(J��30J��(J��(J3�(J��;���%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	����v��$�MYl���b� XP�%	BP�&f	BP�%	BP�%	Bf`�%	BP�w���(J��<���(J��(J���(J��(J��(L�������%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP��~��(J��0J��(J��(J3�(J��(J��?~����P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B~���-�z�5�v�oy����(J��<���(J��(J���(J��(J��(L�������%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP��~��(J��0J��(J��(J3�(J��(J��?~����P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B}����(J��0J��(J��(J3�(J��@��,_Oo��X屪�����P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B^����J��(O3�(J��(J��30J��(J�����?�����x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'~���(J��0J��(J��(J3�(J��(J��3��߷�P�%	BP�%	BP��%	BP�%	BP�%	��P����1z'����(�W,��ph��������qm!D�]��q�ti���{@tX��<����2�]m�dq�WY-,��w2V�ue����:s��Mq�#p�m�N�p<�nv��ò��kI��tgnm�;�����m�wqX�my�<�ݧ"���98'�`*���q���qn�\l�-�q������'��8�o#sW&��.څ�w��=�uӾ�SrM�d��z�:�[\�	%Б�:�g���a�η'L4v�:��)����(J��0J��(H��(J���(J��"��(J��}��<��(J!(J��30J��(H��(J���(J��>�p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg�߿o��(J��J��(L���(J!(J��30J��(K�����P�%	By�%	BP�$BP�%	Bf`�%	BP�	B�b�/�}�L-�9,��-��(J��"��(J3�(J��J��(L���(J�~��(J��<���(J!(J��30J��(H��(JB��߿~ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP������P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	���~�<��L�@��a���XZ����ᘩK��߷�)J����R��u���);��c�JS����Z�ݼ�ef�����)J����R��u���);��c�JR�{��JR��j���(�Ul�g��vn�f �);��c�JR�{��JR��{����C���*bv\i�+�`�Yގ��t�,�2Qp��BF�NJ�I啴Ֆ����1-�ڳ�b�n��)JRv�{���JS��~��R�b�﫲��(�v�e�8f �F��� بNJRv�{��)�u���);��c�?,9)�~��ދ{�KTT���3b��Y�1bݛ���3�!$�^�z�ᘃ1��y��1-;��*u�K]�,ᘃ0�u���);�{��)w����8��݋8f �_��I��W%e�k{�)JRw��c�JR�{��JR�����{��┥'��3� ˶��٘�clާ3���,\ñ�nT�t���mfl�ZS.�a���7{������┥'o��%)N����)JN���y)J{߮�E�ym�7����)JRv����R��{��R�����ǒ�����┥'��消Ȩ"��8f �[�u������ǒ���� p�%.��w�)JOo��%)O����o{v)%m5e��f �A�{�Vp�A������);}��y)Jw��s�S�1n�k���(�v�e�8f �F�{�)JQ�E��~��)J~��߳�R�����y)J^|��k7���Z�m�닜.�g� ��˵�{�цٷc�]�3q���mD���T*����1b_݋9)Jw����)JO~�v<��.���A���uMP��Y�c�Ŝ�;�}�┥'�w�JR�{�w�)JOn��JR��}���oz�H�,rW���1w��g�����)JR{w���R��u�s�R�?|�V�����%Y�1b7{���)I���C�JS����)Be�}�ڳ�bŽ6�j
�4�v���JR{w���R��u���)>����R����|R�����3�Yoy�-��&45��U���a���ݖ^�^�O3ҎY-NqPEV�p�A��v��)JO��v<��.����)>7v,ᘃ1un�'-�)%m5e��)JR}�{��)w����)C�wj��3��|�A���v�X6卙��{��R����|R�����ǒ��{��8�)I���ǒ���{���,UPr�f �@��ݫ8)Jw��s�R��}��y)J]�{�f �A�㺶���Y�H�8f�{��8�)I���ǒ�����┥��v<��< 2���w�w�8æ�ĆWF��=>n�D�d�:�t��۝u��-gp�ao;��p�)㢊�h։�u�ps;7���t�n�)�o6F���v69Xuɖ�^-c��.뭵��	���]�V7f�������kK���ɥ�̹Nv7��{g.	�]i3���nM�̱����۾�m�yY�9��k�S�Xv�L�m�j�	<�/G�j����w��{��{t����G��u�q�c�9E6�`W�eJ3�'Z6��gs��Z��imN;b�Q�����1/{��8f�����JR����JR����3b��>���c��ᘉK�w�┥��v<��;���┥'��v<��;�wk5U�-p��5��R�?w���R����s�R��w���R���{�)JRv���Z���*��b��3�n��A��>�{��)w��|R����{�������N[$RJ1�+��b����g�	/�1�}����1i�z,ᘃ1ov����1w�֜P�T��nv�cv��:�#�9qqƻ�����\�믱%�'8Y`۔U;\�՟�b�{��o�R��]�t<��;�wہ�TFc3b�{�g�����H�[�Cf�ֵ��JR�����@�@	"BxJ�|��S�})��7ۊR�����ǒ��߻��O�$�bZo�W	*u�*�7lY�1R����)JR}��c��#%/������1i�z,ᘃ1wj�]��-VK]��b����g�����R��]�t<��;�wۊR���եA&;(ձ�Vp�A����┥������)J~�����)J��j��3ߙ��4�JX�7QЅ��r�v�s�9�f��`�#>8�.�;/���
�L��y��1.�݋8f"S���qJR���ݏ%)K��w�1-;��h�i�A[,Y�1'{����I�JN���%)K�z�1b]7�p�A��[�	�d�I[MY]�3f ���՜3f#w�x�?�� `�/����)��w��b�����nZ�R�,�g�J]����)>���y)Jw�o�b]�ڳ�b�ou�ʡU7Y��R��]�t<��;߷ۊR��w���R��߻�)JRy��c�޶stEA&B�^�m�J�n�-V/^��4&�8�%7��"鳪��٭7{�JS��}��)I�{ݏ%)K�����3b黱g��ﶭ����e��k���A��wv�ᘃ1���)JO���JR�����)JN���Ҡ�1�ږ;*��3�ݼR����{��)���R���wj��3���D�Ɲ��y��JO���JR�����)JO��v<���n�L�EІ	�-�.�.���|R��i�6��˅���ᘃ1n�x��JR}߻��)w�w|R����mY�1bݍ���aEbt��#�9�Fg�\�"jl���ت�ܘ��$k��v�5I�Xڲ�W3f ���՜3f+���┥���O�������Î �A���R��	k�ڳ�bK���┥���JR�����+1.�v�ᘃ1��D�lr�UU,���)J��v<��;߻ÊR��w���R��߻�)JR}}���jJ�u��H�8f �[��.f �@�}��y)J]����(}�{��f/��l-l��e-��U���1}�{��)w�w|R�����ǒ��{�xqJR�C��3,��s0�2##�'A�4FbA$x-<��lv� �L �(�$0�p�U8�FXRbc��"L�m&_�xL0LJ3	0Je�0I� ��t�PEpY��y��Ѥ7͇�IB =���8xf<p0@�F2<E��6�1Xh���B�8�8�`L!��A��N	�A#��O�R�K�	LBVICL	����֘
8</)��{��敆P����0�v���z�,���p,b5����Iq١�7"9�mt���cA�R߁�XHIHdvp9�¸����(�@��`�sz@�R�@�!+��2��(���{�;�;���	)m�9�5��O^��9m��Ŷ��L66���b����rlv�*v5�����KY)"C�a=6�[d�,�<��<J��@���\	��U\R�m
sM��U�,�q�]��f�ܘ3:�5S����Y�:ݪ�9�̫�a�!4�q�<iSl幦�6�+HXe� 9�E�I*�$��	�in�m�q)f�k��y��i�t��v�6{v�:��� 6�=\��p9���g�[��nk���=�5ѤtVW��첹�gY9��������/>1��<�x8��Pl��TѯH]�Z�����;r���S[E���<8�����v�3���x�{�ڇ1�Em/t��q�l�s�V�u[�4m��-�9��c]�l�ݗiҮ�sZ�`,��'b2�v.���?���\=����:�r�f��f�Zk"L�ll��7=�.�HYN��ӛe��ٳŗ�Ka#���t�z^�OY�[fv��Ɏ�p�]�hV�+^3#W)l*��e��"m�\�d�յmUn6�۝,�^i4������\Ӱm>M;p]��O$tP����,����i3��cX5��Ί]�'�Ɉr���,o=�U8�L��O&Dvx��X��iv6�Q������&錥ʯD�"ek&�լvf1�]��Zx\��0$�v�r ›%�fa@��7bYm��(N��{��|�A0���c2m�j�۶v�b��dE��$ʾ�j4�t�[k=۝h��l"�[U+�����~��F�F	���$ I��'J�^�n�FM�9�6K��U�®:n+�����a��;nsc�(��8e�2g5�Ҩ�39��[�Y.;n��	Wi]�����u�Zz6��c�ں�����h��vvu�4Q�Z�HKl��f�ڛ�m��61.,�Z�8�$N;T;���<�sm�YCF��[-�����V���˹�����;8v��xz���c�S:$p������dࢺC���������}����N�6r�k�ͣ�k���=d��JiJ�ժ��x�����n�\Ձp�*t�sN���]�h������6�5�<&�#�W#d�.e�	ny�C5l�qv�8K��
�G�Yݶ�d��n�d;%�u��u�����x���۶�1�4�N6ݷiUxr�;n�I�eΣm�q�����r^ܒ��ڌ];s(�7� fិ���(_w���
�T՜@q0�vؐ�ڷ\�J ^t���MUť�:gi�J�Dƭ�[b�3f#{��R�����ǒ��{�xp?�\��Zo�p�A���+y2+�;]��JR����G�+�b�����ÊR������JR�{�w�?f)I�����H��\-,�g����qs1%'��ђ�����)JP���곆b���v7�c��(++�s1�A�v���������o�R�?w�Vp�A��{�\�A������99�*��X���A��{}y��1���JR�����)JO���JR�~���1�b��/Sv�4���l&��l������-��]��ۑI�\�!�e����Iq�������ǒ��{�xqJR�뻱g�����f �A��wJ䒩sxo-n�o{JR�����<S�c�JO���%)K����JR������3B�f.�x�����b��K6qJR���ߴ<��.���R�?w���R��~�)JR}{g�m�"��Kb��3�ݼ�A��?w���R��~�)B~�N߿~��qb�|�A�며v�-�b�	���ǒ��{�xqJR��������b��h6>�l�����kuK"֘����Hm793�z�>����dd�I�̸JYj��3�w���1)>���y)J]����(~�{�ᘃ1u}ݍ���$

��\�A��>���y)J]����(~�{��)���S�9�P��w�oz�޵�d�Y%�,�3f#��~��A��gwv�$$=U��{�R����{p�A����q��+��-�b���JR�����)JO����1#3w�sw�V��i+�VJk7�����mG����R��~�8�(;��g��W���ld�T��Q�-֟,L�g���˜d��L�&�77J�ׂ��:K���Ikr�[ae\�A��M݋9)Jw�w�R�����ǒ��{�xs1b]>V��m�Il�Ŝ1)N���R�>����R��~�)JR}w���R��7��]7�2�լ���)C�{ݏ%)N���┥'�{�%)N���R���;���T)e�8f ����o�� ����r�����������%ZI,����/���Z8㈬VUyLRK`l��L`I��M������ukn��,�m8����6	��͇\k���6����4�ڏ�}����޾��ـ[�9�j�^�$����绳��f$�=���U�� [�`�ya�qEȇR<ݹ�V��ݳ 궼�b,��N%$���`�׀l����lt���mC��1(��< �l�:�� �ns ն�?~�9��QX�ƣ�BpQ�k�g:^�up�Ls:�U6�r��#	+՞�ګ�:�ܝ�\��n�W8	zyGkm��:����uf�mcs]���9�@��?�|=���5��7c�q��#��v�[g��nہ�v�i���R�%�K�.��9oi�]���u�a���C�!���0����똣��xn��*���@aӪ�N-�n�ڬ��>T�2����q��~�m�m�F�[6W�׭۝Y¾��26f�q�]v�H�.؝������]�آk@�}-�&�L[%��9Π>�}��Y�z'1����p��=�31&ʯ��޾��l�7����	�7���s�����f v�0v�0��`H��s9ƒN?�=����ݹ���]���_����!����f�z��|^�� [ݼ ]�j�땨�'+�WFxf�Ц��C�6��FЉ�M�#m�~�}w֖��B!��'�{���U���g�@_{� ��{�q	8�MH�#��5[m�9U\H$ٌ�L`I���UUW"�^x���E��� {�� 6ی	$t��$��YW@J3,HWe� �������:��8Ė7�{׀y�=��H&��K-���\V�lI1�zI�@�jڥt����n+X�.�+��U
ݴ���"L�B��#�x�8����R�&^#t�w�o����~�I��L`I#�T�0Ň�.���rY��{ן�6�z�{���{k�;v�y8�܇"�����ـI#�g9UUuw�Ill��ݹSNA�pjI�[�9�n�V [��<�$�}�^����m�[q�e07nD�$�����c�������v�-��1�׫\�UQ��z�@8��<�@����fl�[\�[�.�e���$ٌi%�&w�$M�������$�tS�8^��9&$�]���$���4�[�v�ԒJl�]�_^ҭ/�JO����=}���Kwo���J�I/���J������G#��LI%���}�I%vɉ$���癙ꂻ�>U�w�zo�����;�(F�?9Ƒ;ԒK��bI%��}�Ic�i$�uýI/���s�W�s۷b��z��*^�m�i��.��	�c��gz6�ɞ=3s�՞W��Xkvyت������yޤ�6:ƒKw\;ԒJl�i$��*�' �?D85$��.��Ē[����J�I/���H�U:�q'��&��&$��ܧ�$�Wl�������z}�I��LI%���S��|c�n^aޤ�SfcI$�$��$���4�[����.�q��A�
E�I/��ޤ�6:ƒKw\;ԒJl�i$���B_�/�d�qD�v<uXX3��F#��Q<i�a��Y�S�&�NI���u1cY��G�Eq��Vuu�v����[d9���GU�g9��ۣ������A�����^n�ƻk"����yXՙ�+�6B�V�H�8˦��h�	79��ȋآ��%�֥Z�;6�n|�k��ݦx㤧�bh��-�tI�+����k�?�m{hF7 �Vy�W3�vK�yec6ء8&x����s1�f�_��#���4�[��ޤ�SfcI$����$�,Md�ho����s�I]ܧ�$�Wl��I^�>�$��91$��uXEF�8���;ԒK��bI%{l��&�X�IM��$�Ket�w�X,�ƒIOI��Ic�i$��z�I]�bI/�ZE�MO�q�rO�I"�u�$��p�RI)�1��S�gz�_�Ibۢ�?�rҲ[RVGBڞB�(�ƭlչ囲����8ܒ�EA�ہ���(��'�$�nx��J�I+�g�$�v�&$����S��|$jD��n���������t�ș������I#�cI%7\;Ԓ&�*Fai.)q�� 7�fwe0���
��Z\��q��9� 7�fwe0����ـn�VA���#�ɀ^�V�^ ]�0{���5��&�#�18�B��A��u�9?���ݢ��m��F�|5�(�����mC����V�^b��}��ݘ�7�3�\������8S�"E�I%�����v��l�*� �]�<����q�;����{��_۳�[���%1L�����!��|�,m�&�D�Ac��@��:W�m�Z@��,(RS��Y�"\��� YX�)#%sА]����%���0e�@&� ��i=3B`�D��X�ڑ�H���d�S�WJ��ȏ�
�"�l |ESSJ�����!�� P��t|y�UW����W\]~�6L`�+P)'86Idr`v׀|�׀v� ��]򜟛�Jr4�Mŀ|�׀v� ���`v��ʛ:s��vƜ\�A�x�,��ݙ2��t�D\��5��;<�Ӈ������?m�ݘ�7�1�=r&T�l�)iT|MN)�D��ݳ �������ـn�VA���b�q�0�)�|�� /v� ��0�uX'��g�iI!�^�� ^����F�;��u};�t-rK�P���1��v[z�&T���Ҳ�~ݲ7D<�/![��u�wn�˖�ҭ���qjAm9^���ڰ�	x����m�7e�'�b`uI-�Ol�آ��pi��jG�^�� �[^ ^����
�+�r~lS�m���>V׀�f��^z�����i.)q�~�^��U�� �{V�^U�.V���I� ��������_O��Ol���j�$��"W!_�w�k�͑ts��3�d7fݧ�d����H�cf���W�u����I�kwr֥��$1�ـ�j�)�{Z�۞�ۂ���ձ�M����"ާ�Bk��ڮ#����}[<���X3��.u���ѣ��`����G`�.{cG��g��=S�v(=�/1��c-��MUC����v(�֑�Ʈ�L�z-qz�\���Ꞇ�d
W������`����㵣Zw�t�u%��b�@%��m��C#�k��D����$�Ǡz���>Wk��f��^��V��d��9�E�^�x{l�5wk�.�� �:��S�&����#��f��^we0����аMN&�8�9&��-�=�T�l{f0��@��$�q�we0����ـjݯ �u�:F���`��'�g��&҉��n<7	e�,��q֭����l!��X���ݳ ջ^kڰG���RR(�����_�%�w3�b\�� ��|���^V�V�(��r~$�ɀjݯ ��X���� ���i7.I��+������\��׀uv����L��&�_��y��1��v[-��j%�
}���=��`��[pnc�'cp�r�>�B�Gkݟnu�'9nۍI�2D۟�|@� z�� ջ^V�����+B�58��S�r`�k�*�^� �l�Ҷ�)�R�H�
�׀|��,P��*�00�B��8��o ������$ZQ6ۏ �[^ [l�5n׀Umx���9x�k�p�G [l�5n�`E�[�Il�!ir�U�jnŴ����X�nj{C9#�ћ�d關��WL�j����pI���x[k�>Wk���wW�A1'$�ǀU���mxvـj�׀jݮ&��2g�9NG�^�xvـjݯ �mx�o$\m��> Y��&Ɍ[��l��k�U�°`,@�'�n��ކ��S��X�G&�v��k�>V׀m�m���� P�47nۖ�O;4V�LT2���<�u���볚�WeK�
ʚ�Ɯx[k�:�� .�0[k�m�����2H��mǀu[^ ]��K`E�[B�U�T��-%D�8�� ն��`V׀U�U���0��H��5m� �mxU���f�������$n<���+k���V�x�8)$�*/wӶk�E��,m�Yn�u���\/1Ӓ�А�g��͋�v���S�v}ayW��`��5�;c����N�F7a1p��Z��㮎[&r��̏#sٛb���+�r�Wl����I�z�0E�i��[�;��v.��]9���@���s�pI,�]�5�x�P����)v娢b���؎ݎC��+��-��1��n��i����������;q��(F1�g׳[&��j�7cn\�=g�C�MvјTu%��!�a����?9Ȓr:��� ]�`�k�*�^���5����) ]�?�ʮs�I��>Sסּ�$�T�0Nq��98�)&�v����+k�������JA��HƜxRK`yI-�I&05l��*Ca��l8䋑��xU����V��
�� �:���6�PHm(�f�⳼s�"��t�.p:]��ޘy%��[��y�NFGđ"�< �ـj�^U�?���{Ӏy�?F��B���-����UU�\�9˲,�l)%�	$��$[R'�bbn\�9&�?y`Vׇ������}�ݲ'?�r�%U�-��{?~�8�o� ;����I��|��wȖ:U#l��1���U)>�:�\�0<���+�S�~tN����I��v-��+�zkI�t�c���])�b��W<�;���o�7"ƶm�'��Lݔ�>V׀�����nT�V�ݷ�o{t�g������^ w���,I����2㨅�$���?{Ӏ���Y�~��1fbY������o��Qu@V1���8�17��׀���7�����=�N����E
�4[e���v�?s���O�@��נּI�A�H���z��v����&�SN��e{K��8zr����պ!kg���~C}�8p�!�-X=�|�����f n���G,_�yyE]m�g�?{ӟ��_�IH���`���U�^���58�&�) ^�0wl�߹�/+|��{� �]�n"D7&�������*����r�3��ZS�%e�bY���������lz��S�e���_{��y,K��z {���{ݾ�~����&3��L��]Du=�#��2�<v�:�Li�y���7A��2][e��nl0˻W���[ ��������Py��p�T �L-vY��v��K?fbĤ{߯ ���Ӏ=ݜ����_8�I� 7v����y$�17���8��׀w�l�\�4��Kx�b�����>~�� 7�����b�I����{�[%��o,�WZRG�^�� ^�0wl�*ݯ �x�~Ăi��0q8�������3��&;�/��P�{��ZOP�, �mG�}�Gh ��*�$2Г�=a�t��S�Y�xN�eL,D�WM(p_8�6#	���� �&Y�	HK��	P'��.��CH� �4���"BH_$OX@v��/��v���a	���v��^k4� �t�F0����%ƒx�d���h8YmU[e`���˱u�Μ(Ԏ:5k��h���3X���O�8�!�"�7]UU�P���˱l�*�Du�v���W�:3*KUWq�U\K���EUW 2�(�V�������*��k/ 4������.�Lm����X�t3�zu�Q�YX�j9����r�� &�6��Yv�{ U)��pm����f=v%V���y.xwbkW<1t�y��gbN3ç�%��=�v�:�wOldnn!-3�*Ŷ�y2F��U�^�U�B�vQ�I���
���7>1���>,M��kv8뭃e솞3���ԽG�!�M�2��70�[G`�-�3�o!�6Mcv�Ɲљ942q��6��glv��9����Ӹ�6�l<�kd��q�5�Y�:�����-�k��nR�tH��#]�4)��Z�y��T�!��ʐv��ם1�#���g�k�����Qd����ԏ;p�g�mX�ڞ�H�4c9�Qeu������C�iѭ�s������<�l�ӊ�OA�p�Q۫�r�M9�'���ҬR97!K�����ٲ\.՗-�S�<쪝���E��%Ҥ��n����Ƕ�͙;;�M����A��@��A:���5Z����gO؇>w��9x���=<��۴��ᴒ�c�=�{6u�px�<�����ؔ��Ȏ�F�չM�k,9��)�e� �{U���*�ڡ����:�$wQ�YJ�:�cvڶ�1�@�u�rK�d׮�a���+�Nx	Mvs&��Prޞ�˱&��,�t��� Q����GU�Θ䖪��Ht��K[W%���t��,��MO+C�Am)L�܅���nnJ�m�l�ٸ��r���d'm�`x�L;�cf���[�S��D%0�-���j6 �;O��)E�0� ���� ���sڸ����n9���oi.6�`��r/[V�\%�И��KR&馳u�]�m�	�onZ�fjޣVi��
�x�� �4���>��p������v����8���sŲv�ѹ��PH{Z#�t츠��0�AP�|vaT��ֳ���c�esק��e�ն:ݸ*�q�x�y�;��&���0�M)X�K�ɓn����nx��x�U:�u���sI�t<n4l���n8�y(p��I�vۓ��b[Ӷjr��0S�4]95�.���k�z�M�`{<�J�i��:��ܔ��s�J7&ר݆���N�؋���א=��s+�ڞ��� 3���L�zf痛����w��L�'��k��
G��� 7v�����KI0��ޜ��'�9Tq�(��nL ��0�l�>V׀���bK1&�t���7+$eq�n z�� �[^ ]�`�ـ.�-!c�[���ē�{ޜ �w׀�v�<�f7�� ��j�����H�� /m���`ݳ �]���Ŭm�v(�U����/d�KY�vK�s9z���/Oi�߻���Jx��񋄑�> ��`�ـ|�� /v�wR%���5���q�0��w�l#�T�_��3��5ʯ߿~� 7v��~H7}�����<�BrO�����`�1��RD��`l���q��H�h� /v� ��0�l�����y�}�'���Qɀ�f�=���y��ـv���a�t%C�9�i��:8\�16-�e�yR��g�i�egleۦ��{e�:���$�?����X}��`���?/ɥ��C��� �ـ�fU��o×��|A"�� owo ;���1E�b���1!���ҥ��k��*�;k�*7���r�>!p�G& n�[%�:���&Ɍ�HQ՗V�R�Dq�0
�׀{�����ޘ�ݼt4u���ܥ�B�V"ؑ�zA2�^�4����k��ٛy�����+S��g��҉)#����� [l�ݳ ���wU�Q��E�) [l�����~�� �{�9�3����Ԟ�����5��m��*��=����ޯ������� �؝�H��Q)1���RK`I�r�W
��9I�b��� ��|����{�ӎk#"N6�x����f n��ݜً3��k�ҹ$%q�R�z��p�K]g�sX�KN��VGN�!��d�۵��igEU��k���{޼ �{��k�ـ|�� ������qpRH��ݘ���s������������`vcwRU�񦸧nL�������[��L�#$�8���98��?������ 7v���}���(�ࢋ�h� .�0wl���w��^g{�r�_�P�U�O����[�ÀA��R�;8��OO%�v�\%������v�^���n�<s����K�=fOM�y�7=Y��l�Z��-���b��͟@�1uF���x��
r3����	��9�C뇈�wQ���5�9�����ڧ��nǷkbŘ۴@�,ЇZ�]�b:8�"g��bz�Zf��ǍHRf齕m�m�n+�ko*t�n�(n4!����{����/��%�r�L]�X}q�۰���F��Զo]z�57���r&�Qj"9:m��*�^��vyf0=���{��Q���eu�o ׻���&ϟ���{޼ �{���X���8ږ�,�Y�>~�� [l��ߒ7k�Umx��M*�U|V��ܪ�%$��7g���H��k�*7���r�4 $�I����Ē^����~�� 7wo ;�6?;/�ۭ�k�:��'qCt<�U���ⶓΆ,9��t@4l�]����5��8�wg 7������f$��{߿^�������y���vY�_��ǉbl7����v�}����1f)??/��b.0v� ~�߯ ;���5n׀u[^�l�NA5�#���~K3I�~�x��~�绳��ۀ}lVE�%�Ҏ(�� ��x�Y��������� �wo �{����b��r�m1�F�Hqٽrm���i��v��U� Xy�V�s[Ǆ9��)O�o��������{�}��0���pl~q�^VKL%vY����{�x��������,X���fd��~^��_�c�-�������8}��b_�����l�7u(�`��\�Dr[x�I'����~�� 7{���$��x��
�E��u�,������s�_}>΀I����l��D�_���w���wC�1���i�K�p���礞;N�6I�2s��]qK���M������=x����{��,_�:��N�}I�\�q�R:�-�{�y�X�6y�8_����v�ؖf/�1Hw���[�N&ڎ(�� �W���V׀v� �wo 4>���jҢY���I�{ޜ ��׀���%��-ĒWy��p�J��Y,U���g 7���{=�z���zp��� .�6='�L�f·.&�Ӛ$=40ѣ��jjn�/<�mt=�
Kg�<u���j���o��ـUv�������o�0jS�0\i�F"8�[��V׀�o ;����bX�%�C}���t�r����"JG�_�����ه����H�ޘ�� ����\$`��bI�w}x��^����~�����zp���r��YH�,���������,�wߧ�k�����ݼ�%��yo�_֐��u�8��M��tjE�]�o��0v������z�Den���ݸ��u�C<5�O�E�rgW�g�x�Ų��"ZkJ���
*cH��Z��ո�<������lBV�>����c-�����2ɽltwb"maM2;kMXx��lc9����^S�5�ܞӷ)��A�(ʮ�GjxB0�d
�hf��p��3�N�{��yq�Ɛrj܏�9���֛���i��yx�r���s̍{Y��έ«/%y��>���[ �ٟ���+��z����NY��m�绳��%��a�� 7}��5�ݜ��Y���#���"�;-�����vL`E���[#kU���Pfb���&0"ݖ��[���R^��ZyF$4�'Q�$�*��`yI-�MٌvL`z"�%����x���Nz�˘'�κ���� ��t�%G�f$�9����r���eN�f_������'�c ݓ{e�5��[h�.0v� o����Ŋ	#	C�
 � !�W��{�U�m��>Vן���Ď����܂5m� ��� ��vp��,I��{Ӏ�0��|!�6�j$��*ݯ ������x�b��$�I�~�x�=���',�ʋd������?f,�����}�U�^���./2)�(Nml�Ǜ�eU�,�.����l8qy�r�#l]%_�bK�H�.+%����l�������v[�Il�Z�p���[]�����K6y��p^�� ^�0�+m$4��qɾU����{��u���Ua�t���:�V!Hs�t�LFL�4`i'��8<Պ!�Dt��9�t�1 �$j��B�2Y��D�j�ĵ	�i0�B <D�z�:A؀z���X��%�պ��Ϲx��o �wg+W��.s��:ݖ�I'�����w޸��`n׀j7U�A"rh������_�ff%=�~���ߧ �{�8�ըZ���"��yH�����3�Z���L��X��n��)]�l�[��58�j"90wl�*ݯ �[_�bY����}��>�Y�R5i����`E�-��$�7f0ݘ��s��`����М�RTY$�p�����f n�]��^:4p��r>H�m�f$�~����x��g�W�� q0QNk��5ʻ��ŭ2�\	#r`�ـU�^� ��o ��a��&��0��4)r5g(���[�ezV�$@vӳ���^�i�?�{���?|�I5�rN������:�� .���&0;6[�Y�xSn���,�����zs�ēa��^ n�׀k�vp����	�BR, ��`��&���N�Oy���U���YH�%���Iff7��^��zp�n��I$߷}x����UX�r��r��M��?fb�����۾� �wo �$��\�e$�:�ƫlU��q��Ó=��v:ٓ�ƻ,Fh��m�.��m�);��Ⱥj�#$窚���9кsl6N�����ն���;'Z�YW��tr�����q�;v�`7sܺ���r��ܧ0�wa�[����6�":�]��Fۍ���tP:ܧ(�M�j�W$`����gX=����ocf�
�������Y�p�;:��{�ݔ��m)i��\v���Y�>zi&8�MʆK��4nX�+w�f.*�\lRXՕ7mr���~��wl��fz�Xk*h������H�� 7m��j�;f���Ė~I%���ȓ�ԍ��ۘ�>���`Ir&�Ș�cv�ײF�刍�e���Ė?z�πw��Xnـ��m�"�蹙�DN�%�w��|�fbI������^kڰ��p�s��p䓉��Hc�e�'Auv�ù�í��N�<�s��˘���N@m	H��ـ���ڰ�j�>����!��Qɀ��|��]#���~U[�~��3�}�^���f��� q�.9"�90�������1fcg��� ��� 9yw�q�D�"�'"�;]� .�� w����Ř��o��|���/*��Q$��, �l�?������z�y`�Հ�"�$ꏌ'D�q��nh{+�e��d�^k/Ds���ջ[M�!v_n(�|@I� 7m��j�;]��,���`{}��7Q��I��u�snD��� �����Us�H�ϭ�Y��Tۤ:X��@�����&��NUW$Ɍ	�05�e�f$�T$cv�噘��� 7}��7�p?ؓﯼ���'��ђ�#��1�nɌ	�`z\��Mٌ��fw�OO�I
�)[VFP��%����g����i�9�n��[��!OU�_�w{����nm������_��`�Հv� ݶ`�U�7G9�I����Kn��w޼~ۧ?%��=��1畖Y�����^ w�������_�����z�0O]p`[�y�vL`O\���r&�9��UAH�2���U�k����]�v��A�+v[x�7_ ��������`� ��'x�R~���nn�aۉr����k��{"��f�͎�]f*sÛ�Y*̲����I����'���0	�1�owo�ĳ�%��?~|��R[ke��b`vc ݓ�"`z\����=��G ۘ8�% ��� �Ӥ�{� 7�f�؝�ps�8Ӓ(�� �{V�mx{�`{�V�� <y��7�E�hN,�����x��o ��vp$�$��b]��ѿ?��C�
A�N�q�Fy�����Q��ld^���g.�r� 7f�'۬���曑�ꮋ4��ٺ�8\[SF,]���ˋ��� ����Qqs�`�k�p� vj��n�I�H�9{B���tn�;Nꁱ�kH�xݍ�E��6����ݷ�Ŭ�a�>�'*�6�*׳����skjK�K痊���Ge��:�g-ؤq�i(�{}���w� �T��3�u�gv���x���л��n����|u6v�����ǜVT�\n�l�w޼ �ٌ���RK`E�(��J,Ui�90wl�*�׀|�� .��fcf�6��A�X
:��>�с�$�~�9U�q#�>�$���i���x���ݖ��)����N ~��� n�]���ښ�����#�ݳ 7m�]�������߭�� �۫�fi���[���=�3*=v���!qb��ե��m�}����~�k ��qI��z`wk�:�׀�f�lVF�9��i�IɀUݯ5}��{31Zk������� ����;���L�QN7r<�mx{�`vـUݯ ��E�~��&�m�%���%��33$���x����wg ��^WU��㊨��	"r`v��?,I/�K��~��߿N o��������/��F��Fz2$�0u+�Km$M�<X^���S�Km��GiĮ��%� ��^ն� ��0�l�?��9,�s�8����:�ޜ���&��}0o�0
�����MH�D�q��p~�� }���X���Hav� g_�P�������_g���`]��D�Rp�qI��fWv��mx{�`v��k��	ƭ�V�_���?b�K�b���ߧ���� wm�U֓U��P�bH��Wm���x8��rm*Hp���[�<��=En��q�'8�r<�mx{�`�ݾ�K?�}�|�g��<��Vێ��L^�l�&0;/b`{nD�W8�f��"L�F��� ��׀v^��ܪ�%���0"���=�n	K��NH���Xuڰ]��<4� ��W{����*���k���g?�3��Yq|��, ��ݶ0;/b`OTK(D�c��"��̫_`K�a7fV 8s�����:��p�qtI�7m��R�'Bh���m��� ����bI/���>��ʹi�	��s�L`v^���܉�o�c��U\����^��p��IJI�w��`�j�5wk�� (wh��'9*%$��?�$�>��� ׻����x�ŉc���|�g��/+%�c��"�5n׀�f�v���X6��I�z�&�r
>��'B7i�	���b�<��7i�i86�W�PRk�膑9��r�8z`^
f ��=�����
_�x$��'�a�C��ґ��b�z4ˀ��p��=�ޝ��z��Ȱ��\ڙ�i3 ���9.];�;�۸似׷A���䝆��EmΓ�m�P�Q6����Bj���x^Vv`\��e��
�.L��uB�v��:�.�"q�ʪ�
U�g�а�ԕ���;]��������=���J^.ᤶF1���Kl���Rz8����qmZmm��
�E��e��h݂�L�a���㍂#�`�st������ݹ�]qÜ�gx�-N0m��Ż]����W�s�e���<�T
���)�Hm�����i*�+�S�2v8؋��;��ϲGEۑ��,�m�������vH70�^�M��0��kg�nJ�:K�'m�mCE
��v��ݳY|p�c�9ۗl��1��ѶD������9ه��;�ђ�.�]���������-�%��L���"zY]P�-1(u)�kc�'�jRW�m�G;Ur[k�u�ͦe�m��e��h�����Kk+\���#gp:���:⫴��U�����8��%�A��v�q��ݗa�9.n�r;j�FfQQ�n�]��Dh� �:ι��\�M���Wm�vpvx�@�t��[ngL��wU�������v���k�^uu���%����gon�#t��s�K�!Rð��um�٢���f5�Ň;kd;.S��0��:^���0�C064�[�fȬ[k]�m2��r:�AI���l�!]Ȼfs�L۵�RΥ�4��l��ݬ�^�p�
���l���v�5��H�bIe����W*����랆l���n�y2���ޠ� �b��s6��7[���S����Mz1��� ���cm��_iZ]tA�5�fo���:m��q����l�9�n�g�cr���T��n:����ӣF��bCm����6I�J))�a���z��,rWk�i`F���pp�=�]�3��vn\1��P9������@Umđn�z��`�N��������{��{�w�}v�$}<�:hTU��f���Do4C��wa��wi���ʻ���툃�¶9�ε�����6Ż̝u�;��3�fy���9���:q��<\�sƸ�6pq�:;9��n�[�wѮx�5��7]55���tqn�N�*N�g�Cf�6q�����\\D�9Cch�pU����;�dc���+f�E�Ĝ=/�O[���R#�k��rK8��á2ufv����{6�g!k��Tvz3�M�;1�`��[T����(����
K�}�h�6��g ;���?�n��f���bĳ3�~���7��m�r1:�E�[x�͉��V���UU�U${~��\���I��!dm�����`�k�� ��V���Ӎ�NH�h����,I����w޼�f���$�Ķ�y`�7�D�Rp�s����l�>�Հw]� ջ^ s묰�=�����5���n�˪K�\ⓕ�X��"��%��ww���}~6�[Z? ���Ɂ�V���9]@l��`��@ԲU*-$���7_bI4jݖ�=�c��O�*�����K�T���n2!5�`[��f�v���X����«�n< �Ɍˑ0=�"a�s���'���4��K�@�I� ��V�v�V�����~
���۳-�pbcvs���h�ܑ�b^�[�85֒����Ē|��$Rƿ֮.1��+��?��jݯ ;���>A�?y`|���rB	4D��5n׀�f�v��f���f%��n�<���c��˽r�����U�u��- zJ�
4�,�1�=�P�>�<�u� �mx�eR6p����RL��LmȘ�e��\�9�ܪ�]Ͽ~� ~��h�J�E����f���k�� ��V޾!pԫ���{1�t���^��U�G�<񞓷�7P��l(��j�K9H�.+%���Z��׻��l����[�d�^R��
*�Dq���l�*� ��^V�g=�gt5�y�4ZZYo �ﾶW�[?s�|����}��(����Ĝ�g�G�um��*ݯ �wk�}������Ie�7�N��_�,��Ti��<����v��ڰ�v� uj�l�D��IcTC�V\����2��ўv8+oc���R�s7̷CI$�9��x�v�����v�~��+}8���)*vDՅ��x��g?؛>}�N���?�{��K1%�H�~���Ql���:��Ӏk�vp���7���p>�Ӏw�t��U���q��x[��.�x]��.�x���L�di�Y,�����X�zwޟ�|���_{��LIfb�ff!bHI%�X�M������TQbm��9�.�p��6X������N���g��C���gS�����m�nN6��F�W^�8//:��u���G/@e@��޺�p5v�q�qlgcg��8xո�یu��=��Q8�SQ�������ls'U�#z��pYT�f�,[�.8�^a�v�6�nc�Հ環��1���a;=Rѷ���N�2l��mZǷ$n�e����ezI�v�����ڞK�M���ё��«e��}��>]��
�k�>]���[��7�Ng3�F���:���n׀|���v��噉6u��~V�8\��,��y���>]��
�k�>[���bw�9�F	�'#�>V׀U�^��v`n׀}�,q�q�%5N<z�L�ۘ��v[�Il-�m ����/i�js�.K�Ҏ�YU�-ˡ��*��,Y���͞����#G�un��[��RK`E�-��/I�5Y,����x��g"_ر&ƭ� �mx�uـU�x7�*r!�"8�x����j�>[�����
�55D$��<����ۘ��v[�Il����V���:t�����<������&0*� ���i��䟜`�q�̑��gB�d��p���k1���k�7<�t�Ըdr1�QɀU�^��ڰ�� ����ND܍�"I0����j�>[�� ��`v�ȸ��vD�u�8�7_ �}��¨�b���ܘ��x����Hq�㑧"�>[�� ��`+k�/]� ޵����n8�MG#� .�����j�>׮� ޣ�BQ�.�+�7R�e�MŜF��=uӋn��F�ۂ�a�m%8��(A&��#r`+k�/]� �^���ـT^jj�8� ~'$q��՝�Gu��ݳ �n��$�bM������ī���Y�����Ol�T�l���QjS
G*e�cvY���1�I�}�����|�����+��%OdQ�P�fQaHBG�! ʣ"b�* lХ���W}�y��֤M$���x�ڰ��_ 7�����է��Z9)D�8n5v��bs��5�-�[��;	:�u`ť)�_��O���4J��5alv߀��ߟ ��]x{�`W�`/M���㐜���"�;�X{�`W�`�k�%��٭�yY,������c��&��Ln�����Qwĩ�I� ��� �{V����y%�߻������
)Q�R��ױ0=�� �ٌ�ؘ���\=�Fv�8�sŲvT8-���[E�Dst.\L9��[�%�ꓗ�ֶy�η&˶�H�^z�Ķ��Z���H�7Q�=GY�p,cuEq�4���>K����v.�����}�<r�Pm�K!��n��<��c��u���y�C��l�s��c:�r�5G"�T�a��S̛�g��$,p�It�{d��JO��&�8.�{ϻ�ӷ&|0���l֎��2r[e���;?q���}��47�ֵ,<��B�9ȏ��3�!E#�@�����o ����30�f������Z�TT�M���l�>�j�/^Հwv:�݉�F�Mp��$� ��� ߧu���X�ffd��Y�������m�ĸ9�#"$� �{V����ݳ ��� )ռ��!�!99#R��>�l��?,X�bY�?o�_����π^�� �u.NW�H��)#S�������H6W�����w�ά��m�U�ˇ���qĒjGX{�`W�`�j�;�X]W�>|�lI� �����{!�RX�_P�m>�&,��}9��7��π����I$٬���
)Q�V�8�}��>��k��\�G�}�)>�|H���^:bF+���9���;���}���l�+�>�z�qr'���q`ݳ �n׀U�^޽u��ӕ�2�]+3O/a��9�O]j^ْQ�GF��[�]��FU���Đ�\�Z�-B%d���� ����z���f�v5H�������Wmxz�׀{��>�g<�bl��d�PjYiUV�-���=8���w3s�I�.�1e�F�d����(r��J`&�%%�����p�*	�"����$bÀF!��F&
82ilɅ�-o�w2�2��̰#ı�1�fİ#�Bpc ��ė'�q0Jg�0	İ��7�7,l����8{�EK>�,9����<H��ݛѳ=w�<Cݐ�e�[����<�K�D᠌ a�{[��K\I%&%f�ذ>�_sZl�L@�9�����[,l �d�9�5lHC
��f.Ǌ����)4&�B!)�jA�`	�	�� ����b@c!�b1�d)Dʒ�eRE�,:F!�A�����f���'4�:880���Bv�g�=�$0h�h��zY$��666��Z�1�XLd�;���`����6��F�̲�_�6��(�
x����� k��@�C�S���׀]v���O�9xێ$�Q8�����^uڰ=�s�[��> {�R@^��@��o �}���r&�{r��1���s��%
���߸�7;]b����Ř<���x��%��wE��R�٧[�����<ݽ�������� ��ٳ����~ĳ�~���7O��Rrq����$q����L ݶ`-���j�>�z�qr'��]�c ݓ[������߯�V���;�k�����P��%��b�X��������?�6�<,JbΧM���>��A��#�N(���]� ��+��>����~����l	-KJ�Eظ�^v��n3�v8��f��p���vvrf5�ͨ%�q��k�>�g��� �l�>[��]� ��j�J��K-��v��bl���pW�,�������9_���9&�ݯ ��Xz�׀m�����`��Um���O�}��;ٳ� .�0��xz[�NN�s9��q|�� �s������u[�]v�*�V�~E �"$�O0��&�Q{�f���ݢ�`��rj��<F�9�E��^Ǝ�e"9�:5��n,����7���j�u���t\v��]����8�Y.L��I�n��3`�v-Yr�g���xe5Ӥ7D�y&�4v�9�?��rw�\���ʾ�s�R�
�[���� 2b3\�{����SAr*�렀^v�6d�tZ��Wf|����K�-�+��n�Ŝ�Ij���X����&YD�C�gvS{6:pr���ۮ��k�`m�NQ��-%��h�rt�}0��x������ յ�`����DHP� �n׀]v����������nph�S�	���Հ|��0�9ďo�x�=����6(5l�EU��S�m�`d��ȘnD��(T�USq�,�����Y��y|��� ��u�h��H��c�:C���c��ۉay�i&Yګ�9�躌�F�f�A.W��̕D	�䷀o�u��n�Tۘ�&���V�PAWW�p��������b��7���/�����[�^�V��ⓓ��9��E������g� ;����������>��������J�ev�g��']�x��,��X˵ـovWRG98589�v���X˶m�}�� /��im�V���R;�c�6�gk�e�.B�;b㤘�.2��WP~��������\N6�q||��}�]x_{��$��a�����잊[%�U�����ٳ�ŋ1$ٯwӀog������ٙ����d�)$�����	>��2��U�T��Ș�ٯ��S��b�Q��m�~ǽ���7��X�u׀j�^Qy�� �u<([_ �f���f}������Nߦ���bK;�������@�x������fo.�2��k��*ݥ(MT
:�В)99��̇$q��6����wl�7�Հ^�Vk�bnp9$���� .����~H���{_���� ��dB�H���9��x�ڰ�j�>뮼�����/ Rq��ڜ��?ى/ؖO��ߟ �����]�~�[Q�R��$BU!�qcB���M�w�ܪ���k�5a�����9�]u������}<`�j�>��.T+�\H�����uo`��*��-���l��{dnc�u�&Ԗ�V�{�ݏ�?��q��������[|���/^Հ}�]x{x�G+�'~p����L�z�&}r�"��`DJ��1�����0׵`.�fߒ��bR~{�Ӏ{_� ���j���8���/��?<��x��`�j�-z��'�$m$�x]��٘����=پ|��g �%R�0Y����[�m(�u�BVJ��9oe%ɓn5��08�)L��r�h�l�@e�n;N1����䔯n�K���m;��YǓ��r�dCj�������6q)�g�^����
�מ��x���I�8#{��W�����y�l6�V흜�7Y�ɥ��F/m���3�qӗ���!s�\c&�Ư����'A#2N�f��q��w�b2R�wq>�K&���:����Oٵ�\�UɄ��;k��ձۥcr�e�1UJ]��S��������/^Հ}�]x]�����"��Z������l���Ӏy���7�S ;u�g�"���9�\�l����`O^���R��ƛ��"�GWv�{e0���ݾ�� �|��^��J�x��`�j�>뮼��x��?]�v/cj��܏rYq�yi<�W����b�k��n��79����r%��uǵ�C �{V�]u�wk��]��wO{��T��9ƛ+�W�ݞ��ꙉ&ʶ���`�j�-z�cP��6�n<��x�ڰ��^�|��==8�۶��mRU	S���1%v{� ���|�]�[��u�P���8��j�>]������`[�F�uqȧ��r3��;\�=�9��5W�!����{L{cX������O�$ME�NE�[��U��z�]��*�@>�|a�ț��r(�r`�T~{� ��X��=ě��H����K%�ݞ����s�̐$�JT�ڪ�j�~�^�lD�V���̥�3z�L��1����_�������7���)��Nf$%�/���?L����`�Հw��4\֯�o5�-�/B'l�6%�]:K�:G��OGH��yz���1أuP������~��޻Vz�X˵ـ^��9�BT䳀w���g�{π|����*�^�]e O�5�8��Qŀ]����0"�-���V�jgZ�U�����X�����{�N���s���i��>�������m�C�^DۈDq���*�^�v����+�� ޣ�Bh�W^�ltC��ȉ���mZ�Ns�r]S5���GKJ��$%D�N�X#,�p�n��l��3�9�����`D}QZ�A�����$X[k�>W]�[k�/]� �6��9�i̋�8��������8~������|�}��7gbvEĤG$�4�r`m� ޻VV���k� ���DprqH�'��7�Հ]v�����*�^x�NSA$�)���!LI��6�!2Xbc��NBc%�P=�a�Y! ��BB��^3��C����fE����	��	&��m �-�!0Q�$� �!&��Ɇ��a�!` 1��f��2�	
��� ��	$��xȑ�$̚SX��`�O�qt��$BVe��eI�<L� ����&�]HP�w��{6o[�����ӏ%PmN��f#��w��ՍՍk�.���ܙْ�ŶnA�3շ[��k�H�Z`,!ٻile'\���neLK2�\�\�mj��
J���1�l�
m%�c����E�2�fz0�T���&iy��É6�f�^�9 �j��yL��V�v�l�Y�ڴ�N ��x�@M��52�,dn�8��B6a�]�
e���Bv^�՘Z0��Q��r,�S�t.⫭t���B�7nN���2�Nf��l��1ЅR�yx��2�qUVqӧl#<�"l3U>BG[����v�x�gFڛ�6wa�˻W9���R9P���*��F�X�k$	%nL뵋x�b5�,�ַb��vL�)mu����EM�/"p�\�v�zʬ	��:#nU�d��=�����Z����ͮ
���nqB�!vӻv��(v�\��C5��V؋X�6�8͐�n�n�@yw/:�u��O�{�+�y���y�s�����:��:�m����۶�4�l �TY�6��yYxWk�@����d�������tL�cV9��i�+�xN�9�쮔 �]���-����m���v���X۝q��hwTv02v�����b�7�+˝��#�G0v�]l�G,R'�<��mph�m��4�¹�L;Tpvv܆�\�[g1�� �+�r�Ge-nˤf�V��6g<S����rJ5gu��n�qnyN5nӵ�Q��3U����Vv�a�Q���ucJ�j܁أd�q��N��T�.&��Xƾ�7�*�����]d�j�朙M�p5[UUT��!^��L�VY�O(�4 s �P�d�+���،<�o/9�����N�6��q���vkƦ����a;61��d�y}v'���]�%�X���͛!���}����L(7�ɼ���� ].�ܱ��$������vf��6c��q̦�c<Ps$f�*
N���Ċ�[Um<�ݕ$� m�H܅�[;Fam�'�t�HB�|"(qz�"�/�ߐ���,SY�ڿ�ke�0���)Y�mۆDu9�������N����;\1�d�۝R��[9"��h���l��٭�bqv���wo�'�shGmA�Н]��m�l/A�c˘ݹ<�zA̎����x�ў�k��+��S�A�.,��o"�b�;&�Ӣ6d۶T���oJ�$9� d)����5ͲWl@F�KJ���!h��R�(�9	��w[�&.N�䵡����W<&y�B�tɫ��;]C������{����:]�4N''qP/�����v`m� ޻V�jj��$M1F�� �v�0�K`o�D��r'�*��H���]X/*䵶Ye������n���ē~��>�璘 ?�Q#�Kc�^e�7�"`M����0��s��/��Ӏy�Z���HT�m|{7_ ��/�}=���zp�7_ ހv��7FD�I�8d�6�RM���}�v]�R�RX�⃈����;6�]�#w�)��m�W��L����j�.�Vk��#M��[]m�o ��������Y���_�����y�l�>��ٷ��g���"I�'	D��x��,�ڰ��fV�x�z�nr&��rqY_��ğ�}��>~���5��8�6�Wjj�RG��`+��V���j�;]� ��\�VI�z�Ū.{;�a7f��=)�ΥpWd;g]>�Iu� y����,��o���~[z�Lˑ}ʪ�m�[ ����B����n<z�X�ڰ�� 7v���STA��8~ I�u��*��w]�,AN� `0�e�f�v���c���D��.���-���[ �}�07�"`M�׭�E���9Cn, �l�?߹�~�=����XݱՀn�Oʁ�$�4�Dr�Rvr�!�Y�\b�R���e)4śS��+o�Oњ�{R�k��~~�y`]� ��:�� �������NZ�����|���M�w�y��ޘ�ڰ�F�5$q�4�XݱՀm��ڰ�Հ}����u�h۲�e|$�7���
����9W~�{��E*J/��~�^, �h7�*q�p��NI�o]� �r&}2�`d�^��(*��w����.�B�N�� 7\u��H�ӣZ�M�2'Lt���qт�TaB���n��lu`�f�v���c��\���e�}�Y���&���^�����Հmz�d\i�AȢq`wv��7_fbě�Oy���<�~��Cp�𑋐� ޻V�ڰ�c� 6�0��(A�Ț����X�j�>펬 �l�7�Հq$f	guk6ȅb�89m���0����76oWa�\T+��q�;�.��*�&۫[Wō��s��&k��k���q�P9�A�ۗs��ՐJ1�6�u��M�U.��.�;�F�ְa�'�c�}�[�pK����/;���w��Z8p�u̸���ܱ9_;�쌎(z�8'��*�r(���3�#]�[ ��s���*�����C�����ڞ\^�����tHR=u�v�F�K��y���Y��\�l�ɭ2[#d��*nm����m��� m�`�j�6�V�]I��
6�"r8��5[^�v�k�`v�V��$�
�F��qBI��eȘ�ˉ��Il�Z��>NO�$X�Հ}�XV׀o]� �lU��4�DR8�����ݳ ޻Vkڰ�uKE���>'	�J��j��C	�у��
B]�,6�˞w[4��/D�Q���Bec�z�`�j�-{V�lu`��H���X�m��n�L_f%�]ŀw�:�ݳ �v��s��ܜ�ŀZ������v�z�X{�8Ԝ#���r,���`I��Ș.D��R��!X���#�G����`]� �v�0��k@Ҽr7���?I��A�[Q��l���:�5�٣GWL9.�	v,���GÇ$���j�6�V��v/���N�yk��De������j�>]��U���j�6��g�O9�$H��:��� �mx_����(z�)!#�O�S��I}��?��ݝ�����$��)`�r`�� ޻V�ڰ<���� �g��$��.N	ǀo]� ��X˵ـj�� ��F�� @����]4Q��r����G�7
Wkl�Ԭ\.�䌁Ɯ�b�����X�j�>]�� �l�7�Հ}ݹƤ�9�'�r,������z�X�j�>�O��$����r90m� �\����L�K���R�R�K �I0�`]� �v�0nF%*o0�����!�0��}���Uܽ>�gd�)��"$� ��X˵ـm��M��=�%�������5i	`1x�76�����^�6�k�	4�m5Є��Q��Ɯ�g�O9�$H㋠j���`�f�v�k�`^�^8�d�$nL �l�7�Հmv�����7�,��$�\��� ޻V��X˵ـv����_�9��������j�>]�� ۶`�j�;ݹƜ89$��s�Ȱ�k� 6�o ��u�����$�~BĳWt/�_G�:��p&�F���6���6�����U�Gg]�z��lϲ!�����mͰ39浍d��q�Ը�; �/3ۡ�-�mE����q��wݯ�Ƶ��j�Z��f��v�p[uƩ;J�v'H�i��X�2{X-��;�X��z�SS�cm���n���[hPޒ��\�,s�1�ZJnK1��U� ���蝼ޭ����gQ�	��jٙ��g�ɮ�y�OO�ո6h�d����l��rss�ͺ�4KbJ݈�=a.�L�_�m��l���L��0:�.c�J�J�%�90�`^Հ|�]��l�*/5��r~8DI��X˵ـv�z�Xї��s��[,��?b}��~� �{׀w��KIﯼ��k���IYIk�&����z�X�j�>]����nhlu�c`X!�RD'2�lI�zӡf��5��Sn:��)]���j�W/X\���u��{� �j� ;�� �l7#�HYTv�%|�7_*Y�S��W3�K��7vc}r&}��N�GNq���v`�f�v�k�`v�'�ʒbjrp�Ix�ـo]� ��X�u׀}i8�8��P R)$�7�Հmv������Q�B��NA�&�����sl����u��W�^-�Śժ����R����1
O�@�,k�`u�^ m�`�j�6��X1'�$�E����v�z�X׵`v'Q"n�H�q�ݳ ޾�9w�֌�,$)�� ��D0b,��o�"f10�� |͋�^�y!!�����R]$`�Fa+�J���<׺� *�!��� ���O�/5�z�P�����}Il�|���F�������ڜ���h�5�!��	�y�`l�A�1S��b�ۺS�{��3��  O4c�}J�� Hd�	F��$��IK�4'�|<��pc'P}ޅ6|%�����L�J�Y�bn/��>'��}�C1�$8A����k��H�1���F&��#��n(Y�� r��z���x ���Px

���'�$%t���@>U5�!�U��}��`�u��j�#�d�����X��o���o� ��l���v��k94�$�d��ŀmv������z�X˼4hu@�N7/��J�'g��n�Ψx.P�7S���f��ᎈ�rܭ�4�\�}������~�6�0�{���XwӉ������#�G����`]� ��g<�3g��Y?D�@��8��,k�`u�^���
��N�Ɣd�E�Z�����*�{�W����L��%�d1�I��ĸ�=��7�=�p��Ē#�E����Uv�z�X�j�;ڊ�'"��8q�ȑ���.F^��C�1s��'V�:�#<�Өm�[n��>ǀUmx�ڰ]� �^V�S��pN.%��8��`�� �^U���ֹ4�$�d��ŀZ����xWk�7�Հ}�s���r1�2F7�v�����j�-{V }����^1�rp��#�*�^�v�׵`W�� �B�U&R�_{��b�	buUl��u��4N#`.��;S�;0��%x�{��:�G��i$G��c=VQ5f#�ӪEI�9$�ND�賛�i�k����@:Z���=n����1ۃ]y&L��Yʝ��&e�y��-��5��.�ɶ�%]v��l�[gX��v�сS;��� �U�F��lI����폟��=<�g�K�#�eXj�&���c�v�S�;����n�M�U�t�$�n���۵k΋��K[0R[WM��a���C(�����:���X�j�:�׀UmxE�'R�� p"$� �ڰ���[^�v�hͼ����� �I�j���5����1$��{π{��|w�Ū�$	�NǀUmx�ڰ]� �^V�S��pR.�����b`Ir&��l���ݭ+,��rxK���wz��ʫ�w��fi5��nāE%=5!��&m:�X�m���~,��xV׀o]� �m�7'��#���I_ ��vsRX,HK��]���痙�<�*��w�ʻ�w��ռ\��2rN)r<�k�7�ՀZ�XU���ȆU�7���<z�X�Հu]� -�`D�K����$X�Հu]� -�`�j�- �R4�GѶ�(�"Y D��Bq�c��g��K(��t���\�E9�7��
9$]��< �ـo]� �ڰv'�7��E"|� -�`�j�-{V�v���S��pR.�����j�-{s��> |�A�D7�����V׀]6�j(�9� ��XU��
�׀o]� �m�7'��ڑ�#� �^U���`�� ���a"䌉���ELl�v�n͈�"�;��L�Xݐ���ԑ�Q�3�9�N1��)r<����j�-{V�v��C�*�
8��`�V�v��k�*.�:����"$� �ڰ���[^�v�i�^H���g(�|_�Ӏk���;��|��}�%�7yu�����O�q���}r&�"`yM���V��X�ʵ�y�vv:�Q����<�]��5δ؜h[i�Vmʤ%"�$pL��I0�`�V�v� �ـ]Gs�8�D��ŀZ�XU���f�v������n6�mH���:�׀���������|ޛ��5���jb#"N6�xnـo]� ��XU���"WȘ�R)$�7�D���&��lM��+�Ҫ��_���~A���-p���+�R�cG&�.#5Q��v\I��á�箞j�u�fV�sw����!�	�v�/,�2����`�T\s��ի��n�6��p���v}����pj�ų嫎ݰ#qj�m	������K)d���T�(a��f)�1�9� ��]n��Ż���"�D�:.qt��ĶY�F�+�s�3[Ӭ��k5f� uU����?$�o��v��bJ]�'9/@�:���+��y
��-����[.ɮ�n�$Z�����xnـo]� �X�$b�o3��I�j���v�z�X�j�-؟/$M��P�9,��v��7_ٙ���zo� �����S�#�d�	ɀo]� ��XU���f�:�6���r7k�`Wk�m��7_ ߣ�����y��dQsϴ����s9Ú�^����I��Gn*�^�+#jF7�v� �ـo]����=��, �����$��j$�jG��iCh84��ℰ�0�9#81�)B�2	��J"�88�B@b�*�EW+0����&�l�،��5H��R(��>Wk�-v�Wv� �ـT]u.4���rrGK�05{e�	6c�l��FԌ_��&q%�/��o� [l�>Se�$�e
�_
�Н+.��������䎎�=h�E������f����S�䉹Ȕ�i�� ���|�׀Z�X��xwj|$pL���3Se�$�W�[ �L`uMGs��F�x�Հj�ׁ����"�����o�y����]����7�4�cq`������v��j�>\�:!1D�C�� [l�>Wk�-v�Wv����1�8��"/fux���tC'vnk&�%胛��d(e�.؜�B&{d�8�(��>Wk�-v�Wv� �ـk7�s[Q�h��g ݛ���f$�V�< ���|�׀m6+����L�J)$_V�< �ـ|�׀[7_ ߻dZ�rJ�T��K8��I7�{׀|���vw_���Y�|�b��+���>
�C���� �]����&�l�&�`ݨ	J�Қ��ku�j�q@����.�����N�#Ԭ\.�f�nF������05{e�	6g�\�:�����7~ϋ��nH5$� �ݯ<�{�� ����-{V��Ir�!18�R6&�`uM����&�l��X�j�1 �Qɀ]� ��X��xnـU�x'R�IH������<�Y�{�� {}(;�o�AEE�AEE�QQ_��QQ\AEE�E��TW��TW����TVPTE������"���Ȋ*+��TW�E��TW��QQ_��AEE�E��TWB(���(����(+$�k>P�@�o�0
 ?��d��-'�_Nە@           4        ]<�� � P  � � P DE $�QJ 
! @U IJJ�� ��  ��  �h P   �a �ﲜo.S�ξ��n�����s����K/��t��էɧ}�}���ހG�)�޴�Ǽ �>��I�sJ` '| ��  �� ۟|�O{=*���zS���9:���z�g}�*�  � =P    
S ��S�}��-���=>h� 1� �:;  � PD fP )v@HM @��
DR�  v  &� 1 �&�  N��� hȠu�@ {  E   ��40 =PB ���	��^�о��m��z��\�n-ү�@yL��>�xzιi���|��< ��2��ﶧ�}�^^N���}�Q� ��ny:�y��魯�{ҷ���W�@  �
P
2 w�NZ��nMq=��^�Γ��R޷}eq���[���z�� ��W'�+�m{� O��*�4��x zS�Ϫ{��ګ���3��J�� �����k�NM=n,���} � P  *�6���}㻭/y�ׯ���^�OT�}���b���[�&�˾��� �yK}w�ϧ�^  y��5�ǰ;�}s�L��z�g^�ﳪ��t�� z=�S'vS�g^����n�zt� i�
xJ�  �������*� "x�T�(�$0�A���UI6�TOB B*�Jx�)P  !�)" ��>�����C��������s���{�����Cg������ ��������Q_�EEb*�
���!!���(cO��a]�0�1 Bq��!��]�������	����ٞq�fg9��K�LR������m������e<<�.��O�e'��T��<YO�P�?�W&�E��*�L���7��,Ϳ�[,V������	�D8������Cm��1eZ�yҒ�:��1��]��S5���_*�)�MIG�N*��M4İ�Hy����HI��uUT���I4��8g�G7$&� J�\%�͆Ɯ]�B��>���w���,��j������[̰�{&�7�p�ibo�R�|�L6SY��I\�l(�>�:�V�w�M��P�5�z}�߸A��"A#I`B�C�#R�0�$1!Fb�H$� c���!B��
F37��e����B�0���$���K���1w�%��"�!p׃I-�:��$Z�J��B�
�<F���d`ă2�s�t�c�j�d��ĈGV�LB!\$�ĩ�,h�.LIb��3��E=4�J<����k>�k����7���D!��b�!�xU���i�1��6��$=6C���g�HB\J0����a�a��B��Y
d)��J��@�X B���$
hAjĩ��("Xh)0����"Fy�Ea�bH�Xc#�P�8lnl�%1�q	L&am ��E�
�&��p#.fiu!z&$�(K��K�B�
��#X�XR���!B\��c`X2�lhB�5�q�l��"k
��,	
B�H0`K�J��xH��F6��=称�h�t���BX��f9�3B�/	w�s<�_wH\���$+�����q�9ay�/�&Gf�	tb&c/>�Ba.C!b@`�I�d�FI0��7j`[��c��<���M�9s[fi9�	̬�.���ܞ'�L���3�yr��˜8x�.	0�!Y��!
�y	�졁�v=����#d��'3<g�{���g��Ҝ<P���k)F6�K���]��7�#t��5�5�S7Hc�&�7p�i�(��E�e�e4�4���&4���0�`P�B�-�0��[�)�˚��8�!�!=!X���@�B4H	 �!"�B"��@�E	PC�$"DD ��A�~-!��C��i���F���$`@��*F ��6`BCB&H���>�hG�l�։ �0j����!X�!��
�E�
��	P ��b����ā� 1t-�ۻX��"0
�Gb��c�+��0.��8BC�o!S�9�T�r��I���4�D�X�)��<|H�0���,�#*bk�da\Xщ]���,GR\6%0�<cB4>����H�H,�HJa2Ȑa�B�3XHb¬*¤(��F�A���+	�J`�#��a�F㐴�L��RK<�y2ٯ3O��4���%�Hf�KRRIsX�хX�4�́!p�+�1��p`R"��V�*�"��!E�!X�F"D�H� D0 5b���##Q0,B����*h`�h`'=��x#�0i����.�J�qu\'�<��Ò�(D�Ʀ0�I�jJa���b
`�`h�hl�Ir$���<2}#
'�����6k�J�Jg4��@��x��&D�:��%2�(�e��X"%��tt�-�~�8z�Ĕ��἗NcC������=w����Lr!i��%�\琾p�+�
��M��ݧ��ݫ��7yI3�Ç���}�=C2 � K�&&T�##	V!\bP!F)R"�1aI�VR��%��M̌%#R!LaR4��P"141Hƞ����B�
g.�F�D!�t��F���� T|=��Ç�
*���C	�0<q
�<��S�,x� �x�i����@�i��3N{O) �Ot%�%0�8xz¸�=�����0bB�rx��t�^P��^x�,�%ą�9�\�,f�FD�j��!$@�bH�(��
����!aH�p'6?gٝ��C|��>�q����a9�X��u�Gè��+��'��QO3,:>C��5U���ڏ�޾���)���Dꢇ�����K슝	}�W>�B�B�܉�f>���-Z���Z��	U��{�wΙ�oy"��m�p�M ��n:�Ӥ�r�ԡƋ��Pr���鿥A1����N��G��R�wQ�:��1P��U�x�S�<���d����m*��j��jU��$:?}U�j��'G���!�2���<��� gߓ��V�X������i����GBK�қr� N���S���O�	}VU��T�9��Qy)���'�U�ۺ�}��y[�<�|&i�I<7�Ni�/���,c�a ��H��b�1J����Ǎ#@���	�hR(D�1!����m!B5�JBv���8�e4�
��x��aw��(B�<e���Ӂ�B��È�����0Zf�7�卥h\lۛ�����	L�p��HJ+s.����Z
�iCB2��X1�!B�q�\�@�XP�KJo<�&_9�U�H��ʇ	=��}���cM����9��A�$�X�愦e���}�^8��OO%�G�� a�K�w�.:@�9�@��%�F!�b��AŊ1 Q P5����e3^%|<~=H\u8��X%!�*JS�Sˬ. �HQ�"��ۛ�����y���'�B�d��2^C̣����&,������!Ji���D��h��|g�9��Y'�������%O=�"���(`B�>!��s5a	S���5�������@��B���O��bq4x��1��� F%1���)���#���@��j�`p#\tv�����8��ӈzx1�|}$MS>�-o���GOw�T��cw�N�"1`�!p�p�������) f��jĀ@�8��o�2��s<Jg<�NY�>>İ�^p�����i�]�#H]��;|��(B��dJ�!�����FS8>.o<Li��]�}H'�@�]����8ϼ���G����y�!|O^�y7�.M8���1`1��刄R˾��.�bT�x����y�.�� �
�5!sJ0(ЁN�
:`z1�7�Є�I����������y�<����B�)	rCFT�FD"5=K9�1��	��,@���rz�3��0�	��k��X��(�3~�3��pxIK=�0�6���$I0��BbA(�V��*�8;y�!qu
�P S)�&����Bn33�<H̞�z�Q����H�S��Ra��$��a�pk�#���
a�J�)2�u!pЫg��Oi��8g�1k�׌no
G�_s����&�)II��.lÒ8��
]��XI�}��y�==1>Rw8�a��JL�o��|���IM�o�,k��zsl��C6Z�X[��7\u"Cϼ�|�H�>�L6F�Ä�K�7>�5��;
�0��'��#Ha Fr4�4��	�)�*���)Ye#BH��X�`B%%2���(��b�bP�"4 �!d`r$���D�bB�B����!#N�Ir�!=��t��o%�Vej���%���(D0��U�� ��=!ӑ4�uH_L!�%�%0��rS� `�	L��b}j��P�,�W��Z�����[%��Ow�>��C\aL	p%ψ\%5��aC7��w�{6d9Ͻ��   p  �  \:�u]ۀ���	�\<(k��m�y�m�n�/��2/!OA��C';];�\�3�q�cN�"˞��0Qɒ�g���7K�T�==3rġY�۳9�O=�k���m��u¯=of�/���'C��/j]Џi(�+���7�����v�9 �;tk�tَ���IQC�0�֝�Ǔ3e�2;u�gdRŹn�8�����2�A��1<df_Z
{m+3�d$6K���s��(r<I�Ƽ���|��> ��p�t��)�pL=sT��k�j��K�!��L��9,�զ�qҜ���j�e����	�[�s��yJ�s��<r��B_!!��+�]�½U]��������˃b*��MƇ`�&�l6��:��Jlp�b��h�-�8�
��b]�9�nR�(��R�n@+���r(v�rm Z�x�n�["AǷ:��ϝ����nI�@m��ì�2��q�V�)�Í�b���5�v�^RUe�Z˰�۷1��@���ɤ{uu�r����I*RY��:����m����$��� H�� m�m��&� 'i7\�mڋk�q�h�$��m� "@H�$Ɛt��nm�|�m  	$��K�@Xnm���!��m  h-�$$�J��kh����� m� � 	��K$�A mH������� my3D�hܳ��p�K�v��[,�LEج� ��V�qdU��/��YM�Ӥ�ն�6̈́�   �d��k���^�\xڶU��-�m� �  p�m����N/[�\� ���  �`p�Mۀ�KonE��Wk�    M�I 	&����1������l vŴ8�K.s[4��	�$���6l�.�s�[A�� m�BKm��	7m�ٳ� m��i�1!О��M%�iu���6�m���:u��8M��m�m-��am�����	 �2 )[b[\6�   8�Im�-�m� � 񮳮t�$��� ��q��Um����T��� 8lRJ�� 8p8ɭ��$[@ m������m�t�l ms�6�&� ��>����` '@�:�e��z��mv�յ�� �M���mm�  ^��6ͷ�m&�v�� (-��$�Y0&�8���2��6���>-�8�H��@ ����F�   Ă��`�lH�����[I9�R���&� 8�` 	  ���8k���մ    �3JH �m�%�����j�V� [A  ��   l�  ��t�-�Imxݳl�  $$H plt����Hm � v� �ݰ�M���lH �-�
Q���;m����v �	6� �� ���u�|�zM�pE�m6�$[%�m�l�@86ͱ'v�-q�����8��N��m�     ����@ +jU�꺕eyU�%M $4[i,��  � l-�`   @����\p��m� ��h8k�    ����m�7k�m�n ���-�p	��$d$�����m��@$к���}���  H��"@Eԭ �`�������mն9�հm&�8�6́��Z�8v@#+UU�UKܺ�WX)}��� w/mX�9�{��g�ڴg*LR1�	�UH�� � $H[v�H�(��� [FA�l�#I�t�s��K
3Uj����m[n�fɍZ�\c1ڠ%E��u!ԭm�UR�eT�-�̓wBjڷf�!�I����J���,]<�L� ��Sj8A����G mW[[]��TlrG �U�]���po����mJ��VҭUplJ�[�U [�[v�[@ �,�-]���TuV��Y�@B��jڐ�+j
��6��mn� ڶ�j�m�Pv�vs��j�� �va6�� $��H�`��[���ād�ѵI�-m��t�i6:X7M�%��jړF����9��������΀/+�����iP�8"��I���A��$&�f��H�մ��ƴ��R�x��Vʮ�|���6n�ͷ8$H֊$p���m� ��U]L�5UT��K����-��� ����]UU*��]/,��E��@[@�>  ����8 �l  �m�WvU�W�UTP 8 I 8 �  �: �pp�F�뫪�*��g�� ���6�$  .�   v�&ǥ�p-����GH��6���z$�6�m;����N�q��l86�`m�A�W\�Ͷ�ki�i0  �m�m���n��ŋ�'[odm��tP�@�h� �_�����'mo_f�H�v�I���d�	  ����y�U
�*�TU@����Mf��Xl���m��I%�[l��l '@rIf�*۠lյ^Ck\t@,�瓪;"̀�n*�H��=m�V�V5 s�n�6*��PoavZc [J�嚀.��r޶X mm� ��u�߇_l����,�m�,3m͵�m�A�mm%����)rA m�$<�n�m���M�H�`���� �i3|�7�Aml��F�i��� 7M����i(p  	      �mm� �l  ����H �H�[\&��v��8�ﾻ�6�mm�C�f�HЃ�Ƚn�l��e�(���+��������-�lI��\��75��km�i ���  �� p  �	 �   ��   H $�P H6�����fڛU�6�ۨ�(U�I��d�jCv�m7j�;j��YI�÷nTʵ�S���u.m 6�M�-�-ikɷ0%��[�@� [��`[[l [@�>��m���  �8 H  ���  ����   $���	6�6��$i�$h���J��l�����m��:�N#�C����� �YID�2֮�-UUI��&�%��-� 6Z  �E(p6�wSU�;,���*���m��h6f���e��-�m9a�{a$�K(W T$r�Mv��,�	jր�j�~��9mɧM�A&��Y1>��6������� � i�z^vMM6�� ���J�a�Bs�V�ɴ9�����ۆ=Et�lH�P@���]�'K��J�m:��%V�mQM�����N��*��D�l��T0�I��  -�����۵����@pr�^�$$��hָ�[���&v�*�MK�pnνN	$�m�p�8m��3l�l��p$ �� �im��m�F�$�Wpl'R�	m�����ۖ�]�z�U	��R�p8  6������ĂM� pݢ�KM�[h 6�n� � m!m[%�`�͛b���l z�6������d�   N��  H�l�Ͷ9��tF�i�UvƸWlJ p �$��ݶ��m�u�h��3m�!mmt���P���7i4���@  m&m��H,@����n��Ԧ���` �ki���6�:6����6�@�۪�m l  m��.˳n�廭��  U�YY35*��ےNܲ�@P��j�	V�� ^�J�`0ք���� ��6�p�k� $�rUl٦˛n` �[�i;��6ݜ[V�[]"ޠӔ%���:�M���ۜ$�P��,j]%J�UT���D�V{m�)k$r;r\�n� b)m�*��|�V�*�V�N��r]V�u�cN�7�kp-��d�MU�f���O7+�*ʜ5mԪ*�r� ��B�`.�ej��p��ɵ�n�[I  ��w�c�M��$ 8�l ڴ�m�����2A"�Im i1�     H  �  Ć����	6�m���  pH�@m�-��kmm�D�m�@@H��m� m�e�I@p 6���l           d��\�h�	  -�m�ݭ�}��� -��ր n�pl�m�` $  H�����[c]& p pY��M�l�h6�m�-� m��   �   m�  ˪ș�E�[qҮ�5�iUX5  	   �    � Գ���w���@ [[l �8 � 6�  	 �m�ӿ������d��l:8^�vm˹fY��e�$o/-��QH
�����-�D��O"�����,�� �Dt@�@1�D4E��QJ��(���C�>t�C�y�����>"U�U}S��QHz�/�> �Uנ���߸
�z#�GE
�P�� _�D:q`�Pן"	���Tp)�8���Q}�MX
�S�:�<Ez ��g>���
��q���^ 0�d�@�"#�&�#0NTOD'���Qz����G�	���#�z <�Tx��SU�!��=Q8u����� �`
x �d"���$�A� ���` B#"!��P�'8�E= �]��O�����4�Q��>tQSS����z�5=�}�<�HH���I �1`�$����$%�-!��k!$e�$	-����/A��]���T��P�>G>AO�j��t�P������C��
a� DR
� �>�ݓs�Mkg][��m��nlp�87�hv�t�Y!�<-� ,]��юϬ;��[������)s��Y��=�13��ڌlrU���/(�4n��[ٶ:���x�u6���OG;��p�H�"�,tu�Q;�d��R�4M��hp��kf8&�a�X�A���j�5��qݸ� �<�S�3p'^6�:u�LY�q���\��荹��J�W+�5m�n{�e:��g3�n�9��NMs��j�5�6�٘���LfG�Q��q��T�W���jl��B�Ԣ�]UV�]kpH=��)�C����ꓳҪ�Ĥ��d��@ú�������V�P�(:�%��#MI!����3�l�,�Z�0c�ݔ��r��9s�5sw'FRy��n78ى�l9�mR��<'X��T�4�8-d{;��f5�Gi�z��h��R�ʯ(;g:Efv�R��xX]�q�4g��;8���8X���sL7M�Y��<�`s�$�(c�ԙe��iV���P9��XRy�&ֺ�]�5s�[�r���+�<�=�r��gj��.�岼��A���8��\v�P����ۋ\9֡���n1�����w)��Mnj�ȝ[
�*Ҭ 	ep!X,�RjӕWSl6"����V��R5��c*�7&Gp��b���4�j3�H\��@nYM%!��p\��gtl�J)�S8K�[wX.NKC�M���ݻSo5<[!��mųs�m�]`�P�牫��Zyr�D���#�E��7��F�L=�ɘ'�1��Ar�m�,WI�]�.u�»)�=�*l�T�2����ǐ�@Pl�*�3<���W](lek�c+�7&Y�::�ݻE�n��'�b��t6dx&TΞNeu�uz�ĝk*N�ے�mm�ђR�Ӥ��	wM&��ҭ������� B'�L��e��[zܲ[� 	�XyMـ���.�p/�%32L�m�na0��&��T���R
`�p3��p����DL�~Q#�(�H��l�M�3	�73dɥ�� �2��N��ۆ˅�P��IwW���V�F(�g��������S ԥ��5V��"�.z�ű����:Մ�w7:癸�5�7X{���tlHWn���������1"��,���˻V��Ȓ�f�X�}z����c4l-]���&{wS�o�ێ���t:E�x���,�Rul�����AP��"��G�'o��� �&3Ȼ���y��ySg��9��ʘ���lJ��R:�.7����}��?�I��K���h�>�xO2�����e �)mQ�1�1 �R���"�$F�3:q`���Ňr�3r�>�ؚ}M�8�9�YW� nL@:d��n�s!`n���wI:r�h�ܖ,;�������Ӌ ��-�pD�M�-kc�����[a�7كI�5�a�5qf�B�L�K��t峘����O�ܔ���% 	ɷUw,*����&n�I=�;�� \����0`�/C�x���P��9���b֛) ��H����m�2��Xgt�1aܬ�%���`n�yX�Kiu9HF�6���t�)z�ݿz���R nL@���sJJ)�P$Vc�Vc�V��,Xw+7�1��q���r��
v���'Nj$��k�pҧJ�[2�+�A9�B(�Dn+1�+ ��,;�������lM>��(DJ�GyH�1 �R���ܔ�Ϲ���^7t'NT�J�rX����w�C�el��V�L���7^�33f���ɦ�ҍF78��ܬΜXgt�1aܬ���� I�y�32�̂ nL@:d��n� �ӁsJB9C�h�U#;k��
	�iA��etZ�'�qv�
�Olu�[+��3�y� nL@:d��n�s!`��]N@R���$�1aܯ�I��̎�3:x��٠�>'�w����+1�+3���,Xw+����������z �ݚ��נ�L�.J�Y�B_�]���gy�גN�>ە�4�J%J�6���`bùX��X��Xr��Ji)(�NMآ[(���nB��Kv�K�^ ���3�hMtܡ:r�bU��Ňr�3r�3r���`n���W�F��R���ܔ���% 	�֛|�"@j*$���}��3;����`f>�`]M��%*�̽3&N���@c����n�w��;������m)%���`s&dٓ����@{�@l$2d���v�������t�dЌR�y��kt2�+��ˈ��`X�rôږ�[y�������N��9�Y:�bm6�b�)ۭ��q��n.]ٱ� s=����uv�L�GX{���g%��ݠؗ��Q�|JrsүKs�ֺ���u�As�;.Ԗ��{P�;(u��5r�vb��=\�ql��q���gh*�:��nSs�&x�]���˖�$�nM7K��P���|��#W�/l8X�f{B�]L8��4N1���q"��r��x�#Wi�Fٌ��;��R��@ɈL�����r	҄QQ8�Μ_��H7}�`j��Vc�V�4��t���WW� nL@:d��n�rq`f�æ�N�"�ܖ,;����H�A 7& 7v�]].fU�9w�����@7rR��@Ɉ��V����_S����E(�&�a�lb�7�WN�Z���$u���+�7�*+ � Ҏ�"��O��,Xw.fo�3#���(�����T��&J�O}�w�zA��N>�~���Te3 ;��R��@���f`9�FҒX��Vc�VgN,3�X�Ki.D� ���"��d�>d�=��� ]��of��f��9��AN+3���>V��3r�:�b��&ԌTF��競�ܴp��V�f���+qm�$Y#k�Ja"i�iҔH&�,3�X�% �) �� ����E�9��.�"f���u뙙2fw3#��Ξ,3�X��6��iԦ��.�u���(��K�L��4���@|�w+ ��i��$Q�$VgNrb�$�w% ��s��n��	I�Xgt�1aܬ�ܬΜX������N8���B9$�ך�hb����p�7���o2%��nY]]�3���RK���}����ŀfwK ��m%Ȓ�#��	���s ���%/s�}�UI��q�)B(�(�V溜 ��,;�������lM>��*r�"QD�w�4��ؠ.�u�"Rd�����X>�Ǡ���緒O���t�Ї�QTnKgs�=[��_���`b��`�\�:rH��*CڳQ-��da[�^wI*��LM9�m�ű6Ԩө)�Rq���X��X����;��uv�����tL��q��̙2gs;���Y��w+ ������4ĥBR�+w;���n�w% ��T��ܨ�F5#�1Vw;1�+3�c�V�R��BD���H����6gW��@[�݊�m泉�{ r�;�x�ϋ<c��i�%��W�O��|�q.萛����uF,��u����Y�yq�g��Sv�%�%0	����x��6��Dܑ�d�/J�I��Lcn$�I;�m�f��ݞ�v5��cwls��s\�a��̪�F;=�[�gQM��m<Vî��H��ԣ���M�$�vE!�N�`�4�8܈�9n(mu��獈��3��f�d�/��.����.f�6folT1��.�̺M�cgmQ<=(8�y�٪3���V�������'�?6߿�����J@:��ܔ��nU��]_9Q(�,�ܬU����}����Ł���M�%N�J�i�`b���ܔ�ndܔ��ڕwt��:���B����}����Ł������[���9��@�9AE`]��@y�I�Y������(��z6���~�f�w�N'$��E\V�s�-;�m�8�	t:�5��}����3�y������w%{�ϻA����=Z����ʉ�`�V*���z�D�
k���Pg�>�;y!���1�+ ��m�J!"M�U���n�s �n��9-�l\��J5J8�ΜX��X�;�����������'N���U�x �) �K@7rR��F���������=r�Z�L�㞲Z�ϋ6��Ú����F޽����A�-��]T��N/��[�;1�+3�c�V�M��$�R��8��ܯߒ7}<X��V,;��ug1���J	�L��{:Pq��j��3�Ld>���H�"����HF����@�G�H��@�,
I	����~�HIX�&6�c��e�� �L`B�*�1� D�}G�!��<i��{1��a �EQ�FP`F"\D��BpB4 Ea@�P��n鵖�>�3�7�X��QW�UQ���!�=RmANa�'� ת08�2�I%�㮮��;���Z�5J���2��(9��2{���Y��n��/(���('ӗ���"&G�22���ؠ96d�?�ft�@]����w���������\�f����Q�h�u�nͱp����AM��I2ISMRSm�����/��w�|��`I�R��@7rW���Uw��=Ǣ�rE$�	��VgN(��z�^�Pq���^�3�K�ǘ�:���D�`w?��`b��vc�VgN,�\:n�*u*T��nϐ��(��z�gJ
X�6�$�gffM̓%�͓��(��w=H��)�xV��@7rR�̂��@:���?���.Λ�����y6mUZ�c�$������Z�N�T���;��~T�GD�|��Ł�Ӌgs�3r�
���>�Q26�)93��9- ��H�A|�K32�r	ԁ$,�u�����+3�gN,�[B����F�R�#��[��Rw�� �� q�hf�L��$�	DQ8�ΜX�8�1Vw;1�+uUPWUu�j���j�?o��\;���<[
��$�Ru=��@{���=k�6����E�.��Z�-�Y���(��t8�f;cGIXڐ�V��:0��Y�6����TI�<;��g�F�ѻ��w���.z��1źR60 :!.LU3��g��k��.y�e�"�s��R�UX��5\�lwk�yМ��c����N�x;CW<�Kr��h������q����|?-sQE/)W3��R��+q��\_������R�I-�u��"-n�u�8k'NDF�wt�`bùX��X�8�7up黤�ԁ*(ۅ��f��q���Δ�Ξd��2L��`�`������<&�4���,ͼ|�����o�ׂ�A�A�A�A����8 ����ӂ�A�A�A�A�>��^>A����>��3?Y-�t�p��x ����ӂ�A�A�A�A����8 ��������lll~�~�|����?�g�M�72�������lll~��?N>A�����~�x ���߯ �`�`�`��߹�pA�666>�o�������tզT�:��3�vOA'm9��z�r������Z&��ś�$n�>A�����~�x ���߯ �`�`�`��߹�p ��� �`�`���s�pA�6667�����Y�C3r\�f���� � � � ����x ���Q������g �`�`�`����� �`�`�`��}?~�|����A��g�\�����7n�Y�nm���lll{��N>A����s����lA�A� �~ϧ�ׂ�A�A�A�A�w���� � � � �Ӽ�.~�pݓvI�36pA�666?}��� �`�`�`��}?~�|�����o�ׂ�A�A�A�A����8 �����焦l�7eۙ���A�A�A�A�>��^>A�������� � � � ���~�|�����~���� � � � ���������yh'��]��Ăg]�gX:�ٹ�����%��$���D.n����6� ���� �`�`�`��߹�pA�666?}��� �`�`�`��}?~�|�����g��왙�d��5�&��`�`�`�`���s�pA�666?}��� �`�`�`��}?~�|�����o�ׂ�A�A�A�A������i�&�]�\ݜ|�����~���� � � � ��O߯ �b(��Px��~QN���A�9����A�666?�w�� �`�`�`��çl��34ۆ䛻8 ��������lll~�~�|�����~���� � � � ���~�|���������[�L˲\�f���� � � � ����x �?�b�{���I�k$�3�����s�fe�Ԝ�n�e�������g���F��4��{)������K+eM���\`݊��\������nd�% �)�����	ԩRngN,Xw+1�+3��'t*p%H(��@:��ܔ�nd̂wW&�uu)IB�)������t※�҃IZa�MJ[)UlP��}J�'QE`}�8�3:q`bùX��Xf�W?�9Q��$�'٠:��p�L���1���r&k�VV#/J�Ix�*TL����!`ft��Ňr�3r�3:q`u*�ބp�n�	 �t�) ��H�A ��)TS/R��T6�&F�X��X�8�3:q`bùX���H䔤Q�їyH�A �� 3e ���n缬�b~�u*T�Dۅ��Ӌ�6R���s �s�_
��\���Dg��z�ݶn��	f:�r;]�6��[=����u��#,6�<8؋<)�=I=tG�����ݠ㓫�m�3)���ٝ�d�4n�v����v���	ZhM�n���#!Od�yC��Mi��i�6�v0*\qN�i7ZN�I�L��Яc'�zP���`�F�`'R�����#���hLcB��μ��ݛ�Z`|�5'0�rL�t�nm��˒����a�[�N��8��p�tN�g-!;����)���R
&�|��+1�+��Ł�ӋwW$��D��)I�@7rR�d̂��@��m�*T�DTTI��t����Ł��y���X�k���DȚ�(�����^�� �=h�J@u̅��6��G8F�0�*��`f>�`ft����ŀun�e8�RI�M��\��-��y�q2����S6�0�ir���d�g��۪~m������̂��@:���ʙ���|y����&"^���ҭ&LB`f�K(d$�\�9��@[�݊�7^��6&'�N�	 ��3�,�v{�[��Vo��t�M�t�9D��]]��t�Z���s �nd�rN��N�"�����}���:q`ft��ś���6����T܄Uv㞖��Ͱ�W���{���|Ʒ6�[\6��7R�cnR�IԤED�XgN,ΜX�yX��X�k�>�M�#*DL�@]��\�$�fF�����׳Ł�7N�$��a$,�ܬ'��{ySEX�
�����rI��<X`�#�J�q��*I���� �� �w% 5��2�32�"Q�Tn+3�gN,�ܬ�ܬ����&GDq4㍂u/]�nŬ���q��ڰ�8���␂���ϋ�哩@"m��7}<X��X��z�A�����;ɶ���(� �n�f�s;�����O�Εɝ�ռ&˨�:�!8����~�>ΜY�L�y(��O�v;�@�`��N�<)NK�f^��3�uq@ft�@]�k�Ze�x��I@ @@��"����?o�9���'O��BSn�ʒ�!`ft�����Kw�>u����:q`up>IrD8�T�&�����j�"[Iyj��y�g@m�qt�����R�$.���7Q���w�,���׳�&d�p���;�s�]ӼGI:�����}��U���#7�Ł����ŝ�����RFut^����
�"^���※�ҎI2g||�2;���͍���(��p��~���nuq@c�tPq���L�(���(���m���J%H(����7����UT�'����gJ2f��f�_���}�G�F
�1H?	�$Bq�"0��e����)0�=���@�#B�R��X���k8��*D��a�� !�B0 �`��@��	�@`�a+$�Ё�D�+G��!*@j���m%	R!d�`D�@�_��!>���_>$$c1"@"���0R0a		1b�H F	�9�b!� D
�	�)��B�,���!(�b��` �!1O�,�JF@�"��w�w�n>���}��[J��T�͓>�M��;7�F�J�H�m��<������$����`�9�^ĩ%�T[tm���������m��f��Dv�a���c[�<��(�s����Ș��MP'��eW�L�[mբl���a�9�p�4�ъ��S3݊�Rk&�=����0ݓU����d�yz`N�ci�I��!�#ƃ��nիó��0�I��"b]���Z�mF�����+��탩d��<�N��/G �.���nkC;�o=<[�'A۝#<�\�=�Z�Z��s���.�Z�B�g&5��i����>�^��jt�\1�U ��wku.�\�,���K��ؼ�k�B��)T�AUn�J�ٞ��V���f1�6"\j��OT�n���np㓘r&-��/���_2��n��q�&]�\m��]9��v�q��#F�4�����/�rsb�B�[3dVm�J���m��tb{gu�vK�$�$��GUҪ�R�5вnO6^��*U^�Uu����/�w]ɰ��ۮ�[gZ7-ȸ����I�]�e}P\�����r���:�4���d��m;G+۞�Vq��^��ú:�j�.s���Ѱ�L�Hr�m[P�9	l[4ɨ볧�C�,�ji"�e��	8j�V��ٌ���g'8l['Psldn�`(�M*�W�J�ìg|�O=���9��]��
Y��m;�/N� [W������[v1�.M��E��m�A;l0���M͌lu����[k��nG$��<�8��F@GL�JD��������m��r-\p$c�����yg�^U�X���L��[�#ɵ�9%`�*��` yk�cM�8�s�V����M9�l��ol�w��>|ۜf�r�E"me���j�z������Ƃ����I>��-�������ygf��l����ۊ�j��]�6�v�&^aΥ��e�m�ˮ��\�Y7f�ꢶ�jx�a[c"�gkdϻ��>��S�V����@O���`��<=�ɜ�wt���ɲ�y0�y��;R���K�k����,n5!�r��moE�v]<�uP ���c����q<@�+mE��m۫�!�n�@1.��ZlYsi�}�o�v'�uL�m���p�`nL^=<�d{�`�u�B�[�+V�҈���^�;U%� ����B��eXrp���KW�t[��ugۧawL�ےܹ��L0��pܐ�
���w�|����^�����S��듥���������ұ�P�^����������ΕB���$�����z��Ҁ��ӓ7ꯐ��`��~�I�2*$����t�I&N�gO��4�n�s&��#�:�K�!7J2��HX��,�6h��fJ#v=�3}>(Q�j��"��a$,=_�R[��`n�yXgN,=��n��X�\*�RR:M���ܔ���������و7�����֪�j1h˱�P���'�J�i랝�mg�����>﾿V3J[F����+3���=����VV�lO�N��@�F�3:qv�/�&d*O.̘�^�b��#5���z�2M�����BT���P��Ew�G3�dw=����f��WQ�p�!���=Kv{���~�3:qa�{��=[�&�N�JdTI������ml���)����⩸+�- �H�m��T��v��6�v�q��t9�b�?��w�>Q���Wk̮�����t�Z���w% 	F��$���FB�ś����#u�=y�@]��^L��f��~w��çy�OJ���v=�>��z5c2fI	����fv�� �ޚ�Pk�lĨy�x�LD����Fm{�@n�|P�l���~��{����$�@�F�ޘ���������rR���o���Z�VW`燋Ec�V�8��`q�.��<�q<�2�ɿ=Ͼ���5�G��> �������������A�����;�N��t�C�ܖc�W�ԑ��@ft�@{�\���:㓨QRE`n�yX�8��I��`n�yX�k�t�MҔ├����W�������Kı?g��Ȝ�bX�'��{x�D�,="���U\e�7g�yeC'8��Oh��I3!��7$����%�bX�g�܉Ȗ%�a���|���O�X�%�������bX�'����O"X�%��{�4�.���K�z��:!��ـ�#)f�i)�>!1v:D������d�ք�3;����K������<�bX����ND�,K�{���{"X�'s��"r%�bX��w����4˻nf�nf�'�,K��;۩�?�]��,N���Ӊ�Kı?g��Ȝ�bX�'��{x�D�eL�bt��ə�eɺM�6��۩Ȗ%�b}��~�O"X�%��}�Ȝ�c��Dȟ}��^'�,K��?~���bX�%����f]�3I��s6q<�bY� dN�nD�Kı>�~�O"X�%��w�S�,K� e��qL�8��N2�:xT�!f�vK�7r'"X�%����'�,K������yı,O���Ӊ�Kı/�gv�"X�%���}�a����0�:v��ºnk9c��WQ������͒��=�=�T�9��ք�C��2b�[��z1�U���̶qqr�in���Ӏ�FD�L
�Ǭ�3n�[s�lhv8]�I`���h��t9CG�|���	� �&-� 1�sv�	�͇�%�.��)�;b��nn\�b�+��c6���.Q#\vP�kT� �z!Z�=ǽ�ظk:n�ca�[�u+�'H`|�;esf�-��K�S,͙M����}ı,�]ND�,K�{��'�,KĿ}���"�}��,K������%�bX��'����ff�Lݺ��bX�'����O!� �r&D�/{���"X�%������yı,s�����eL�b_��g훚L�6�&��'�,KĽ�~ڜ�bX�'��{x�E8�(@�#���d�'fuqL�ı,K�/����+we�rn���K��@ȟ}�߯Ȗ%�`���]ND�,K�{��'�,K�"g{���"X�%�ߧy\�٦��s6Ss6�<�bX����ND�,K���{����}ı,K��mND�,K�w��O"X�%��f�ݚfᛰ�OP�c	�)vx����/�s�����2���nB�v�{��o��|�C�"���~�ŉbX���?�Ȗ%�b}�gr�"X�%�������Ȗ%��~�u9ı,Kӽ���w0�&�������%�bX�g�ܩ�C���� u�ND�7����<�bX�s���"X�%���gȟ�  ��lK��d��f�vK�3r�"X�%������yı,s����c�Pa�2'�~����%�bX����Ȗ%�b^��$�ҙr��nwoȖ%��FA�~���bX�'�~����%�bX�g�ܩȖ%����v'{����yı,O���]٦\�r��۩Ȗ%�b{�y���%�bX�g�ܩȖ%�b{�����Kİ}���r%�bX�{�����C.i�NU����t��6q=�k�M�tKO���-2f����/8M���ݓ3M�nI����%�bX����Ȗ%�b{�����Kİ}���~U�DȖ%��߹�q<�bX�%������·v[4��ʜ�bX�'��{x�C�ș��?~���bX�'�~����%�bX�g�ܩȟ���,O{'ye��tۻnf�nf�'�,K��?~���bX�'����O"X�DT�1Cʏ�����L���~ʜ�bX�'������%�bX��~���e��[A,^��oq���"}��?N'�,KĽ�~ڜ�bX�'��{x�D�,�����MND�,K�?~��̻�f�v�s6q<�bX�%�����Kı=�{���%�bX>�{59ı,O}�;8�D��oq������`E���c���ڰ�W4N�kNˠGsC��WX]t�i7d��n��Kı=�{���%�bX>�{59ı,O}�;8��2%�b^�?mND�,K�>��\�S.K��n��yı,{����bX�'����O"X�%�~�;�9ı,O}���<��)���Ŀ��7d˖�Cp��59ı,N���Ӊ�Kı/�gv�"X�%����'�,K���٩Ȗ%�bw$���76L�6�&��'�,KĿ}�ڜ�bX�'��{x�D�,K��f�"X�S`���p�<�������%�bX�����f���)�n���Kı=�{���%�bX>�{59ı,O}�;8�D�,K��wjr%�bX�����w����)s74���RK���veEj�2O��Iv���L�n�`&�JY�c�����{��7?~��S�,K�����Kı/�gv�"X�%����'�,K����\�l�]�׻���oq�{�y���%�bX�ﳻS�,K����oȖ%�`�����O��n&ı/����˗n�ٻ.\͜O"X�%��?g�T�Kı=�{���%�bX>�{u9ı,O}�;8�D�,K��s'�f�6Jnf�ND�,K�w��O"X�%��w�S�,K�����Kı/�gv�"X�%�z{ܒ�Je�.������%�bX>�{u9ı,O}�;8�D�,K��wjr%�bX�����yı�{�w��~��C�#b\\��6ɆA����ngV�彻�\�9��;n`���{v�u�붪3����ݥ�;aAT�Ô��WjW�δ�M�����{r���N��̳�i]��7��^�v���Ok�����ͤ��Y{"��.��ڙ��\5D�wv�������+���2����W@�ɱ��۬�/*#g�����ʛF��I����~{��O��Vl��/SЦz��Y�rk�	���D�W�Os�%b+rF��p�Ȓ�=�/w���d�>���8�D�,K��wjr%�bX�����ObdK��?~���bX�'����p�3M�nI����Kı>ϳ�S��G"dK�����ڙİ{���S�,K�����8�D7���{����X�s
��g{�o%�b{�����Kİ}��jr%����>��?N'�,K��w?eNoq������߿ ��f֖�K=��d�0�	���eC'8��Y�\Ryı,O���T�K��?�������<�bX�'����s�e�t۷m���S�,K�����Kİ�${���SȖ%�b}���x�D�,K��n�"X�%���.��[qٵ����IV;2����s^'�6�e�=�n��wU.��l��Մ[~{���D�,N�s�T�Kı/�����%�bX>�{t?�I�L�bX�}���Ȗ%�bw��-�8L�4ۥ�37*r%�bX��{��y��z��&��:�O"X=�?]ND�,K�����yı,K��ݩȟ�r�D�/���K��m�]w2]��'�3*dL�?o��S�*dLʙ﷝���L�� �
��Nr�~���S�*dLʙ3��ۼO"fTș�3���fn�n]̻0��u<�D̩�>�y�x�D̩�3*g�gv��Tș�2&g���ș�2�n����]O<��3*dK�}��O\���j������{��Q>߳�S�*dLʙ��߿~��{2�Ḍ���u<�D̩�>�y�x���)�w�Os�����Z�:nT�����f�I!5\�\��I�'vy���i��{��?9�����0���Ow��{��Sݑ3>��w��Lʙ2����O<��3*dO��v^�
�*%�'9S"fUt�z��;(D;(wN����$R��,���'�3*dL�>�{u<�D̩�>�y�x�D̩�3*}�gr��Tș�2&g���ȟ��(9�ș��������,=]�/w���w�O�����O"fTș�>߳�S�*d`xI�Q�$\3o���B1��R$@!�	!0��|ŉ�"���"$B"�"?
� �i\M@�EA!b�*D�H�$�`@�	F��r�_H����)��A�HA"@IL��f��0��.��u��0���O$g�� ��adX�gތ�� � �����I��#��p�� @���b�:�������@SDT�C�F�(��UG��p��ß��eO�f{�ۼO"fTș�o]O<���;���͝Z5a��w��-L���;����2&eL����ۼO"fTș�}���y�L��S"}���<��S"fT��r���s�.�vfnT�ʙ2�D�����y2�Ḑ�Hs���2&eL���?K��&eL��S��;�<�D̩�=ϝ���Rf �95�u�/k��J�p��礏�9=l��+l2���~s��~s����뻻�{2�Ḍ���u<�D̩�=�y�x�D̩�3*}�gr���߾�ș�2&gn�<��S"fT�����왐��E���=��)�w���|����Lʙ2���w*y�L��S"f{�wx�D̩�3(�����ʟ���S"S���p�3v\7I���<��S"fT��?eO<��3*dL�~��ș���iȜ������ʙ2�D�����O"fTș�=��[۷K�6�d�&��O<��3/������x�D̩�3(���]O<��3*dO~�v^'�3*d
VL�>߳�S�*dLʙ�k�>��t6M5|�~or��{�w���yS"fTȞ���O"fTș�>߳�S�*dLʙ3߻���&e�;ܧ�����~�lv�Tkl��D�v9k4��.}ZcVvM6�t��j5�ٷn�nf�O<��3*dO~�v^'�3*dLʟo�ܩ�2&eL������y2�Ḍ���S�*dLʙ:w���έ��������{��S����ڞyS"fTș����'�3*dL�>�{u<�D̩�=�y�x�D̩�ܧ����ߜ/,F^��w���w�2�D����y2�Ḍ�y٩�2&eL�������&eL��S>�;�<�D̩�3���nxa��M�ni�O"fT���7h����S�,K�������%�bX�ﳻS�,K��=����%�bX��>�37$�n�vR����Kı<�{���%�bX�ﳻS�,K��=����%�bX>�{59ı,
�@}ωtLw؎L�������n�a$nW۞�j6�w���'v��n2닋fz1��g�5� 9̧\H8��{M!�9ᴺ����k�3�������Mq������Mb#nz��..gY�q��ṳ���:�$
 ������;qե��.o9�,Ӳ��n��lӫ\m�]v3KŊ�����/+�<+���X�;��V���?0j3Q���6LB��*\�7I���i�Cmw1��c��n��L���Mݿ'bX�%�}����"X�%��{�s��Kİ}��jr%�bX�{���yı,Oa�����ݙrm&��ND�,K����Ȗ%�`�����Kı<�{���%�bX�ﳻS�,K���/r�n�6sfY����%�bX>�{59ı,O=���<�bX�%�����Kı=�~�q<�bX�'�K�%�칆��m73f�"X�%����'�,KĿ}�ڜ�bX�'����'�,K���٩Ȗ%�bw�{�fLٓM�7e�����Kı/�gv�"X�%��{�s��Kİ}��jr%�bX�{���yı,OfI߸�:jC���OS��q�mY���8��<���izub�˛���S�,Kľ}��Ȗ%�`�����Kı=�~��yı,K��ݩȖ%�b{��p��m�nSp���O"X�%��w�S��p t�bX�'����O"X�%�}�~ڜ�bX�%���x�D�,K�}�fnIl�2���ND�,K߷��'�,KĿ}�ڜ�bX�%���x�D�,K�����bX�%�O���sd��Jn�woȖ%�'�^��$�O>�w�H$���blD�O~߻x�D�,K�g�/viw7̛I��S�,Kľ}��Ȗ%�`���S�,K�������Kı/�gv���7���{����>�.Q�Cl��u����YI�L̑�NB��Mӱ֨��T���sM��4ۻ�O"X�%��{�ND�,K߷��'�,KĿ}�ڜ�bX�'����'�,K���v�ݙ�n̦�swS�,K����oȖ%�b_���ND�,K����Ȗ%�`���S�,K��N��̙�M7dݖff�'�,KĿ}�ڜ�bX�'����'�,bx�ʊx��*p�%���f�"X�%�߷��O"X�%���幓��3&i3�ݩȖ%�b{����yı,{����bX�'��{x�D�,K��wjr%�bX��}�.g�t۔��ws��Kİ}��jr%�bX�{���yı,K��ݩȖ%�b{����yı,O�ߦL�vn�3t&f��b1�:�-��[	�ͭ��*�k��Y�ڶZ�58��Z�~oq�������{x�D�,K��wjr%�bX��w8��2%�`��MND�,K��l��%�-7I����Kı/�gv�"X�%��{�s��Kİ}��jr%�bX�{���yı,Oa��٥�ܙ���]ݩȖ%�b{����yı,{����bX�'��{x�D�,K��wjr%�bX�t��}��WP���w���oq��Ϸf�"X�%����'�,KĿ}�ڜ�bX��I�lO��;�O7���{������ez�tt���"X�%����'�,KĿ}�ڜ�bX�'����'�,K���٩��7���{�>߻}z���y�]�]����I�㕍���բ]չ�פ�$T��9�i���vM6�����%�bX�ﳻS�,K��=����%�bX>�{4? �șı=�~�O"X�%������N0̙��73v�"X�%��{�s��?G"dK���jr%�bX����^'�,KĿ}�ڜ��*dK������n�rI����%�bX?~��S�,K�������Kı/�gv�"X�%�|���'�,K��M��#[Nl�ֽ�7���{���~�v�<�bX�%�����Kı/�w���%�bX>�{59ı,O0�wf��n��n�woȖ%�b_���ND�,K����Ȗ%�`�����Kı<�{���%�bX�0@'��Uh��Q1;|�Θ�����=���n�6�n�ȕ�Mۆ��qh����i�n�U��وܯ�1>�0 :�dKx�Q�6���%;v���
xA]s��]r��B��2�R6�m1�Q�sv��v8��0O,ri^���y��Ls����{n^��r*h9�(lnЇlАѭ�J�p�O7���[���k��)�m5�ap�B������A`�cSP�<��V�[FR�s��[	s����۬�䳒�c.���&E���|��{��7�����~x�%�bX>�{59ı,O=���<�bX�%�����Kı<�[;�w�v�nٷwx�D�,K��f�"X�%����oȖ%�b_���ND�,K��{�O"X�%�����s�30ݙM��l��Kı=�~��yı,K��ݩȖ%�b{����yı,{����bX�'zw�fd��i�&�nfm�yı,K��ݩȖ%�b{����yı,{����bX��2'�s����%�bX��O�nd�sɚK�s7jr%�bX��w8�D�,K��f�"X�%����'�,KĿ}�ڜ�bX�'s�����n
���+�buK�x(�'P�����剚�]��=�tvsw��Kİ}��jr%�bX���v�<�bX�%������"dKķ��L�8��N2��"&B%ȉ%\ݺ��bX�'�oݼO!�D�E�Y�,K��6�"X�%�}���'�,K��;۩Ȗ%�by����7%ݖ������%�bX�ﳻS�,Kľ}��Ȗ?�a�2�����Kı>����yı.����;�8fR���{��7���=����%�bX>�{u9ı,O=���<�bX�%�����Kı<�[/v]�wa�v۹���%�bX>�{u9ı,?"1��~�x�ı,K���jr%�bX��w8�D��oq�����n�sR٦ܱ����k�ĵ��=p��Xxg�>�v�kZ��'#:]�r�M��S�,K����oȖ%�b_���ND�,K����Ȗ%�`�����Kı;ӽ�3&nSM4�m�ͼO"X�%�~�;�9ı,K����<�bX����ND�,K߷��'�?�*dK���-̜.a��l�73v�"X�%�}�����%�bX>�{u9ǂ�`�A��t�9��?^'�,KĿ�g�Ȗ%�b{��r��7r��m&f�Ȗ%��@�?o��S�,K����׉�Kı/�gv�"X��,Ȩ��e���N2q�@oC�L<K�isv�r%�bX���v�<�bX����?mO"X�%�}�����%�bX>�{u9ı,Os�̲v͐˗�6n�=p<^�ս����M�tKO�c��3KE��'8L7�76Kt܆�7v��ı,K���jr%�bX��w8�D�,K��n���&D�,O~�߯Ȗ{��7�߸��X�i�2���D�,Os߻�O!��F�bX=���Ȗ%�b}����O"X�%�~�;�9ı,O:o��ݗd��[�e���yı,s����bX�'��{x�D����"dK���Ȗ%�b}�w�q<�bX�'��rK��s6m�m6��ND�,�"�2'�s����%�bX����S�,K��=����%�`b.��=��{u9ı,N���\ɛ�ݓM6�����%�bX�ﳻS�,K��*�������Kİ~�߮�"X�%����'��oq����o߼�풀��k�$"MPM����rR�ö���q[9"�j4��7e�d��ڜ�bX�'����'�,K��;۩Ȗ%�by�����QI�L�bX����S�,K���e����3]̗w8�D�,K��n�!��WblK�����yı,K��mND�,K����Ȗ!���}v�>�;#p�xh��7�������oȖ%�b_���ND������>ϻ�8�D�,K����r%�bX��|}�w6K��)�MݼO"X�,���~ڜ�bX�%���oȖ%�`�����K��&D������%�bX�}/J~ͺ\��sss.���Kı/�w���%�bX>�{u9ı,O~߻x�D�,K��wjr%�bX����އ��@di*�"�x��8�$�
T��e%)+@�PB�X���a�XE�`���3�uR@[i�sL� W��'�9��hH�#@#�>��	$�oft�`�*�JB�1 ��H�0�x^�����S��u�Z���ܸ�nkW��=[��;9��8ˁ�У�$��EaMιc �d��C��G�K�e��چm[m���N��l1Y9�a�'dɕ8�T؛8Xx��@�T��t���N��U(I7c���;jh�Ĥiڃ���ݲ��֧��FN���5��2\�YX��1�KC��7v��MS֕�� \��׬*Q���F^���R�5�-�3U5m0��O�V켧�z�l�s�&�e�C-UF��7KQ�Yv��t��kYp�Lt��(tی��
�+!�I�[S����i�� *^Z���m�+P����d�r���Xm���R�mJˎ�Y�V8e ��np�:��u�bQ�,�i��#�n����ɺh����k83���V�T�j�
�ࢩ�P�M�b��dɜ����FN:�TGnONj� ��1��I[8�1�Z�vviUxvR�m�@���lݓV4l9�[sm t�6�[[c����G�X:g\�:�l����=�sc*{!�KcW�]ێ1�(�2���aRmVc�b�,�(�Ѯy@�[�� q��5Х�v�f;�v:�� ��A\�A�In��e�ЯW��%�F���;�Q*ƺiIn�
�X�v�:'��h��1
���� scK�:0u�=�cJ�Sel�Zq��h.Is�E�{;l���p�(�3Usi䫝)���2��em�E�i�\�t���^���!�[ ؝�h�^���ur-S�d�x��t��88\��lp���96��Ꜫ�N��d1��l�v.�0�ۣn����@[����<k�a�h�^U.��ז�7\e��N�q��'X�W�$�[`���d+�ch+�˹��K�U;`{L�H�"،k�sl�1WC�\8����)rˌ J��T�����Et���y������������(�� (�8�Q:'�����B��-�,�)�$���ڨ=��X �5H������e�B.�������X+��m�*Es���ꦷmk;p�;��v���ε�%��J��b��Z_Z೺��`���d;f6�9�ƺ�g^s���'%��D�9��lM<.�h�Td1�y��'&��,��r:�-��"�0p{]��OU[������V���6ckkh����k�:^,iX��Ֆ�P=h6�n;���bfZ���{����k�o���ާbX�%��?~���bX�'�oݼO"X�%�~�;�?*"O"dK��>���yı,N�������p۴�mͺ��bX�'��{x�D�,K��wjr%�bX��w8�D�,K��n�"~\��,O߿O�\ɛ��&�m�����Kı/{���"X�%��{�s��Kİ}���r%�bX�{���yı,O�w.8[�n��2nf�ND�,� �ȟo���O"X�%��~�u9ı,O=���<�bX�fD��?mND�,K�����͛�n�s%��'�,K��;۩Ȗ%�by�����Kı/�gv�"X�%��{�s��Kİ}~��7-p��-Kxx�&�YȒU��ժ����m4��#_���|�>	����\ݺ�D�,K߷����%�bX�ﳻS�,K��=������Ȗ%��;�YP��N2q��j�S1 ���I����Kı/�gv�!�����P�+C�My"X��w�q<�bX������Kı<�{���%��oq�8�㾱q2,�T{�oq�ı=�~�q<�bX����ND���ș߷����%�bX����S��{��7���_��f{4p1����̖%�`�����Kı<�{���%�bX�ﳻS�,K�L�������%�bX�;w	s�3&�i�ۛu9ı,O=���<�bX���{�v'�,K��>���yı,s�/w��7���{�����K�F6��P�:x%Ɗʶ�s\%r�b�j�q�����O�s'�t��w���oq����ݩȖ%�b{����yı,s���<��,K߷����%�bX��~˙3��3v]&M�ݩȖ%�b{����y�#��,���Ȗ%�b{���x�D�,K��wjr'�TȖ'�;���7$�f�K��O"X�%��~�u9ı,O=���<�c�P8�$D
�%<NDȗ�gv�"X�%��{��Ȗ%�c�]�O�m�7g����{��7�w1=���^'�,KĽ�~ڜ�bX�'����'�,K��;۩Ȗ%�b^�����4��r������%�bX�ﳻS�,K��=����%�bX>�{59ı,O=���<�bX�<n�����j��S.�k=f+�G6a׮�4�&�h����+\<\t���f��]ݩȖ%�b{����yı,{����bX�'��{x��L�bX����S�,K���������3v���w78�D�,K��f�!�9"X����^'�,KĽ�~ڜ�bX�'����'�?�D2�D�:v�Ys�7�n�i��59ı,O~�߯Ȗ%�b_���ND���Dȟg���O"X�%����59ı,N����:�N�X�����{��v�w���?mND�,K������Kİ}��jr%�`~��� ��O�O�D��}x�D�,K���.d�0�6�,��ڜ�bX�'����'�,K���٩Ȗ%�by�����Kı/�gv�����?���`�9#e��s9x���E��6�6ϭ��tl6��u#K�];t��p�%B6)��?���rb��hpu,�Ð�*"$t�2P\n�y&L�;�gt��%�{�����`]]"�I���(������G��g���� w�m*��i8�jI`b��`ft���r���}�`{G�y8�ȩ'�V^Z��@uܔ����D�[ⱃ�I��$�6��f�r�����n�j�1���x�D��Al�\�2���v���8�;��d�F0RTKV�g�'��� �(0�f�l=�'@r�����v�6��W![�iv9�_ �c��������l�t���0H��;yDgm9��C�Rɜ��Y�ז�Xe��l��͌{t��)R��Ц"�8�#ps�������:�k��d˺{k�@��qW����ع�.\]�����#t5�:77*�F���͍��٠-�6=��O����M�5JJ%H�qXgt������$j��3:x�>��z�o2�7�y��D(��P�ܖ.��3:qg~��k� }�����IJT�4St6�z��fm�`=�z�r. =��7��us�.��D)tD�@}q��2L��w��1�y��8��i7$�8��
ɳ̉.*ae���nOg�l�w1ez�0�p��ka���(�+�1f�36q����f^L�\l{�@���z%�<���12D�����eI$9w��y�@}{����2�2�=�s��&&LL(x�o-'����)�"���h͉	��tHQ�,=��f�yX��Ձ�7����������T�Ȕn+3�����׽����,���|�~}{{�R����.�sRZ�.���5�WH�rZ�r��Г�j�F�QnW�QJJ7%X�y��8�>�ܽ�����Ձվ�&�#�I(R;3�J�נ.�iP���̓2�4@y臏!C�*K�&J6=�.�iQ�ɮD��N<oE��� -X�F� �����"������}V��;3�����}ԵQ̌�n8��X��@{ﹻ��=�z�ȸ����ˮ����!�b�֑��H���)-��4\m�ۧ9��pRӤ!��g��e��]�H�3�}��ml��7�܎Dʕ
dD�%���י�2N��4>oEw��y2N�wO8�'2%��7}�`b��`ft���r�3ky���n���%Q�,9&|�ފ3���נ�I�6	*��_��7����Rn��r��H�̂���=�z��=�Oe�;���7ۋ���e-���WE��gY��X�[v�s���5`m�ݻR�ۓ3�������{1 ��}Ϲ�h�x�
�uz��7U%E`�����ؠ>��(�7^���3$��?=���㑧%�˽��������foK�z�'t9$�r(92fOy��y�@y�A�d�3���;��C�T��*m���k�̼�2e��5��׳�-�/£yܿ�I����6ͳ32����0Z�j.�q�w7���S�;knv������Kv���p2옐�����lb7a8�ŋh-َ��m�ᇚ����p:�Y��"���$��ft�5Zۤ��q��{b�֣J(3[����Z6�nk� $��݊�3��ӣg�m�MŖs�� �{y:]�`^Y��m�z�ʵ�GZ�� e�ql�!���};u��}��ś4P�@�ɳ�,�ۓR�˖�[e�k�a����]mIZ�k0����:	c�m�>���oy�@}{:y$�o�/#��ռ����!D�$LL�oy�^I��ܼ�‼���ٯ332N��QI�ɇ)�������`}��Xgt�1f��9���hq����Xc�Vw�4���&fI�:���W(�@M��ID�Xgt�1f�3:q`}��X�S]N�PNA�$MJt���P�f��\7u�jv}[Zɚ�w�g��w{��N0�r�M�$�[�vgN,��+ �ޖ`�.N8���Q�rI���uS�)긠� �T�\���4���y�;���:�D�)ԅEM�X��V��,������;7�Ł��֛$e)2$ۊ�.�f���ؠ>��(<�y�Fm{�@o.���҈���u134����dɯ:����z �ݚ�37F�Dr��`ks7pv㛂���n�.��ԙx+���s�7��H���uwϏ+���Ⴍ�'�� :�J@ɈOe�	���Ԫ!�J���Xc�W��UI�,[�vgN,����Bn&�J&e��vh{͊5�%ko����0�l��	i`�B�%#%��iK	�2�)	(V�!,<��Lz AA����"��"ے;!aJR�1%��m� w�@�m�S�pv�B6J�,�Im����X��#粦c�F*cj�1�����BQrH-"]n"dd�����a�k/�J�#+��K�^�� ��_�SD8�������!���x�� q��_NӪ� &ww��O{���vUNS�)�q6Ԓ����U-{�v溜�}��3;���S��9#�I�K�11@]��@y�2K�$�f׼����`b��`}�GR��)��Fy���jݻ]�&��s�?����	�XSF=�L�΢�S�IR�HTTۇ�f�yXf����I�2_8^t�@v��w�3R�FD�qXf����F��;7�Ł�>��U_��#��!���S�%Q����Z�dw% �bx槈���Jq�S��Ps&d��:��/����I=���$@T�)PS-�� ��3�TCR�GC��>�ܬ���t�Z�d��8�*r������1vy��V�qu�X�s���s�bӷ^t���V)�_����;���o��vmx�� I�؀t�Z�dw% �ڣ��
S��m�%��7�������3}<X��V��,���i�Iˏ11@}{:P\n���3���4>oG�p�6A�r&T�S"�Q%̒{��z ����b��&d��\P�˼.SyR�%܈�z �ݚ��ɲ3z>3���נ>V�4��3��g];�t��ex���\X9���N��t�����6�]��7!b�U��%@�$��8�\v����rTOq�:E�; �mk/E���۬��L&�$v�ې���|�� ���G]��P��G����۬�;��������=+�9W��l\L9�▔�n`�r�v�ǥ݇�v0H�uv&��.��M*o�{�޼��U�풂z�s6ZK�k�lY(�TrH��{vw���m����{�7�But�u)Ȓ���{����Ł�����/���5gr��O.<ĸ�3�Y���܂��׳��^�f^ffh��p?��)rS��D�@fǼ����I�7������Z��R�q�RP�V�_�RY��`j��>͜Xc�V�-Tu8�FJqFDL�����,��Ł���כ6Ջu@��S�6q�H�&��i6�-鵜��]I�TC�-�������)�&(�'J�נ���$��[�vq�?Q%Ju!QSn�����}@m�B��@�J)ffM�(#7�����>��(�bN��*2Tq!��foK����y��y�@f�<*Q
S�%Q�,?����׽�`f�x�>�ܬ?�R[���:�ަ�҈R��ԡ8��A�ﹻ��tw���%�:�a�k�P�����r��[Ð�o�U펷W�U5{#�:Y.�n]n:b} ��H�1 �����n�< {��S�*Rn6�J��37���;���t���}��;���8�N(�s����}��9��J@{%��=B�G)(��%(�>͜X\n� ]���g���7M�u��*ȥ�DI@}q��2g�ޟ����`}�8�;Z�s�m�@AI9Qi�L��͎��m��x�1ms٭H�����E�mO����uuR���Cn/�7{��ś���:q`}��X�����%A*�I`:{-�2���{1~���'7ަ�҈�s�R��3}<X��Y���ޖ����u���T�5RQ3w% �b��h'�~��}ݪy S�G��}��I䞭��T��mT�9�foK����?������u�$�뷹	�!�Iw�v�v�,qw:v�Ҋ�5�.��mkX.���T!D��JJr�M�ܟ�}�`}�8�.�u��M�J��zh�q�̊5�IG�����}��>��`[�lV3s3(���(Q
(�;� ^�yXۮ��5���X[��]Q�)ʊ$6���X�y��8��W��6{��ޮ�M�ID�J�rX��@7�]�H�L@W�p�w~�Ϲ�\�ԥ�ݧF��]'����z���ˠ��=	�ֹN{v�]��M�ӢS'Vw��j[3��D�l0��g�Msz;k����0Ke��-��kb��,�`;G-��F�`e��mR��Zp�9x�IɷF!.�g-v��o/;����,�[�t��Ū��ͺ��R.r��Ѹs�&8\]7J+�4j��ku��i+����sKM��܍�U��+��J�usv\Qmt���\�(�4Dz�W�R�t�Q��H��O���\��t�Z ��NNg2��]�3�f���\��t���+�2d�s�(���y�L�&^�/7����أə2w���̎�6�}l�$�ٷ6�3w�~@_�E3�?~��g� ��H�f ;9{EK$����RG`}�8�3r���X�������E����H(����r�ӷm�]����a��]�����j8���;��z�JW`���HTTۆ�����}���ŝ����Ł��u�Q�G�����$���y�U��*�˿�g �����}��ͭ�:wDRQ$����t�{�G�Un߽Hｈ�{ܙ�.[�7a�Iws�~TO�\�����~��& �)���ժT�K��&d�>��zə�%��ɒ��zl}�����Ҁ3qB�*#`f^MM%��Mˑىcs���q�uc�gm@��t�����ָYN��6�����%�:�!����R�\+�����^!4���y�&L�^l�@n�yXٽ,���s$�����33ד�w�F����&a/&e�,��3y�$��髚���@j̐��*S�U6�`f>�`f��1gs�>͜XY��]Q�%EH��`^l�d�%�ɛg}�3z|Pq������?~�I�P�*��#�룥�T욺3���l��Q�.n�ں�wgE���efbӒ�s �n�}�����,�����q��*)Bq��8�;������4���rfwF!�zNRL��!`n�yXgt����RZ��v溜�]O��j2���z ��f���ؠ.�t��̓2f�����uߕ�{E��8��q69%���h� �n��& %0��z �f!��B��c9��x5n�֭��W�h�mӴ�鍕�eh%C��|�N��n� }{�̓3|Ꮭ�@z��6z���**��p�3r��٠-�v(��+�d�;��f)�L�B$F����1gs�>ΜX��X��:N�E ITI%���Ե�tP�<Pq��L��'{��5g���Q�!QJ���6q`f>�`^l���'f�@C�Ha08F|T��[bR4�
$$� KT鞔#��D4�Ċ���F,HP	��	�!OS)%�`�Yo�2&e!!3� Bi)V64�K-*R�%�JZqb&�)	�BS4��'���¬$)(F��!*��Y	F�{�p��E0��|�m���&�n9�����[6�&��+�.m�j�������=�
ґ�ny�v�M�y�.��k�8���c.��ױ�L�8*}2�2�yݶ k���Y�ȉ�'��-��n��\nm�V�l�d���k<TM�^[p.Pг���g�U:�q�K5\�l��mkp�Ѷm۩��S�F\mAc���e���������a;p��rl*��R'7k���	�'�@��m�$�u<����f1����8\��3֍�][����mٻIl��@ܘ��;�nzv��<p][�ڇl+��M5KvL�SS�R�Vm@�+K�K�:^FH����۰fR�U�$J;l#=.'&T�b�/-Vg� �*�D�S�.Cac��MF$zn�(D�����۬iF6��q٬�[i(��-/6���v����3=�@z3�K�\BY�2���k	�l�2]��7j�vw����ڴ�5kn���sv����Wi���,]��0�;�L�媗�iUxuW<팈Y7RF�A����s�kʹh��EF�ڬ.�,�n���c����u�����JN^�B��8���hx�Mǒ��,&DQ;��-��U=����`�%�q����Q̫*�*�[l�"���3�xA{\(Ų�Jԥq�u�Ғ�K��N��i��Vi�b�!sfj&UU#����j��m/C����v�ʝ�Y"Z��s�e�v���d��a(`�WCsn�7\ta6�n��={2I*�d�tM��[/N���s��������\�7+D�F�R��ch�5l��k!ևf���Z8��f+J�5@mwP ��kXSeLv�2PO�X���@Q�nĮ藖���E��j�/lj���!��Wn�ؙwnc�s�r��[l�ع�8�ڍ]G`�]�%�[��aݧ���*���$*�k�eƵ��v�vl �d���Pg��;T��#�ۨ��Z��m���UW�j���Ԥ�����ܨ��%�	w_C�gD�u�MT�U@# �<f�}�~ww����v8�뱃^�p����B	n�W!�����R��.{q2v�w5Xˮ��c��h'�k��D-�0��H�Pa ���{��\ӆ�v\h��\kPr�l1�bE�h����nb�UI��x��e���Pa�G.I������N��(��7<��^�pv�P)�W]m�����/\��%��s:��)�=�c�8h+&x�u��p���7R� �kp�mɫYY�[rm�w��Ȯ�&�	nH�t��\�\��z	��7^�>�٠-�69��&o�36x�<���?T%&�j��Ȭ��,݊�'J�׮d�2gp�O�B"@RTn&�$�5o��͜X��X��,���s$�qJ�$����Ҁ��נ�٠�d�3�gtP�d=I�T�EM�X��Xߖ�>V�����Ł���MI$�D�H'�ɓ�,öMe�bJ88a�!w���A%kS�z�~��M�N��*J$"Dn/�7}�`[��P{:y2fd�����j�!<](�ImTNKw;��t̝8�3#5��vk̓$�j��")<'��!��^Zw�� ��H�1 ��h��WT�u*7B��}��2�f���ؠ��ϙ��Ό\����/,�3��R nL@:{- �� :�r�?�W�o�А" ܃�H��jT�T#p��s�a�a_&���H��a�?�ݮ��6p%F�n��`������Ł�>��UU��@n����S�K�)	)72��̂�� ܘ�t�Z��>H�ހ��RT�**��qX��Vw�4�2v{{͊�7^��Y.�KD�/.�DK�y2fN���@c��Pq���L��2������;�'�O/5 �D�1f�3r�>�ܬ3�X����F���D��'Z]��gAw4�d䆖Q!��=s]`ٵ������/�R(���8�u����}��3;���;��uIuuF&���"�3�ם�3�h|��7^����F.Q�IO0A2��z ����b�2d�n�x�7_�������9*7t�fh{݊�gJ�7^��2e,��I���7����c����$�������rb��h��誜w9�O$�s�n�]ѻ�?�7|��`֞U�1ڥĬ�!�X�����m��{~� �����̂�7*����!Q!��fwK�5oy���,��+�~����w��t�Q5Q9�7����Ҏfd�������4�w6��t�Q19B���8�>�ܬ3�X�y�Q�.�����9�D�@}q��3&O��?���@]��@BfL���] B�pN�b\�����:z��G��レ�;d����^�rޭ΢c��6n#rv�c�����nɭ�5��h�$KZݸ���,�^���s�c�R�ʷ-KuqM�1�����iGp���;'>JLJ� �V�`L9�X�����X�Ν�m��+�v�$d9g�'�t�j휗�7����1�D.)k-�����1y�8�v#���\�3�f۩;<\Du�;5�iJ��x�}I4Q��JIB�NT%&�&��H�7�����̂���F԰��Q��jI`b��`ft���r������*�Jt�M�8��g�]�H���t�Zt�*���HTTۅ��>�`���ś���:q`f�ğTE8Ț������t�Z�dw% =Ͼ��W����YyB�d�����ܳ���]�bE��:n�kd7M/��\mY3sLBtfg@���@û�� ��@=��m;��BF�8)��t��~�+�W�)/T��nO~�v�I<���$��~�`F$���4����Xc�V ܘ�t�Z��@JἜ��3�w�����H�1 ��s ����>�j�Ҍ�����,�vs ��) 7���ʮV]�]��/ll�F�)�QEj̯<��U�z����	I�-���.x�[jg�������`�r��zX�y���&���f������) uɈOe��Ł�[}Q�:������������%	32t�]��@e�k�����R�$�9,Y��͜X��Xgt�3ky���t�!EaW��ndܔ�:���%�o���}�k�,�he1�e�
�:q띄�]�klu���jϮz�n���y'5�� ��H�L@:rZ�� ��ЩI���(�+ �;�����_y�͞(�1�̒fL�k����`��M�I`j��;3g����}����Үp��#m���a���3F�}�͏y��ݚ�u&d��DA�Tb����s9$��5Ԥ�N�**m���r��zX�y�f�,�I�8�d�GMԙ� ݙ���5�ձq��d.�d]�m�^�G��������E9N�8!����`b��`}�8�>�ܬ�y�;������Oe�:� ��) u���߫�$oWy���q��A��ޞ,���^�@:{- o��'/�\/��3�����\��t�Z}�&O��� pj�"����Q3/@rb��h� ��) ��%�+����4�\ �z7T�s]�=X��s��<��M���9��ˋb�����G*Ex��P8��`ݵ��g���q[	�)X�85L\�Ŏĕ<��Kszz�'睺�9Ƨ�\\[W�x�u�.��0a��{d���@n�~O�ყݹ�q�;�r�n���Yr��%h�tLJ�9Im6�I��{�vH� �ab���$!j�n����`��z�V��P�&�z.�[H�\�s��v�6��R��	�M���q7C�|��;3g���fd�8��@v��D�ʉ��]�9yyh� ��) uɈOc�;�mu9*S�
 ۅ��>�`^�����/&L�Dk�z(ޟ,��ꈧJpCn+ �7���7���l���r�7M�&�N�9��f���ؠ<��2�$əf��,����>��`w4�>9$�*i�ut�l���m���ч5��]�����6M��Q�`�����f�,��+ �7���7��m����$���!`}��yQC�$V��\j�A

_P}��@c��P^N��I�w�W'ꄤ�RQ$V�ޖ,�vz������~�>�j�:�$����A̛ɒIF�������@}q����K��JT�*�N8��g]�H�f =���� .������́�Ϋ�"������zw��+������҇�����D]��t��B�6����R �وOe�:� ��n���e�:����V�oKo;����<�;��ʈ[;���.^�3v�]ٚ7����t�UX�0�:�@�$_����~�=�JqU� AX�S��c�!H\�0"R,b1�� �' 	��!-�2$�!�.*��me0�����(ؠ0Dd $$U�@�1.1��ĀB��VXTIZZ�0.0�1��@$=�,#�,K,dR2A↑5�*�*��$����#���~E~
��4��%eIK�cH�$�rҰ�C�~U�~���b��>OPC�)_��O�S��H��+ �ޖmo4ۺ�����(�'J�נ�6h9�2I�3z(A�^�S����J���>�`f��1f�>͜X�-�J��$��rԂ�{Y���ډ�-�C���u׸�u��ӡ!(�JS��(�?ID�Xٽ,Y�ד���/2I�6=�3�8�IQ8���,Y���gc�V�oK��JT�*�NH��'J�7^�d���������v�"mz��J�Tۅ�ߪ�n�yXot���ZfU���˶a�Q,�S�#qXٽ,�׽���<Xc�V,}B�SrD⍶��Ű��,�J�+@	vH�3��؞u���N�K�D���9�$�,�vٳ��}��>��`n��6(r�A���'J�3$���w= ^oMoy�\�&I��/W�STH%B��~��zX�y�f�,���S�ҔiO�8^e ���t�Z�r���sӐ�0�8���,Y��URW�\|�w= }y�@	�7̙2P�	U9R�f*��ψr���ݸ!˝�vClZ�{]i�jv쩚�Ey֯g��7�z��݅�5��r򹛀�u�g+�#�!�t�t�&6�g�iuq�m˷	����i�Z���0!e�<�഻t�\�!��VS����	u�,��uyHٷ\I����~|q����4�i�nsi�������:q��Cƺqj��Cٴ�9[�t�l�n;�����C'l:��"9�m��չ"-7��6�ܜFv�����ĒʒECpq��O����}���ś���6	���(�"TӅ��) u�����{�@n��W8O�:%8"7�}���ś���6q`}��X���j��S�Q�`b{- ��w% �1�l���ȩJq�Pn;3gc�V�oKo; ���s)JNF���	M�tn�knra�gH�^�3m��Y�����1�k����"~�	�Xc�V�oKo;��ŀpm.�ߥ(ҟ��Ȭ�ޚ��32VɓD���N���@rӐ�0��M��`b��`}�4�ə$�y�@��@}�1>��D���Rpq�f�,��+ �7���7���lS���T�SN��� u�����{�@v\�ww��Y���+�Y��kLp촴vmhʹ6!w�w]�\��c7k�[]X��Ͷ��~����ד�$������j�x38[p�wl����I����~DE�{�g�u���>��~H�;�6�D�"q䈘�/6x�.�u这$Ɂ.�UG}=,]�v��}R����J�&fI�'���zh{݊��Ҁ�FR�}�R�FT�9�}���ŝ�@}y:Pq��2e�&�\��5	9.��e����m���-�II�E�nJ�F:�)D�Ru �lnO�վ�>͜X��Xٽ,����r��JN�;����#u���3}�`b��~�H����GNA)��,��+ �;����������Ł��ğPL�rdrb%�92fN���@c�tP{��r@��AUhb��-:�਄�D�@�sw��'�v��$��F�)$�1gs�>͜X��Xٽ,[���"M��H���P�Md'k:7:ݓ�t=�\k1�/2��YZ��ʂ�REIA8��gc�V�oKw;Po>�I�Q��,���^�@:{-׹��8�����C�Xٽ,Y���~�K7��5���;��*@��M��@:{-׹]�H=�S��@9����ܦ��$vٳ��}��>�٠-�6(h�&g}~�N�xu̅t�Žd�s��:�Ms���/F�m<Kk�Z3;���i���Ɛ��g��=�8�g.Gf�[՞�h��<��l�b�β��a�gc�mխ��jG46���[2�d����˾@�;��A ������f �<4Y�ӝ��p�b���l���plG[��&v����^ח��dخ�9:�����1���g��������g�G��w=hH�F��s��鵜˒b�VR��,9�<�)��Zy����zX�y�� �}�`gWD�����"D��V�oK��[�vk�+�}��ͭ�黤��!T���ś����>�ܬ�ޖuo4ۺ��REIA8���+��׳��@m���3�A��ᙔ��) uɈOe�{��0�i.䍡�&$�D��s�u�%yX�{�/V���ցL��:^��9�C�!Ȭ��,�vc�V����v-��T�H8���ś��e�L�dʊנ/#5��͚�N�ꎯ6F�6H��9#�3_yXc�V�oKo;��&>duQ�Tw���) u���%��ܧ�=H����DH���>��`b��`}�yXc�V���)Jm)(�N���`�n�K����j��n���K3�iw(A�r�l�(ڥ$�,�v�����>��7�:��m�&�J�$���@v�� �{��:������y��RD�DtI��>�`f��D�D�"�/���Q<����8k�V*2�S�ңq)IȬ�وNK@u��A�}Osޤ��=Fr@��j�ܖ,�v�����>�`f�������P�D���I�F�)�46"�'/5`�<I�	�����t�nRu"���`}�yX�yXٽ,��ulk�%7F�7oe ���;$�]��}ʢ{�ğ�S$�T�A��7�,��������������Iӎ&ڥ$���b���5���z�gL�C;%��TY��`}���m�(�J�$��v]�w% ���t�Z�%+*��Mv��qc�+a�
�md���̝tn�'�v�;*Fn
6���{T|�uܔ�:������v�v� x7��~�*7)8���>��~Hս�`n��>�ܬǵȕ G�F�RK��h�e :�J@rb���F�ܤ�D'�������>�`gt�1f�>��&�2JnR�
�r�w% ���t�Z��Rxs�w	ra���R�1�2TZ�^yD���!F �B# @EdX�X�D�RB2��X���B1�����B� F#FD�$`!	aY		D�"	�e	X!܉�~c�+�{}�iJF��X��e/���
[a	Hn���AW�$'e�$���`�e� @.\E^�῎ ~��ŌBc�`$!$3Z�iI��������U.��ÙܷJi�vm`�v�t�=yjbz\�׸[�'I�pC�7:�eݺ�k	B���v�(<s�[�i���lw<úMa�J^0���q��|�';��)��5��|�mS:� �n:We]��S:	�u�m���Z�������y��X��Y+v��#sU�e:�ϧf+e*mt����og L���iLNqQƌݫn1�Nکu�mw�I�򣯄j㱙���]��<6��<6���0Ҧִ�!m�]�f�:�{:������L��5���dRت�2�l�Ӕ�;v-XU���˪^T��t*bd�ڥ�Qu��2@�<���,� 6Hi�L�B�fyvAܹ�5j@�f�n�u�5A���.Cp���k*��m�u�yQv��m�7%nv&�՝rsHv�8ꎜь��� Dv�a�����	�<.��r��n��mmL\
ch|�4���\��P�8ɇغ��{]�뛋w3�z�r�������R�sW/�8z�[#+�l�E��� fQ��݃�������[��2s��s�K	�;%��E��I��M��:=�^�w=9]�g�Xl�,{�I��y{e���I�f���9UeZU����)���������K��k��
�-mn�Z�W�?2���p���g�����=uU*����U������6��U6x-º�<KM�$�;�Q1���4nM�ͧ�dN���/��ڸ7*cM֗�3��s$����KUf�r��l�.L/�Y�2D�,���:!�^8Ha<t�&�kg����{WUUef��<Fy'��b��*���p�>�]��������|��d6E��Z^zQ�^�a��8;iq���F�Z�=��q����v��tp.�Ӌaˑ���j���"����Khl F�+v섴6�؀���e��m�Y�kVcY0[�T���ʚNBV��������USs��㝕3���ܪl���>�"#��=Q�꿑QODh/WQ>TNb8~H/�:� ������d�6]�d�F������������t��I''C�:�V�xv����I3r�Z:i�ѵ�:,s܆��'=)��8{;`C<`�4Ct6�3Ͱ$]��������\����g�綺�b#>��ظ�S(a��	�r�Y�'n��-�@����]W�����t���D6�-�]�;h�kp@�>�8�U�rݜ!�֮Ñj��M�4�����������lm0]F��6���X�][��ECHA�������iۋs��n�J�* G�NK@u��@7rRwj	Ӻ�$M5JI,Y����+1�+ �7���[�6�N�IPRZ��R�������C��@mo�hA�M��M1�$Vc�V�oKw;�{��86�S�ңr��"&^�>�٠92e��������n�6���}�%t��GV�Ak���Ե=�k(�x�^y�Wj��\][-���|*����뽔�n�ײXm=��E �H��9#�>Ǽ�S%l�ɣRI&�#bi��͚��b����UI��&?2:n"8*��`f�z�^�@:{-�{)���U���Dd��>��`b��`}�yX{�͞�;�xN���9"i�RI`b͖�뽔��) u���]�U��K��؝����Y��<y�2n+;�sW=֝n��t<]X�[�z�!a��o�����>�ܬ�ޞ������u����H��"�3r�W�߿$��`j�y�c�V����Tܤ�r+�O=���'���98%��	��7��׼���u'Rp��n�����뽔�n�׳�^�\��N�����
���L�fGs�y�4w�4�գ�""�����.{�}��툩d.�L/�N�r.)��{Pi	D��A1�GI�����Vc�V׳rb��Rtܪ��>���$D���lW2fI��3�h��Vc�V��t7NT�IG`Ɉ��H�J@d��e���(�J�$�)%��Rޞ�7_��>�w�q
�_UP�}�w�I�=�m�Ji��#�H��ܬ7�X�����X����B7*�T���˝�m:g��ԈnL�x�]{�p]����{mq)ʔJjR��H�7�X�����X��Xs��N����'$�-�v+��3���@fGs����m=�l�A8@n!����������L�$������2�H�F�0��GQTN+1�+ ����,�ܬ�������FAA��7�P�������n�L̒�B�����_����iH�e�3v�]YqA����l��O*�1��v���ٻb����5�-�Y��Cc���7F'#v�Q!�ꛄ�ϟ6~;�;l�T�Sgh�LO%q�@]e�-���9��H�x����N��ֲ���Obnm�&ބ%�U3��1�>5�m�y8��G�}�d�v�7n��8a��ݝ�/ca����(q�议|����7	�s�z"�%��̛��7v��Us�l���n�����31��5�qd���P�M�5)�NT�I�9> ��K5�+1�+ ��i��n�D�S�J��X��_��H�~��zXgt�RA�7���Ji��#�H���+ {& ��ے��N\�p��FE`���3;�������Rݞ����'Rp��m9%�fwb��H�J@d���g�wV]l�BhUͳ�9�m�]�nM	mzV^�a�{*8譖�zz]5��r�M|�?_�i ��H였��r���e�&�ۛy$���o����&w{���7��������|�j%yH였t�Z=U���@=�z��5tۧ*F$Ȝ�,�vk�V����f�K��j�D�T�J
��nJ@{�{��tg��NK@~��^�c]��02�$��Mf�F1�$k:�43�����U��1�3���`��H�J@d� ܙ��l�z�i �WR�?T�1FTa$V��K ��k�Vc�V�-���T�RA��<L� ]��y�F2ei�*�����L��60��U� ^���(ů
b`�*Sq5�k�Vc�V��,3�Xi�&�2:RQEQ8���H였t�Z��H��*������r>x���Xns�f��u�l�f�����#�n����9z�A���m��1 ��ے�w% �vU�T��F$Ȝ�,�vk�V����gwKt�j�R�����ݹ)�rR rL@��8�˻������(����ɒg����頓�~��N���#"B1`�FbBF#0`F"$HE���)`, H����0b��
B�~^�f�@�'��OT��?^I!����餻e�s�fR rL@����H���o�w���~�?�,Xn���=tWh��n���-�n�uֺ��$d��JSZ.��\T�URI��zX��XgN,;zXu=�N��N)���Kq�R�d�1 7���7I�ʻ�	�J#��'�����3;��foK1�+kv$�D�8D�H���1ɈOe��)������vz�u�NA&I$�1f�3r�>Ν(�vh���d�0�I��w4��8�HU�/;`�Tm�Q��Y��b�fSq�=���u�Ud
ه����mtmv�e���0�]�g�p�Xb;�����t�q�6,���|M�+��%e����ݽt�,Fv����E�K[B\�� ��.�*\�x�	��#�Y�J�K-r�8Ԗ-��rod�XѝL�T�(l3�I�H
Y���m��%/���CT��y��o۹�n�-�pj����U��.Em�l��6��c��g�����:�%k=t�)��?���@û nL�����@祗W�g-8�jJ���r���`b��`f>�`մ��T�JQ��$V����@7rR���[�wU��S�'Q�����,�ܬ��+~�Ԗ�,=K��	�)85�w% :�J@Ɉ����=�������\OB����o=dh���Uf�����%�S��vn[�YK8���q]������� }���\��=[�.n�0ݙvٹ�y$����4T:���Jd��$8fo�@}�����@^aΚwM��$��%�foK1�+�}��3;�����M\#D��%Qfb���w% 6b of 	��4��4�!�(r+�}��3���fwKu�+ �ҷ�N�$��9 8n�n{\��'5�ylFXz�'w>�ڤ��q=qJS�(Q�%E`���3;����������}�k�JT���m91 7& ܔ�n� �L@��͑�I�	��$�3_r�3r���@�-O��� 0%�X@��> D!+����@ 2# 0H���*�upt"0!PcB!�%���#RPR4EXXR#Q�@6H�H$����đV561C���+	��P8>$H�R(�H1I��E��=��� �^�X�bF0�#4�B H� !!���B@j�Q��`�.Jq�f���7n&����?!��:�b�#cX�$��od�HYdH��I�eɊ��y�� ��UD*�߁��|Ez�W�����%EP��<�:��d�������Mzl�:%<@�(�R�^%�9�I�'��;�h�vh�ܬ�cO�J�"�D�V�����ݹ) ��H�۲g��Wm�R�������+WKm�F�ͯv��b���Cŧ��^�H�|��߭�����������ޖ���M\#D�%

G`n��`f>�`���ŝ��UUU�#��co�)'Q�C� 7oޤ 䘀t�Zv������ �#*@�+ ��,�v���䟾?) ��QW���y�`V��F�J�(�FԒXf��7_r�>�ܬ;�X�����D�6��u�G���c0���q\Eь魸@�eb˵\��]7c�(��}��y��7^�/wg��/���z��ty�M�Ԩ�7���������o��`��V��W����ti�D��ʊ%qX�ޖ��������������:i�6�BF�������������>�`�����ɦ��l���TJE`n��`}��Xv��1a�o$��H%A����g��3wr��E�bl�*��E�WLr��/)���Ԇf����6�I���6'�M�q�n`���壍��g��� �a��ѱ�ܘ�7S����.��BCY^p-��6��-�Y��F�x���l���Ӡ��c&��F�'m�I�CBHGOd��B;B��\;;���ŝ��n���5[<5���m�r@���8�\�����}�}���L!wv��Ҕ�srL���1s�V3��uɹ�����lI�(��n�@��$_����V��,Xo+q�+ ������*:$��3�b�6R]�H�A N:�L/9*8�uQ�`bùX��X��Xgt��msb�������H�J@ɈL������؝J����Vc�V��,Xw+�}���j�GA2J���&�i`z{�贉iհل�O+�J�[1d����nH�9QD��V��,1o+1�+�}���ӝ4�u!#ISno$��oݼ�>���E>:��2I.WE}[����w�4���l��Q)������>�`���3�9�m�JH:$���) 7& �e �)�=|%/S�1FA�H� ����f.�`]���q��32d�wt(x�]فMM��^:K����-Q��D3ѫ9*�j�!��S��H99Q���$�u{���}���}��3;��nk��%%RUU�u�yH�J@7rR nL@��`n�&��JTN+1�.I'�����2��.�?ا@4�N8�������`f���H�9D�e]� ���IH�J@7rR7NtӺmԄ�%M�,Xw+1�+�}��3;����U�ꊜ��Aڸ�U��]&��v��]Rt�VM܍�XsnR�DM�)F�J@U�X��Xc�V��,1o+����T���2�fe :�J@Ɉ��H�r�9Q���@��JH�3�Xu��ܔ��) N:�L/0*�uJI`�yX��X��X?߄h*u>��{��O��㹒줡��E`f>�`}��Xgt�ż����<?�6ܤԑH��*��FS�b�gSi��P�[=&�ʸ�N^�Zb���9M�ӔB*�����V��,1o+1�+����9D����rb n�R���w%/}Ͼ�7���nQ$BU��7WyX��Y�ߩ,��+ ������&ںQ:�/(�eVe �) ��H�1 7]���v���)!��:$���}��.�f�.�u���zRMi�d�	�x�����<gm�X�d{&泖��dǅ�'mz������\R���]�w7���?y۟��gCo�ؗ�Q�ᠴ�8�eG		����cpkv�m�������H��쳗s���k۬�g>ycT��,�=�H���<9S��^�K��s[��h�Ў�:�@N �vy�e�hvEN�3n{I��8X�U塖�.fn�	⢏��Q�����̹��-ܣ9�9؆��;���T'e��ձ�JCJbج���涄'E�2�&�u��ܔ��) vk���F�6���ņ�3r�>�ܬ3�X`���IIT���/�@7rR�� ܘ�t��`}��W'ؤIB*��`}��Xrb�6R���y�Ww9ue2R�Dn+ ��,7�������>�`un�.QT���m�Ӡud�z�^g�a�4x^ղ[�F�̂�7TR1*��`b�yX��Xc�_߿~�����;���WJ:r%������o2�#h�څ
��LT��oޤ�{�����]��I�IC�XgN,3�X��Vc�V*6�S�4� Ӓ+ ̓ZIH�J@uܔ������Q:��RK���}���r���`W���T�LnQ#�&�n�sv���Βts����Ns�2hö:M[MUX�RQM�7�����V����fwK���kb�N1�H�q"7�� ܘ�t͔�n��n&�SLN!J�F���`b�yY��(!A@�O�(����?[y�o'M�	�)�F�2���ܔ��) 7& 7M��wDu$#i�+1�+�}��3;����`j6��()I�28�P4�&j� V�����sf����WV�卹�ېdCRP�V����fwK���}��86���4� �I nL@:f�@7rR��g/iu9�Q:��RK���}���r���`u-�N��Rq��p�z&fI�'����z �ݚ	I$�B �b�uQ
';���l��' ءQ"7��>�`ɈL��ܔ�{�Fd:����:�C���vzi;GRh�'�㕺DZ)���M�M18�*%��fwK��נ.�u��o�3:x�7u���Iө	*7%���`f>�`ft��3;���o��'R26��3.J@72�1 �R ��e��	2Rd�9��Ӌ ��,;������peu7�h����,�vh	�d�,�;��ݎ$���EE�DEE�Q_�""����DTW��Q_�EE�DEE�E��QX��������������"*+�����DTW���DTW��Q_�EE���DTW��Q_AQ_��PVI��{)�"@�v` �����Zw�    �                    >IE$��J*$� �JQ@�	Q  �Q@ P(� 
H�T�
"�
�`  �   (PPa�Nz�_{�/}��=j�z�^��������})�=���,���۴��C�z\[����s�_W��ӓ��}� ����K��>�g    �Z@=��y���t���o,��  =�@   ( ̀
{¦[��A���ɧ[�˹zn{��O,}���^�ﻄ� �`o^��}� ןnU9�� �� ��D^�q�tӗ.Ǽ������Z���㳯��� x   Q 
  � {������緧�=^��x  �h)6   6   �` ,�  &��� @ % �J� D�l�   �l ( P �  P  Y� @ DPS�@D
 �o�w�
���{��;���w���ͼ�)��\��;�����w}|  O�R���^� �,�uNX�&�m��y�gХ�C�;��;��.�:�/��� � �  � U �`W>�}��t�:�������� >�헋tӓ_Zri��}���� i�ӓ�2z� ���og�{+� �W�'��}�}/y�+��s�� }�=}��}g��^��+������M�%J�2�UO�PS�UJ�   <z�T��R 2 Ob�J{J*D� �U?�	S�T�J� h ��II4���"��������o���o�fvw;�\�s����Cr���Ȁ��T���*+�T@TW�QX������y����\&�n�m�\J����#B$���e	B2f���0���Y̦���s,!-e�md.��$�	Yd���"ĂFH��*K[��<8<��W)�F��J�:Gf�N]���O�yr��Oxp��.�K�CRf�@ăYR�S)r,�g<�3���VaR1�2�%1� ��g��c3�۹ςV���bhˆ��3|�(ir��<�'��+.,*8q��B%�T�aL!X]�e�.��O���Le�\߂\�]��y�e³g6\Զa�a�`��e<�%	B_/̹w���.��nx@� ��|��`1)��j��XhCS�G�1c,#!�]|p�ыf��sI���!s�*��8ixwg���!�D��1�āgx���<���a�k�)w�����<�0�N2�xI8d�2�@�`B�(�0`��*B��a	$L�)���
�1#���L�=90��}>�O|�6�,�Y�����%�ٜ<0��ewSK�BH7
�CT�Y}>!�<��=���1�ׅ1%�4ҍu�х3RS5!L�!�ǻ�����{�14�=,`Xc��XJh@�B��$4!LM6!F!��̗0�IR,�!6$�g���"�CЅ��B�Hp8�|�Y�7iąHP�q�}>nN%��s|S4/��fa�xx����}�s�Iq!ՅT�4����{�X�Jf�<��s��C�
css��L�S=�S�y<���=��6�H9N��/<��<�E������J@~����~�~�	���6le���<��O|����)�!�Y'�~�,N=����Ǚ���W.��&�}���~_�jz,_��S4qw�o��O��j�8��[2�~����$�;L_��?7�{3���߿ s��>���y���I$���>�.�эFSK�O}��>�ĂD�ID��!L��\SS hfL9
aL0�<7�H�����8��Mc\YNBp4�7f]�3@�p��6I&f,n�bB��0a37��H2�8cla�pЉ�"o=�S7�L���L��Z�.s�����"Ddu��%�P�b�d�.D��	ƭ�� �P��SYG%��FO�O<�z��X�x"P��!��B��5�%��ЈشH�,&���D�R40X��$���0��$
`�V#�F�u#\��t�'�.y����g��CBo+*]�p�p̘�a<�^��.R[���a�B�'<���np�`B��q�!��yJJ|��	+��J��˘�K����BJ�$����3 K�C�x��.O���ݴ���9#�|眇�%!�K��9�zC��M�0�XbƁ\�7u4�M��9�.o$x�'���%����7}'���l7��`T��ԅS��G|�����B��y=7ݧ�I.-JF��,�|iC�/m��&��$X�2`n�o	M�80��zºf���.�����8˞�ɾee���7RHذ!G���fO_�<n��6�K}7t<����+@�`5�D����H�J�	`|$
,`$�2�����:X��!M3������<������� D�p%��n�_<=��}{���X�3.%��<8�HRجJ>��
�F�)�0Ԥ+ ���
�Jm�s@�!2R%���Q�<���'�}H$�3 �p�e�"�1�Lb��� @ab���=�3�g�ĉ1aX���^D j�@*D 8��P�	 �0!����@�h���˾�O1�.�p�!�%�#!YH_}e��%X�!Le1��F$r42�d `D�!Lh��X��)$B�1��g,H$X<�&�5���y1����C��S�Ջ� ��	i��YHQ��!��.�4����oa
x�,�L!���~O����`�]����Ҟ0)�@��o���*�!�� B沙�9�V�������ĬXc�0�y��H�o	��
ń����=��
�B��3gM�HS3Ni<����048���������>�������a/�<���8�o���oa�)�Ĺ'�.:C���ߠ\��7�#�<=HS���	�ώ@�)"A�I
�<m��͜��	q�ō�cFR"FB�Be I����1�p����g	sRf���a*J�"�����Ƨ�4�� Ђ�q(���5��Ť!�Ӛa��5�N>7cHP�cn�s�B!#L4��`�]�$�0Ji�q<4�x��'��4)���|�\4�c���-��p��k��p|p�LJaM7�h�p��=i�$�h]7>	��Ōi�#(�St�>,B�hp$L�섒��M79��Jc��n��J�uԍJld!�B���F�p��H+HX�#�jC)禐�% �@�����xK����Xܜ�ݒ��6���ap�M˧��G��p�|�>{t��@�
�Ŗ$#Yfi�a��@��o\8B��5�<�y�����|	s�$�VY�HfL�Si�a�&�2�)o<�L�RƄie�*C<�f��G����L�.�q�)�L�s}�2�2f�hփ!�
�B�K�ְc쒸jB�i=C�� F1#������S@�!R��İ0�5� V7��! ��p"T 7�
B̹�,J$OBHT�6����<��	�Ä)����m�I,����3VS�3%1&��f�����L����<a���=	.n��o�y=��,.HL������as#V8�y�
o!�H��d��d�!y�	t!���0�E���H�LIm.�ؐ٦˙Ja�篆���s|��!s$&��2F�6���0��q�y��.a�hJ��p��B�B0��́����e�	B@��3�c����a�$��J��1��f��(JC!P!�(�d."F�
A�¤H��K�3��H!��!.0�$�e�#�"B$"�@c�S!HRV	f����Ip.$24���ɤ�4�wv5!���4�p����ׇ��3�6����o��_`�y�!���	=�J]��OJ��&r{�����H|S��ꑉ�:ØN��N{�����ul���8y�߾��@�A�� ������D(��0B�)B���� �F��k�E`0�Z@+�ha3�l��1Q %`� ��4aT��@	 E�	1��)(E���"S,&[B�@J� ���!���@"�X����H!�9�����X$�kh���,J��!0T#)c ��k�"�%cH�B��i�i��B2���5��"	1q\1Xa���1 U"�X�$a��'.p��)Y��Cn�!LucaW��1�1�a�,XjB�u̙��5�#�8o(��&��
p%3\!��Ɓ ��L�l4���\�!fi�
$���#@�s1\1���p �3Nd��f��!%���"ILCX�!8�֌��4�)�
�SM����w8h�!p�97/SH�`e�8��\Ӄ
�p�%M�%���Ƅ�	t���2�!c�,�)�a��#[-���*F�� Vfd�l2SNrݼ3		�$"B&B�#��a�*@��D����<��<�n{��iK��=琍�9=��{�CԌHR:���ėb�
��ߤ/��p߷�'�$+�
b�$�p����`Ɔ02YrK�O$��s�А#a��e�|o��I9�!�)
,}����`���D����Ȑ����ꐫ�>~I��     ���l ��  $�Xն�j�\fk�8؝Gl�q]��n�m;qu7겔��Xpp�x�K�mW3�Gq�gs��������Rc#���3E�p��
88U8.��3�
�۪z�g�,72��+-2��x�{v5v��WR�]L�ʜb�.�v�j4���x��A͐A�蕮�X6�m�H ���jݜ(md�p!�!�m׺Բ������~|�]���[  �y�M�.��qn�af�u� H �b�q�i�ASe�U-��iIE�J�d
�ulm�+U��Q�M�k���wM��� ��� �m����	�A��T� cƢpҭ�U3�9%Y��U�	q�+v���YZ��������T[sc��v��eU[��*�ન)j?�>w���=�-��u��郛T�L�޺F�����$ {��M�K�-�[���)E�ȗ�m%lK�pU-�J�UV]̨�p��I� p���ɶ�$�Vt�F:�UU��힎eP�ܜ��mN^�`8����K�UF�-� �JHh��` ���j�.  m�� 	$ kXm�����Ƶ�����n]��`�M� ���z�4�H��/-�UT��  I6�T��N�cr�mm$   �����I��UUU�T�@H-�� -���~�D�im[D�D0
L	#m��  ��M�[@ �c�n�����[A,�k��� 8Ӏڳl	6�@���{a��$� q���v؀m)b*ܶ��W[¯WR�mTR=;s$�UU@#��
�y�9y��Ryꪮ���YV�1�j��U'�Z����lŴ^�|o��������ö��r��pt�
^�vUaų,�s��m� ��f�}v�}�(��I'[C������m�5�m�$lm%�1e�` �חC������k�ƲJ� $����Wl� Hn�v�}��n��'I�������x��Q���B]���h#3
�7UV���S��U���[8x���{�e�b�     p 6���t݀*S���0����(�\ m$h���lk�[{m�M��Ø��8-�+�Ԏ ɛq��N�G����j�,aq��e�ۉ ���E�Pg\�!GmF��uA�܌���A�1���5:�5��aƁ��`%`���[@��G hm���$�@h�&������hƥV�]"��I�S�ꮕ٪Y� *��ZI�\H� m��Bc �39� V��uUrܘZ]�7�����٫�`*�1Hn� �[�TW4�m�o�Hl�@�K&���c��6�*�@�q�ɦ֒-�8n�$�l�V!m[C����h�޷��%��V!��.����8&նw$8w�n�������m���n��n�r�u� �i-�H�pHD�U�� L�F��9��UJ�B����T�Z�vZ�*�����6�mZn�9��i˪���vX�Ҁ�O.Ϡ)Y��T�P:
�8*(����6�Znz��۳�h�,�CNSms������D��*]���Z��d������咎v����V�e�m�:8&���ۍɜ�L����ne�� ����6��l��v9!o�@ H9  �I����*�V�;!ۤz�,��y,��:].� �kh$ ���8��Am��nm�  �ְ.�6�b� I��` � V�{6�*� �E�A�Xl�9�s�j��r���\��r���#f��1,�U/k4�.mխ��햅�#m�� 6�-�GpH�e��m��l��[JKԫ�Ӝp����J����m{k8@�9V��`.�W����O����b���-�坕�=���TK2+f[@l�mB�H	2sniյ�aۢ�)<��j`W�1'o�G��ckƞ�-�'am����t+>�����ƶ�ت2-Լ��NҏUr��>hss�,�+�TYp9]6�[�m��
[Bڶ� ��6r�6���n�lv�ul� 8 knٶ�l�e�m�h�B8��d�v�pps��)�m[쏾��k�kk��E%t�   K���ʢ�E\���S,�>�,���N,̭ܮ�UT�.�^���t�R��,�jU�Bl)��*�)�p�i
g5[m��m��|��@ l 6���	 	 	 �    6�   ��Y&���)@��j�m���f��n�p��Қ�m�am ��:d�i��cj�@ַ2 �m�訶u( =J�';z�4�um�bi��cmm�i$�a���0�۶�$m����m�׬��ha3��V�ڇ�Sm[Oe�d67�5��[�����l-�    	 ж�@�`h � �[@  	 �6�    -��Ā h   Hp-�� Â@         �  �H     �i7`�l8�� 
��I�2se���Kz�)q��ࢳ���j�����"�%� �@	6�@H�m�:�&�j�"��5r� ��df����� �6�k�  @U��@,�@U��l-�S[&8$��@T�F�����HKh�n�*u�-�$ ۶�sl�Sd0H  2j��D�]���m$I]�P��@�4�B��ڶ�^Om��jD� hH �   ��  � h�	    p hhڶ �� 7m��   H  �:[@    m��ۀ �`p -�	    �  @  lH ۾�| I���   	�� $ m�!m ��m��\�a1�-mWUU: A�H�_.h�l��m!���	m�N't�7D��l -�8'B��,��o�-� �춀 	d�/׾�����I9qkU����
�hٮ��}��6��l [\����� H�6n���Z��mn�  Hk@2=�+�T�/m��UU��v�9A��%���[gv僪���yiITp��l�E� 	-��I& �Ѷ� $  6� m 8   p H [[l m�pi����      �m$ �h �m�ڑ���>�}�� h�@  ��` ��   -�(rNC�m�� �9��v�-m���\9eт궫�Z��Y���R�͔6���L� [@  ��[V��l�`    �b��%���]ZZ �ր��Z�8�  ��z�/T��RԫWU�jU�k���p 6��Q���l�AE���'��:*�ݪTbU��lH��` �m�`�ɭ�]'i0���měl	l  ��`HH  � ��H�m�   6�-�j�:U��uu++<�ٗ�*Fٴ�M��&�f��[�Ų$8�۴� m�-�� m��` ��ۤ�Ӷp�7a��h  �  	 8�]�m��,�� 7m��p>�����PY �e�M��ۅ�j�i��	 ��8a���&�m -�[��I$[�����葁X��l�;�(����Rev�z�v@-� 6�   	:� N�BF�r�h� H  ʶ���im%(��5W@Uc,I��*���$�Cm��m����NIe*��	�U��7 �:�0�m�j�-���6�Zꀮ��m0���� �     @V��s3�[��ggf�5s-@U�V�t3(��آ���
>
���Gen]�薨 �^���e�s�M�n^�rFէ7Y��+(����%[mͧ�j��]���ص�k�յX Uy�v�����m�i�h/O4�D�����R �;vH^��E�G���> V���rQ"F�'K�� �m�m�   =i[� �`�E�"v�l��k� �l@���p  m�V�N.yM�U*���˾y~.�T8�[p  	����$�m����R��uu�����($��2�R񓭪�ڞYy���W����n����U�H��ܭJ�֨ViC��������]��BjݺKaya��#�*k["�6�3b�-�l��nj�[��퀓��`,6���*�UU��nn�kv��	#U��P� kdbztK�u� *M��+��Fݲ@��,��� �n-��� ��k��`ȽQ�V��ǧM�[:�H�]�Ԁҩ���Pi��-�6�8�  �l[� ��      � �[��ɍ� � m�����$pÉֹ��oAR�쓦������f]ɦ��m7O��T��R*,� �!��Q�U��� ' "��> 	�� ���M@1���@[�z@5C@~⺁�2� �D8��C���'�=�>���������(�C�@�
��P�-O �/TS�0p��N1W� �~�z���@_�S���< b't 0u=
	�1Fu: @ ��E�= ��!�	�$BH@ �B1@DH�`@ BX�T�P��|!�E" x0���AO
	�W��� |*	��Z����Qh��!�u���_@zDo8
�=�x/���s�Z|�z=��EV�z�� ��Ț`�/P�S��ON�˨|l�K)K J��[k-���+1�P8u@}W�>���#ϑ\h,(
��`z|�H�������i$�@A�re����*�]ln��kB`����1zɪϧO/8vm�Vwf�/J�t<kR7V�l^��qf[e�7��\1�O���-�uX�h'$[,�-���n�Y��gs�����m��#J@tQT�"���JI;5cY3�k���:Vgf�Z��9�1H��{�9a�*�^�Ž�ic�ӷ+zgPFݙKk6l�d�e�]mt��S\f��F���F׊�`;k�'��X�&�d䝻q��c*�D�w�Jy6�aqv�i^�;����	�y8vU�h��=��{��&�ч]vn�V.�r��a���r�Y��Ǖ�6e}�ˬq�s�X�{BQ���r��mх,�X� d����Ws���F���F�n�43TW��lp.�]v�n�e뀊Z��6��t]�-��nI��=*�>յM���r4r7��U�4��{�wU�����;<��N��nx\�r�L�Z�0� Z�86��kn����d����r��r��k��4�.pi��vۑ�jU�8i��5*�j檍J�Sr�bmp $-ڶ�dڥ��n��V�EJ��g;��m#�g�nqi�mh,[�6��[��x�(;�kPڤ)��)��*mm�Ҁ�T�6�� ��]Wh:��-�6������6�7� u�q�\�l��8��m���b�a�X��bP'�T�4UW6R^
嶺@�L��jJOg��m��m���ֺ��y-���8�]�����%�)�<9� ���B�9���ʜ�.�D���g��Ve�3/3�0r�t��#��� 㵸\��A��!nEK�v6�*���7��b��닋���pRY�*�R����r��Й�8wRۗ�6��g<n͓Y�d�+�ni]t[%m���lPU-���IV�>m;7(b��X"���۷Hm�!�`���G=�J�QkE�U��̨�����8j�d�U�\��L��sw%�.i� ���45"1B �����@�E=�>����Qt�WN 5F ���ܛdٶf�u�b�iP�%,����ҹ<7c����n6\q��,ۣ�l�:6����v�۷]�q�m��+�.wB@O\�mn�q�#�.C����tt�!ٲӰ\� n�
�[q[����G$[&6�����<��evܧ�����1�����N��4cF�'1�c�wE��8�;�։���`eSFl��v˻nl�(T_��p�>�>m���`{������An �('vx�g�{l�8U��1�x,16Q8d*�^�w��w�㙙����@���65#�1�Z�� 7y�3�>}x:|�W��;�6���$R7$��f�ɉ�Jcz �����>(�^7$�M�Jh�W��� ��h�.P�x��Q�Hh�W�.hc�&&�D�7���d�j�ۤuΘ�c��Y,�L=�!&4�� �*p=�.H�Ԏ!�L�� �)�_u�޶h�)�yzנZ��I�Ƣ�.�R���I=���H����� ��E����s��g$�����$����n�hIdĜ��JhLo@�	˚�V�^��T]Z�U����H9�� {�x���:�oG����h�R= ���4�MS�9���f^5��"{ d�]�Z����m0���@���o�)b
�Z��֤k�������q4	Lo@�;��]>(�\�n29$z���9^�@���������H��.|iF�#��*����'o�w94S��X�� y�����v�h�)�r���crb��
�Ve�Hށ�h8��/@���@r6D�m"H����q4	Lo@jF��J�՘^f�v����*&�
���lnm���s���W8.҇H���m9���"iŠ_YM���
���:��@��Ճ�iAujv`��Ή�H��V ��,��h�[Ѷ�$�%�H�z]ΰu�aЗo_\���mRqP��48c�8����/�����{'A=PqF���h��Os3��5w^��cƮX�1�F�@y��%1���#q� �z%�4���Yό���N�u�7M�k���x�S-�Vv2���ۗ,m�3�=mt���[�l����Hށ�h8���8nD(�&E#�*�@�����h�W� �["cR'�4�z�ƴ8��7�5�	��~*�:(��WV`z">�0���
�נwYM�mX����x��bWf�m��11=O�� �vF �ۜ�x����T�߬/��J]��^ҫ�.��q�u�8�W$�u�Ԓ8�&IwM��C�L�Ԫm��]�h��zL�0q���-��'J���lpP�c7���Z�.^+p��&��������=�=k1���#���v�'F�n6�Q���`@�@���v-V�F38��C&�'���Mn\����΍�Нu�ɝ93�t���5���i�*���#!�?������}�6g]��n�ć��vn;z��hla8�e4YAw��LR�*�4�.:��F9"��/��@�s@������ģ�D8c�8��wۿ�C�&�+���o@�r�t�W��c��R����mz]���)�yTw��&�⌌�C@��o@eƴ	.5�<�hSM8�j'2dR=���j�/����mz�33����<qG'�!�,Qd-˭��f�]�����I�u�/hM/0�Q4�q'#ME"��}e4+k�/>�@�<�x�u��p2(�ZI�{���z聏��> M9�����ڴ��h�ڱ���	H�%!�~Vנ^}V��Қ���/Z�kiDI!�G��g�����-��@����mz��j��Pȉ?�#�@�>�@����z����쩹$Q)����Ǔ�8��n�:�ʄn�4A��.�F;^�vآ��q!�77�"�/����z����^��U��M&HG!�y^�~�����H�O� ��V �v��ѮI7Q�xӏ@��z/Z�k�+�J�z+9�wy9$����I;��v&6��NF�(�Z/uz�)�~W��/;V��y��Ҁ��
e�q4�����WF��?~�ֈ�)��a�s���Tu1��x��c�7:'�DĆ�L�mO3��
N
����Zց+�zMV�5���DI"��u�~��H���h_�Ɓ��^����lO��JE����̽KV��@��o@j-��p����1Hh����w{��v���$����z(4߷��Q�B!���B9��&z�u~�|`]� ���uV��u2�A����=t�8̱�5�5��t�q����5#��W!�kQ�\nV6����K�h8�ԭ�k�^��vwUp���u����L�JGo_/���wW�{�;7Y�b$��4�M�V��o@�bhR׏rDĚiH�%!�~VנU�^��;V�}e4z����qFIwuu�5�� ������|`/��6{�����>��v�=sy+��������r.jm���x����[ρ�q�9����6<˳�kҪ[fJ���NQ��,�W�m�4n-�2Y�ϗ���[[`��u�Pr��^x��t���jX�i�nb��:9iNN��R�:�̠Gl��p,dYY\��$C���2�D�Ӎ���*��5��]n7]~�﷧��nh��u�i��&&(�{����>�w{�q�5L�6V���S-ݻ�u�t�pؕ�pv5��q��vuL���5z������@y��:�o@eƴ	�]�����"�/����z���wJhUL&'�HG!�~Z�`kZ��)kw�����j�T�MĔ�q��U�{�U�_YM�]k�-vȘ�y I���X۶��b"&;{8���V ����m�ϧڦ���=�n����\��iɛ5�aC$��v�2Eg�H�������uUf �v���� {Z�L�����=����iE
C@���ϒ(�@ �(�g{�����{4�)�wZ�7��D��E#�,�ց�bh8���	&]�uB�6�,hiǠ{�S@����ֽ�����° �)?��Ԇ�}q4�m��5#zI���r�v�5��iЎ���뢒*��s��ͳ�7�3Fn9$:v0�������lO�����o@�14�M�)ˢ�b��cN=���wJh�S@��נZ�Ȇ�yI��#�=����'}��rzr|#�3� Ԕ�V��������x�|���T�t�B�$H,-��ꯤS�	�	X�#q�}}S�E����>,����֐��A� @=�h)?�<~���=�����o�@�<�x�?��Ԙdm�h}��﷌��� ku�B���;�+"�45�H�$�~]k�>ϝ�?�u�����fbf;�%��Uuj���]������뛧��C���g=OR�-Ź��ݚ��'1���G�?���@�t��}e4˭zwF�i��Z)U���=3>�<�~0]�V ��z���M���?���/����u�@�����s@�����Ƥ��?.��wW�{��h<�fg�C�1� 7��������r�[RbSiǠ^}V��=�s@�����P��>rH��H�&�OS�JJ���rD��n��c��6�6`㩉�0��E2'15"�?{��}n��ֽ�����I�ț�m�3@��}�uE���:.�@�����ʄ��P�*��:v���Ο,w^F}n��jkP������/>k@�bh.�@���I�m�Q��DŠw>�@��s@���@������Idx�����575cmngB2���6mep��s��y�����H&3�bNs5ֻݱ�o1���i�Wy�ԗ�f��ݧ���vvb�pX�Ggu�n�G7.���ѡcSl�J�`�t�ϗ�����1��+��� ��ݠO=[2ږ1n�c�������,Һ[�a��+�[��D�X��s�������n�p�B�-�m���{�������TͳSn�ki3�%2�.�Y�v�]�;��]�Tn�irL
�&��.�x��@�~���>�o@eƴ	R7�u4/��,���H6�h����U�r�@����˕��#�9�&����T��8�ԭ�q̡'�y��$z.���b_w��@��Wuz��أ��ڏln=�@�������cC��4�����q��VA�����E�<AKj�۫�7Z�T�e��G�
0��X[���n�b"? ��� ���=y�%�Ǡ^}V�bA����l�>Z�gLLBCn�E%
␮AUk 5�^ �v�*g�b`o���}���@�]tm�DF�I�,�����-��ց�#zR�piL&'����ֽ������F����˰��U�{=lV&�<��y$[������!��y*P�R5�&�sm����-��������^���}��H�����R/�uw�_[��~]k�/>�@��v;#p����"iŠ_[��~�w����(��#U}�w���ՠ~�{��5�l�,I��?.[�>f&�$��'G}�H��U���X�Q�z�Қٟٙ�mߏ��U,lw��� �`�`�`��~��8 ��{����?Т�*�r�yh6\�n�q�]m��x� 乽�dF*i┹���sg��A�A�A�A���?�"b�`�`�߻�Â�A�A�A�A�?~��|�������ӂ�A�A�A�A�����37n̻.M�%�8 ����|������߳��A�A�A�A��y�pA�666?w��8 ����߉�r]36]ݙ�� �`�`�`��w�����lll}��~�|�������>A����w�� �`�`�`��~���,&e۶�ff� �`�`�`��������lll~�y�pA�666=���8 �@`9���8 �߷��d���sp����� � � � �������lll{�xpA�666>�~�>A������ׂ�A�A�A�A������\�3wY�hXM�˹
"6�YN��q\�ɶ�P�2݃�J�At���������� � � � ����>A���߷�� �`�`�`������� � � � ��y�pA�666>�w�g�ۻ).Y�ini�� � � � ����x �o^>A�����ӂ�A�A�A�A������
|�� �l{����[7n\�ݻ�wv�A�666>����|�����w�� �`�`�`�߻�Â�A�A�A�A�����A�666=�y�3�L������� � � � ��y�pA�666=���8 �~�߯ �`�`��������x ������.n�v\��]��� � � � �������lll}�~�|�������� �`�`�`������� � � � ��zv����ɻ	����Ĭ�F�6dV���,�w�V�}�	K�.K�瓳�L��7�g�cy���*ul���n�]�ٸS��qѣz�'=g�S��]cp4��^�xWS���N{y{"n@P��a���q�Kqm�6���nö�k�ƻq3q9�S��8S-��.���*d�n:Ԓ��Nz��h��V�^"��L�]eƴ,��&���g~"��f��O����w�w2�pq���<��v�4��5�p�ƥ'�6�ɫ:u�7rf���Ӣ�A�A�A�A���?��� � � � ��{��A�666?}��|����~��>A��������3wmٚi��x �o^>A�����Â�A�A�A�A������ � � � ����x �߷��ٙ���fnn�v�A�66 _��?����Ϫ�?W�h���ؔ��3@���~��s�-��M��}��=K�{��(�#X���w\k@����kZ���r�囁d4u,ݛ{��,�1ggvvZ�u	e����R�Ŧ��T�I��o�bhu�h���:�ށ$˺|^av�f۷vrI����x ~��g��~���Vg�|`-���f ��Q��s$�rE�w�S@�2ק�X����@���hTZ2`�1���@�bށ�14���N���#�Y9��c�@�zS@�>�@�t����k�<�]�Q���H�>�[��Egv�بm&;h͐�k��:��:�i�"ci�q���ㆁ�fu�|�zύ��_��}gƁy�g�8�*����V��m�鈙��U�{Հo���@�>�@��V��Ģ$��Nf�hn��m�d�LL�T����Zց����;�^�&��"��(����Iq�tw����_�@��u�$��G�2%�������s@�Ϊ�ץ4A�;$�E����(����i��l�
��K�&��Ҥ�~�年8�x���/�^�nh��^���������ZTddA) ۑ�~�i�rG���|��^Ft$|�/�d$C����j=�Y�w>�DD�f*���0���`ֺ.�UJ�ꮮ������M��=}��~�k��=��
|' �$�:D�E@�����o��rI����3e�&l�t���k��=3>�����|������ ���H�$iH�?�"�u���k��nĜM�k�뷷g��N��j/�{�w���(�(�#x���W������mz"#�?Ps�d`�z�\Z�E]��.����:bb��=}��{�U�ٙ������'��dȲ%���w,~�f���Հ}���5��ʺ-ET�*��Ļ�8�5�.���fD�Bn��˺�⋊��UՕWf��N�zbb7����wW����~��I4�F;*F�}���@�) �I"��� ��p�S8 z�
��BF2�(��HH25م>d%�\eP��pĹ3.e�`�����A�Q��B�B%
Z��+
BI!,,��j@�F��$�)�4�W!o�@"$�s��b��`T�F2�ZE��H�$�	!!�S�C�#F%H�%!E��āhB��(J�����
�X���*V��#�D��HR�I
x]�BSR,e�B����J�#
++K	(�(Ɛ(KF��a!d	X0"ڿ!0�PXA�*�b$H�, �P#X"�BR!A���,HA#RT
T�+)J��"J�IP%bD�"@�e�m*B1bA�	$	 �=��{��� ��_U�[�ζ�����a��
Rkv�#��M������Q�n��Q���7[{^Âg�5���E�N�u�y�N��p�z�&��:�s6��n�n�N�x�{:$m��"�qum[8������)(�K���'V
x����H�o���D�Cn�]���U�x7Kl;pY	�ଋ�ݱ�0p*�0ji�Q�v��]���p���"`qn�Z��q��ywK-R��y8�n_!���1��W�S�ޣ���{"v5�=3�����NL�6��<�;|����n�ԫ/[�8�sĔ�te�۔-J�t�υ�-�����셬T�˅˘����xi����$s��W��s�d�&8k��v���v�v�յHgGR^�촓+��s�.��y�mu��mtlK�@,v�-��dM��kgaseu���F��T.�l�I#�w"R� -&�8�0\l�TA��@�Y=�^�6�me��ݵ�>^�m�6�ջ�[����N�������lM��6� ��RZ؍h�ٕv�&�ɧI��D�p��^Α�Y��&4���:���u��.�ղ�ۮ9��:�h5�l��55l���ȳ���d���/�m�"p8@6:�gp�
�3�V�RW�w]{|���o��9�$,��_>Q���8Mv�9d�;�3V]Z@��Z[�����Ѫ����k�`Ba��f�.y�� �]k�vgx鳇b�۳�뫄�e{	h6e�9� ���2�+�Z�N�,���R�`��kCm���v����; ��m$��WGp����O2c��h��w$�4�`��_ɹ4�u�� �R�k��h��Km(���ϷE�\��*b�\h�6��6�a�V�a����p�*Ym�۔�UV�nu6����yN]�nD�zA�e�]��	�l�V�q[p��v)RtTi�q�I9�5K���ٕ`%���j����3$��&�(�W�P�#��Hj����?-�'
*�;5��{u��$��h�0X�ۦ킐��7F���l�Z��ǝ��7<˹��R͹�v�E���D���O�S��[Y��a8�Y��ϱ�sF����mNNݰ�;Pp��V�g:�I۷U�,hx�96�JY��c��R�&��-��_��*���q����7W^[-�D���g��
y�Dmt4TI4����l��%���ﻻ���r��<�.�P�Y����6u���o���4<av��R��w���#4��BD��>��O�{�k ߶��?�k����}B-UuuwV������L��"b���� }G�X�Z�tD�CڇT��b�*.�]��0���zfj���X���h��^�LD��G�Hh}���ú���,��L'�8����dM�Q�G�~���>���w��/Y�w5k�?{�Y��$�8)�b���;��c�2�n�tQ�d�7)�D�vN-S��~Z��M�&4G�)_��~����7i7^���A����<�yE\TYP*�S����~��@Gj4d} %�f^נz�V��ֽ�ZTk&4�Lq�w�h]-�7�	4	�@����a�����@���m��+����;������RG6�Z.����/5k�?W���m�ϧڦ���>�g�":�e�\���f�$�n.N}�3�H��R�]�ȉ#�;�)�^jנ~���333�~��W�	#1�����.�n�ε�]6��m��11��U��(���G�)���h]�Oؿ�33>��-jנ{�&�o&4G�ӆ�ʿ������-uסؽn��Z��`��y$q�������?wJhVנ\T���&���M��b�u+�:�[4��;�m��g���n�3i����u��k|�}��[�>n5�JV�	�@�Ԣ��150�8���ZWj�;�)�Zկ@�ۀL�IY�h��t��#t��|�k@�~�t�@�<Fԋ@�t��ի^�����"��D(�����lw,��"��wvT%v`�7XL��o��;��-�Қ�Ԟ�"���$mm3ٮ!s��!���k�S:�R������-�$��Q#��R=�}V�k�h��:�k�=�J�k�bȲ%� i�脇���R}X���uX��1H"�M�ҚV����M ��hZҬQs$#�/0��7�|�M �s@�14U\C�Ƥq��JhLB}��z��M�S2/���v!����k$�/\��Z��=���]J��t̈́*�N-[.-\��z��.��9\In�=����^sɍ`�v�)�S丹K�tN7e�t�5������ ��D���:	�M+3c��3�χl�]���0��KZ:��MUS<;A	�ȯca�Kb�S<9�n!d{����ێI���m�[q����<VpQ��[2I���ݻ���7�4$zl\�Qgl����8���땓��[9������&FE�r)#����>^�=�Қ���DD�L���s�0��qh�j�QtU�`��3�f"R���@�����]��%0q�X������bh+z鉠}%7�(�x�p��G�~�)�Umz{�4�Z�wDв�2	D�5#���xDL=y��R��k�����i��Kn���^ZQqS��Şi��,���v]\�t�Y0(���%I(쬼�t��#t��|�k@"�@�֕b '2L��h�k�ɉQ�%uw, ��wm�鈘�D�Q�ˡ�wUvQj

���7��, ��xtL�M�� � m7V�
J���ժ�V�?G�3v�� ���7N�`z&'�3��y`�uR�\]RQ<LRI�wt��y�^���V�˭z�ꇱ8��@bX�BBY���4p+&��DO0��j�	�����-��N9�m�ŉ8~���=�v���]11�6���Չ+�t����TU���?:mg�}1TwW����M�t�F�j����J�E�]ݬ��גO��{9 �0D`�M�����rC�|�
�ռY�$Q�!Zb��&�� �鵁阘�W>�рy{�����&'0�f�W�٠Z�Z��Z��h{/2�䄄F5#k�ٶZ�%��̻��v�b^�v�Q	L�xf3O�I5�nM�j�=�j�-�s��>V���Z��4!�)qRUk �|�g$wwd`����mg�'�Cu��h�����E����{�R[��ց��zzA�e�^*Ut�*ʫ����u`�ܰ��k$� 1�
~'�~���'~�����kM��x�q��V��t����s@R�X�&w���ڻ��wt*���AV4��h�K;�ۗX����n,��[�����}u��E�rE�>�O�wu��/��]1��]� 寪��m+��T�.�\`��3�R;i>���o��3�1鈪<�ԗ��h��v]����K�X�M�=13>������;����C�1�0iǡ�b��~��@�빠Z�W���hCp�9"iU�]kXL�o�G�;�>���m�����߿w�9��n��9]EWa�g�=sغ�.��	x�{h"�;��g���vr�c�B'�v�sg/RϮ�s[�)��'7-�T^2!og�\�{8훮�҆�@�+��l��հҎ�@�d�7m�km��"p�&k�9�؇:�M��Df�5�ˋ0������|�v���v�b�ںO��ۤ�������d�rH��#FX�p⣘������8;��5�x�����@5�X)��peT���{���F�<t#v߿�������Λ]33�>�� �ά)E�ʥj��+������&R>��_�?�w��Xo�0�]V]�J�EU]*��Wu�~t��5�kLL�����u`�uHP�E�ڋݬ��M�q�6�# {I���Dz&f���,���U
,����U�v��yDD����}�ܰ[��L�DLB��q]UN���8��sdv�8�:z3�Z�������l�۬�L�N�i�V�de�@��$<�{Հ~t��7�ֿ�#��d`._�_�L��Jm�2�����{x�����������G���X�����k���H>�|�PiȆ�M'�y���7u�a阏LLU{�w� �W����j�B4�pǋ"IŠwu��/5���6�:fS��X�uaJʹ�V�.*���Z� 虏�����r�7u�f�����}e��H�p�4�F��hꓵ������ 6���iӮk.�T�w{����v
�J���.�����oխ`��=11����ɮ���uHP�j��X�2�	&&�$w�]K�ͭo�{ؑ�:�LY�rHI���o���Mq��� ��� �l �Փ�(1��|!&	�`X�`�$� E���H�F�4��$bH�ٖBR6�t_\��I#$ OD�#�0ID#$dD�&�!$I �� �HEH! �@������'�S�G@5!�#��`E�4`�8��)��cNtCE"� uGA����QJ"�����<P�3LLODB���`��4����
슫������]Z�� ���`�t�;��h�\ڠ"d�E�NM���-�������r��x�����+^�P�ݍ(oi���m�a7C�e�b!�gix�b����:�aUU���]��Xo�0�M�D��>��?��hW�?�pɄ�Bcƈ��;��hy[4�ڴ^���Ď��f5��U]+����� ����6��JMm��߷4���B$Go$RM����u�n���ؘ���f
w������+�I#�A����^���s@�ˬ�?Wj�/�m�� \�o=���O&�<��ͽ:�m��=ni�˷g"��M�LY����mH�m�s@��٠~�ՠw>�@��ITLQ&�E#��U�l�?Wj�;�U�wu��?*��1��Li94��Z�@�;����m�����h�mcIš�V����I[��RIW�l��$�ݭ�I.��v8d�C!1�Q�~��K��5$�~V�ߒK��ޤ�����ۊ��4Z��J
�E�H� ���S�ܹ�@�-�M�z�nsZ�#�]�Ԓ;C�ԍ��鋣I�w�4�/D�y����LM�-��V������S\���v�h�8�t�<Q-����].�:f7l�l���֫1ݻ$��M��&��q�ҍ��������`@�6Çz�t�8�
v�s.��'#��q������Tݢ]�p�7gu�L."���i�5̂y����xK��-Onv��s�N6ݜf�=���צF��Z_�o��雳���	]��Iz��_��%�SuX�I��?~I%�v�K֪�,1!�7��OߒK��ޤ�����$��I%Yz�ߒJ�BŹ�I2�ޤ�����$��I%Yz�ߒK��ޤ���+J8
B9�9��$���RIWWY��Iy�[Ԓ]gU��IT��+��OȜr�J���ߒK��ޤ��:�ߒIw]���]���RI�)$1���E�e�N�g��G���W�d���}�K*m&t�F .cc\�X�_������� �w]~��Ku��T�����$��Uw$uS�2� ?oߧ�������A��a�$��[?~I/7kz�K��[1�C<J'��$���RIVz���Iy�[ԒW�i��Is�$x�1Ħ<���ԕ�m�׺�^n��$��8�I|�u�I%�|���!�7��OߒK��ޤ��:�ߒIw]�������������f*�%qq��(�ݶƤ�:�Dۇ��c��^Cj;+��8�O�w���c�r]D�7#�I|�����K��5$�g��g��\��7�$��b�(�9����$���RIVz���Iy�[ԒU�}??��S�~�����..�k| ?�}��������r�!�"*���<�Go���]��I%��̱$�8I�''��%��oRK�uz�l����1|�}����"c��I#ȓ�@��� 蘕���嫺����?@����Y���Gn�����۝+�9��Ab��]��Ǣ�ț��Ct�%����������������{���PFߖ�ˏ�č���L2bRM���z"5ou`�r�������˫
 $�<�94/Z��)��#�女U��4mlI-�iL���r=.&�w.hQ�4>������̷o@������"s�4޶hs����.��^���X�pj9,��!��Xٵ6$�5�ȍR�u�:�3�r�=�vh�-��F�L��1L��'�*����>_7X�mzf#�w��\�u�$�*­R��Wx���;�Gz�� ��h��o�ؐ}��E�7	$yr����@;�4	C�:�o@z���.�V�һX)n�^ ��׀|�n�:e>��jӫ����B
�"�+��5��=�����ܰ�{���4AP����\(/��G�o�K�H�7�cUIVꪕ.��E%'1c&og���7[;n��f��]���c��,d��v�G�8���s��MY-ˑ�M]����`v9ț��l�;E��ڠ�rˍ��H�MY�7�����P	�m�z��Sٞ��Uʸ^7[�qpp�� �cu�;c6��I����{4z��D���rv@���4	]�bY�n���ww�L��)�bCm�'U�Rn71�h��)�C���j�0�eN�{|�o�V�Д7&�'������րw.h�s@U�*�ٻ���UeU�`�k:e ������<�k߳3*�b�E�MD4�6�'�٠4+�W-�q4��(sqvX\\]���D���u�����ف�1阉�o޼�.�+m8&����<�k�/;V�{������/c�I O���!�⫇ʇ���qW��������(^�����j>|�蔌Dm`)'�>�wu�G[~��D���޼Σ��WH�V����*Wk 7u�\}3$K��"ۼ ���kY�	1�ͨ����J���O߳@��������Ԯ��+�]��YWw��+k{� ��V {������[�k&������u�zan�_�9�x����=߿�)���=Mv+�nn�jC&�u��OnIؘ�rm�����4,�T�ӌ,j���f^�w.h��urހԋ�-|в�L���2I�^V��ֽ��Z�[4ʮe�D܉H��Iɠyzנw>�N���ٟff��|���h��ē�6�xګ�v�� ��� k���t�L������V�q#&"7$��qh�l�9y[4/Z�wJh�䝉��鍃��F��pqZWpm�n����Õ�\>��d��/���|�z:�v�ۮ�6�O����:�o@�14�s@�M�V]�co$��jI�yz׿bE���@;��hr�4��$-�#�j,��=~v� �����4��[�X_i
�$rDF�������w�M�U�l���{��1}	A�:���y�^|в�L��
d�94
�u��}0�����~0 ��{��P�]�#���T4f���l�R�
�ns�	�/^��L���+d�����7�l��n�b"? ��������AwbUU�]`�kY�D�U~��Mw� �|�g�f%!�C�UЈ�E�]�$*������k�=	j��U��yx�E��2bNM����>_7X�����Kw���_h�q���H�5$�<�k�9zנ|��j�x*"%}Y$�r$bH�1��!b�)E�b0b���@���#=��{e%�R�0$��#(Q�#$i(��������DO��# �
(��@X���a�`DHD"F@ ,H,XF@#) E�B@ ��bń`0c"�b��!֥� �0#!�[5HJ���98���'jъH��f�Б$!I;ӿ?�?�������:��i��`��ѼZ����g�̜��ǰ6��cN�sZ	Ӹ{f��s�6�nϟ5to;���VQ�X�����=X�vm��ڷ�p�t�"-�U�%u�)1�m�v�В�%`�S�*(
�&N<'L����@T���T���`\<��	�=�O2�Z�Q'���m���I2�X�+�d=VW!�vÞnC=[�b��c]��K��m��˭�U+�7�/��3�7t�\�ls�A�8�wB:�r��/�+rc\�b�x����	�'�s��̽ڸ	��u�95���קvv���YT�8gR����p���e�N���v�ע.�J�x\��!���4��U�s��P9U�Q͕kHt�A��c6:�C;�,�8ᝤ÷���8s�we�u��řc�,�s�1�o2��ؼ�v�g���l�	z�.)�y�0,GR��3�c��i�N��5��-�JCc'sc���uÓ��@�Ù;-W1.�=�ݻ6F��<kG �PU ��n��$�RM�6���jؒG&h��[ӯZ$�X.V�X%ж%�vuqG[6MrݭdM�f����vmg�u��&%�=UF��V� n�J6*�
U�[�i ,b Sl�V���jy��H烧��dݍq��m�T��t�� �77Y����*ԻN���
VM�͖J H��jmYN�X-u*,���g�s���z�	ڎ�<����I�K�,��]��5g��2)m��I�A6nUy�[ex;ez�+Cr�d�V�S��m.�r��^5��V';�m U[q:'�;-o'cg0
1�³�+�U�y�c�<#�tu"0D�<�G(n(��<��:Zyw���u����:*�*�LNGnZBz��WV���!�M!� �+A�Gp4r������ب-�y���Su���8��l�V�Wd�V��W��L���=��B��W��_���*�v[!�}��#�ݶL۵\3vtLV�֔�CT��l��P�SN ���q�:�R�!6�;`����'q�si�AȎ�j#��\�0k�Z�i�#�r@�6۶D9gVĎ�qg�j�Z�HR��sbK��nգ�;Ev�v�=l�x!oН��)HU�� rG6�
cv��؛gD#.�֞A�{y��i7����q�-��nf�0�����|��QT�9{�����N�[h-�M
�K��޼C�]#c�����/��܍�5BI�~���l�ծ�& սՀ}ԙ��+�$��2�/@;�4�G4�[�:LM�?�c�5G���zn)Z������� �׽x��zwJh�l�?*����8�cIɡ�b��|�oۚ�[4
���|��!)0M�i8�鉠˚\ۚW-��Q���W�ջv;uǞ ���(8����k����c��`@�N���>R��C�p+oͱ'�٠5͹�urށ�bh\6���e��[���v����'��&&`��!Pj�u�kv� ���=)���S����I#��@��|�w[0�F�u���� �ڡeUU��@^^f^��bhr��-�\��~��Y�S�$��' ���^��^���U�v\|�㑎Ll���TT�w�Ĕ#�ury�d��ݜ5�\m�ӌ�)�LM��"�M�Z�/Z�^��g�w�Mʫ��<�I#�*)U����Ι�H�}���׀j���$��X�Av�)*��7��9$����&�W�������$�������#d@D�I��&h�l�$�����c��:�m̿�(�'&��v��ֽ׮�{����'\�@�҉(`�K#��&ۮՎ��9��[�A���&n�d3�j�Mi��TuY����:�o@�bhr�+��������?蓒=�Jh�l�*��@����ٙ�����2(��X�� ����n�虔�O����-�R�	�H���h|�`�n���`�" ��"I�"B/���� L�G���g�����yyv/���qȒcN=W-��րs���z��Q0������è�UuWw4�X�
���l�^�=q��Yc���)"�\㪤G� I�&�p̹��{ı,O���jr%�bX�����yı,N��܉Ȗ%�b}�����%�bX��}��ݛe�nn�nfl�Ȗ%�b_{�w��? ��,O��ۑ9�ĆDȝϿ~�'�,K����֧"X�%��{;��wsm&L�.f�Ȗ%�bw>��ND�,K����'�,��2'��~�9ı,K����'�,K��gs�.��pɷ7�܉Ȗ%�b}�����%�bX���eND�,K�߻�O"X�%�����9ı,O{�ܴ�&:W)����Ȗ%�b{۽�9ı,K�~��<�bX�'��w"r%�bX�g��q<�bX�$/WXN�ې0�K�vn�\��e�mZ�Uͳ�uJ܆{@]��,�"v]���;ݰr�\k���k�v����nn�u���0r����ݷ���C��״cv�p����
�IE���� yB����Rj��=��m��L�;��D�&�k=��9$�s�u�)xM��i��)����4��]H�-��GQ������@�ܗ%.\C�������|�Z�\��vx<��cm�9n�;hܨ���r��Ͱ[���,i���a�%�~'��u�b}����yı,O��܉Ȗ%�b}�����=��,K����9ı,O߻y2M�p���ܙ���%�bX�g{���P#�2%������yı,N���T�Kı=�{�ȟ�{��w�������gvh+;�Ȗ%�bw;��q<�bX�'ݻ�S�,h�lO{�u9��{��I�O�����˚��I���y�T�Kı>���q<�bX�'���D�Kı>�{��yı,N�������[��oq���{߻�Ȗ%�a�T����r'�,K��}��q<�bX�'{w��"X�{��?�����:��E�Y�{Wc\��6lnۓ�^|�c9�nr�ɍ��K5쓵��O"X�%���w"r%�bX���q<�bX�'{w���� �&ı,N����'�,K������-�%�͹�n��ND�,K����'���DȖ&v�eND�,K��{�O"X�%���w"r'���,N������J�6����yı,O߮��9ı,K���<�bX�'s�܉Ȗ%�b{�����%�bX>��Y�&��,&빛jr%�g�DϾ��x�D�,K����ND�,K����'�,K����Ȝ�bX�'{���Y�l���������%�bX�g{��,K��G�����{ı,N��͑9ı,K���<�bX�<���������62Q�]��);vt��+�\p#��|�\��c๻rT֡ⳅ�2�33r'�,K��>��8�D�,K���"r%�bX��{��yı,O��܉Ȗ%�by��d�s$��l�̹���%�bX�w���,Kľ���Ȗ%�b}���ND�,K����'�?�Aʙ��0���vͶ]���]��"r%�bX��~�'�,K��;�Ȝ�c��1�/�p�&��}��q<�bX�'�xT�Kı=�gp黹6\��a�����%�bX�g{��,K��=�s��Kı>��ʜ�bX�%���x�D�,K���L�t�6�ỻ�9ı,Os��8�D�,K���S�,Kľ���Ȗ%�bw;�Ȝ�bX�������+T����Kl�n�]�NJc�D:�.���̚��O11)��pv�nn�q<�bX�'{w��"X�%�}���'�,K��w��9ı,Os��8�D�,KܿK/]�nm�f�ʜ�bX�%���x�C�� ��ؖ&��ۑ9ı,O��߳��Kı;3�����r�D�?~��|�ݒn�-�����yı,O����ND�,K����'�,K�����r%�bX��{��yı,Os�,��.m�˻�ffnD�Kı=�{��yı,߻���bX�%���x�D�,)��H�ϻ��,K��=�gK�sn�s2��Ȗ%�bY߻���bX�%���x�D�,K��w"r%�bX���q<�bX�{����M:���d9�s����k�2���N���Y�t��d;m�C&p[SngR����Kı/�����%�bX=ϻu9ı,Os��8�D�,K�~�br%�bX�糸t�ٗrLٔ����yı,�ݺ��bX�'��{�O"X�%�ٟv�r%�bX��{��y�2%������wIp�nnI��S�,K��>��8�D�,K�{���K�ș������%�bX?���Ȗ%�b}��2�xf����ۛ��O"X�%���v��Kı/�����%�bX=���r%�`~@	�;�~��O"X�%��^�/�ۅ�tٻ��"X�%�}���'�,K��w�S�,K��=�s��Kı;��ڜ�bX�'�
A9����}�羦׭����
6�mN#�M�
�ݺ���k%m֌%+���۵�	���ցmNqg�+��/���N����i�=,��ޛ#���ۊl��pώv$vٵT!Z(
�[��:܋�W�m��9h���L�J&������t�Ș5=˃�*��W��xlUǩK*gA�<��q�i�3�4���֖p�>���>d��m������9frΞvuڥc��ĮhM.]���[�MZ��.�-�j*��~oq�����w�S�,K��=�s��Kı;���ND�,K�߻�O"X�%���M�n��qQEE������ow�{���~�L�b~���*r%�bX�����O"X�%���n�"X�%��v�:nl�	����˛�O"X�%���w*r%�bX��{��yı,�ݺ��bX�'��{�O"X�%�}�~�j�M��Ow��7���%���x�D�,K��n�"X�%��{��Ȗ%�bw>��ND�,K��w��2�6�in��<�bX�s��ND�,K����'�,K��}�ʜ�bX�%���x�D�,K��~���)��F��yZ�]O��G�Pr=��KRWE:��*pե&�鷛�$�۩Ȗ%�b{�����%�bX�ϻ��,Kľ���Ȗ%�`�>���Kı>�{�a<7fa����7w8�D�,K��w*rLQ+�2%�}���'�,K��}۩Ȗ%�b{�����%�bX�϶���]�]�w.nD�Kı/�����%�bX=ϻu9ı,Os��8�D�,K��w"r%�bX��׷�v�77p��ݻ���%�bX=ϻu9ı,O���8�D�,K��w"r%�bX�����yı,Os�,웗0�f��۹�S�,K��=�s��Kİ����~�Ȗ%�b_�w��<�bX�s��ND�,K�&{߯�o���q�(�uޙ{n�@��1О�V��&��Rd�M��LTl�=�bX�'���9ı,K�~��<�bX�s��ND�,K���Ϟ���7���{��_�u��pU9ı,K�~��<���r&D�?e����Kı;�~���{"X�'���9ı,O�����̷M�f]��'�,K��_����bX�'��{�O"X�}M!�HBN��5�S���ƪ	OK�� Ke��7rYi�fuҪ�@���0�� D
D�u�g!D�X@����L=�:)N G�_�q =N�A=A�$�Q|�<=J
(�zX���}�"r%�bX�����yı,�^����7,��s7*r%�g�� ��?s�����%�bX�߮�J��bX�%��wx�D�,K��w*r%�bX����g�inə��nnnq<�bX�'~��Ȗ%�a������~��'�,K������9ı,O���8�D�,K=߿�)���<�S�\�g�s�lf�5��J���a����L�PT*YI꺭�ܻ�S�,Kľ���Ȗ%�bw>��ND�,K����� ��Ȗ%��;���"X�%����?\�n�sw��ۻ�O"X�%���;�9ı,O���8�D�,K��w*r%�bX�����y��L�b}���fbK%'����oq��_�����%�bX��gv�"X�%�}���'�,K��}�ʜ�bX�'���鹳2I����˛�O"X�~BD����S�,KĿ~���yı,N��܉Ȗ%��8,t�/6'w�w8�D�,Kهs��n���f攻��9ı,K�{��yı,N��܉Ȗ%�b}�w���%�bX��gv�"X�%��w�s�sn���݃�F�W�nϊ�<�9$���{C��乤�z9���2s����t�iww|ObX�%��;�r'"X�%��}��Ȗ%�b^߻���bX�%����<�bX�{oy���ْf鹻�9ı,O���8�C��"dK���n'"X�%�~����<�bX�'s�܉Ȗ%�bw���Y���wr����yı,K���'"X�%�}�{�O"X�dL��?~܉Ȗ%�bw;��p���2%�`�/ad�\�6�K�����bY�@ș��߷��Kı?gnD�Kı>ϻ��yİ?�Y�3�����Kı?~�����&�6��ۛ�O"X�%�����9ı,?�#������%�bX������Kı/��w��Kı8b��=��m��Rpۇ&����-t0�k�nţ;*��Jx�G[�x���fQ�p�rv�g�d�m+�^��g��Z��*���i�^.[��mg�x��mk �('FzK��*��݀G3͍�y�e�C��e��ΕT��x���nθ74Xٰ5��	�6��z��=<�=�X�^��� �ևtv�u�:X�f�}�{�������ի\fd�5teg[e�V�ѻv�Ϣ��]���Յ������E�I7E�����,K��?w�q<�bX�%����Ȗ%�b_{���Y�L�bX����'����oq�߯�����{i�J��O"X�%�{{���Kı/��w��Kı;���ND�,K����'�? �n&ı?�ٟۦ��p�攷wq9ı,K�߿���Kı;���ND���DɄw��gؖ%�b_�����Kı=�gp黹i�.�-��'�,K?�D����T�Kı=Ͽ~�'�,KĽ�wjr%�bX��~��<�bX�/{{������\37r�"X�%��{��Ȗ%�a�R9���؞D�,K��oȖ%�bw;�ʜ�bX�=�����(jF���OJ�@��woip&�J�B�Z�kh��磵U%	�#pu�!���O"X�%�{�wjr%�bX��~��<�bX�'s��P�y"X�'������%�bX?e�/����77v�"X�%�}����kՁ!�6:�R���9"X��gr�"X�%��w��Ȗ%�b^�����{��7���o�}�A�:��'�,K��}�ʜ�bX�'��{�O"X�%�{�wjr%�bX�߾���~oq��������f��Yi�,K?������yı,K���jr%�bX�߾��<�bX�'s��T�Kı>�ߌ����MͶnf\��yı,K߳�S�,Kľ��w��Kı;�gr�"X�%��{��Ȗ%�b}�.wi�wwY��I㷇���17�< [$�5	�=X�
b8jK�7sI�i��җ3v�"X�%�}���Ȗ%�bw>��ND�,K����'�,KĽ�;�9ı,Os��:nnJn��p����yı,N��ܩȖ%�by�����%�bX����'"X�%�}���Ȗ%�b����s4���t˻�9ı,O3��8�D�,K����Ȗ<�F��ؗ=����%�bX��s�S�,K��~�g���!n�w-���'�,KĽ���r%�bX��~��<�bX�'s�ܩȖ%�by�����%�bX>���2nnI1����'"X�%�}���Ȗ%�a�V?��~ʞD�,K�����yı,K���'"X�%��E��������?��6d���v�V���Yg�kc�w<k�c�	Q�Lqtݧ��zg3�ul�f��w���oq������S�,K��=�s��Kı/o{���bX�%�߻�O"X�%��v�܅ɻ�7rݙ��S�,K��=�s��?�9"X����q9ı,K����O"X�%���w*r'�eL�b}����7TTg��{��7���������bX�%�߻�O"X�ș�~��S�,K��>��8�D�,K��>�j�v�q�S������d���w��Kı;۽�9ı,O3��8�D�,/��0)��8�s"\��n'"X�%�����˶Mɹ�����Ȗ%�bw���Ȗ%�a�G�����{ı,K������bX�%���x�D�,K��p���8�j��k�WH�]��3��X�nE�l��[�#e��'h��n��i�w��,K�����yı,K���'"X�%�}�����o�6%�b_�T�Kı?\�2ݤ-��廹���%�bX����ND�,K��{�O"X�%����"X�%��{��Ȑ_�&`�Ӱ�e���˕6	 ��~�	 �'�_�lD�����'�,KĽ���r%�bX������e��ۻ3ssw��Kı;��T�Kı=�{��yı,K���'"X���>�����KǍ����'/V)��c��{��7��|���'�,KĽ�wjr%�bX��~��<�bX�'{{ʜ�bX�{��z�����>�y7u5ۗ�a��4dz�6��㮚�:�*Y�h�b��B�[OU���5gQO+�b4`��śWm�1=`n�KVM��n�{�n��[q�u���X�
�֭�M��mY	�'=��n6�gv�u�7m�X��0��5�7=��.a����'N�5��;��"\l�Ǥ���h�!'0�r�{Amc`�I��@�9��6�-ܗw{�u8�2����V�th�.�d6���ۣ��C����y��:�����������b2n\���v%�bX���۱9ı,K�wx�D�,K���T�Kı/�����%�bX��^�wt۲d�sJ]�؜�bX�%�߻�O"X�%���w*r%�bX��{��yı,K��v'"~*dK��~��fɹ7s0��n�<�bX�'���r'"X�%�|���'�,�T!�2%����ND�,K����'�,K��os��[�[��e�Ȝ�bY�W�TZ~����O"X�%����br%�bX�߾��<�bX�'s��D�Kı=�ݹ�e�H[�n۹����%�bX����ND�,K����'�,K��w��9ı,K����<�g���{����|���Z�\����\�۱l;�n@R�k�a�ⳙ4q([�p�ڦ�{�����!xf\$���33v'�,KĽ���x�D�,K���D�Kı/�w���%�bX����ND�,K�߳q�� �+W�w���oq��_�l��u��)�"r%�~����yı,K��۱9ı,K��wx�G��7��������G-�9���bX�%���<�bX�%�{��,KĿ}�w��Kı;���ND7���{�_��?n�&�:�k��{�K?�?�(lM���݉Ȗ%�b_߿oȖ%�bw;�Ȝ�bX,ș��w��Kı;0�fwt��a&改��9ı,K��wx�D�,K���s��r'�,KĿoȖ%�b^���9ı,x��?O�MkӺ�ƶ�9�r�z�v˶ln��K<����:���]�ɑ�ɸ���\��'�,K��w��9ı,K�{��yı,K��v'"X�%�~���Ȗ%�b���s.ɛ�3!sL�܉Ȗ%�b_;���~QA�DȖ%��۱9ı,K����<�bX�'s�܉Ȗ%�b{߻s˖m�L�wr�nn�<�bX�%�{��,Kľ��w��K@U "X �PMQN��QNț��nD�Kı/w��<�bX��~�rf\�72�f\܉Ȗ%�b_}����%�bX���r'"X�%�|���'�,K��w��9ı,N�~�\�0���33sw��Kı;���ND�,K�QO�QJ�����'�,K�����Ȝ�bX�%�߻�{�{��7�����Җ�I��Sm����YMF�gK��յ�ݣe���wC�.9��Cf���L��2ff�ND�,K��{�O"X�%���w"r%�bX��~��?
�ObdK����nD�Kı=�צg촗wm�wl���yı,N�{���B9"X���x�D�,K�~���,Kľ{��ȟ�0�;�ow�{�_泞8�pj�����%�b_����yı,N�{��,�T!�2%��߷��Kı?g�ۑ9ı,Os�O��7n����ww��Kı;���ND�,K��{�O"X�%���w"r%�``�8�"�� ����"s�w��<�bX�/~��]�wm���.nD�Kı/�����%�bX���r'"X�%�}���'�,K��w��9�7�����߽�V"��65콚���;\�i���x�1��E���%ѓ����-й��.���Ȗ%�bw;�Ȝ�bX�%��wx�D�,K�����DȖ%�{�����%�bX?e�/�3s+�e�Ȝ�bX�����oؖ%�b~�����Kı/�����%�bX���r'"�T��7�����Z���Z�{�7���%������,KĿ{��Ȗ%�bw;�Ȝ�bX�%��wx�D�,K����.m&��2\ݵ9ı,K����<�bX�'s�܉Ȗ%�b_{�w��K���"�"~���jr%�bX��צg�٦�wl���yı,N�{��,Kľ���Ȗ%�bw���9ı,K����<�bX�'��p�#A$!}�x�Ò>����sM�$ K&|�S˧<+e$���8��p�?"�׊�H	&-�Y 8�R8��D`�	a���pb?�6!���rD>X�`@ �	s��wwwww2L�:K���<1G���e�5�^z�M��-�^������'d
ݗ�3z�Z�Uw,������lF]� ���q�\Y�v�q;��t���ig% M�N�p��g<: v|�"gTge\&b�k���6ҭ���g��m���v�A�m�<�S�hH�]H�8����̪[�5��9��;k�h�g	��-%х��l��P�����ZS��v��n�����������s�l���[#hq�v$����)n6˃�Qgkm;;cl�����^�k[�mD��G$n�۱��.	ٔv�I��μl�KtE�㬁�V�B	��.^���2�w=]����n��\�'K!��܄��l�)�-���<F�4�ŵ�����ASPgln���]AhF]��eR���ct�۱��݋PVe�]��2�Z^X;=��Ns�6�e�ё���s�h��N�]�hgk����<jr�i�y�]�jRe�Z� �x8��D��Q'�����u�Irn5���g�lKj�VT	N�iS02�lKm�@�f��D"[�V�u	�B+s4I���N� ��RU�l������Cm��˘ƪ�҂ĢF7��V(k�8[hu*L쵰UK�8b `:��]�f�&ܫwXn��m����[��v���Ӟmɱ��5�q�V��	/2�:�m��חzl�J���S��K]J��c��Ɛ�:���;l;^�'F�ŕ�&�+n�U�J�qQ8�¡��y���sR�H&���mn9�<�ø@��h.�pv�Z0Wm���� ��h�\�ڬ��]�������nM]�� �;x�:��kb��TvE�v��< �6-Z[,v��Ş���r8���k��J-�]K�NPf+��ـyh����.��mk��uƸ��`㭛j�=�ŐkGjN���]�jZ�l�6��cv��Y�v�>�˺�`��]�����^�qӣ�7w{��=�����F(*t �@�0V������5A�@}=�~qn���ۮ�v�U�:�nb�͡�Jm:`� ��D��t�bɺ�qu��pMP���mn���U�Yps��ֶ�/���;Wm�O�^1cH�D�\�u���ZP����V5v(�Q��9�n�v�d^P�:��j��<��=��aD�wU6Gp;j�	�p#�m�f��K�v�����v�J��um��n���<�]j���ͳs���|�������uu�gm�7�R����G��F.�:]�q5��G��l�+7Y{q���;����%�b_>����%�bX���r�"X�%�~����'�_�lK�����Ȝ�bX�'s�����a��m�0���O"X�%���w*r%�bX��{��yı,N�{��,Kľ���'�?(��S"X��~��[4ݻr�4˻�9ı,N�~�'�,K��w��9ı,K�{��yı,N�s�S�,K��v��I�36�����yĳ�@��?o���9ı,K��߷��Kı;���ND�,��7����O"X�%��^��l�Yt)����Ȗ%�b_��w��Kİ��������,KĿ~���yı,N��s�,K���w�����m���Z��H��$��c���f��,�����n�5?����'ϋכs3K�����n��D�,K�?��*r%�bX�����yı,N��s�Ry"X�%����O"X�%������B�f'9i=�7���{������y|+�6%���y�9ı,K�wx�D�,K���T�O� ��,N���3�ͳL6�����yı,O��?eND�,K����'�,K��w��9ı,K�~��?7���{�����~�֞�i�4��,KĿ{�w��Kı;��؜�bX�%�wx�D�,� L�u�u)�&0��L:b�ʲ.-]�f3w��Kı;��؜�bX�%�wx�D�,K���D�Kı/����yı,O�����mͻ��V#vOanm�.�\��
ఏ=��N:S�[�%�X�T���wy����%�b챼{ı,K�����yı,K��v'"X�%�~����{"X�'��։�&0��Lo>T/�R�U@�Z�����%�bX����ND�,K����'�,K��w��9ı,K�~��<��*�L�`������2鐅˛�9ı,K߻�x�D�,K���Ȗ=X�>,��"r%��wx�D�,K�����Kı;���/w3snW,�����yĳ���?~��9ı,K����'�,K��w;�9İ?
��؛�����~oq������L���E�bs���,Kľw��Ȗ%�b^�;�9ı,K��wx�D�,K���W�oq����~����Uj��k]F�n�kɒ�%�G	�iGc��uᇱ�պj����L�%�f�p�w<ObX�%��?g�Ȗ%�b_{�w��Kı;���ND�,K����'�,K������i����6��ʜ�bX�%��wx�C��DȖ'�����"X�%������yı,N�s�S�?���,{�����,۫���{�7���{����~ʜ�bX�'��{�O"X�%�~�wjr%�bX�����yı,_�ۜ�ܺfK.�wr�"X�%��{��Ȗ%�b_��ڜ�bX�%��wx�D�,@��|�y7�y�9ı,O�w��|�ɷ,��n���Ȗ%�b^�;�9ı,K�~��<�bX�'s�ܩȖ%�b_;�w��Kı=�������a��6�3vltܾ���N�e�ģ��X��s�:�]�F`
���	wf�B��ڜ�bX�%�߻�O"X�%���w*r%�bX�����yı,K��v�"X�%�߾�a~��প�����{��7�����F�h����^ wo^ o��:""!#��Wء�rCbq���M ��虘����� k�V �%�T�A(�1I&�u�4��h_U��fb^��4������s�Y�@7�w�tL>������^��"b��_��fgrK�6�۸[sa�����(�;m]�k�u���\t�A��� �r�k��=`����E�m���.�X�bIehw@�8�-�Uf��!{;�6��S���h �Iˢ�Gm��w]�1�o�����2�ש$��s#6"�6
X01���zѐ�F(s����Ks!m^���_>p=��؎靱�!-� �.�y��B�6��v��ì��cv�utv���:�z�NKTA�{]��X#m�K�͛���Ůuz0��p�����~�V�|�41� ��;�j��3L&!<iǠ�Y�z� �[4W��?^��o�0Q1�4��@�h��S�>�z�x�H�����f����W���f��X�*��bi�8�h�k�5=u�6� 5��*6��T!fa���6�5�,㭎�v�rn��R�W-�۷FD��ɛh�k���}?�נ�hc����-�O]���lܛ0����O{�� *}�=�`c�:��S���ۼ��DsG$��f����W�������fI��G1bnM�[�%1� ��F9�}�{wr&�LBxӏ@�z� �l��f���z�B�HܐmȚ�,s�I�g1�S=mI��89�&�\Q����ǘ)��E#��f�u�4W��9^�@��?���1��c#�@:��7�Jczn5�w9w�h�#ӎ5$�+k�*�^���?�8�DDF���3?bu� o�� �5��/�܏@��zW�h�f����E�n�# �n=mk@9�4��1�7�n_��H�I��t�^�Zy��s���v� q��e�j7cG<B�IUF�y1��J>l�%+zLo@��h��S�щ�s6��9[^�H/W ����$�߳(����ۜ���e�K+������r�� ���:�V���T,��W%]Z�Wu��31���z�$������}��o$�B*V=  &0Em��3�O=ϰ��Ct��y?�q��f��ڴ
�W�r����e�UWtZ̊2�*j��fN���9�b�.; �f#���]����{�����Ƀi8�RI�������*�^����޳@��ʢ,l$BNO]`�u��u�3�a!�$Ῑ�)�E	�q������u��*�^�|�rI#Ds�@�x�`=u��1k�� k�E� dbyō�4�)�Uz�����f�e�1[��%��s�u=v`�n�b�$��'7�BZ�HX�sjX��l��w:TXge�ɪFIy�:j�w�d��$����v���t��9f=]N�ۜ@p/lF8���#����U�ɔؒ�єC�� Pg��+�aunƶ���R�����ݩ�q��7c. ʜ�.ٵ�:��/O{y���|,u��v^��ny������������ E�ԭȻ;c�͠3r�v5�:8,�uIa&ݺ0k�̈́�.�R�?˻� �6� n���"c��_�{��Q�QuJ��v�� �V�W4	M���}._���D�j���^�hm�����ľWW�|�����"șffh]���-��� ds@�SV�*���� k�� ���L�b"g���|��^����N�J�=������n�1�2��5�غ1Irm�*���9�W8�X�<�;�Җ�4��h�h#�W}�5�z��/6�[w-�)����N��w�/A4����A�À��@����� |���m�z&f5h����.)T]�(�����0�n�艈KWwV s}x箱U��j��
�j����D�LW������X ޻�7]� �u�,��1��R)��mzoY�wYM����K��)��LNa����dԍ�p���Jt��Ў�֚�����{�2�`�����UsWw_ {���7]�@��z�����⸁ȉ��34	M�7�u+z ����fbG*��@HM�#Hp�>__������&�|�O �B{�1=���j�S�bI$Ȥ �$�� dXp�&$����u��#c!@�	
#hF,E�B� �$H��mq"5�2aa���0b�5�D$ �GFcX�QCB$�z�=�Q!�JJ���e%�bB	IBVT� ��@�< @ BI��0������BA�Q�%ŉB��e%H����B	""`0  H�"� ����D!2�'�>*�B(��E�Q �b@�`DbD�F,B!F,$H$bBXD�)�!24������xp��A�ੀ4S��	��C>����h�M�K����DMB`�z ��x ޻��l�阕�ϫ ��AțBJc��)&�[�h�S@��z}l��VI�?�2F&��=�ڵ����3![gs�p�T��N戢����a�LXۓ@�ҚW�����鈘����׀w{ՕUw
�E�ܪ�0���$ϯ ;�^ ��07�A��RG�u�4�Y��b!'�|`����:LGQE�*�����������z�����S�s?��}f�ޱ�WD��'$�7�l�=1[�_�7�^ =�x��O��j�&��]/dãmqͻ��r�y�����|��w[��ݹ��BE��#D�y_���נ˚ܹ�w8�ɭ��6+��TwX���D��L�EP7�^ �{� �|�g�"R;i�]ڸ�I%1�Y�@;���=�j���J���@=�}4^s��!�yŉ�x����o� �>� �ۼ ׮�NU�rLjb��@�z���л{���׀=�k q?L��K��N@2�S�a-vY{�I�M�ˎMZ �j��,�\�=����&:�`leL�2i9����6���0(^:6].+�W	tͧ�ӳ�N?�7���踪�<��Ǟ#ڹȅ.�z��I�E����B�7j�p��m�FD��t���`�]�� ܛEك�7�'+�[�k�؃t:v�PO=u�Z��oWa[h�q蹟b�$t=:4e�gs��w���|n�V���7m{a푹`�k���dԑ�ܣ���` ��N:9��q��Rb�]րs޼ ׮��]DDG�s���Q6�bmI��&�u�4
���9^�@/���cx�Ț*J����]`��æba#����~��E��15r ӏC�g�Juϫ ;{� 5���X�[N,E�UV��U� ?��鉙O�_�>]~z+���G#$����L�����&��n���8Л��v���	�}Sf�����%1�X��@:��^��W��~@}o�@�����G��X��䓷��94b�'S��Ds���= ���h�f��*�Sr`�s����`=u��w��f&f;�^����;��,{�M6�qH�z���Ļ{� ;�^ ������KD6�O��jL��4޳@��������@�Vr���8�(�:�H��ml�I[�x������nɵn�4_�����qjȇ��rO�|���^�@�~����ϯ k��jB-]R�E���5=u�0�w>� |�����LL$�⫢�XU+E@�� ;�o$������ *���>�䓷ֽ��G#��Jb��9&��3��'ϯ ��� ��� =n�~J6�҂,.��B����f阗\�� }~�h^�@�u��N)$m8�0H	�9���^������s��'fo-�L�e��L�Nc�-�����@:���j�/ulL�ci���G�[�鉔����9��jz� ��q���i)25$��f�z�a����}׀o��5I\]�4�UWw�阘\�8����ۼ�S('�A"��"1�&�Y�U�u �Dĉ��9]u�z&Wwu� |��ݳ 6����&�ΰY��Ȍ�ۭ����&6����0�V��}�����+�m�����?~��41�\MS����S%�,NI�z��)�r�^�[l��\;"�G��X����ـjz�DL�""��{׀���4����Hӑ!��NC@�z� b�F9�1w�#vU���M*��Z�� m��=1舊�w��=�{# �����3Q�ϳ8���B�f1\�c�9�ج6ӭۖ852�����qi��ԣ�0mŘ�8��6�Gf��&��o��|~|eW�)�X�b'�\Ϝ\���棞آ{]���TӵB�qJ�#�ɴ����p�6�Q� �T�s��gF��D�Z��h�둞�8���63�X:lh�8뙻[���i��x��΃��u63u�6����k�����:��)��a��y��F�4l��g�
��i�v��L�PT*ub]T��]+����^�����k�������w}��8���i�&��y��T5��`��^ o��~���*�(H	'0�����zz٠�f�z�� �Wcw"Pnc���@/[4޶h����?�>��}ί����%1LX��@=�f���h\��\�%zT����3��7v���z�C���f���f��l%��m�t�nNb���tOK�_6�~���0|�n��w����x�wU,��d���m��<�k��nd�o��@?z٠^���[�A��84�q��� >z������5�Հ~�ZBtB�	]�һ�D����uܴ^���f�ޱ�VF�oR]�f�ҷ�Jcz �������o��jծ35re��[�3�3�}Fs��J*�a����x��}�Db��M���˺��^�V =n�^�����ՀqWcv%��Ĝz�� {���5n��5=u��ιu��ڸI\R��Uwx ���kZ����fd����
E�(?\̽����l����2%����Ĝ���X�� ����"c�U��^��U,��qwH��uk ��������/}��=_U�_XVI��kκ2Pn�ۜ����D�Y/;;9�;,�\i; ԍ�D�o�ƤR= ��hz٠u}V��z���f+��I1b�wx�k��JC�|`.}X�]�3�#���/��0r$��h�>4�7��hc�T�����`��ʫ���ou`�׀=w�Q蘟�3�8�� ���U֔X�Z.�ח���h1�7�%rށ�����*�k�l�nx�˽t�����`�T8�\�.���g��8�
*�K�U.b�����u�`�n��\���+Ϝ��bo#x�7&���z/Z�W��^�@�ŭ��c�E"�.�� ��u�jz������׀U����S���)��G�ɍ�1�S�%rށ$ʳ���J#��z��h��@��^�>�w��'Ŀ4�� ���B�J�R�];_ ����nl�kc)���n�~�Þ�s1�Q�4(E��!$BT|��H���"X�"E!��,��%KIB��0"
R����X���$ZB��FRP2����� ��FT�`�D`ĄaD�"@�e��! �$+,l���(��0@�)bP!,��B��H��$a	R P%%JT�D,�B��`� D�$T��H��ĉ�@a�H$C��<��D�!y��A$Q!$UB�lU� [*B	A*��Čh°Xabő�@�H��)*Q��A���4-bJ��BV�	�B!Ng��~���ګj���Ϯ�9u�g�s������u�e�Z!�L�E綆ڕͺ�^�&�;j�����Cd��6���|���u*�V���G�m�����}7]VB�{v������a��r��FS��5�Wj\�JIs�Ae9\�Z��h����Y���ʍD;�RZ�ة�:�u������}�"���u��$�Lq����3�$��B/ki3��c��.��\�,�����H��u�ְ(��%-n��.m�p,v}54�Ol9��n��c�8v{p�'���]� T�����$ӹW��̔q�\�z��M�Jd.^;��ÎL(:իg���aY7;�V�mm�a�,.���I�j�:Rͻ������i��VaoS�5�������1zۗZ]��&��'��n���:�C�BLG)Y�i��ӟ@v׷�\�9v�X�������7�6:�əN7CO���!�*����N����-���AGLCZ]$dwH�Q������N�ޛ6��Rt��8�#��z&IZ��t�m�Ͷ��ui�` �M��V��up�۰ON��WT��m��`� ;k�`��D9�\Yێ����Tc�n]�q��#���@�cj  �Z��r6��)2���UUEJ �Um���;`]Xk[��v��`����g�Pg�5b֦L"��(������mq��a`��UQ�C�o�����Vݶn�d�-�ؐe�g�������.rY��ˣ��n�C�N�/[��V�tʴ99��Ԥ�.Uxܹ9�s ��%4�l"�w˖���$Α635	�%��n�Œ�p�{m2����`9��k�w�]�W����ض]ɮͧv)�y�;�-��K�-�l�-u��S�E����e�k*�c����1@!ͮ2'//�-۾6�\�L���^�k�=�$�綼�m�%[�]$�I�.���Asp�Dͻ:��c�t@+ӻX�=Hut��yem"Ӏ֛t����X����� �*�z	�"�hQS����\���&�0��$۔��2c�3��1-i��5Vޞ�1��|[�x�L<ܦI��1�ֻ�� y�ԦG���[]��m/M�`L�`�c8z��v���5Ȧ@� te��5�5̩��5�+��hܕ3��/��;��rU�Z�ۈ�2�VEİmv�B���6K-Vwr�3�v��r�m��r���nI���պ�T�v�tj4�Ͷ}���{ȥ4���ݞm���.�.�74�0r����9�֬��,�䙰��M͙���3����ƞL�	G$��~�=��z�l�{��?/#�@H�1H�G�~^n�u���]�&�g��D�""j�O/EW��*�uqWWX��^ }��D�%��� �>���N��t��Ҹ��Wx���۬����3)[��@�y_�qH,M�o(��<���=313�>�������x�I�)�F�&��6��{\�`Շ;d�$ghB��S��:9wFd6���;]\@��� ��4H��ѽ�����m�᛻ws�I���U?��+������ɷY鉄��ڡcS�)$�~�h�ՠy[^�z�4z��\��<�$�ɠwZցԭ�+�"��(\�	�)qhVנ�f�w[4W��?{u�#��Q���A�"X��qm�z���dۗ�����u,싛n�!#�2'�u�hwY�r�^��[^�y�d��F%��NM ��y�	s��>]�X�7x�Q���q,M�o(��=_U�~Vק�����'�q979�y$�[��.wV��1̘�S#q�����s@'G4��"�eiU��S�H�z���g�=�h��h��������D�'01��y���S�ۮȖ��rq���
u���6�kT�5ɍLmF��@;�f�����^�~��ޱ�W�$��1��sֳ�bf!#�ϫ >����]�4[$x���('!�~W���٠�@�빠��e�d���L�ǁ�2�s���� o^F�Q331�ޯ@��[Ȣs�dǉI4��h
���cz��Ni�̼�^���;�K�j�pڭ!�d�V
�9�qr�al]̑Cqh���l��U�m�����hS�W4ts@�E����fuqJ�º��~O]gLBA��x ��wYM��ŢL"�K�H���w]��3	5�Հ|���ݺb/���"��M ��4���?+k�^�@��o����dq94	�&�ԭ�1� �s@}�������Wg�&�'�=3v�V�9uӉ��u'5G�8���n��m�����k��9��b���L�=#�� ���DѦލV8Ct2"�yl����e�V\g���66`�٣�=H	ڞ�wF;A��n��ٕ�[7F?�����1��v�y�Pʗ':�;t-��������F6­����c�1ى�g�j����FV������������R��5'I��Hl۷<rkh�[r)w7��m�X�>-�iӱ�,��4.�.'�I�_���� �9��4	\��j���y�s �F��^�@=z��e4_7Y�12��\��-WV"����~f�:ִ	\��u1���Pcr0�ǉI4�h��z���>�Ļ���=��[�<���K��%1�����4	ֵ�|ϼ|�C1e�k�s�e��x��S�ڇ�hw;���z�f�X��aŰɋ���2��7��%rހ��$�؋�f)�"x�@-�5fg�L���31A��� k�u�|���>��T*�Cq�E��$�9zנr�^�b\��= ���@��u"C�2H�p�K�:�ށ���1�W-�]��c����E#�<�W�}���~�������W�_5]Q��	Ē@��v#t<u]��0�oݺ�c��2iY�u<)7�$c��@:��/Z�W��<�W�$^x�ϙ1���]�hO߯@����7��hgZ��H�E���W��<�\�_����/
�=OE{�&}�M�U�z�Lׂq�cF9"��Lo@#�'Zց+��	&]����XE1��z��z�h�k�z٠{�+RG���dc!ϪQS`7f��Z�p$W]�n��M:�m٦��z6��p#��9&��YM��z�[4׬�9r:�"c�F�pNC@��zܹ��4�Z�5U2�1��do$q��l�^�@���@��^�k���$c�$�C�fe-���5s��>_7X� ���h�I$# �1�F"~h�!I!# ���B2 �H	0�B`��a1a��E��F!$u]0!������_���@��|ҹ��x�'&��z� �|�`�����xDL��w~����C\�1�%�]��N�1r�=�`���jH-�ɳ��5�lո�.��8���|��٠��@��T�x9�	c�G�w[4׬�<��@��^���؋�j<k���3@9�hJށ+��E��cySō�?��hVנr��@:�4׬�?.GR$Lppn����%rށ*-�#�R��O���FQ��l����/]*���n�e�2+^l�L�vW!):�"%�rP�-���:Z�������/�n�C�ۭ����7�7W�8v筴tl�lHO
�W;K��Ɲ�m��dT��x�f�Ի�մ9�@m��P���<�э�nt�9��<zd��$F�Bn�6��\����q�J�����d��Vzux]���=�5\�X�ţ�f2~~AP�O=�_sswf����ik��1�Nn���qX�cj��h������.�%�5���{�z{��<��@�ֽ�$x��D$�@�:���[�%E���/�8���M��ܚ��h^�@�mzoY�{:��q�x4�H�š舘]\���u�z��b"S��Z[�f�"qDc�)�u�h�f��ڴ
�W�<���8�$��N�8}�\u�{m�z�:�Q�G�1��㝯��E�1�lX���O�� �>�r�P��4�¼0M��ww�O�����>�|Ѡ�U�נ�� ��h�#�(�R�	$Z+����@:��Wj�*K���9�'�H�Vנz���h�W�^tU�PRGD����f��ڴW��9[^�圹�7'򌙀Ҋ#�G�ǆ���cv�N��!wj�g�:4Bs��u͍ٔo&��:�V���z+k��f���[�ǊCȢ��Z+��W41�6��s�oǯ+�1G�@:�4�Y���ن�f���!z1�a@��A���*��,�@H�1H��'KLD�!��<�aa�`i��2����8#:!YUk ��0hUl�Ek@�0��DH��a�s�CªA<9��������i��B0BR$�$1 DN����'�AX�F,���"&R@�`E�T�X�"D�a��!��	D��"dC-��)��DO>V�t/����*�uD~�ZA(Ș����TT�����@��wtM,�Ƣ`�]�zfR�}x��X���~n�z�¼��$YrM��Z+��z٠z� �ˊ�I!1J��{c�7O($n��%�8�`�(g�6e���F��O&(I"�9^�@;�� ׮��\������IE]�]��Y���4	Lo@�cz�7�^tU�PR)1��1�&���z���W����@�<猸��Q�H���>O]`�]�~@w>�19?�0�΂`�����?g$��fr8�x�G6���@-�4
�����@�܊�#q�m����[��e2N��\ts t7t1]{GA��d��FU�29��rh�f�_u����L��k��v�(袡Z*.�Vf�=��Z �s@9�I1��$�G�@��Z}�h�f�_u��GP$"�͓$����,s@�hq� �K��I!Ɣ�jI4�٠�f�߳��I>����&)�P�B*� $%����������In͸*܃!KZ�K5HQ(T�N��I�-�:�����_a%�a�)�6�js�T�w��[���&I�܁nv�Y8s��+\��vý����ɲc�;�\5�*�.A�]�6�F�2u��UU�N]u�OI���o��"�K)�{rQTO���kkn�J1����Li��];����nw&�[6n��p�sh�'m�w����W�|?'���um����ړ�v�C]�6�h,��6v��t�:���b���\+�� ������X ��x��x��p@8�x�7&�˺� ��4�٠�f�ďg���j(	�.�EU]`k���w�LL�Gk��>V���[���ŉ��4���G4�o@�hL����%BHܚ}�hwW��f�_[4��ʛ���f��S�m�0!��Zv�������؇k���]��<D��i�dq�?��r�^�[�h^�@���1@��$z/Z��= �C��@��O2N~��@/_��Wuz�K��do#�a���� ��N�h\k@>c����$#�L�19&�w[4��h��@/���[3�D�8�,JI��ύ ��h�Y������3��G!#J%#�!�8B;tŮX˺Kym9hۋ�JBZ�Fc^�ɪ��&��������� �l�/��@����(�&,Rɠ�� b��\���:L���C0Y��'&�^�h�SG������f}1Q33���u����7v�*�1'#��G&�}e4��@/u�z٠yTv\�9�@&8)!�[��+�������l�>���V)�RI��<��	�x��)d��5ht�:��d�7MwXv�����]��j�� ds@�q4��n���H�)�'$��f�}e4�٠�����Ĝ8�,����@\�c� ���u���2!<dq`�4+���]�}�{��'?��O�k�(�o��NI>���s2�\�ۙK�2�4�s@�;�M ys@�=���M-A ػe݁�=c�PvP�v���:�`�qhw�S��I�:7;;��e�|�f�9���4����匏��@nI&�޲�}l��f�^�4*�ˑ�1�	ت���w�u�	�^�]�@<U̲'�I ڒM ��h�@�ֽ ��h�Sn(�&<������G4�o@\�K43��g+�IF6��rx��	$�E$�5�8������Si�M��Z�h,���FA�8.!�Z�mC�{f��sT3��;tJw۱f1;g�����EG'ktwd�-vݻv՘��O<�@�iU87]�jws�Ua�������[3���0����:Y���;�vĕ��9�����5�Wmg�ˬ����l۳כ%٤�г�V�o���{�����@���/��oۻ��륛��"���XW�#����St�j2�ۋ��2�0>d��$mƀjF�bnO��~�f�^�4��h���k""6����9��h����h�=m#ncf)rh�@;�f��&e.��X�>�wn�(p��**��̫��	���Z��� ���ю�C�x7$�@�v� ��4�Y��� �쮩�cQ��瘋�c�8烞6�-����`�̚�]�ɵv���2ai���NC����@/u� {��1�v�r�9w]������2���I;���t �D?�8�"%DDfo� �� �� �6�T"��ȅ��4��@�YM �l�^�@�򼱷�ŉI4	�&�1s@9�h�hz-y��M�!��4��@-�h���׊�2D�A��Ă����m��w���:�j�t���жz9��q�	��b�nM �l����������ie�8<o"R8�hW4q4�-��h�X����l�M�)�~]k����� �GU�n����O����ʢ�ȱ�y1b�	�h�Z��f�{���)�~\�;��ȇ#���yz ���9�+��}QoC��߶���Vװ�GG+v:.=W��aM ����hɴ��t]O�{6���e�|�hq4�-�4��yc�&0q��dnM����?.���f�{���mX=�O�)y^+0�>����hH��{�Oq�l��F8��}��٘�����O����'}��rL�C�:�O/���d��Hԓ@=�f��@��ހ1s@�1�����j�j��FQ������uW'.�Np�FK��Z�f�6U/b)��5�m�������u�@-�h���?*��<O"-]Wk ����DL�ϯ }x���?*�X5�Bd$�ȤzoY��f�k����]+�di���i(J��9&�� �� �6� -�4��x1;�C�ɊI4kZ�+�m���X����131+�� *+��P�� *+EQ_�E�(
�����?�Eb��+�� *+�q@TW�"����@TV�������
���(
����*+��@TW�EQ_�E}E�1AY&SY��by�vـpP��3'� ad/�	 �l4     $   2�      4    PJ����� *�E*� �  �      
(
�(��   V  j  
��P�� �ϵn��_}�ŝ������o�>��9>�\_u���Y�}����8 	�l���|��w�ڽ�s����%�t�Ε��6�jv�c��%`��| {  �  |��n� �@  E �̀�{t����׋���I������:���_o}o�%���xr����o��ͽ�sd�w� y�1o�����}k�����E� }9U�,���w/j��9�v�< ��  �P*�(Rɠ%^�S����m�m���y�����*��}oW��ɜ�}���W��n��k�w����w�}ϝ�*p >�����]��ޓ�iV]�W�J9�̹�����۷�v^����y�H 
 "(�� {��7v��k��n[{��@ :���� ; h" ����)�
" ��   6�p��@`�@ "th4b 9�  ��f &�)���   m@  
 
V@4 &�M���
Pm�t��> |Gr��[�;������N��==��C���Yw�}엖��  ���t�{��|��>���W��;ϼsǎi�;�ۀ=>�}��z�S��j������_ 4�Sb�(�0S�FS5R�   <z�R�~���� Ob�CTJ@  S�S%<ԩR� �""CRRHL�hx�%�������P������v#i}��BQ�z������
 ��DPTW����������QO�����?�R��O��=0�S0�"H����|�fdu��8C��&o<��zl)�M�m,^�*�M*B��V,Y�/
R'��}��R��e�2�2\�����RX��!�r^By��d
s��U���\�I�=!s�
��
��/��p���a����,o�T�A&e���*��)5}�YUPM*A58���BD!|��V_���r`Sp%��'����2�Y3�#�>�>%ͼ���Hz����!��\��4��F}�_09�#x@��Yp�.]��(����J$����+�����!B�o �ȼr�2��d���zx�7É�\�9�	����������
�o���\}���sX^ӛ{������i�B�Au�B�T
J��4�^����)9�7(��hB%"OB$������ӵ��a1�`�ET)�~^V�M)�����+�O�A5I	ߣ�9/"���%JbK�.C4)���BK�!�ŋ"`HT�>S�*����E5��M�|R��F��Q~ϕ���h�+)o�B�z0l��&�
���0�}�D�ϒ\a���!�J_k/8@��\�0"I�����S��}�"L�E���y�y��%�hp��M��y�慯��_�����B<�
j�T��_Ԑ�W�ܻ��zp#�`K�G;�~��ԗy���eY��Nӌ����dx�K��3�{|=�T�3t�����)�7�O|�BQ��s� F{a@�0�d'�ԓ7͂���Y��N,a���#��=����_Isy秉ce�LОg�k���}3=�w��B!SN�ϠH�*^��g��7�x��B37��L�����7���Z̰ؐ�c
c
c6L5����#=��)<����^ar��+/1�9�{���� �i���Nd�RX�fL����>������1�j
aI3J��c�ā����!���1eŹ���[���(Ktv����+
�zi���,j���}�5,X1�!F8�
cΆ�X$�L#�KaHf�����L"GH� H��"0*a6@�"\�\Hi���=%�xF$5�4����\�ac��b!�#���b<�r�b�����Xĉ�xr��!����XL�\�"H���
�`�B5ą0%�8Ns�����Ba8i<=	L���%����9�=e����HbA��@!���,	(B�d�L� ��g��I��L"o���yd�$SX�Ғ������
��p._<!B_~�!�)�d.2�
c�=}o�=Sy7П�v5�Ԅ.��D�+�C�W���Ç F1��`���8j@�����@� �	r/Ǉ���)�I��Ȑb� �5�Ir�233����.O=��L�&� c����^$�(B%�H�2��,H1HH(Į+<�q0=�!R%"_�t>CR�B Nzp��$Ф��4�L)�����t<�fBp�G#IJZH�l*@�x�"h�d� �����&�������b`zp��̆'�Sr$�aHA���B��0��62�3��s��0e�B�X`K!f0�HJ��R��^C7���p���.;G�����^)"EJ����/���!M$UP�"�M��rʦ�
i,��"�!�D��E�"�H���
��"$J��1�"愌��FH@5[ld
)��#0��`E��4�R$�Ĉ`A�`E�h�i��J�l��8o�SOPp4 �\�@�!\c�C4"��!�
%00��o���������(B�"L���q���`E�<O
�O<�.˩�B45���F�wOSG�.�R	'+d�c@�j�H>.�	�� $X��G\p!LBR%rhE (`�p�1�41ˡ�hF�2��MB5"���
c��!���B)C7FT�!Ն���v�,
��JK����H��H��8�(`�D�L����(�1B)�.�H1ơ�KC�V$0��0 D�Sp ����Hb� +� �pā\cLH��� `�!H`Ĭq"0"�#��č,%0a\H���5�3Yt6wzJ�k��\�r�O��=�/eU�{潗�n;���:y�i�z�kų(���O��A�WU���}�i狯9�y�|'���3O}�����"�:Uc[�Y��*�3/�}{����ݾ��Ao�.��W���������+����_5��vo�|I!���=o<��0�YR-�TϮɷ6�H�L�ݕ|%��9�����J�5��f��	�\��A�Ͻ���� k.@��H��1��H%�Ѕ29��QcK��"Bn��!0�8P��ɓ|�,��3t�ԁ	sy1�bB�f B�D�,�\0��bI��� �a� ��CI#WX�_F99���%�����
P�Z
�`V�c������/�z�(bd�_�ax�[nJR��a}ILӌ���J�)	B�+� �
#饳4��Z�n��H��������~� �A��%��H�@%�f�\��L��Q!R�`D0"CB4c��)>C�H
PC##\ؖ	"��`}k�R
l,d��L IL	`H%"I����k��I`X����D��	h#&��(`H�� �)�I�Dj�(�1�F(D*E"�W�U��%���@�"�H@���#���$�:����.�!� ��B4 ĊF4��1B5aR
^��F?)�p#Hd)1�J�"���0b�	�, �� �. �+X�j���A�@"�B)"B%d�	0�� �rHXG ��IHD$_�4�A0�P�4 X��$C���Ka8F��2�LQa0HŋV**��x|A�)���B�+��Ġ�`� ���!p�N>�A��	�4�щ\�2�ՌpٷCH�<vV�8aRFT"� �H�Y�>�qԅ�@�V-x�
�B�1�#�F�
��B1�"��(a$
A)��=�]3��W�����=dhqb��"|�x��"@`Z� `b��0�	r�C&9�4���,��
��D��V2�����*Q.�Ћ\�fAԅ��8Yg���"$B+�Q=���� ��_P(�B ��}�)��.®04�
�fA�!M��=#V!!|fd׍��q�8xċrM6�4�y�jD��'��J�/���B������Z�H4�<�4�Ĕ��aM���4aF\��|���C4�<�[d�c�(>�[0�+��ԋ<��3D��GyMd��lcs$!�4��iD�N]�O��x20*��H��Ҕ�4�wd���i�\�Zq�>W+���`
1X�,�a��Z��Db��
$"@��B�*�B0�,����`�}���RS!�T ��H�$$ld�la%M���L��8�3w��BxØbB8���d�R��D�
rHS��lq�n�F�0�RBH2IwNF���k�$��K�N�v���ɿ��aB�  �[@ ���   -�  #4�k�$�gf/*Kv�va�UjǴY�x���'��vӠ7���=ns��1
��ʗn�/<���j�W�a�aSB��r���������Q�qCZ�����c�`��J���j ���l��mqcS�Ⱥ^@Ļ��7)�������6�i���� �2� m�    ��n���/^ ���ݴ��� HM1&H�@2N�)���"��I$��! �d wZ��t�n�n��	�D�l $p  
Sm��^�B�۰  p��m�m��9�ua�� 6��H[I-�m���m�d&�  $  -���K��6� @�@  ���-���  �� [z�UU�6*�\���NӦ��D�-�� C��������� � �m� �'mp$~}�m��� qm�c[��/i�/-P�P
�U����dЃ2�e�W�g*���Y���m� 6�IV�Ԭ��(g3)+�Z�z�Rl�t�  �D. :�b�]���˝\fݱO�d���W:��h6M��;�R����Q [r&�7f�����/	�@�	�/N'��m׬ۋ&m ir9�,b�a�j��v�Kj�� j���x����Y媦��lX܍@V1Oc0��Y.m�mܞ��YM�n���-7`[Cu�N!U�Ҋ��c��2c�%��Z�P*�� �  5�t[�KoT������ jT�;.ƶ��j��p^�i6�]��#��͇2�gb^��`*�BN��w��R��)�z���<
�UU�U�d�cp$iyn �p��% v��{[�ꧬēV�[=�n6�b�m�/;u�b�-�[��  @-�^k�I6�HZl$ $�hj�N��q�Fs�p;4*�T�u�|7|5�۔��m�,�ۍJ8�-U����;@�Rv�f�`7k�*�����S`U^�A6&]�(*�ml^�F�����@��wW�H��UUUC�UU�/��8�96U�p5��0�l�S�p�]��Q;N�#Cc���r�Ni�[]I����UT��n4�V�K��e�W{U]Z�OD���L�2�xĸ����r���m[��$�z� t�4ڬ��V�j��A�6@9�#�Pv��k��YR�k\�cDp:�]��5+� U��[`�R�֭��<*Cl3��=���`�����m�������]�6ͤ����l$���TUmYI�eZU����[,V�[C��n�6��I5+$<n�"��lۮ8%�:�8;6�ɒ�`����U]K�[J��';Z�:
��m�:H$-�����`m��IրU[m��V�Y���lm��m o^lit�$v�Y�fگSʭ��p�wf���qX���&�sv��  崐��!�vZ�`��;���d�KՄ�m����ž��i:�kv���o\�hڳ��[@8   ^�P��m����o��6ض�鰐�i[��Av��J�l���m�i�^��m��$�D��ä۶i�l�۵�&�]d�]����Eݗn^� Y�ګ���n�����m� Hpsm.M�I̐��� ���E��8l�U��m���m��}'W��-���p   sn�6�`Ȗ�HqK�!����X�iv�����~o�J|��e8�� 
V�:.��^��K��� 4����Id��[[-lͺM� 6�t��	$�-88ΛV["Lp��"@�`m���#m&m��m�����BF��  m���9#�� �`,6�#U�j�"�����jڠ:�UWf� w-Tk��oX��͓�[��ZÄ܈��p-�6	u��
�,���;kj��"[�ڕvڶ���j�6v�ă�-h�m���[vm�oW� Ā 8 pH�� $[R-� m�M�]�W�W�����eI&� Y��d�� $��m��ml -�  H�	$  m6�`6�h�U�LRL9:-�-���9��I�M��H�2�i ����}4�o� �Z������s�  �a�Ĝp  m&�H �E7m� m� p  �`�[A�$�d��$ �lޑ�l�L<��BKK5m�m��l�g}��|    ��n@6؛\� l   m m�6�A�AV�aq�h����8��E9��$�l����  ���` hm� H7m�A u�� [F�@N�6�m�]��			n�� �m�� �l ��6�l�$�K/��u�M�X�]6 H �[]	9�m� �I�`#Y�m�� �e�jN�kd�F�j���m�޻a�fY6Pq  8 �b۶�n���'Y0�+Yk$` ��闰ܪKR���2�?��O��kl��d��Z4�E�ܥ�I���
�ԣNrG��ж�: �0I"/Z �m�g H  m�ض���m��q,�-4����ä� � � �� 6�[)�� H �sm�kV��@n�;j��l�P��8���m��-�U���m&$$Imn�[[V�  ��  ��o +m��#[�h m�m�l ����C�  m�   � ��l � $  � 	       $jj � 	 ��  Kn�l    �     8m�  �cI���"������mz�@   �   Ŵ -7b�m�a�lk� �M,���:���� �8l�` 6�-��L ��   Jm ��}� $   i��X`�4Y  �`%�` � �&��`��Q����    ��  �l  m�,������ۀ��m�V��    �` 8h8Hf�0-�-�   �i�� #Z� � 5Lm�  �� m� � �S`ݶ5�� $ ��ٶ6�� 4P[N �pɻv�q�gn�Ywl ��[�Ip$i�7Hr��Kkk�l�USeZ@"������j�t�U��p �n�yh}���jF��eu�����s� �� 9�oYm�-��k�m�U�1��
U�Q��gi-�!�[A�ׇ�M�I ��J��6͵�.�z݁m�wM��@-����-[]<��f�hڶ�� �ݭ�Y'^rړm�� �M��@ ^Idb�<[����d$-4�P���]����ԇ �����  Б���LlH��ݫT��R� R����8   �%H �sl�ݴ�[@k{i6K(���i�m��	6��	*���Z�X�� �hm�x�h�6���Y��kdvp n٩d����mUR��j�e��S%("U|��}���$mm���i-�u�`�P����  ky��-�-�q��k�����&�!#���K#�f�kM& �u�K:���n�jN ] T���R�)�� �%l��X�H-����l[[��� [@      [@ nM&-���D����m�fӦ�Ӎ��N� �m�� 	��@��=����U�ʯ-��WT��Utl����R@⪬���J��4��Z��6�K�[�6�ss��m����R�etm*� Ul��b�h����]v;[p]-A�J�T�� 6� m�tͰ�����WD�.0��m��H�    � �v�[    �au� �@6� �m ��id��d�   � 	 �     [dȽm�i6y@        m m�    m� ��    ��kpH��  m��۰ � 	 B�8   �-��`m��l    �  >�  �$6�Rf��[�� @   	��6���� Hj�88��m ���}�� .�8[@-�m�am m��� ��H   �-�  [@   $6ٲ�@ �I.f\��m��� ��� l���H8 I��� 	ӂ��   6���  �    �6Zm� �-ִ���u-��h    ��lm��m7F�yk��]&�m��`,0M� ��ݸT�kj\�ڀU�:%�x�@U�m���@X;m��G[Ub�%Cmv��䀒n�-˷M̓n���PD*���"����<GAD��` 	���/+T�G�㠂�G������5� #QQ��p�P|5QB�Nj"����THN� *x�B�k��b���Az�z�!�UO �F(<@�T�: ��(Ċ@Rt�a"����U_�T: ���T"�_�Q}PN A@F�B0�@acB$ f"N���"��T爨GAꎠ=D��(|����	�+�@�(�z|�{{�C�*�����^�Az���h��Ϣ �!�߸	��=����20��JG�8=@S���8"�8A�tQ�x�>U��*�QF��EEpG��8EIj�X"�G��&�[D���rN:���m�����m���[i�Gj��f�H ���<��v ��E��`��tb@����|�;�,����yRMhb�����/]QAtY&��!��K�A=)2������I̦nH�.3��)�,�kj���Y�:��{C�Xx;�Q]U�s�%��O.�t�Mס{S����!�Ɩ.�W�<c�ɵ�!� ���χu�`��yn�p���v�s�8\ �ѻF�u���|�O�;u2�;��{[N�ӌ�t�f�mi6���g��<�Ͷr��R�؍�J�S*�36��X���.�7VF�ljX�-�I.�4�e��	���E�n�OHR����uӇ�[�&j�sDí��t��JKӤ����p�<K(�6�P�F�KJ��#۳�=��T9�7���7`֙T���ٍ&�[;V��k��5X�JK��U��D�q�Zi����i��b�˻�Ѹ��ݲ�"�� �s��	`�7ddɶ�c"8�����,O���gXy!�n�mٜ��(.��MZca�S�v��v�'J��(�Nى֙v��U��E�#i6hҌ�J�R�*�+UUqŵ�ր[@�[%����H����K�nYق�U.�4�R�51�-��i�ݰH$��Nel�� k[�$�d`%��B�͌7td�]�ݫ���i�b ��;V�a���s����Hz[�v�^�S����b^������j�)s�1ڤ��H���'�c�tM����n��l���u�PnƹnvpYvf
ܚ�	z��pd�85�+��&Bq��ΤA��X�uǜ��ךլ�m��q��LC���U���f� �Mp��(U�*�U@ml� -���k$��Hd�Z�UU��]�HK������r=p��T�UUEV�u]����4��dI�uP�z���1��5o� ���",�F1TP��T?�u5 �(?Ƞ���x U^�Db/۝�f��'�L5��v���'\�W<�d�m�)�g�a�Zۮ�,�`���k\��nDz8x�lh�ҥch�S�Z����g��Z[��	��n!�P5�9^�����������G5l�X����:ѡ���h�=R���"�@k =���=FgDp;x��Uz�_F}�O:���:��8�x8�g�nz��f�L�M&�n\��x��D|9�0��Oc�l&vp��<�����w �	�w�� �����\4�0�������K����h�Tӑ��!����/��#���+9�`gV��ۚ��r��E�F�
ň`v�ft������ ;�1U��v�$�6`3��N��������2դ�	؝CN������ ��gٵ`�f�L���a.EMJj��u��͖{���6�su���"��WX�f�V��N���	��v�/z, �tx6J�����ف>�����C��z z��;w�g$�gG�M� ވ�+L�:�N��l`Kޘ�=�o(0=����呅I4�2JleS� �ٮ�D�ٯ�z?����,V��X�J�L	�����^��������$u��ࣱ�\�-����qV摈G.���:�5U+!3��/H6Ѧ�P`Kޘ�=�o(0�T��Z`�m� �� }�7�0��0�"�cN؝��:v�Xٚ��=,���HP@��X�2'Mj�.��w��N��	���e�n�V��wm�o807yA�/zc �Ș�(�� 1eЫ-bCw���0l��=�K�%>��J�n	r��R�i7F���Gwe�l(-�l֞��3�7���7XHl�63iv*��閛4��X���	��n����e������5�l�?�W����?��	�F�V��X�I��	��n�/z, �tx��N�髫L�3 �c����mXۚ�&-��E$�q��TO{����'���vfL�l����0%�L`�o(0;yM�m���}�l�7 =�sr"#��2PM�6��;�e۳�����#\��f�q+49n���v��{��B��NoU��κ�$���SI�r�o(0;yA�/zc ��]�� i���[M�w8`����G�M� �J�&�n���Zl��U�t�����&���w4V��N��U4ʧV���$�6���|X>ͫ�Qp(IE����m��ĺ�<���$v��P��!e�d�����ז׶��\p��uyGbnv-�n/�7jqnmی�żv�m�4�f�\��=꺄�N7�YƋq��;�L���������9�N�
���V]�g�kE��^��m�8��C�p	nH��㞩��͞�ul�Y�p����ͺ@�?�͎o��)nq��l�I�������FQ�����L��+�M���ˣG
��r�7"AƤ�̻Ev� ube+m��p�;y� �� }:<H�j��2�L�3 ����Ӣ`M��"��]�E��-*`Kޘ�=:&�P�;ze`�D�[�ڷct���Ӣ`M�oGL	{�bɃ��7v+T�;i�o8`��Kދ >��W=(�Z�i�H��ګ�g�sۮ��ۮ�K��7��sm<�n.�:�F��E[m]������Kދ >�7�0dQ
շCut�2�s�I�~���pD�Ax�
���/}i�:(0;z:`wr�*U�����1&��0&���މ��].��V�l�m�_�g�t~0oG�N� �8�ګ�N�0V,C���7�`�o(0߇���ݵ��k�܏g�.��	sV�f�#Q�U�Y�1ɶ���5��.��\X�"�oD�=:&�P`v��[��IMQNJh%�`{u�(Q����S׀oOe`������ݴ�S4�ne�`}�͛�fڲbyjQ�M�oy��O=���$�{�SpTR�(U��+`{z:`މ�{z&�p��D��n�ҫtݴ� &�L��0&�����L�a��]W[�ctF�5�80۱۶U�8�ͳ�Q�/m$:���y���,��7���m���0=���ގ���`{���b�Vb+$���K`{z:`މ�}��}2ws�NiL�I#hj���7��L��0oD���K`K�,�e�IT�i�jâS>��`��a<�>��8��}D��wӒN��&+�'j�X�m� �dxں^��+ >ޏ :H��I�mպ�����n�7�쌄Îu$�nj�$���X�-���m��S���xں^��)�{z&�0	:]����U�]9�=��W�	(���o; �w;�.��"����%V鍧X��x�0=����0'U���2�!f$�=�&�:[w�������"V��Ս��o �WK�=�=�|�<����y˅Z���\\^/]����GW!�tq��y7P.�+c�9O�����-y3]c/<�O�a=�rvgY��j4�8(�bW�Ŷd7HN�-˵���N�!qՕ��:��g�c	�g]�gs& ��ڹV�t�d��m(p�j���m��u�=������Ȍ�Zd��1-�� 3K�<�'-�P*yP*
��H�q3�J�.�Yz7V������{\�i���W���s7Ngmvr�v�POKӮ���b�Г�š��e���&hOe`����G�M�_H�鈴��۬^���0&�w���K�2�2�T�CN[� �ۮ��c���
g2?���68�Wi�t��N��m�&�w���0�� ��P�&��5R�����`tBJ#�7����`o��`|�k��Wn�����X�<`.-�k���]��%i%=v��n�m��M���[�6ـKދ 7dx�p�U}a��� �(�i6ZFn���I'�����E����ؠ���1��E�/-U��),I�7��A�/zc ݑ0$��*�"��VZV�ݑ�׽ }�<�]/ ��:v��M]$�l�Հ}��`rQ
'ݼ��[�`g�mX
w:�ID��mP!��jS�M�',g[x]Ε�h�r���۬��2<�D婍$�!�� o������wt�����&�5jӦt��������vI=��m����� %J�bt��ԡ�r�́��j��}�V|���Ӫ���-3���'��>ȿ��I	�\7�RO�81H@d"	�0�O�K�IF� �D� �T� ��PS N :!�_�?��Ͼ�I;�����H��-]պci���WO+ �w;�Vl�rS��Ł�Wt̩�l��N�����G�{��g���Ł��ڰ?(I(�;��|���i��ק8�#����Npѵ�%�_n^��m
2_��MM��M ԍ��7�?o?Ł�c����mr�@�w;��S*���$mJ�X�m���d���gs�7���6��+T[�"���� �� }�<o8`��o)b��:`ҵHT�,`�o(07yA�ԫ��
'E@8���g$�{����˚jYW���I0=�������zc �2���ߓ$���&Բ��2XT�%[W�)��R�2�k��tˣ���vI��s�����X�b����ޘ�=�&�t� ��բ�t�+�t��0�z, ����l�P`N2K,�ċHT�I������7�����}{�`E]W)ZC��)[o �WK�=�%�={��D��,��̴+�J�Yi[���w�`{WK�&��-�m�Cv���]�1[�B6|]�l`a6(�=��v}S9��;vp*[N�s
'�d�ƳÝƝ��X���}F�]�g��a:!1��M�^���b����q��m���o���Ǘ7	9�9)���PRM;v�$�r�m�+K';iݷg�gV|qp���MG<i��{2F�;ņc�9�Sm������a�df1�������	+�)1��ܻn���wN}���%bS�Ϋ���Ǝ�$��#غ�i��������c ����llP`tγ f*�Y��
���{�`{s��=�A���E�}�ƚ�i�mU�t��o �WK`{�� ���D�:�BZ.�X��V+�V��E��0��/ 'tj�[�4�պm�� 7z&��0=�%�="��s�*��<.�%�5�ਚ]X͌<�-���'Jt���m�/&x�WF�����Ͷ����0;yA���D����Yx+�M��n��c�ġ(��u�`��`���)���sE*��3-��T��ϋ �f�:&�QF��;5�m�j��2�L.�0l� ;�<w8`H�w"R��:BWx�-$�;�&�P`zE6k�9DD��t�d��h��:I�T�1-��i$��p������
\�=6�I	�*�9���Ӧ�m��~0�p�	�< ��v)�˂��N������?6G��;�0w��ʧEJ��r�`��`����(I*J&(��;�=,n�,xƶI�j��2�!f$�;�&�P`zE6G�n������M��	���:B�������`�����/���+��n]���n�܌e��by8��uk-`�������MT��J���WhDπ�y��	�< ���	��m�*-�-Zhh�L�	�< ���	��}#�܉JQn�	]�@�i&��0'r��(0	�&�(���U�А$ZI�;��A�/d�+ﾳ�D�%J�yr��`��1$0="�^Ɍ��`N� ސ)U�L[)U�v��m��Ak\-����5��g���ӵ[����Uչc����m���y`oG�N����[�JշE�*tݤ� v�x�P`zr�^ɏn���.Yx+(�)"����A���	{&0ޏ ��
�t˻n�j�0�8`�E���_���{��閯�C^Ɍ��`N��8`o��&��c�-�����錘Z玸�jw4=]U� �&�E�u�>|ȇ��l8۫ct�g�4YNd���J��]�Wg��G�\�^�����..ĺ;��	���^8w[�[����[�=5V6���t
�ZC���
l��@��n7�]ƩP6l�
i�lC.�����UT�v%&�MmhΝ:�j�U��t�wwi�7l[1�;]iyxW\<n���jx�;��W*�c��2�Y�	�kk�����ks�r��OG�N����Xz��X��~K��j�.��HI&�P`zr�^Ȱ���
�(�"S)!һ���?�������� � � � �Ͽ~�>A�������>A����{�ӂ�A�A�A�A��v~�\�f��]7v��>A����}��pA�6667�w��A�666?��~�|�������ӂ�A�A�A�A�����wKp�i�s78 �߻�x ���?N>A��������� � � � �Ͽ~�>A����M�~�76�ݙ�+��@��k3���^�qsd'mj�Z॒�`�[��gMg�}�����wz����{�ӂ�A�A�A�A��y�pA�666?��߳��A�A�A�A������A�A�A�A�����rL��[wI�.l���lll}��~�|������"UP�T8<D$lly���pA�6667�~�>A����{�ӂ�A�A�A�A�~��L�.�7.nM�nl���lllg߿g �`�`�`�{�o �`�`�`������� � � � ����8 ��g��l�v[��i�w8 �߻�x ��w�� �`�`�`��������ll?���������A�A�A�A��o����ۙI�!�77x ��w�� �`�`�`��������lllg���|��������|�����s33ff��Y���Š\k�ЫӮn����ˣ<�G7e�J��&\��rnd�.�����lllP?���߼��}�����w��pA�6667�w��A�666?��?N>A�����w��3a��i4�ۻ8 ���g"?Ȩ�C ��A�A����x ��������lll}��~�|����~���˗t����3s��A�A�A�A������A�A�A�A��y�pA�6 ��D=C���<���?s��� � � � ��w�pA�666?}���	rm����nn�A�666?��?N>A����{�ӂ�A�A�A�A�������lllo�~�>A�����s�nL�t�m�&ٙ���A�A�A�A�������lllo��x ���߷��A�A�A�P��y�y$������\og�����]�^3Z���8��]u<�X�96���N7W���v�WLѭ�?$��y��u��ztG����3k��H�r���
d��}��d��Łۯ� �f��=�=�Jm�n�Mcm����=����Q������o~v �j6jV�(uCU.�,:�v�ټ�=��1$��D$������E0B! ?���?��rI?���h����R��ܶX�5�������O?� �s���~�$��j��[t���ͽ;V�])[���Wq6[7Xt\�	ѿ]_����V�uv�*tē N�x�zXn=?(�J?%�?o~v�t��&�r"�T��n��c��B��ݯ� ��v��w�"&L�}5EUKL��hrU2��k��7ٮ΅
d��vf�,�ժ�Ii����D�2â!L�o; ��v�������Ł�G�̕Ls�S%�`��`r��;>ݯ� �f���A���B A"B$"D��H�Ba I$aD�B0 0"!H+j���aD��B	��HFB, D�)*�,��$��e��B �a���$,�&� �֭��x,�1!	��A E� �l:��jDLd��K���I�[
5$F�� �0F�"���[ H�f�p%����V!H ��/ !�O`�h��'�a �E@���H0�U�H"�B0bDO�g1D#=�Ex�!��P�h��H�D!J�2�3;��۴�6���Q�&-�l�����m�E]�"�Y���et���b�)u�I�r��fۘx.���D�2\��Eu�r���E�[+�7F�i;+�l��� T�S��Zɳs�Z��\YgRA���D�6ڒ���$��!UȸT��.�m���Z����c�0�� �����nO���T�8��׌�K�.�L��jV����ƌm���I��� �c�m��ѥ������|�@㓵�n��bwQ�A�y�s�$���q���LWm\�<㮫��2m�����$���l8�9�ݹ�P����d�f��ۃm���)��[�m��"
䞅zu]�9]���]Vz� R�P�9�<1ڝ�,��3qG:�A�z���ɯS��;]��v�&fF6��8.�%�v��e��$.ۈ9���3�a���!��&��8�3�WM�RK p(G!I�-��78Ed�B�o��ݭ�@u�du��l���k��]&��h�H�h�e	sl�Z���2	WK��� c�,d�����ܦ0�ԯ+���������U��B�m86]�v�h�(�iY[�@��v2�qV��f0�@P�YV��@VYZ���r���� �n�m�N�v��T����Ò�P�VR'6���P�㈖�j�U�Z� ���|d����5��Wd�bX��PA,uלG.�;����6^G���Jkt�ɖ+�HK��{9��,8`{�@��wB�UR�JBSDWe��հ��6�vK���lg��E�]Rc9H�r�s�c�fz��SIWO/n�D��&C�6��gEg@�]�EYױv �;�b�p����n�Ų�6^��� ��j����f8,���]UR���V�*�P[*�*�Un8�Uz��gn�m�m7Y&[Cv��l��һ�c�h.lb�
�T���
�i5���ʧ -��=��ʹk[-��g|�:���c�.[Ҡ�p���tC�$4ED�a�&�fm�f���w0��rGRq�NBMcsVm��M�v�v;e�La�w3��Wn��I���^��C���ѷ���`��m��n��o�8�A�q%�*��,��p^��G�݉���m���4�V��8��Z��l�ҙ �m�=��З�Y�c��p�H+��%P���rñc��\z�u��w>�4��M�*���蜳�ɡn���=�����o��'j�0�V�crۙe&���+,=�]���)`tg2��=���>|�i�N��lm��~�ۏK �f�I%���r�uT�d1�T�l�=����D(��D(�����ߝ���K脦C�w&U1T�R��ܶXgs����~J*�w?Ł���,{%�U4驚UI�USv�L�w;�_���{7���[=J��jB����7`n���L���y�oG�uoL��\�f�p��Rv�s	v9�['���uA;��n�lR�P�Ⱦ|T.�-�e���/� ��0މ�7�rT��KcN�D�2�7ٮ�6!�J)(U_U:y07�A����$E�RE^*E��oD���NP�	�<该:v�N�n�o ��	�����c ��0
�*^fTG�Y���INP`K�1�v�v�=,��Ʀ�p��*�P&�[&�m��n����-�r�]�h��:�h�L����VZ���I+H`K�1�v�L	ܠ��s����R�Ӣ�+�MZM`oD���NP`K�1�*����;�_�����uce;m����>���ДBj��o~� �f�ٯf�UL�E媼��CӔ�L`���e0:�j��144]�`}ր7�Ɂ��NP`&B�B�ۜ�Cǁm�%і�Qfp�h͔��R�s�6n���լ<����=��o���w(0=9A�/d��_JT�Ĕ�SC�.��7����2{��`t��X{5�(��]�2UqS:���M��_ϳj�I)�sy����՚�T�R�J��r�a�OVoU�no;}�K�%���*wߋ���ʦ�0�Wt�I� ����t����/z,�zZTe![��ةZ�մ=���&��US�S�����msv�!m����.�e�J�H�i&�P`zr�^�������T�!�.�unę�}9��/zc ��yA��%K0-'t���v��Kދ ;z<o8`Np�7� իO�;N�S�� v�L	�������L���v�X��B�k`M��(0%�L`��`z҄�	!D(_�U�M���v�.�u���W�t���{=�6��7Q����2�8�R����U;Z0#�@�d�u�&e�h��z1p(�^�ƞ$�)-\�N�����Nv`XV[r�O�ga�+����[l��m�Kla��j�R��z��-iqoN�����.nPS�q���Z8x��-�	��/U*�V�@[+m3;P�5�&X�z�U��^s���3[�36�v$�y5sn��[��-6�v�ݳ�\�7
�W�FKѡF�uCU.�>~�gٵ`����J"c��|Xr�b�b�j�KM�l�6}�W�$�Csy����>�zX�:�v��-U�:j�k ;z<o80=9A�/zcw(����*�"���yA���	{�oD�ގU�i��MX�0�8`���ޏ ��r�e�I���t���h��띤6���RT��G!����]ǒ�k�w|ӬBm�!44]�|��� v�v��	/�39�`f��2ʪi9T�S%�`���I*��_g>,}�����QTgW���&��S@�����X��,铳y�gs��]�e�Ɛ�[M��p�	� {ۮ��P��o� �[�ULU-T�t�$�7�`�&�P`n�m����qy+i:u�i){Tm��]�
�l��l�\��ջt�n����6���#3`�&�P`n��"`MTIV�N�Uce;m�9�=���������<z9E���-:��e��k��3ۮ�	*�>ICf�:8`rU��[�5i��-!�M�0�w(0�U��~�����n��'@��k 7dx�p`n���˒�.�U��I>����.�˺�D�r�n���
���뤄ΛiӢ�cwBt�7�N�v8`�E��< �"��1��˴��݊	{&0�w(>J&C��2Jb�j�KM6�`���7dL	���݊ӕJ�ň/�i�T݇L�w;�_��KP�TN�ss��I;�}/e̛�Ʌ��V�`M��P`z&�"f�߹�Ｌ`k2j��$���ɸ��k�w�Q�^��3������݇�7[�fb�A�M�쉁7�rU��[������z< ݑ����=�z_(��7hޑ�T��AL�݀fw;s�tB��Un�� ���;쭭MM��)�˗M�t��� ���K� n������tƓ�4�0��z�t���y�{^�DD(J~�
�e�n�P���z���D�ɉ�y�{Fm�{7H�\닋Jmlk�Ė6�_]��\y3[>݌#�����knp�ZY�Hno���)p�<�%�L���fc��}�3��}v��̈a�c�V�q6�;f��{:�@�*��z�Q�7���!��z먺س8����f�9W�wez3�����RI�pS�<���n�Mֹ��W:�Kn�O���~��6ܝ<����[g�"n+Є�۰��������N�&�͑ͅz�+v.]uV�������7��`�νe��Z��tēx�#�>���*���?�<�	����l�UݶR����A�n�LvD���;%UIM��iҚ�X~���ŀno; ��]�(�v�mu"z&Zc��C�i���vB�����Ł�k����(�=��,(��U:����]\rʵs��\r��c�=��6��:���YUN�Md�� ��vۏKv8U}a/���yz����ۗM�n=,P��B�Ir�e��������z��+�"�MLi;I����ŀg�]���	U��;?s�X���(YW��T�C�zc ݚ�����ξ,�Z�&�s3HT�I� ݑ�������~0�����~����u�(�6k@�����k	��@���qs!��Yۑ֛5$�׻�ϥ�ܥ%E����{���0�迪�DB����ߝ�����&�)�-:��ؠ���1�nȘ�A���΋ʋ��Lj�CE�`}�, ݑ�p��@$ @�d@$`@ 0#	�$�	 B,B�X�B,"�`A���E$B)�� ��=uV��@�S�I�A�|FD<���`D E���h� �b�"	���Ƞ-4@5�WA���. ��*UE�(|��"�TMs�C���uE>U'���ﳒN�>,�7IsUN�MN[��3��<����0��`r�S��i�E4���=�zX�||NwU��L��`d�rjf���4��\��ɛ<7b�(ꉍ�u��P-�yDӞn#�f��sb��4��i� ݎ�Ȱvk�Q�g>,�ˠm�t�T��6��ɌvD�݊ؠ�햢�n��
�5i5��<v8a꫾�?_{� ����줨�O�v(07b�od�
V}��&lw.�V[en�BL�7c���c ݑ0=�A���L(ً�̵v�@�W�Z�&i���������-֋&�v�Zhh��oz, ݑ�=�A��2\�Wy��v%@�ZX�7dLlP`n��t��E)Вt�	�64���v8`���� *H$����4����A���-�nȘؠ�=%O��Wj��*Đ��ޘ�7d�I<����'��{9$ @�$մH1
�)E�Q3�ɤ:m˻-̱��u�V��$����&un�#�b�S��:sϤ�w���{Z	�[k"tWN�a���c83��mZ��Ō���bvMgU=�8�]+�˛k`�{u��GC��|\:`+��{�i��T��^�
���aY�*�1�$��h�5��V5 	��#g����#�p/9���M)99����,���r��sC�`�b�.ڭ����>O��Q�2r]nNI��O@g����J�r�vto��=Eӆ��Tēz�w�������y˴]�e%E�����8`lp`� ���\�����.�,��C��D�7z&�(0>���閭44Zf n�x��0=�A���.ZʼH���H�� ��ؠ�����3m����AIڛ���2`5� 
6�6VX{f�gtupѝ����k]����$$��ؠ�7z&��`I�rՅ1�`�������P�KU����7~�`��`}�z0	�>���J�$0މ�n�LlP`{b�l�Sĕ��J���0ڻޘ����8@��`v�.�v���]�����8`lp�ޏ 7z<�WO}MP�	�h�QC����Z˷unLbF�ݷ,J<�]X���	)�]�'n��l���T�g�oy��ޏ 7z<�ܥ*��t�V��0މ�n�LlP`{b���-���J�۫-�������N&�0�F��w���rI>��))����R����o �c�~���]ݝ��www{��wvT�/1��g�W�1^$���߶8{�wgtt�����E�]��������g����ݫ���ԷZ�l���g�n.�����vM�H�k��s֞����W���몷������ww{��ww{V����=뻻�j�a���Y[�������� ?~�c�����!��wd��yww~��� �
j���i/z���(�����p������0 ����~~ ~�}��/b�`zxZ>L�U{;�>�fd��N�ff}����2BK��77�ݼ�����e�e��f�x�z�����ݑ{�ww9En�����ϻ��}��sd�d�iS<n���0j��[%ƺ�g�u�[s��$�<��5��Պ�� ~��}�? ����?{oNJ=ꙓ��;���k�)��M1J���^����Q[���lp������� ��~ߟ�������>�m�j����z��'www�"����b����ܝ*���U�j�$��]ݝ��www{�/z���(�����p����e����=����| �߿o�����>[m����-�}�xo-��E:+��m�~n��N��^-��u ����b�c� �tq�u����n�v����q�]��ѵ�/�n�,��i�6.�S1�^�1ι��ns�.LQ���FzB�Uŕ���:�=C\)��m�������ʶC�2Ptl�)��F��m�
��M��@��=�9��R�ae{:{m=�l��a<�����@Qe���.V�"^5��=����|��̻\�`L��aTZ�IP��`^���Wi,r�뭴kl�C)s�m�7�������G�����{�wd��;���ދ޻�ފ���QiwyIU�%n�����޻�'GI�������� ��}�������ˋ�e�8Q�]ݓ������d^����Q[����������]�4�A�~ ��޻���+www�=��}��~�c����xN�	�;�o�	��0�2�vG�E'�7v��v��m��it�����P�+�ݫl��g��g��6�/WjӵIi�v���� �镀�&�0	$,1/��v�RI}WUv�&�07b� �_T��MݪV:bI� n����v~S9���3w�X��7�!K����ZI�{�Lؠ����nȘoK�-&ʻ�M�&���ott�7dL_I��3�RWk1*VF�ӏk�� p�N����1�sKĻ�h�=����L-�,I��i��L� ݑ0=}&07b�_L˗b�t�ժ�"Ҧ�"`�g(07�:`}���Z��
Li� ��1�g%�����V����t�t��
�x�,ēg(06tt�;dL:""gs��v�mêEL��6�wGL�D�&Ș9A�+��./%v.��aӪ�ś�l���76	غ!�v�nm���]t�u�L��묭�6�l��vȘ�A����N�o쥔U�����I0�v(06tt�7dLoKaxQiwyIU�$�݊�0� �0'E�R���e�;-3 ��+ 7dx^ȹ&�E�<��(��wy9$��za۵��]�UbE�LvD���1��::`I0��T+	fRT�[�N�n��C.���ȶ-���yB��uňMu%mQi�B�o ���0�2�vG�HH^4� mU��n�{^�ЦL��V���=��gJ�I|�T�$�Ύ�쉀}�<v8`���6��v�v�SV9���=������`{3mX:忋E�Z��H��� �H��A��͵`��1%�B� A" D@�$��"��	@���BHH1�ஐ�c,E �b�"�	!��D;�O��jh�Ԋ��H#1 �@�J}���=qT؈������SĀO	R0BWC�>$�`F!K�x �@�� B"�* ����
����"|{�{��
ЂA�Ib��R0��j����n�[sPjڻu�=qb��)�:��g�'<IGSuq���m�����q����b�v�2�5�E�s�$�<�v�Ӕ��m.y+ap1�4��َ-I ۪�ヱ�Zz�q�';��1Ե��L�R�7j\�Ub��;�n��ײ�U]����DW�wn�W�;XGG�	� �lF�/�f�+���9���L�N�q�
�"�IQ�5�c��kv�%3�h�[�X�ܺ�,q�v�Ι��<�g��9ݶr�����9��q��mDl�㮜u�ܝgd��v69!�]X}B��pt�ŧ��P� �&��9����ld���NC��"���� U^ֳ�8sq�iϓ-����AŚ.���^M���v�P�#r8ګ]�G�����͜�&玴�WXòL����u�W5�s�g^ƘץƖ�u���C3���¤��n�:2��b�2j@�pkQ���-����m��$sS�d���i-I��5C���Wse Κڞ]��<�R��܆�D"��<meW��v�C��w)Ö�ef�r���L������ձ��9m�@�B
��7�-������\]�R	���2IzҀ��@�V�Tej��ͻnr�v� �	��ˬ!]���U�샭D�S�,T�[PkF��U��3�ӷ,D���pA�%�A�l�T�V�V�N��%ޡ��ګnW��m)�gk'��,�SH袳m��:v�&�,bMw-�d�[����NЧEa��2���u3��v�#�w�d����6���ʹ�S�Hj���,cv\�P�C^f�eM�Wq=��N#���ғ���v�7S�J͎�>�v��Wi�n��͊�zW��h�p�Xm��Uu$6�yIٺ�����X
���*�ym"���6��e�l 4�I�K�M��ji]ڷ*���� �4W��6mtT:���-����
���!�nvz�sY�f�d͐���H�i�P5���#ɫ����=�.�Lٺ�jB�M�.���r�����cArq�w4Ź���u��5��X�u"D�,�"N��c��k/pɝO��c�ˮ��6��Ϧ�"*m��pw��m�����I���c<�G(�K���,l���ڴV��W�5�v��d@vV���zC���\�g:A�n�^@�S�ũ#F���"�^�nd��)6�A��d�j��b�N����9cR1vz��3hf�ٻ�:�4��' 4�5�ww=&i������=*�Ġ�A���� ݑ0�ti@H�L�i���0�2�vD�;dLؠ���T�X��ڵV$ZT�7dL�D�݊�0>��-�-?�V�RcM�{"�7b�gGLvD�����V`%�yJ��K�A�����"`v���������k��]���Ē6l�B��n�l����Ǟ�N�8(���a���e۲�I$x�?:`�&�$��P`ND�Ӷ�ЬtƓ���o��Q�H�P�ѕ[s`{���=����Qd��b(�]պ���M�n{� ���GL^ɌoKa���Ee�RUy�07yA�����jL`�&ti\�+t�V�-3 ��+ ���X�#�7y� ��q�J�����u���������K��U5c�w3��f�ms��scLtq��6߇�}����<w�=����V�K�B�?�n���ʧV��w��L�|X�֬�jE�HIv����V��i6��P`l��UUKﾯ�={Rc �H�nj�昤�4�m����6����<w�0��Q�m'v��R-b��jL`�&�(07d��6��Кn��j���n�.�j���hU����Ά�gk\�4ȗ��qqv�+��Ɍ�P`l����E�}�/(�6S�T݉5�n��nڰ>��`z}�W�"!L����U-2J�#�i�v���Q�VtDB��M��`fk���͢����2�-*`{p�l�����_W��ꢇA	����y�v�K�f�1b��b��"`n�gGLm�`rQ���&�]US&�	r����Q<>�&6��78��ȸ��qݘJXe�L	ؘ6�o�;��l镀}��`l� :t�4�@�P��m��6��I%'����s�������F�j�����u�}��`{u�����|X�֬ܝ��L�T]�X�0�w�::a���g����@%�l�v�����7y������	1�vȘ���WW}}��w��u΀�ā����(q�y�92���lQ��N��u��([�Z���ѥ�6�nE��s'6�[(Պ��;Ia�p�����M�^9�0WJe�:݋C��e8����b#9�\p U���Ӯ�$�Eb3���b�P��q/m���]�h
7`d�H9e69\�8q���9mp���*�C3�v�;s:�ڄ�,��O׾��4��lEg����Ʈklnҳ�F�GV�1�O.�FӘncj��iX�+t�-0h��t�V��E��?W꯬;��K�K�s.Z��[Vޣv��D(���`fk����ڿ�BS'��檕K�:�%$15���n������ڍڰ1{$�iMIJ�j��(Q�e�`w����, ��N�����4�e��͵`r����7;���$_�.բۺ/�V$�n�7'��N�z��'�uѻ-ɱ�M�l�uZ�JjM1�5`}�[�`��`{����(���(��A�����t��)�#S3M�+`�&����w��0=�����ȩ�>���d�!�vn����~_�������K`�&tY�j���3-�d�,:!(S���=�������_D)wMwn�H�-��*ݛ�%
w;��fk����+ >�R�Ҷ��6�	6&��^�d`�n��2�$nwi��jk������9�e1�줊i� v���p�6t�興�C�GuX���Tڐ�S�I07yA�����	1�vȟ���(K�(UA߻�ӖЂ�!��l�7�~�`}�7j�""%!����=,�R�M�-X��N�=W��y`�y���l镀t똊.��n����n�=���;>;zՁ��ذ��IQ��ؓtJ�6~�Ղ6���q��f�[V8�vn^���P�4�s�� �����7y� ��+ �Q"���y�y�g�նUݶ���l镟�$���GuX�s�=�z_(J""d�ޣ��Zc�rԍ�ڰ=�wU�g�S���0=0�fY���������vȘ�P`l���ꯨ����J��ߪ�7�l��e&��$��P`l���æ0�߿K��N��v�n�mE����]�8-�7U�ݗ���vn3����Kj�q�Vi�tv-!�������;dLw(0���n�j�N��u�}���G`}���=����Q	L��=j�)Х����n�s��f=,脢&s�����X��]![e+�Mդ��c����ڰ>�3já%	)���`n󪓔Զ)�l2���ڰ:=�ޯ�7;���c���0�#x]b|�S4�:���o��^2�r��P�wNS���t3�Yr�n�r&�)��dÈq��&7�G;ۗ=��6������ד$Mȕ9r͗Cn2�u&-C�lD�Dd듀�ճ��I��MKe^��t������7B���lwA����IZ���a��Yy�{<�hx�ý>m��eٸ��`����FY�͘���i�\T�,sD��R���ݺ�盢�LeU�*�%Y��Ѭ��!\�.�q�-*�0���vȘ�P`l���D��'LcI�IM`l� ��A�������$:Ya��䌥X�Lw(06tt��a�l��t�yk	QB�J�::`}���G�}��mu$�'l�fR�,�Lv1�vȘ�P`l�`b�Ҩ-Q.��j��L�i�&�y��*��B�ܜ�	/5=l�6z%�Yb��Y���B�0����0=���N����@�;�I���'7���5E]�f��$�����G��$�J�X�ʻ����0�?:`{���D��r���!e݊���Պ��Lv1�M�0>�zXtDDOn����Q�.i��TUS����	�<߫d��=��}�ͫ��~}ߡ���l���P���I����A5��ϙ�6uݠ�̜s,��~����Y3�ة�i6�	�����N镀}��l��t�/�(��I+H`N�}
d�ѽV����H{u�`Ū�ye��:n�u�}��l��~�P:�@���8*�J'�@���W=�F�`[J[d$%)m	IXC�̖��R���E#="��dh�E�#42���'ނ z��uEz"���Ծ���w}��w��V�-�TRtH�f�*Jua�"g��&ȿ	�0=�t�Ύ�]#%���MSvُK�~I%������#�� &��	��SWm&�t;�ŻN��d�;�V��L�cM��o��[1*BJ�b*��CL�'t��>�tX��|�"��|X9��a,r�8++J��:c �"`{�A�;���(IL��7�m�c�r*����=���>�p�'t��>�tX��w!L:)�:�݇BIO�o��z�$�}���$���������Ll�b�ETP�%i	�0=�t�6D��r�WgJUj��Ec��n����r�b�N�I�K'i�Z�[��7�R>��m�UUt���nj��m��&Ș�P`N��;�c�2Հ�f�*Ju`��|�L��|X�֬�6L���-��1�ZM�w8`�ea��w�� =���;�J͒�jI�L���(S۽�=�o� M��~����V.E� �C�]\�[V�FmX��������|X������%*""V�L�4U9:���N��k�Mg����g�ۍ9��;j��H7bv�<��½r���;z��\v뱸��e�;�Z2��ڻ5nJ��x]<�k�%
�F�;��S��+�4�u��u�Bڕlc���fY����5[n
g6GO�c@\'PU90��m�2�ۋ<����v�;W4(�f��Z��2M�6u:�5�m�Ɵ���{��ώ��4�ʁ�N��ذK�bŻ5�9V��hݲ�ç2G5]c�}�>�}�W;6��vRC\���<�镀N��#�m�`��̅4!:)5N����tt����݇L`z'��Y����U_��4ۚj����Ձ��ͫ�Of��n�� ��Um9�3T;Y��/rT��t���0'uE������v��� v�x���wGL_WL`m_O�3���+�q�⣧<ю�Wb�!5n�j^;%���C5\�N�T�m�	���o ����'fڰ=8�k�/���`n�]HUMQ#`�M�s6��}�/�B��~�|����>�2�����v1!���u�o#��	�<=��g���zOe` �i��vRCXߪ��������Z�73mX~��oU�o�I�*
Xe*Ř�`{�:`N���â�	�< ��bC.�T;���[����Є�ۑ-/�ޟ}���<�5ɵv��l(tӴ��='���:, �#�;ze`�]bR��wj�:n�u�za������S
�J��f�)M9���3ٶ��(Ws�t����l	�@����Pb�ē�GL�06Vt���`vk�[HT�D��ڰ>��V�G�=��7y���VDB�Ξ�*��ٹ�\�/[0��N��I�W^���!��f�ؽ]St�V2����m��s��> l��0;dt��a �/`����+`:&oGL�0>�Y�}�)��;����C*i�2������GLJΖ�6tL��ȨEAB���S�GLJΖ�=�������P�%ni3Z��.�%y����-�l��03۶�K��]SE:ne���(���/\�@<A-�GV��51Hqk����-s��L�E)�? go;=�j��nڰ>��^68t�n�	�������GLJΖ�6tO�}�Va'�WV�Aj�ISg���}Ը`n��7�2���U��ĭ[�n��>�Y�`��`g�mXtDD�{�V��G�$�i?��&����;ze`n��6��
���f�h�e^wex)Z:�Z��:P6[�=�a��$^��z�,mn�'�G1�'���g9㛜�I�gXm�M�I��Г0���r=�m�^�K���tV���64F���,��]�i����즦���w6��U{	1k�Ji������o&�=gII�:Ӌ��m��a7�ѻV��9�l�-�k�,�S� 	7v�ɒY�on>w���M|�U����;"S�t�;Fg[�3s�o^G�rf�:�a)a���{�V���c�C�t����z{�X�L�莋 �� :JJ:@�:i�u�zH��L`u�L`v�t�}�W�]���ם�@՗N��u�o�<���?$�BS;�֬wu�=�۩T�Ț�i��N�:/Д$����;{���0=0�	�J�����ui$����6GLJΖ�6tL���&�qTəjS��i˒B��04�k���i�x�N�O"6��ޫ���w�ܭ�D�k�J����t����lgD��镀m�Q�tեj�N��XҗI�[
!(l9����޵`g�mXr.T���1��Ċi� l��ގ��:`zVt��L�2�Tˤ�2���	(�������`v��j��#��뾓 t��`�:(tӺj��nڰ?%	$�%	$��������3ٶ��q��Hʔܒ�(*i?:�ݰ8���z�:lm:2]:�C��&��h�.�CTU�:j�u�}�`Ώ ���������ʵe/��Q�b���w�	(��szՁ��j��hͫ}
�XZ�Q�WKLގ��:eUW ��Q/�5�Q�":BP��Q�U�go;�ʹ�S4؋�J��:`za���+ ;z!�n��C�����ڰ?B�J?(I(��ߟ���֬��m����Bz:�"RdjKF�q]�����u�7;�_GEk�sK��."��J����73]��͵`o�mt(Q��'� OO
�+�@�i��i�����0=0�	}������'r��!�K��ӧ4Ձ��j��hͫ?B��=;�V��� ��N�� n��R��T��æ0	������? �[����w������YJ��T+1c ��0;z:`M���GE�n�Tb):��ۿ������mLgv�NhК���4m���rlP�b�e��	
��I����l���]��%��y���cj��%0`�V����zyoU�nf�=�j�BIBJd7;�F��S%UU����X;��;WK�>�e`r.T��le��ĝ�k ;�<�t��%���J�W-��]AT��f�b�Ę����:`z�t���rH�ȋ���'�5��@�= ������KBR��R%m����]ה��p*�3_B�`�4��hF᠐��"FPRdQ;Ͻ<��w6�@V�2k���G��b�ɹ��'*.I���	�@ �EҌ��[�%�@z	��ke\�L�]����r��:�[��,�=�T H��t�Ӳ7a4�g%��L�:Y��VR��XD��Nt�O�����o'��(�muXN F.�m����C�:�p9(����t�v�b�[�F�mˍ���E�aϜ��f���5�ٷ0���2b����ǵ���Ξ6������t�[��LZ,�Hl�>y�5e�j�tɄ��+Τ8zH��������<m�(i�u�]� n�,XTX6�F.,�vE������S�E1l�9:�ƃm�ݸ�Zu5[��;�gk85+]жg����u���4���]Z$3�5�Z.�mI�vv�;p�k�]fm��Cp*��&��I�96� \i���4�,��:ݲ�I8� �ap��,\�p�^�ي��(�uPq��uk���7&���B3cll��	�;F�9�P�v�8S=���1<�D" *�l�m���K��vۜ�h�y:�O���HE��p�uq��e�V�9����� @T�[O�ݔ�ӕ�v[Ú�cWH�R�*����Tm�$崶����N�ݠ �e:8)�\��j]��U�X.� 'l�s��j�ܴ4P�[RM�*��� �#�mmZӡ!�BCj�m�v�mK��UJd�o@�v�G\�1n4�nm��S�i�=[q�$�m�O7ZmZ�@ ���'PS�pt��ki[F��]�vU=i�<K�WT�5;ݺ5Y�,�x�h(y�s��Շ�d��A��yyj�nd�B�Qv�.љjۧ�6��\�ێh�i�KRS*��kZ)�1,�,�m q)]��^RS[t�H �U[��-��"۶���n۶�4�km  3'B�R�wI�K��s���m�e8	��.M��4������p��%��@sk7K����I�̔������J��A��(�tC��ɣQH���� �@��"�s�;'�3L�vm�H%�l붝;
Ln֞GBu��L��K�Nid9x�qy������ӝ*Gn��F��%�k�Y�����jt��-�W����<��D����xIm��[�q�nz϶��V�����x9P*��Ěv1��TYM�գ�;\]Ι�i�*#������Pq	���ke��zNΫ(�n"��]]�P3�`�Rڮ�}��r-�	�ۍ�x�P��mv��gm���c��u��h�7=Y��7-룒���9������ڰ���B������ $��N�aM��:bI��GmXfk�3՛6ۻj�!(Jɹ��R[��Yi��M`�� �]/ ���ҳ��;b�WJ��ʄ�ui�a�D%;�zlwu��U�6�B��ww���޶6�i��S��I2����s���� �]/ ��*�h0��=��"�u�3rBk��gTU(��笕�*�2�w��{����|HӤ2���5M|�V���5��͟Т��6{�X�_��:��N�H����D���Wܾ�6I��`n���Y���	%2wj�J��s,��ʦ�ʟ����ҳ��t��B���e*V�+`{�t����l{���$�q�M�v�MU0M���*�Sҳ��۝-���W�߼�|����!f
�fh}]���9U�$>z9�qLr΄�N캵E)r&��hji������Vl�f��
>��*ޛs��.�m�=Y�`zH��Y��wD���U]�'�EM62J`�[���j��hͫ<�
�W�]ں^��-�Nյv$���ڰ�	(�r{�`����Vl�t(I~Jg�߼��'�͓Ld�jJ�,V�;�&nt������-�����P]{E�W^�}(�H�84옒��[�U��Sc.������o�\��6�l�ļ쟭��#��gK`:&�̟
�-}t�-,V���ҳ��nk�3՛7�d;ut�N�&��i�'X����}�`�K�>�2��"�B�vS��:Zw�m�E�v��`}���Ȅ�.:�_w���s�R���`��$��%�=�:`l��x���:�)��ht�4U�ݔ��ӷ"��"�WKm�N��H�uZ<�$$))VX$؋��t�X�]/ 7�?W���x_���N�ұ$:L��$��ϻy���ؗ����<�bX�'{����Kı<����y�(eG{����c�t�V�1�u�=�7��bX�����<�bX�'�ov��KȊC"dO{���Ȗ%�b}�f~ʜ�bX�'{���,�v[�&l���yı,O���Ȗ%�by�{���%�bX��fw*r%�bX����<�bX�%��.gY�.�0�n��Ȗ%�by��É�Kİ�*��ܙ�*yı,K����<�bX�'�ov��Kı4 т�@AH ?w���u�2��ܙ��a��,n���FS�R���$^�����qp7G5�mv컐���8^F�L����/��y5ۍ�WS�rY��ٞ4��
ďU�$Bt��OtvK�ni��we�=��d:��QW��y�"殷�u�v��lc.����OC��m���cM��O�Z%�^Xe �ܻɧ3�I���ͦ9�V���n��[�S��6�9iT16kU�d��%MΝ�����#������묭����oq��N�ٟ��"X�%�~���Ȗ%�b}��lND�,K���O"X�%���w8fYv͖�4�fnT�Kı/�}��yı,O���Ȗ%�bw��É�Kı=���T�K�I}����M0�H۫��
HRAb}��lND�,K���O"X�%��vgr�"X�%�����Ȗ%���읶S
��$�&����$)���Ȗ%�b{�s��"X�%�����Ȗ%�b}��lND�,K���f�ٻl��Lɹ�q<�bX�'�ٝʜ�bX�%��wx�D�,Kﷻbr%�bX�����yĒ��B�9�)�L��74L�ST���;N����Y�x8�����k#�͵l�����mܛ.��fCsmO"X�%�w���yı,O���Ȗ%�bw��É�Kı=���T�Kı>��L<ݖm�nl��sw��Kı>�{�'!��� WblK�w�O"X�%��vgr�"X�%�~���Ȗ%�b_�r��C.��.��Ȗ%�by��É�Kı=���T�Kı/�}��yı,O���Ȗ%�b_����76Ct��ffi��%�bX��fw*r%�bX����<�bX�'�ov��Kı<�{���%�bX�}gs�e�d��3I�f�ND�,K����'�,K����؜�bX�'��|8�D�,K����ND��oq�߽��ﶘ����ܓ�J�s�l�1<%F�����U�˧q������4ͅ���yı,O���Ȗ%�by��É�Kı=���T�Kı/�}��yı,O�t�M�3vYfl�%ͱ9ı,O;��q<�bX�'�ٝʜ�bX�%�ﻼO"X�%���ݱ9ı,K����M7m�2i��3N'�,K���3�S�,KĿ}�w��K���4�,Mϻ��,K����É�K7�����/?m��&3��Ow��"X�'�}�8�D�,K����9ı,O;��q<�bX�'��;�9ı,N��n��6e�L���<�bX�'��w"r%�bX�w���yı,Os�w*r%�bX�}�|�y�q�����L���J��f����(�:!� LV�uٷȌ1�&(�ʍ�3μ�I��swr'�,K�����O"X�%��w;�9ı,O���q<�bX�'��w"r%�bX��;t�͐�-4ٙ�q<�bX�'����@?��-��
�-��$$!^f89�PA?�dK���p̲�[fi6�ڜ�bX�'{��q<�bX�'�ov��Kı/��w��Kı=��mND�,K�{Λ..�&ٛwsx�D�,�
��Cb~���؜�bX�%����x�D�,K��v��K�����T�F" |J���+y����%�bX�N�ܓL��e���.m�Ȗ%�b_;��Ȗ%�b{��ڜ�bX�%�ﻼO"X�%���ݱ9ı�{��w�����6�����������q�7D덤�Q����!Ѳsd��ބ/���/��|����sd�����>�bX�'�?�ND�,K����'�,K����؜�bX�%���<�bX�'�l��wM�6]ͳ&]͵9ı,K��wx�D�,Kﷻbr%�bX������%�bX��s��"~r�D�?~���)̲��S����)!I
H[����Kı/��w��Kı=��mND�,K����'�,KĿ[�됷Zi�wv��Kı/��w��Kı=��mND�,K����'�,K�̉���؜�bX�%�{�i�3l3KM7n��Ȗ%�b{��ڜ�bX�%�ﻼO"X�%���ݱ9ı,K�{��yı,�}����jF�E<:��#t=��K%M��GL�YЇ\���R9� 3pw��N{���r��vwMַ'N\T��8��\�Rjwk:l�Ng�6y6󖶧]����{V�3�43�1���K��ٸ$���:�I�0�Ā�jܮ�z�vwne����{�<�P.�T'-�oM�tB���;p�6:YT
��|�%��f�ղ[����r��л�dIogӒd�%�I/oRRr�Lݮv�j�qk���<�n^	э��0{�7���{������O"X�%���ݱ9ı,K�{��=��,K�۟�ND�,K����32�M�K3e���yı,O���Ȗ%�b_;��Ȗ%�b{��ڜ�bX�%�ﻼO"X�%����4��2Y�M��؜�bX�%���<�bX�'���Ȗ?�!�2%�{�x�D�,K���br%�bX��gN�m���p�37ww��Kı=��mND�,K����'�,K����؜�bX�%��������{��7����73e��Nڜ�bX�%�ﻼO"X�%����"�_߼��ؖ%�b_�oȖ%�b{��ڜ�bX�'���6ʷ%kS2����q�ۭ���b!à9װو��f��	F����_=ߛŉbX�}���,Kľw��'�,K�����9ı,K��wx�D�,K�ol3�B�B�e�ݱ9ı,K����<���h
� � �|����Ȗ'��?Z��bX�%��oȖ%�b}��lND���,K���4͙���SM˻���%�bX�~��jr%�bX�߾��<�c��Dȝ����,Kľ����yı,O����r۶m�L�m͵9ĳ�?���6&�����yı,O߷�lND�,K��{�O"X�%��w;jr%�bX���iTQTԃRS6��)!I
HY��br%�bX��{��yı,O{��S�,Kľ���Ȗ%�`�����^X$c��C7	u���mvjI�v�������nJ�e��_�{��_w�GlK,Λeͱ<�bX�%�߿oȖ%�b{��ڜ�bX�%��wx�D�,Kﷻbr%�bX�����f���p�s.��Ȗ%�b{��ڜ�bX�%��wx�D�,Kﷻbr%�bX��{��y�TȖ'��ۚf��d72�d��S�,KĿ~���yı,O���Ȗ1�x {*a)�����VT�+B��(@!+YB		X�\cF$�BQ�bЉH���Ic �����*�!)
�h�(Jb���	£BA�0# ����$��T�C�E�ͬ D ����0 A���	�@�@�0�����D�H8��eS��E}�Tr$[HB��$"�"��!"�H���감�0�$�B�6���"��>��H#�B��eaRT�`P!�+��@b0HH>"�(�8��PE�����@��Ax��蘒��L���{���%�bX�ws��"X�%�~����.if�̚f���'�,K����؜�bX�'���O"X�%��w;jr%�`~fDϿw��<�bX�%������[�4˻�br%�bX�{��q<�bX�'���Ȗ%�b^��w��Kı>�{�'"X�%����v���kC�{9��\m��ɶ��`#]st��y4�f��r��e��^qvw����,K��v��Kı/~����%�bX�}���,K���Ȗ%�b}���73.ٶY7dۛjr%�bX��}��yı,O���Ȗ%�bw��É�Kı=��mND�,K������M,͗ww��Kı>�{�'"X�%��{�'�,K�����9ı,K߾��<���¢��溁���$��$Ӓ��K< dO�~����%�bX�~��jr%�bX��}��yı,O���Ȗ%�by�����Km�Mɹ�q<�bX�'���Ȗ%�a�G?w���{ı,N�m�Ȗ%�bw��Þ���7���{�߿^���u�ܹԓs-v��8ݦB�K�Dn@�ؒ�}Mf઒hz��������oq����n'�,K����؜�bX�'~�|8�D�,K��v��Kı/��txR�H��*�����{��7����X�����blK�����Ȗ%�bw�s���Kı/~�w��O�\��,K��-3�Ji�wv��Kı?w��'�,K�����9ı,K�~��<�bX�'�ov��Kı/~��M�4�6�i�s4�yĳ�`dO�s?Z��bX�%������%�bX�}���,K����Ȗ%��{���}�T�ڶ�w��7��b_���Ȗ%�a��{�~�Ȗ%�bw���O"X�%��w;jr%�bX��
`�!'
���{ε��HBݳ�&�ܼ%v)6piO	�[�YS<�Ύە6���n���Gl��=���A��?��j�9��mڃc)��#�������skB�Uҏ�:ؠ�Xc�{O��Fr�Y@�jX�-��郠k���#l�Sז&��<9u�u��a��#�hvx-1�)����n��68�{tU����\]h3kZ�ݜ�A�w������=�;��׺��f��uЬn�[6��#�q!��;8��
s���9�6���ߛ�oq����w�؜�bX�'��|8�D�,K��v���DȖ%�{�����Kı;?i�	�]�e���.m�Ȗ%�b}߻���%�bX��s��"X�%�{��x�D�,Kﷻbr%�bX���l��ͥ�ri�.�O"X�%��w;jr%�bX���w��K�2&D�w�؜�bX�'�߿xq<��oq�߿���W/XXܺ`�|�bX�%����<�bX�'�ov��Kı>�{���%�bX��s��'���{��?~�en4��W�w�Kı>�{�'"X�%��=����ؖ%�b}�s��Ȗ%�b_���Ȗ%�b{;��e��Rd5�;���Qn:��YQ�G5GY����A���m�E� f�vɦ]���,K����Ȗ%�b{��ڜ�bX�%����<�bX�'�ov��Kı/}��vi�Y�e4���8�D�,K��v��)��1T���QLr&ı/~��O"X�%����9ı,O���q<�bX�'�]���e�6�L�m͵9ı,K�~��<�bX�'�ov��K�B"w�xq<�bX�'߷?Z��bX�%���e�35�%��swx�D�,�EBD�y�lND�,K���É�Kı=��mND�,K�߻�O"X�%����,�eݖY�&�slND�,K���'�,K�����9ı,K�~��<�bX�'�ov��Kı<�~��A�(Pl���ڥ5�ӵ���ʶ�'Y��ymq��d#������wϏ|>Q�N�e����%�bX�~��jr%�bX������%�bX�}���	�L�b��ݽ�_��$)!f����)�Y�˗smND�,K��wx�C��"dK���br%�bX��w��Ȗ%�b{��ڜ����TȖ%����@[�r������{��7�������bX�'}�|8�D��Pb1S�k��9��<�9ı,K����O"X�%�g�̦u�[�M2��؜�bY� ��?}���Ȗ%�b}�s��Ȗ%�b^��w��Kı3�!Y
HRB��e��jF��i��Ӊ�Kı=��mND�,K�E�����=�bX�'{����Kı;�{���%�bX�ߏ����d�	hT�n�����쐦nkS;�.`�[Y�Zۂ�&���v�w��ŉb_����yı,O���Ȗ%�bw��É�Kı=��mND�,K�������fX\ٛ��O"X�%���ݱ9�Q�L�b~���'�,K�����S�,KĽ���ȟ�S"X�����n�e͓d��'"X�%���߼8�D�,K��v��Kı/~����%�bX�}���,K��>;{nn�-��Mɹ�q<�bY�"����g�S�,KĿ�����%�bX�}���,KT�$U�( EWd'�o��|B��������2�4�2nm�Ȗ%�b^��w��Kİ�P�{��byı,O~����%�bX��s��"X�%��w{���=��:]��*t9[������2��x�qf�wl��D���{��|��(���>�bX�'����'"X�%��{�'�,K�����9ı,K��wx�D�,Kϻr�l6vɦ]���,K���Ȗ%�b{��ڜ�bX�%�ﻼO"X�%���ݱ9ı,K��v�홥����33N'�,K�����9ı,K��wx�D��_�Pi�6'����'"X�%������Ȗ%�b}��;�2ݳl�f�nm�Ȗ%�b_�����%�bX�}���,K���Ȗ%��,ȟ~�~�9ı,K����q���e�����<�bX�'�ov��Kİ�PX����N'�,K�����S�,KĿ}�w��Kı<�$�30Y��sa��ST��i�κ�Gi�\A��ky�/I�"^n8u�lN۳��ĹZ}��wc9�蓣!����l]*�X���/)�n���;��ϓ|��];��1��q��z�M���LӰc�\*�)��^eB����ꘌl�r^�x䋎E`��{2Ks�,u򖭵۝�lsۇwO�`l�g7&�&���,�g��Mu���w�8b�:qgFc���jqc��d��.���E�!�4�'d���ՍSs-��4�eݱ>�bX�'{��'�,K�����9ı,K��wx�D�,Kﷻbr%�bX�g�oe�ܥ�ri�73N'�,K�����9�F9"X��{�x�D�,K���br%�bX�����y �,K������#v˦w��7���%��wx�D�,Kﷻbr%�bX�w���yı,O{��S�,K�q����d��E�H��w���oqﷻbr%�bX�w���yı,O{��S�,K�2&w���O"X�%�gYY�a�,�e�ݱ9ı,O;�vq<�bX�'���Ȗ%�b_�����%�bX�}���,T�����5�TU1L�`��lT�k��3�Kƒ!m�vz��
N���q�Q��U�L�m��M�����Kı=��mND�,K����'�,K������g�2%�b~��?N'�,K��nٟ��vͲɚM���"X�%�{���'��r�"X�}��ND�,K�}�'�,K�����9ı,K�׽n34�l�6]��'�,K����"r%�bX�����y��2&D����S�,KĿ�����%�bX�N�p�0�m��훻�,K?�FD���ޜO"X�%����֧"X�%�{���'�,K�2'{�<�Ȗ%�b{�?_���R۹�nM�Ӊ�Kı=��mND�,K�ﻼO"X�%����D�Kı;�{���%�b]���~�����뵲�)t�J��Y��έ��AZ{vqYm��V�(_���>|���sI3&�ڞD�,K��oȖ%�b}�s�9ı,N���p<B�B�ΐ�����:����UMS���7x$�H�����K���Ȗ%�b{��ڜ�bX�%��wx�D���2%�gY�-ٳe̓L���9ı,N����Ȗ%�b{��ڜ�`*=TB0Ef��Ib_��w��Kı>�{�'"X�%�{�{��fi�t�i�s4�yı,O{��S�,Kľ���Ȗ%�b}��lND�,���O�����_��$)!wKSS��5,%�۪��bX�%��wx�D�,K�=�?m��Kı;���O"X�%��u���oq���~����m1L�i`�֕��vzL�׶cFb�nq��/��=�妳4n��l�Y�.��Ȗ%�b}��lND�,K���O"X�%��w;jr%�bX��}��yı,O�w�i�M�d���v��Kı;�{����G"dK�۟�ND�,K��oȖ%�b}��lND�G*dK�����3r�ͳrnf�O"X�%����֧"X�%�{���'�,K����؜�bX�'}�|8�D�,K�߿�����Y�]0{�oq���|02&~�oȖ%�bw��lND�,K���O"X��=`��qW�D����S�,K����/Lٻ3w3.fٻ�7x�D�,Kﷻbr%�bX�����yı,O{��S�,KĽ���Ȗ%�b_���r�n1�n,�ʸ���1��Ԝ�2
��l��*=-ms�lN�%Q��7������Ȗ%�b{��ڜ�bX�%��wx��&D�,N�m�Ȗ%�b^��~.��7n�7.f�O"X�%��w;jr�șĿ�����%�bX�����,K���Ȗ%�b}����BivJM�6�ڜ�bX�%��wx�D�,Kﷻbr%��2&D����8�D�,K�۟�ND�,K��s��e�fYf컻�O"X�%���ݱ9ı,N���q<�bX�'���Ȗ%�b^���Ȗ%�b};��L�7aff�l��'"X�%����'�,K�����9ı,K����yı,O���Ȗ%�bxs HA�c��c���(D#a�XBX0�!X��	HQ�@��� IJH0$@�)��1HB,�`B$�RVV$aډh�%B�J�BP;�E4�1 Ab
�@�,��@P� *8�� Ab0�E��Xb0`P�$B)�,$,	 � �1b�b�0X|O���J_O��˃.4����!�w��#�# �� @@ @b_�-�$A"�`���`LP(�'�@�S�
�$`�`b��$���H�s߽�wwwE�[EU��gI�,[Lb��u�	m{Q۱͠&�esm�����!K7d^]�]���+ծ�2H�����vP���(sHtD/;*�wD��ʄ@��]0�6�63��jsݚ&��F�e��&Շ�3��:�vg˚�\�]����e����O���6��C@g�
Ƹ�";1n��&����v��>i���P$g*��	���O@h�5	�k�;a5;�]���w<�p��;Z�p��e�m�J�9V,��4�[��tn�Z����M��C�[��V�(\�[M�y;ff��ݎ��2�`4 �Zڨ
�6��5���3id��^Bq�ݗ<��5�ٕu=d��lEn���S�5 ���s���MZr�Q7iկmA���e�ĸtr�݋0�:L\:{&�k�!eiN�Y`LY�MZ�S`��3q� �:+������ڕ�\�$jN����퓒;v�.�Kz=�Y�l�ঁ!iҗm�[l��]:v�㵬Oe�rm�+nйIN{�9���|K|M�r�cll��G$�\�7k����Y SS���j���%Z셷K����G�*��'�v����M�6�-� 6� $$Hkd`H�z�[]/Z	�m� �] S�m�!��i�-�ۖذb�bY�5� [RI]�&�lf�v��׍[4ڠ%��h��aɥ��۝��4�v�Bu<��6�A�@���
�g�Su;F��#Y7�t��@ɵ^�7d2��	Vl��=@a�9 ���%���$��n�mS�s=�f�k��vw�����3.�q�C5�6*�nܷ�6:`J�;&�i���F��c����`�E=FgBaz����[.�̫Ƥ�T� URC��)WhZ��
�-;; ��myt���:MԁPm 6�Ͷ:��H���������U�c��FY��m�d�U\�v�;eH���ژe��e��f��舞
��(zuV��(��@;�q�w{����P���:d-�z��V�y����Y8�+��՚�8�9	�4S]�	�i�V6�qveGq�c���ce�k7�ڹ9��ɋsRN��ٿ�������B:r�s0�����0ݞ2s]rm���m�%s��ݺy�{Z8YZ,�^ƫx)��RE�[�v�G[���,�����0������l��K��T� ��0�Jr��d�V������|��\�)�[��:�����	V�H�u�`�!M�6F�oU+���t|�݉��X�;��ߩ�,K����S�,KĽ���'�,K����؜�bX�'{�|8�D��oq�߿����Adn�t�����%�b^���Ȗ%�b}��lND�,K���O"X�%��w;jr'�Eʙ��߹�vf�f\�.���%�bX�����,K���Ȗ%�b{��ڜ�bX�%��wx�D�,K�N�2]�ܹrM2��ڜ�bX�'��|8�D�,K��v��Kı/�}��yİ?�L���?Z��bX�%�������a������%�bX��s��"X�%��"������Kı;��֧"X�%��{��'�,K��;�6Ĺ3���=>Ϸ8����ȞJ����j�a����S���LuͯGT��"�����ı/�}��yı,O���Ȗ%�by�y���%�bX��s��"X�%�{�s��2�,�vnn�Ȗ%�b}��mNC����AW��6%���9�8�D�,K�֧۟"X�%�~���ȟ�TȖ'g����K��4Ͳ�ڜ�bX�'��s��yı,O{��S�,KĿ}�w��Kı>�s��"X�%����6��r�ͳv\���%�g�2'߹��ND�,K����O"X�%��۝�9ı,O;�vq<�bX�'�m�d��ݲ���{��7���������%�bX�}��S�,K���gȖ%�b{���ND�,K��{�]�&�G8N^v�Vqg��wZb!àl��&�Qճ�����R����yı,N����,K���gȖ%�bw;���P�DȖ%�{���'�,KĽ��?;��],�d��"r%�bX�w���y��L�b~���*r%�bX�����<�bX�'{�l�Ȗ%�b^���ni�p�i�3vq<�bX�'s�ܩȖ%�b_~����%�ʽU�L$M���l�Ȗ%�by�y���%�bX�l�Z�ha(l�L+!I
O�	2&}���'�,K����6D�Kı<����yı,N�s�S�,KĽ��݅�.�2������yı,N����,K��#�s��O"X�%���w*r%�bX����<��oq��~ܻo�X���T[�b��Bx2٬��mQ���	��Zu�缷Ϗ�����3w.l��Kı=����Ȗ%�bw�{*r%�bX����<�bX�'{�l�Ȗ%�b{��v�33]�3lݗ6q<�bX�'{w��!��G"dK����O"X�%����l�Ȗ%�by���Kı;�މY �7l��{�oq����}�'�,K��{͑9ı,O;�vq<�bX�'{w��"X�%��{���]5(��-|�~oq���;�ݻ���~�dND�,K������%�bX���ʜ�bX�&@[bg�}��yı,K��;���34�i���Ȗ%�by�{���%�bX������Kı/����yı,Mݶ��$)!IeƷ5.&�[$=�Ơ���M��nbc�ݬ�9�;i^����tS�/C�7a�f��	��33N'�,K��n�T�Kı/�}��yı,N����,K�����Kı=��$��n�0��$)!I
}���'��H�L�b~���"r%�bX���?N'�,K��n�T�O쩑)
{:��T��*E-����)!I
b~���"r%�bX�}�vq<�bX�'{w��"X�%�}���Ȗ6��ہt��*��K/��E���7�<�8`�T�Ҷ�j�v6Zf��0_I����`tp�5~�������[�vW���Z2U������;5v1r<�yJ�Ss�p���Cմ��x-����-r�m��woX��^^����6��ږy���,�n�']!��U���;@4&���鵖2����I�����0z+D<����U�P:��۝;��m�][d5a���厽4����%�4[i�^��f߸:_�vx�6ۛ���$�b�Ew�{���Ӿ��,�7e�/a�k,�Ͳb�ݴ�V�d��e��>����E�]��vˊ�6��OɁ�����	�\�B��iZN���xlp�>��n� ���d�i�IՃ�m6`�:`l���`v�Ӣ+2��5V��V��g8`Ώ ��s��`n�]N�������XΉ���:`l��м�㹸{�]��g̹��$�ܙ��v��e�.�E�q@�n����lx�U|�~�P`v�遳�Ή���-�2�MS��,��j(�P��;������0�*X�4�
��L���6tLؠ��+ �W)\t*i�i�%vف����;��`t�X�p�&�r��ڵjݍ�7�v��l�����G� 7�<�e;�Vt�`S��`���Nz��*�ѳLo���Lm����d��\i3�ݲ�e�H`{�t������W�&s��L�����T�:UI�STՁ�φ;�`n��0;�U�0$���X�k�3����q�	_XP
()AMC���~�>�3��`f��(�MPLKe6݇�������6s� N�������a��X�	�:`l�;��;c�����Ucv�b�e�U�L�����oAH�M:Ֆ�j��,�C/RN�I���u�l� ����� �&V��R�M�]�@�m�;�`v��06r��+��N�i	'bj�xlp�>�e`K�� $�)���'V��ف��(�ww��έ�fk�"���(I#F1�D�B@�##��B0 FB�R@�@!�V�a!`B,*B1p������0�d(5��,��m:M��*��*����l{�`v��GL�UU{����>�����"6I+��ҷcu=]��ذu�Լ���mm���sO.��1�T+J��~Lؠ��H遷�c ��e�]^*���!bI���06�L`�z+�V����U�ň`{dt�۝1�n�Lؠ��R�V�MRN��n���`�D��l���r��Z�Z.�Pf��7z&lP`{dt�����«�QC�`*TE���}������0u�JR���Ռ��������:Y�(��L�\]8p�s`oUv8N޶s����]"�w/V��Il�`i8K�Ν9��'{O<�<uќ�s�1�U&�	�w����V���\[�kWf�,2f���T	Mڎ-��%�Ч�(�{ge

3r �շ,MT�n�k^gj@��DڸȺ�
�>+vccr�c�6l(�Q�o��i0�J��O+u[���,Rϰ���k��л�2�]$&um�C��6��ui�7 ���}�mX�z~�@��v��s$nT�H*�X����遳��D���J�J�1$� ����0;b��#�w*��V 2��hn�a�&s7���ϋ�͵aВJs���v��J�jBb[6���0=�:`l���0.�u�|�.K���ј%��*ۦ��'b�lu��Y�A��$$닱A�ncM�6߿c�ݯ� ���߹�lR���O&\ɦ컧$����� S� (�������>��$P`{dt��ːX�����t;���0�2����c�iݴ7hI:�ě�;b��#���lw�`K",�t$X*�X����遳:[ �����n����e�ʶ&Y�v�h�M[�*�gLKӬEӜ�u����R�)'umRT�'X���w��;b��#�w*�Z�WF*�lw��;c��ɕ�l]/?��o��`�M5!1-��v�>,��j�d&A�$V$���a!"D���H$��#1 ��,bB,b���:H!�\�Nt��c"�@�H�1HG�'�!�a�Db��x�����}RYVF%�T 0�@ �+P�)V"Bc=��V	H�LHb��B�/��1,B,FEA����g��a�V��_��9,(@`�����@^D�<j�`F$U��'�Z �@���)
2�hJ�JJ�2�Z�IVIVH�@�XHP�%HF!ec�j$�D�<(FF,B� < ��A�_@@�@�T��ר�t�УQ���Ws�} {{����x%�[�TST�t��>��[�`���;c�ܥ(��h���M��`�͛�DNgs��|X��'skvͳ`z��ver��)�{띳��9{vqYW�2F��B꛵��@�u��쉁��:`lΖ��)5m;bN�16���nɕ�{k6l��w�D(��˙%9Cd��m6`��V�t� ݑ��� >:K�umRT�'X���	���I����H��"�"H<TG%{u�+w�sT��5(��-̀{ۮ���B�����fwZ�=��?6߿s��]1TM�tj�f�j�4�����R6^�:�ך^2���s%l�Y�pf�c֐�`v�쎘3���3\�R�-̪)�r:e��nھ�2gV��gs�3����&�r��R��wI�-��;�z�vG�v�vL�yr�:ljڻN���x�����,{vՇ�P�Nsޛ��Ԛ�lbN�16���nɕ�{����I���I� ��,RAU���ÿ�/�5ѫ�y4nn��S��k�OB�\E�����.���g����x��;[M{R�M�����4�u��Ω��k'T
l�v�^˱�v�M�Ufg��q<l�S�2,���&�Ov�!:��I���ہ�Ǝ+b���|��K*�g��;\g��Ī_�0��ncDj��۬�/@+\�����wQ�9d)M���[7�����{�u��������#���*Nθ�蝮�K��'�;s��7��5�Y�UJls%9Cd�U.�8�󿵫�t� ݑ��� >'J�umRI�USV��f�(J&C3�����=�:`wr����V+.�T+J��G`g��g�P���wZ�3�zl��X]����,Ę�A���ff͇�L�o;w��KD�2������06gK`�&lP`z���ݵ��5�w箒�965m9ŧa'Qq���6�vNm��oE��K�P]0�06gK`�&lP`n�遽����K��h������
& � >�*~�UH M�������V�t�ld��m�BIզbI���:`lΖ�7dL�H��;���Ҷ�0�2����� ��里݉���J�2����ޛ�$�3���>,{v������������a�8�Ka�p��:�NZˣ�9����n�t:+���ݎh�V�.�T+J����`v�쎘3��HEWuw��_֐�`v�쎘3�����0���ZI̲��#�X�֬mf͉�Ȉ��Q�.JaA����3y�`ztݢf��Z�M;I��t� ݑ��� ݓ+ �]6;jڻN���x�#�=;���;��b�x�H�;Cuusp�c�\h2�nV홄���mnZ���̱����V�W͎ؠ�ݑ�ft��"`*Ev���Yv��:`tΖ�7dxNp��Jj��V�%N��u�tΖ�7dL���ݑ�{��*�
ˣ
Ҷ�"`t�얬*J!G\yDFBIBK��w6�ƴI3M��#ct݁��K�3���ս6��vb�T�TS�-5Y�ʷ�z�yQ[�a*�:"9�L�ٺB�!k��[t�؝'n�>�=��t]-�M��A�/�����E��U�f*`lΖ�=:&lP`v�t��]�۶�݉�44� >��0���s����ld��i��ui���;c���+ غ^���ϻ����r�S�6H5R���ͺ`lΖ�=$Lؠ��V�}\�.�^���jw\�J7j��d&�XΫ/Mպ'6#�t2��J�v�.�k��'�7o�u��Y�u��E������q6�ͺ�=���םn5�*��J�]���Wv� �{W�2s�&��Ʀ�����)�9]�i���~|I���s������v���U��۰&�Y�g��(�T�HK�խ�r����'���Ǌ���"g��羻�rh]�2��q@�\[�d������"..�\^��ڹ�c�qm�VZ���:e��@��^ }:<=�O�(J>��޵`n��&�T�T�I�V�=:&lP`v�t�ٝ-�zT��.�"���.�Lؠ��fڳ�(Q
g:���=�����+T���������遳:[ ���� ��$��ݺum�:�6.��=:&lP`v�t�6L�f����,��g��]RQ��[a�r�/��u�e��<uh���N���ߟs]��ץ��͵о�έ�;9��ff�2ff�777y$���g=W�
��(K�!
R��kzՁ�[�`n�`*Euu��H�U��!����b�x����� ;�(Л�5IR�fb���lӢ`v�oGL�q��+lV]6Ӽ �txlp�;ze`K�?����T|�N��[�{r�s\i9�j�r�Q�/9��_n^��b\�(2�M��$�:1-�-����Ł���ft���0;�������E��b�0;z:`lΖ�=:&lP�:��J����j�ZbN������v\y$��DD%	B��~,�u�yH6;M%l�hi� }�<=�K�fڰ�9�zl�g2Z�i�I:�ն���}�2������v{{��ə�R��L8�u�]0.:{3��cjX�*v�̘�drl�;$��l�:$X*�X��7��L�����`v� J��7WIӻI��t�䣈�P��3{�`ns���ٶ��q�Ю�6M��� >ޏ �zDDϳzՁ�[�`b�[D�ӑ�.���(������oZ�=��6�D~Yn��vٮW'Jdi�˫V,C���ft����A�O���@�n�S9��������D��&-�t�n/:��0E�^�6�,�L�����`v�����m��'bt;�ޏ �l��3��;b"-U�"��Vb-$��l��3��oD�:t�t��,+i���z{��:�<������ҔIZe��T��T�۝1��vE�'d�s�$�AQ_��AQ_�DPTW�dPTV�����
���(*+���AQ_�EC��PTV ("��
����
���(*+�T�����(*+�蠨�������
���(*+�(����"������������)��'\���4( ���0���    �  *��@        �zT�RB�((�   
  @P�UH (          %AI%@  
�   ��    (a k)JSE����4	��J �}2waq��rt�nM }>��.��]������`   j�,��`" ���u�rk�{�=  �    �� PU�
��
`�'�b:vu*ɡ`�n �&��#�[�i`��C'��<� f{�8ZG݇'�3��{���A��X�C"���u귀| $P  @	� ��U�݃�]N����.�@Pw��\�U��,f�ۉҬ h2wbq��z�yh�o�Ϊ� �Ү.��=�Sv:}9C �}*ũz��ˋJ���Wχπ���� 3���L�YW�b�12�����>�냓Tbwo��Ҙ JVN]��8 �rҖ3J����$���aVM.�x��V� 8��C��ze�/= >�@
�( *��A� ��K���^��4������@)�����QM60h�ΚP i@�� ��@  �M�ҔM Q��iH��JQ�� 
lf�i� �R���� Ħ�4��@�viҔ PT�ʔ��!����OBDԥ
d��`S��IQ��L���D�*��Q*�L@ hEO�	L�*J�2�""CRRTi�2h؟%������������j�������g���_�b
���PU�?�E�(*�����+PT�����͎�4(f��.,.�(Ć2cG����!���)!�&�Q�L1��B�b�D��HN]�5 �e�e���!�+aL�1�1 ˄�2!32o!2���#�
� �)��� �Io����Ux�q�t]�J����M�h��\lN��3'��;�p���w90c��*���}'q%�o������Sj�.��j+D������&���w���H�..i�N�`�-����ˈC��b�w��~�}Q���1wy�{~�5ʇ����9À�)�jTMA1�}Knb^�\|��ώ]|�&ң�j��m8�R\�\���Gb�;��(�-�޳\ˢ���]��S͜h}�r郘A�E˼Bip���n�2N!>�n��L7�Kg�&��8�_fn�bD��d/
���I	4
9!�@�5X$@� ����=X ĉC�h`���"(0/��тDO{��+�B� �1�]
�<	r�HCX]H������X��CXX$8s�1�D(lB�6��Cd����%5�0X�b1$5:'́!/�=����Hً��0�!cI	��8��<YK\�P��� �@��L����|��hP��c��74"� 28�����0K���G�5!���h0`@�.,*�P���C@�SB P"Q��F�04��H0�LD�p5cC�W�}�.�]�|�sp���I.0�ׄ9¼B!cQ�e��F,B$Hē��RR�@�F��/	9��E�AI.m�X�A�@`���
$��T��PR0
���A��h�<i��@���D���B��q<�>󌾜<ND�R�,J4�2	���'"@>��(�MV�T��E�u%�K�̄��M���-"q��	�J�b�>�
`&�6yvaH|󺇜�!�� b���A�"�`$Z�H����0b8�E�j$R����.o<f��|��|�bB}�M>4��J�0垲�{���͋#HxJLH��{��=a�<OhH3Bk4��SSq%��!a����!B`D�4��3FˮdI�	���r��E�m=��}<4�4�e����$X�)-�xhF">�)��*���o� �Kk�00��(���1`%UxE
�E�YO�.jp�jD�@<T�����L4x�)���h`B�����<�K"Ӌ�i�}d1H�J`K�
&)���&$*D K�˚@�Q��E#dJ0*��B�F5"R�HV��_�p�+�*F�5$���jf��M��`���a��&�p�S{ϰd�4D��[�4s[����ni�.k��J̑��h[=PĢN`F5RV1K�7�w���CX�A�H���ǿ>�k��<�
�t��qoM�u4&_���}�ӱMx��|XGd$0��T���so<�#C5%H�$0V4]�	t��	�Jp��1�|�>G����;���F,RG֨j� C�t�j�}"�ք��=�a�� �R�xa)�s��D���!1B�"aa%HÚ��k,����XZ�\��d��"L�i�fr8.�]�Ȅ�\��X��$�8մ�y�<H����ġ�>*����!	1RW�1e�~m�arF!�/��[�l��Oa��T)�ɩ����ĵu(X��Z�k�jF(��E羸V5`D%Ic%��Q�"�AX��Ȱ*X�`�"D`�"T ���1cU�GxƦ
hp��G0H%BF�ı:"*H��8���a% S�P""�#p	L�R8�1�2�"T"p!]�4��0�%p�	V`4X�(@1"� 	V%L"U� W �T�@"�H�X� �`Ł@�T�S%BE`Q Pc\VH�B#�R-`@ W%@�@#VV	F�A �pM�l�5caB	�� �=��3b2Ɛ`w2c�8=gr���\$5 ���!��@�"E)�J��P�#"B�$� B�,!���I�A*1`�b��0�$
� "$R��$�a�$j`�H��jD��Ha�F��i �1B�Px�b�|4�iBQ#�BpaR�y�ȡ�L�!(@h� Dh
�`+��b@��H�)�+X��Y�ԋ$H�� �b�b�R��wÆ��>�{���Xz�*`� ���*h�
��Yh�F�VH"Ё�T�L4�a��Z!���H��8�B/0�#�k�8l	
�,���4��
渚8�W7yiIC�0���Ck�7G���yjH2�aF�f�ݤ��L؜� NJ��#d#dq�X2�`fP�L�x�3�CAe�k����l���L���N�ɨk���r/	!v<�CNl�+ƻ6��CI\���$hб�l�0�0!!�jpI	\48Ƙc���I��%��5�2<(aC$�8K�<�X�I�!m a��-�朁��� �ȱV���I�%�gH�ݮ�!�Zf�ɻu�Ұ��F���My� Bᆼ�԰���%7dg,���8`H22&�2�VNg!HX�7�n�L	p���E"��HXC��iSm%��,shX0��Z.N,���t��H���)�3ymX##X��sm.�:m���f����+-K1Д�1��# I
!����ws\�%����*iD!C��B����)8�$���0h!�Zs�ʄ��	 E��1hHrP0�ل6p�Ʉ�
�b�X��BBS %2I#1#��Sb�b�`0O9{��`<>����y�.$.$��篶i�C�3=���m�M�y!!.r���$��:�T5�d���l��.ph�d�΀��xB��
����F[U+��8�\�nm���>Csko��pӄ�C�$E!RI�P�B�	%��0�`Ub�8�f����G�@�bF�B䉰�Ф�-p P!M�%0և##Lhi͌��`W#	LuH�u�W �Hm�
�e���5Ȱ�H�I�F<Hņ5.�:��_V�;w�9�<��h������&���f���R�R� �<p65!xhW�%y�.1���$1%�\4�IpM%���
i���ǋ��bB#
�����:���!��<i�P�p�B�
`��B(��m���(A��PH��D��D�`B�E�#�����t������  �         6� �l             �     �ѭ��m�Z� .�j����ZV�(읰-��      6�!�kn�`���mv�Bݭ��R�.���e]$�� ���   AmI6��  ںl��V֩�inԎP'���:�Tڶ�� �W"sv��z����UVҬ�R��>|� ��@�9�t ��T��ѷU���� �����i��*�Rn.��v�8`
�mp�f�:��H  �tR�L\�k��H79���gZ�e�I�ͳn�y(	\��:LU:8�J�dj�T�ʬ��UQ� h6۳l[D���r�jv�m��Éo������X*�Ή�B������N[��A6-�C�m��!��UIz��9�adȥrmJ+��qfWe�Uye�iO96#�bvm���9�P!J��Y�7&�`̙�x8��U�:ڴ��e��zܩ.�� 6�d��Md(mf�*
����`,�J��&��  v�K�ôml�m�b��mmAN��r�� [<����t����8	�+�� kH`I��$�d�]��6�r@�g>U�Y*��궠�) 5R�t�Ԯ�KK2l�s���ԗR�W,8MUS�&��A�h^C��k��[�km���ۗ0�n�K+j�jU���ć����ZVcԲ�q�p�E�-A�M5�@ p����qvu|}��.���g6����x�$1Z-����Zޜ��y�:-����b���mɣS�O78uU�+`�������N����'�u�"Z��k t�������˞��Q��I/J�����Qew:��5U�cB��������S��w��q�@.�P���%�oJ7Cr񶬴���t��z����n����kn�t�q�=�*pc�]��wb5XJ��XҶu�:�������$ ��V�w����m�@  �8-��m��m[   ^��m��7[�ݩ�n� �uljlL��%���m�mH[A�'��E��l      ��� ]�p6� m� sEr@H�����   m�l�l���l  �  6� m�� ���Hp       � 	�� m�,��m ��8R�N�[K�l 6� ����Ͷm����       h 8�b��g�ym  p   �C��� ��n�m��M��p$   	m�[@[@       8@    @ ���`l-�  p  �mh;Z��m[@$	�H�[\��b@�l $�� �cE��m��P.�	 t�ۍ` iIg�eZH*�Z��٫m�״��i��  'I�� 8���5���޶�m��lH�-� $�7j�@��i�	86�-� �m-��pm%�n`-   k*� ��GMoF     �n�$�iW[N � -��JvV-�L�����,���e�� �oP-�ͳI��!k����I�V���h �^� H tZ �R�H6�a�ml�[l L�Ru�m�m:cm�X���[@dP �m{M�i%� $:��l   
]���  �m��  n�H�-0   ���0�E�[nY�u��nP������.�S���[�ƕ�t9y����	mu� ��M��p� 4Ӱx<[V�m lmb�86�[H0 �`I�[@H��m�m��4����-��  �y�]]�m�mQvD�`��۰,���ۉ_�w��l�fI����N�%���%�	n/h۱ �J�M���`o[Mj�l�j�Б�� 8��}��\�� ��zvI�[7��*����w�8�۲�[��JS�Hݍ��+S���4���v.���*�cR�m��@��a�,'C]�-4� �]Jݤm�-�l�nh�U��m�	f� ӖY�5�&�6I��c��,�ћ^�����!Cg3@m��a}mU�UV�4�g@�_Z��� 	6�%^U�؇WWUJ����@��  �[�\q�e�8Ӗj�����s��[pd��2I��6mP!�T=�e�V�����yC��2���5P :�2@ H�l�m��#EI�%���@9 Im[%�@��	����U2PԖX����-� ���s�A����&�9ש�n�   -���&ٶIf�����ʹ����!�k����"�Ҥ$�km���  ��l��E�I�z���km�m�� l .��L� s��(��ʲ�T�'q�6��l�6�H A�Ŷ���68n� 	��[���6�M,��k6�F�I( 6ہ��qmq� l�[ X��$ Hrt`�bC���-�8m�Hz���2  ֱ�[d���     �M��� ��V� ,�6�  pd�8�npp�6l�  l	m�v����l��N m�����O{�� -� $ o ��ۤ� �%6�n��-�hhI� �Rm&�A�m� Xe���    hku�  m u� �   j۶�Ëhm�2��  Y)� [@ 	��%� [V���m�A��	�7m�� � ��     8� $l� 	l �    -��8[@-���� p�6ض��������� $m�  h��x6�m� l ��� ��۶� m��`$� �  �i8�	 ���� �l�l �t� � 6�   ��  �ll8 ��_` H�   m�n��� p � H� @ 86�m�� �ն���h �mi7d���5� :@ � �[p a��  p8 n��� ���$ ��m۲�mm      [Kh$�m� �` �`�[@�  h �kmm��l p  6��̓��   � �mk ��i�l���n� ��    m�[N  ����[p8 m������mp H�  %.pkX�l�`l m�  6ٶ� �   mi�   l�9%�km�6�`ݶ6�v��	�  �  [@�B� �ۖ��oW��l m   �m�!"A!m6��pp/]-�� �$�p�m i+`I�z�m��� @6ۉ�I[v��V� m��]6p�lh6� -��&�qm��C�V���� �i���]*�Ǯ�v3J��L��V�2�G�.��^�&�ONlp66�ƛ��e�!��R�����j�X��� 7I��ZΣ��`�o-�5�m�@��Y�zn�x  -]��L��В޻r��kv�m����l���r�UV����U�P�z�m�� m���l%�Amq���H�k6�5��U[J����T9��V���d�4z�*^YUJ:@�X�mu��h6� )@��6�퐚�vYbne`*�����=�ŷ�(C���IR��!j5If�^� 6U�s�*� Um�UR�P������ ��M���l�Y`��	 "M�ێ ւ�   m�l�A�a��m�m&ٰl�]m��  hp� J�٭fՖ�Zi00` m���`  $��l$h $[D�m�nݵ�m ��j�m�e$;lӶ� H  	  m��  ��� $     ݫa  X�ؒM��`l�L�v4�86�޻`  q���l[@�l  ���m�8��z+E%���I 	�m��  �V�� ǃ�km�l5녴    lI�|��u�m�%�-�mI,��� �� 7j:�}�k�ݤ*�(��\d��(VUP �۶� ���@�_/�N��` �:^���UV�����=UV�K�[U][P@����Y��}upضT�UT��h5ey�$�ڱUU@  m'հ$,4��0Zk��6Ͱu�@�\s����a���Y{l�#e�K�!�|�򪪥P젫e�eV�}t9݊�j���*�����)��E?У�T��A@04R�� ��AE7��J&�
t �5yR��"��	���� �P��8(`���T��GQ�xx�A��x�����^��CO<=���,7��S�<�D=�=DN��!C�AT8���A� *) (�J#�T�8
@z��� V�!�� J8�S��@�Q ��^h�Ra!�B0��	����!� ��#��^(* z!�PP��z���xD��(}訸�<�S�Cک��N��z�u�&@��Tt�Dp�>��LE���O��"A(���w|;�Dw�C�S���6HI�K0��	h�E�$��2�ŌC�}S�#�!�� !��Q�AH(� ��p:�AD�@4���E}?�+ $D"��� �A�����Ͼ���������7vKh �� �&�[�`�UX����lr�T�ʪ֌{U�U*��l�������������"�0'^�:Mƴ/^t��Y�\dl��n�����i�u:3UQ�=���j5<����R���pGJ�mU@.2R+pD ��sm����.J����.��b��9ml�lg��k��y�0uGk2u�ݟ�W��or��zggu��)�#�ef�p�f�KUR��Z4�ݰlN�Iڧc#UUU�	�2�@��
�0U+�ВRNz9Zhƪ���j�ۅ���v�OIʬ�lJ�P��]qm�����I����tn�m�"���h-��� M�L,�$�n�Y�sv$�YӀd�M#� �X��Uڋ�J�:�	��5���뢶ܫ=��Kv�R;.�r�*�� �a7'k	�[{�p�N�nf���k�I9�t񽇸�n��|0K�m�ZG^�E�]s��V�7g��vyK�%���'gB3�q���n�=��\&��-�z�I�VM͛vm��ʌn9t����@Csl��e˕Z@���탭�au��s�]�IKj�gjں�6t��)n�9�Z�S �<�#n�m��3��r�R+mV�tm�KTU���j۔�1u@G�����u��� 	��T`�AUA�@�l�y%�%@ծQ���f�� N��shv���;@<�S��)E�8�­�LԪ��T�6����tYD��\�A�VյV����@�W9�����xn��s�iظ���6����N�l���;8���6,dܩ�&�nenk��mW��}�%x��ظ�=#m�Ā�d��쏮wDfx۴�X�E��i�z�`:�^Vqث��ʸ�V�ub���gl�<��[x��O���%�u�����i����۳j�=�v�Uo]R���N]�y= tv-�inݹ"�&N���j�@���&��+��.��Y�������/㘠��� ��DX ��*��4D���q<}�@~�=�2�f�ͻK�J�y#\���ٹ�6�6-�:7i�j�d�u�{qInr�u�Ͱ�ΐ���۶�����g�����e��\��(u:���tF�s�J�v��ݸ�^���6�8��E�䚣a�ۑ�gv`MM	�\4�87 <$t��a�#C�un&\�j�\c[��c�8ѷ5�k\F��٩��l0�&l�ݳeT�A<�wK�p�(Р��
H!H�<��a\;aA6{q��g�d�D6�Ĥ�e%i*,G>���	 �'��lA<�{�p?�
�?DȖ%��~��ND�,K������I\�[����131z?zL\��E#�2%��}����%�bX������Kı/�����%�bX=�/GG+c�V�F�����������'�,K���y�Ȗ%�b_=�w��Kı;���ND�,K���ev���]��n.������{�ND�,K��{�O"X�%�ܽ�br%�`vdO����O"X�%���N�B�d��Zbf&bf'�����%�bX����'"X�%��{�s��Kı;;�br%�bX�������K��͜<�'���g���x��I����a����)3������s���{ı,O�~�ND�,K����Ȗ%�bvw���Kı/����p��L�ŝ���X�@��Yd�Ȗ%�b{����y� RAF1D>�P󂀞*?bW؞ı/o�n'"X�%�|�{�O"Y�������b�131w��"��v�.&f�Ȗ%�b^��q9ı,K����<�bX�'r���Ȗ%�b{�}��yı,O�I�����t�n̻����bX�%���x�D�,K�{���Kı=Ͼ�q<�bX�%��w�,Kľ�񙙝%̅��dv۸�bf&bf/G�I�LLKè���y�O"X�%�{{���Kı/�w���%�bX���e�,��K�qº׊0 �:G�t��l���t^�m��DM,��Ia��9�����ı,OsﻜO"X�%�{{���Kı/�w���%�bX����'L��L��_O1��[VUGie��Ȗ%�b^��q9ı,K����<�bX�'r���Ȗ%�b{�}��y*dK��ݷd��3L����Kı/�w���%�bX����'"X�X���@�HAH"�w��r&��o|�'�,Kľ��q9ı,O{����IeMV�In�ቘ�������ND�,K����Ȗ%�b^��q9ı,K����<�bX�~�⇤p�Yd,�b�131w>����%�bX����ND�,K��{�O"X�%�ܽ�br%�bX���߾?��u��.�ٌ�Żz�cu��v�]��.�#�gu�Q�\��w��B�˃wp�d���'�,KĿ��ۉȖ%�b_>�w��Kı;���ND�,K����Ȗ%�b}:M����ۻٛ���Ȗ%�b_>�w��?
G"dK�_߳�,K��;����%�bX����ND�,K���ffuIe��#����131z?zL[ı,OsﻜO"X��2&D����r%�bX�ϻ��yı,O���a��9���������o��w8�D�,K����Ȗ%�b_>�w��K��(�C�E��DS�
~��';|�19ı,O}���-�wm75�͹��O"X�%�{{���Kı/�w���%�bX����'"X�%��}�s��K�q��������r�0Y:���A�����]��@o��	���d~}�ww���실�ݙ�f��yı,K����<�bX�'s�ܩȖ%�b{�}��~I�L�bX����q9ı,O߿���KeQV��qp��L��^���9ı,Os�w8�D�,K����Ȗ%�b_��w��Kİ}�d�C�5++,��LZbf&bf.�}��Kı/o{���bX�%���x�D�,K���T�Kı=����OH�m�B�n.���Y�%���q9ı,K����<�bX�'s�ܩȖ%�b{�}��yı,O�I��������n�n�r%�bX�ϻ��yı,?����T�%�bX�g{�8�@�N�{��|!�0"����3�ܞ٘n��mf\6.�������==�����t���Ǎ�5ò����q�tr�.8-�v���9!����״�Ąiy�l眔òV���W�]Ir��=;�\q�.��T�0k���dd���p�g;H�Ni7fzB8�p E�ص�&Y��VyNv'�<n�-�D^��&���0S[v��BL<�.0��9���s�Qu�m����������.�Ht�bd�̝<��N��vk��V�!9���n]��*�aQHGRI�:��=���@/m�ffg�� m���b�q`�IƛMǠqw���@>�@�����P��ds�&���f�}�f�Wmz{^���nG�L���I4��h
�+�=K��TDL��.K4m0I��$��,cNM���+���٠�@��^��{1Ƞ6��5���$A���d�<�s�@������.�6�jF��'�$��#b��W���^�4��4
�k�9�x�m"H�2d����N���=D� 	*�#�L�K��H2�f��^���W����;ۄm�9$��#rhݶhvנqw��-�@>�q���6Ґ�6��Cي��=��= �hݶh�$PP��'m7���W�8�������m�?&�@��C}�}��U�&a浩�+s6,�wV��Ǚ�chT��s�#�]�Ul(:oS&��[f�}�f���^���נuUۍ�S$j`��m���߳1"��=��= �h�`�ǪI"�*,.�4�J�Wr�Dt�gL���(�CTD�g���$�o$���I1�Ȇؤz{^�r�4��4���r��7[HR<H`�z�l��l�:�k�8������"c�E&ciC$�����s��x�j78��8�`6e఻]?��wv^ү����c�����4
�k�8����٠s��n�� �n9&�Wmz)r� \�hy,ߢ&b*�ofV��I�6��@�����f�w�����gZ���ds�&���g踉��i��ɼ�rW�F�dEDD��ĳ/f������R)J�%�.�3@?rY�9�v���u$�@%��p�n�d��Rc�A(�(Ɇx8�(0;n�j\��8sH���1U�"`ܚ]��]�z{l��l�;��x�i1�Ȇؤz{^�&""�"�9���7�W%z�����IH�bhn= �hݶh]��]�z{p��1Ȝ�s�M ���������@9m��;�6�	�'0Q�$�Wmz{^�^՚��� �n&bf9�[L�+"�7C�gy�W��}]^;$9,��Ed�8�4{x并'��^��q��;6P˞K�eV\Ys���{^��6�>�XZ	4=U����Z�9:��Ȟ΀ݺ�sk���Oe���:Xn˄�bsI#�N�Kks��۝l<4�ղ.`�DW���I6d��jV���N1�,�y�rgb��Xl��& {n'�&�����C�q� B�fyn��˛�l�6�%Gi�}:x)2�������nQ��;Ki�d�
D��H�i�����z{l��l�*�@�Q�BD�9�Gq��@>�@������@�/j�70q�LjI�v٠U�^�߱.u�- ��w��$���$�0nM����>ՠ�� ���@�~�)=$�:�	 �_~��?f,��{��wޚWmz���;�
7:TpG5��;]g����ݸ�1�y�PmF�tFz�����r�ye ����o�߿o��l�:�k�f|����@��Fߦ73v��]��I'����*#{�-���ɠq����w���8��7$�bR��$�:�k�8����٠r٠s�\�AɁ�4�z;^�r�4�[4���e,.5	d�Ĥz�l�=���b�}��_y�\�z�33��!k=����뗅��Vv�g�f��8��.��/|����nl�q�ě�R8�5$�����Wmz;^�^�4�Lx�̒ck]�h
�+�1Turw�7���f��vc��m�Sؤz;^�_��K�I�	u�d��Gۑd1s�t��i�"�����<P�D� �p�*y��)HI�u{�B��x��T� O�Q�O.|�< B#�*:
��<��T}-�T�31ELGQ�f���޺����.�i%"ŉ�8�>��w���wޞ���@��z~������;�9[���ye�T�É���������\LDDEQJ�w����_��9$�����@W�'���0��u�]Z��Nd��8]�{d�� ��������+�+bR�;�DDL�W�����"fg����	���� ��~��y'������v���M̫�.�/@���\D�LUm柢&"*�sy�*mۈ���Ux8��2����/*�/C�DU&�h����R���]�z]�n$�q8�x9&�}��y$����$��~�rJ����T�?fb��女�{<	<z�I1���&���^���N� so4�u���Y�q.�.���(n��Xg�ɽ��ڇEqQ�;y�]6�v��i��֥"ȹ����?��r�4�[4���^��n��R,H`�z�l��l�:�k�8�����I�f69����<��z|W�z;^�r�4���Jࣉ�1FԒh]��\�z�l��l�9�.H����' �n=���@9m��-�Wmz?.��E6�M���gV6^v���yu���&�X��{l`M��հ[�]�����ܖ�D] c��u@\k+%[C$i^��q@��t�)�WZ�P]��I�ƶW�U�[ 9�wnBT6,�C���7+��;ccFu�\µ���Ƹ�r�Լ�pl�-���ŵE�^Ze�vq�E2��nE?�'ώ٠!�(��M�l-{)7w���R��4MU�廡�V{[.ӳ���Oa9�S����n�zơ"X�P�%#�����}�f���^���נuU���M��'��hܶh]��\�z�l�/m0I��1ɍ,`ܚWmz;^�r�4�[4��	㰑�B&�#�8����٠r٠U�^���7���JE��@/m��-�]��\�z�u\d����݄R�ݨ����&�칁ud�Ƅ��oHgk,V+l[	�#mH�(8ܟ s���*�@��k��ٟ =}�r��m��M��6�34\����D�P��^�~�@u�-�$Pr`G�m7�W-z�h�f*���Rn�B-B��$K���Z�l��٠uvנr�ՠu^���m��O$��,�:�+�<��h�Y�9���`��ԻM��c%���S凇����΍��m�X�tf�)��=Lj�/e�Ͳ���Wʴ�,��Y�8涂�?BF��G��Z�l��٠uvנw���74H�!�8��{��y$�{��'�>AS���yǠr�V�޻�1��jI�A����٠Umz+�Zm�@�_pM��n&�ڒM�k�=��~��'_�o4��h�[p��˫���Wc/�� ��.��ʛ�etiGi���4�4P��E�� 4P3���?~�_�m��4�[4
��@�Qܸ�$K�Ĥzm�@>�@���.v����7n(��&�}�f�U��\�zm�@�Ǐ\d��o��*�����@-�hs?~�s~��%�9�x�$n �$z;^�v�4�[4�k�:��,x�N���;��f3hs����A���+V�x]�r�gtn�p�^Y@����o�l��l�:��@��k�9�q&7[C�~o�M ������.v� �o���&�q6��4��@궽���@;m��-�k�X�Q�`�R$��8����٠r١�ي�{�@�x~�cP�7�8G��m�@>�@궽���@�?f/ߠ�{j��+\A�-��M�[Mzύ˺x�u��Y���;q��'=�ή��\�vu쒠V��6`�n��[4���'-��ֆF��uڲ�ʹ4s1u�j�ɶ�Sn�;Z݇���\��\P�⍌s�w-�/[���@Y,�!����=*j8�>5�z^�)��7A�z8n��g�q�։���ީ�3��<P<��T�Ҧ�E�I*��$f,Y�6M���f�ԝa�ٍ{�q@"�Yk�g�h�#O��X�M��(brN�__�u$�@�{���@&�h���2�1	��@궽���@;m��-���Ą��$n �$zWo��v�4�[4�k�;�to�I1!�q�m�@>�@궽b����;_�&7��M�5���ʶ����� �h�+�CvpV��Kl�ҸM;p�2�1R�t�H��X"\�9��v���c��W�¦���r� �?�����*�Yr���[�h}��y���Y��D̩���LÏx�f�.O4����;���c�B8��@;m��-�{����:�|�+�X�M��(eeU�f�~�Y�u$�@�{��LL�6����4���c�8��	��@궽���@;m��-����s$��MlV�b �Z�[��.v�@Y�E>68�a&HOf��	ᬑ�d�d��Wo��v�4�[4�k�;m�<n0��ȸ���/@9%�����a��@u����8���u�I���m�E����@��ޚD��X�����_Ñ�������}��n���fL�)$�t��zW'z�,�u^��@N�8�Q�`�R$��8���+�z|��߷�O��?~��|����������w�+�L5��Z�We�a���ϧg9��)�c�]�Ҽ��|l�����ݷw8 ��߿o �`�`�`�}������lll{��~�>A���������A�A�A�ı����r�$,)n[ubY�bX��������Ƞ� � � �?~��|������g �`�`�`�{������lll~����L�nnf�&f3w��A�A�A�A�~��8 �����>A����A� ������� � � � ߻���|�����~��?d���n�ɻ��� � آ� ��w�pA�6667��~�>A��������� � �(~�@� �(�D� `b&�������'�A����>A��������3rLݺa�e��>A��������� � � ��~��x ���߳��A�A�A�A�>�����lll�������xą�����l��>R&������������cb���������⊽�i�sw��A�A�A�A�w��x ���߳��A�A�A�A�>����
�9����x ��~�3?��ۙ��r���>A��������������>A��������� � � � �~��x � �������nnJ]�7nm���� � � � ��w�pA�6667��~�>A��A�A�����A�666=�߿g �`�`�`���o��eٻi�7s7fn� �`�`�� ����x ��߿o �`�`�`�����pA�66���g �`�`�`�}��6�fMɳ.[���� � � � �~��x � �~��8 �����>A��������� � � � �|�a�i  C���D,A�x`$H�HA�>H��|T��#$�h@"F
Aa-���� DHؚ�g��B+��$�@8�@��|AH1 ��OP$^K�#k+<Q=���YH��u�Oc//�"B�\�.#D��,�a)g	 A $B)� !��$X��@ �@ �Ŋ@�FG��H�+"0�`A�IXR&#(@��0��Py � 0F ``�=$���$�I$�f hG�\bA kB�"�#JS������?`��m Ӛ�nl�l�<=�1R���郞�x�]�+ӻ�a�z��@��v�ݷ��6�&��h���F�kmn�޲���r;l��eMa��<peCf�C����!�)��n]u�譶�
^�Qޓid+9��v9��v�Vk�:1�Н��9��'\�ݤ���������cu4t'i��`��F{p��WF��[�]�i�m������o@^z��UR���WG�`��k�@R��y������E���
�0U*���H!Y�%] $-$���\2���s-!�H9�2����9��n���m�ԏY�y�p�<�mu�O+V�TC�5��;-��PW0�n$�@9�VC�J�k���k��b�nIY�	bth��f�`ym�4P��}�9�'V�۪��6�'�zO0?:���ے޳���	�J�Ƈ��ɮUsz܆y�k�v�3��t�[���خ��; ՗��s�v[����-�����q�CHm�@�{���f�m�Km��%��h$M��I�];:v�Yf�Fz�˶�]]Y���V�r=W,�M��fv��C�+r��ڢ�u�v9���68�� �1ڮ�ɢ�k5�޺n�fNÂ��՜8�jDF@�-�@AOm�T��Y�F�(�耓;2�P�ж�[!�nm�!�հ-���[JKHMԨ	��r��Q,gn�^�<�[;puHm �\F� !K���b�V΢j V+����)Tujt��2�S������u��Ӈ]n�i4[@�`����g.�6w�l>
�㛳�v���S�@��]��y7 ^��(���8J�6&����c����u�;�MѺ�2�T��@:��=�g=8M��ℯ� [Vk��ef�(�Mn�6Gc:����#[��H	 _��z�\nD7k-lU���뭷f�Į1�e:��t��]�v���;�ۜ��`k�L:5Ɋ�}q�Y�2�Nuq�ٝt�mrd��������> y(��}�@"j���'�>�]�I���ws6�M�l�z���]���M��񶬨5�:��'���<d8�n����lb��y�V�((��f�zz�P=��Ju�ɠ�bj5�DXs��Ά9�6ܺ��X�a'I��ܽïk[b�E�m9t����w���2�$���լA7Gl[�9Ks�q������[l��^9�ӭ�x��7b�)Y�Z�-E��]����� �]����w|���������N�lT�B�d���"�v�3���|<��d��wq|��s�L��&f3x��'� � � � �;���|������g �`�`�`�{������߿o �`�`�`��߹,�?\���ٙ3w8 �����>D�Q���A� � ��o �`�`�`�~����A�666=����|�!`�`�`��߿y3&e�n��t�.npA�6667�߿o �`�`�`�}������/�D��g$�����z�$��i��"�M~�K�����7z�ܯA�ESM怹`]ݲ���d�ҒM���~ξ�?�;�zhܶh�n�nBH����3M�է�7)�N�.�&)�6�Є��k�����"$�"qƢN?������f�}�g�AU�������j$Ƣ�BI4����f�ر��t>���8��M���@/-�Q�FA���hܶh]��\�z{l�9�\k��D�M�ܚ]��\�z{l����s���;��㑸d�c��\�z{l��l�*�@�:�*r\�7,�$�ʝ��ʘ:;on7�����%�����[�h�<��Q�;��o��l��l�*�@��k�;�q&7[I&@D�ɠr٠U�^���נ�����߿bE��~I�p�RL�6�@�{���鈉�����s@>�@��,Q'�'#Q'���נ�4�[4;��T�Gh5	d��BH����{4�k�8����:�m�G#ȤPp��&�$E�[КB�ݝ����ѝCu�����l3ح����A(��hܶh[^������ =�zho�cX�!$�ܚ��늣��� m���K5�L��?5"��H6I�����4�蘚���h�w�rKJ�������¯/A��ESm�{��RJ�=3~?f{?fdS��@�wc~mj����K4�>���﾿ �?�@Jh;Tċ�榧��� Ʊ�	�s�g#x-Gg�l��zs�ڎxzE���pVʿ7�4���/���qs����f|��}�{��$��8�Q'���+�陈�.���4��f��%z�*���R,��5�����M ���<��������v�$�Q��(��hy.wޚ������נ�� �j��8FHD��ܚ]��^�z �,��K4��&�*bf#���M��.�k�y�tE����2����*��z]��;f���{,��`�(��Û�����+�Ӳ�"���t���Z�j�b�l�3٢l���<�Z��� j�g��8iwCə��!�a6�em� <qe�p�tz�u��T1��W��5��V�nm>��Nކg\+���?'�@ذ��a��KvЖ\�d�˺��L]	��3����X�l�	s��Aa�\���m%�����k�j��Wb�4��%�-͗4�6�����trY���}3���n��Ү.��܀�0N= ��o��fbA���@���8�����I���6�"��@>�@������@9m�y��D<Na�F��h]��\�z{l��l�-�,Q'��ډ��.v� ��hܶhvנ}�����eV�̔�s�z���i�/V�V��6���P�Z�=M�,d��Ě�z{l��l�*�@��k��A��8�IDܓ@>�_���l����;^�^�7��|��c��47&��}�qs���@>�@�{	֠�P��#�������� ��A�DӴ��	��\]����`�z{l��l�*�@��k�>�Q����f��HHJ8"Żr]=nW��m�,s��������������6�"���wޚ]��\�z{l�;��m�!�s�4��@U�^�GW'z �y���h	_Bʉ51G�Ȓ���.v� �i��칉b�39�z�~��@��=��֪b�B8��٠r٠uvס�ٟ�_o��{��iģ��(��hܶhVנqs��m�@.Z�J)������nm��a2h��yL�V�h8�Ό�M �-��J�i2�ͷ��נqs��m�@>�@�,0N��86I���נ�� ������߳/�����܁ �8�6�@?y,��"�Sn��N�u����kN(����������}���@�����I=���䞊��/��9���'{`&�1�/�4��@궽���@9%���f���DL�R���]�Sq��G>��@nֳ4ɐ\��";V89�n�v��l� Qn��@@�������~`;m��-�Wmz(���"�G	 �z�l��l�:�k�8�����3�A��=�8�sr(���o4�J�s3U��ހso4�+ǎ&� �ɠuvנqs��-�@>�@��X'Z��Y��H�W�^�y%���f���^��pD���������H�!5�L֎�u�t�gt!�69�m<��uû\�Bܽ�����c��;`��C0��T�����,���z����t�V3��n3ͤ��g���U��l�<N��G$,Y��dM���a�)�ۓ�jЦ�:��6�b���,�n�s��ٞNjx%'t�ЋW-r�Z�3[��WR�tt��¶�n"��wn�e�f��n���@�#�?����"���u�ܕ�0�bݝ���[9瘋:��d�vۋ�[���ױXyK���;'�r�hܶh]��\�zz�$��kN$�(���l�:�k�8����٠w���u,x�H���������W���U�� �7�oab�aG"J&���b�����ޚ�-�Wmz(���"�F�"�= �hܶh]��\�z�����3;�y���x�HI$r91t�u'��۝{]۝=2;���!�4[(�$��i��&��> �}�uvנqs���@��8��47&����7�.��Y�'�ė8k�{4����}�f�~����`����Pō�H��N��Y�����h
�w�rKJ�mL���@;m��-�U��{3_o��k�$���ē�,�y���f��[n���ހrK4w�?]�2pj�z�&ĝ.ʤ��/��e��c,��Nu���6�a�U��A�˪�������r� �}3�����@����(���r$�n=���@;m��-�U����%�Q(���z�l��l�`����Č$��!��@~�O nt���MXh4`bl��%E�XE�p��d�Ѕ�m*ODO@2�cF�J�AO pV(h��C�4W�TWE5H(��*'ʏ�
��|��ꀞ �:���v����@/.V'i��&��U�o4M��=^�z�,�=֕ȱ��!�@궽�}� _{�@>�@:Ze�q�5�"�J���
Z�����;j�-ƺ�ݎ�s�m���L֦!��H����@;m��-�ٟ ����/�����܁ �8��٠r٠u[^���׿��bLoͬm�E��M �}�u[^��uv����4�n����#JI4���.v� �h?ٙ����>�,S&H�!IǠqs��-�@>�@궽��b�)b�B�D�����w�SnA�/�7V���N(��N�"&,3�D�4��o߿l��l�:��@��k�˕�ě�$j2G&�}�f��mz;^�v�4.��X�ɎI��ɠu[^���נ�� �����:���6�#�8����٠r٠u[^��ۣxڙ�$'�v՚�sy�M��=^�z�L�I3R�E,Ub���홆��:Y1�m7;h��U���0/E�i;`�-���E�n;�Vx�һ.�ь�k'27l`��=���p�J]�m���K��~A�)R�<�j����6LX�-�y0P;���ZэfJ�e�:��if��Be���L�6�vWf�
��;3���Iع�!=d���玭��]�rl�iC���\����{E�c��OUr�̻r�~@�SӘ[�䲛�t���@��^/��-ɻ'����cmqԆ�[�r��	bocq��������4�k�8����٠w���u,n(��RI�u[^���נ�� ����}�X�	$"���.v� �hܶhVנs�'P�JD����r= �hܶhVנqs������N@rG#�@>�@궽���@;m��r��i���ڛ��z$�����S���W1֗m�>p���H+\��\�ֲ��m�}�������@;m��-��a�j���6S3%��I=����� ��G��a}=4�ޚU���7����b���f�}�f��mz;^��ۂcu��I1̄rhw�k�u[^���T �{٠^vm�51~��$�:�Z;^�s�� ������|�i<����B9E#g5���{�vJ��=��:4mr�غD��29�dN/�����v٠r٠s�ՠs�'P�K&)1���z��4�[4uڴ.v� �;��ĥUKl��[��t�=�Y�0X@�".DaDL<�v� ���}�cX�P�@ ۓ@�]�@��k�v٠r٠^v&��,�7"qh\�z��4�[4uڴq��S��xH7B�����6��.̘}ۍ�''��xn�g�S�la-VoS#r���v٠r٠s�ՠqs��V���md�Ls!���f�@�{���&�@Q�6�b�Q~��$�:�Z;^�s�� �����ʔX�L�jLs"yZ��;�M�~�Y�s�f&&o3��;�V��ibQ&LncI1����hܶh�h\�z�uU�DS��N�xt�;Vv�Of�[u�!U\꧌�<b����+�\�9�f�<��f�@�{����@ro4��X�95 rh�h\�z��4�[4�a�h��Acr'�}�٠�@>�l�9�j�;�toS"rcĜ���4�v��v� �;f��n	���I$�G&�}�f�λV�s��@9�f����}|P��\��P3���6��+�뎆B�%��z��0#hx��q!�#�ޱ�(��yk�n�vp1m�a���ZYp\NT�\g�@�Ƥ������l5��d�]O�N}�u$�z�9�퓩y�f��`�rXv�rtc'���gmJ�[YH�v�s�%�J���xI3��mm�܊f'J��˽�|-�Vtlt8�
3GZ�
ll��tyqKA�g�1/�L�\U��uݎ:<%3�sC�\u�Ӱ-�0og�m�틔Gkt�$[��m���m)$��Z�v� �m��-���*Mb�2dd��e^V�{ܳ~������h���=֒�9��J$ɍ�!crM �m��-�:�Z�;f�w����N@rG#�@>�l�9�j���4=�v��@;�䱬p�Rdrw��v��$���|�G]�jI%�;g�$���׿�k.�q���m�y^���v��e΄6B�oT��s�+��)��Ú(��$�;}>�$��TԒK�vϾI.�kz�K���7���91�NO�I#����J��bˉ,��w���m�OzMI$��l�����q��#�jI%�;g�$�[��I$��l��:�SRI\�tn�����$�|�����I%�;g�$��=I$��l��\�U6�s"��1�ԒK��|�K��5���}��6��{�km�.��yRU�YĔ�u�W`�r#î�X';N1��3	 ;�:���Dc/\��r��� ~�~٭��;�^q��s�s[m���^q���ʱ8���HH�z�I}�g�$�S�=I$�����$��RI.w�,k ݢ$��o�=�5���~���jIfb3طv9���m���^q���Q1���"��I$��l���v��$���|���߽�5$����xڙsǉ9>�$�v��$���|�I[dԒK�vϾI.v%�F��Cf�HI�8"Żr\1�0kn`�v�[;��Ѻ��ܗa����#����I$�����$��MI$�����%S�=I%��tn���JI>�$��ɩ$�9�>�$�v�������� ����(���k��I$�����%S�=K�k����$�^����}���B:�UI`�Q�y���IO9�'�$�;�O�I$��jI�ř�����7~4Tsw~�w�-�_{ٖ�ۛ�53� ��}�~~ }�_���_���O�I*���I%���DI��)�c=����p�F�M��q2�T��m�wGfR+<�/3'G4rV�YZ�� �~�� �s�}�IT�O��3��K����$����k]U�E�vۭ��{��9�3�?�~�z�Is����[f��ۣxڙs����9ZU���h�fbb�M����h�`��mBH���8�?�fEW����� ��f��13�7Zλ�m�DM��RI��� �>��>����s���=�՚��b� @#x+�j`0�G�`	b		 0Q�8)�%�`c� �F8E�Ⱥ'&)�j�� �H�	(K�-�<C��Bx=�x�Lv#��F` .EXE@i�Q�@�z�w����b�5�e�l�� $ "j�)��@�Ո� @����vۻ����8Im]6�l	�{C��U��q�`���*�ԩfY^W���� F�E���8�̊.�`D"�A�]nL8
���w���X�ӷC�M�#�/[�=����]ֶ[R5��`�&X6�[��؝�Pp�A�mn�-t �V�(WxW��O�O`ت஋F8nN�ݮֺ;&�����Wl����%n��g�v�k��#�Wu�l��I���ٳ �-�ܲK��6텶YA�i� ��pm@����UT���������Dr�T܂�H$&�H5Ul�&�$ݮ�[�V3rܬ�Q�M���t� VI��gNޥv��V�klb�P��!�i(�':��Bl ��9�kg�k���[٪2,��J�r\�s<�����[�"қ�7i��f��&'SF�v��`}e��Z�l�(ZW)a۶b��7F���mHJ�V�i`w&8���1 Nz�@'�y���y�ڵ��&8��26�Y1ve���h�r�۝Tl�uJ��8�ڭU��w�K�%�t�����0�*z��Rs�<VN�W����Q��դ�7c��]���8���g�kS������Q���N�����S6�kE�#��'"����U����U3a@���#YW3�(���ʫK�2pV)�P�Ep��.�R�<�H/����:EQ�by�^�<�[tn9 ��Mk9�2uB^emSUJ��u�
8�Z5�R�mH�q�P*����ZZrҀ`�m��������mU�&��X��#���$��^��D9]>�ó[o[yZ^ݚ����i'#�q�Q�v2e���kZ�c{Vw�������ط�Uu��JF�V���F��9ϪR�-��׳ۡ��f[j��\5�*����5[&��d:Ym㶶J�j�� �Id6��cư�S�S�mmɉ02�scV�dPy����m[J�E��V�$�N�QO��MS@�U>G�<Q8�t�?���}�پ�ɗlٳsvfm5�J�%n�l�{tn�#���Z�w^ۜ��nw�:�A/rXҼs���f%z��6ݦ�v]�VI!��Gb�hn;]�b���xĠ;���=�Ї=��n��Ng	�vt��R�Z6�Υm+�Y�d�Yv3�v�Xv��S�W:�8zݧj��<N
�^����jx2:U㳸uZ��]�gu��1]�G6�l�Z�s�ۥ�[���V6TT*[[N�:���3����{��?��]Xm�yuw������Z��g�D�DLq�����_�1(���b7$�9ZU���h$�@=�Y�&b"*�]�y�Ĝ�9�(��wޚ�l�s�h�ՠuv�cX�XԀwy�fb*�o4�N�V�h8�����h��h��B1��4�Z�V�h�,�If��>�]�������]�ab��Mtg����c=�a$]��nN��_�{�~|��]q9�g����?����@;m�W-zm�&7ۗw7\�w6�I=���pQ�C��J�""&\G��y�z�w�r��~��u�o�"h�FԒM ������^���Z�[4�T�q� ��q���8�k�;]�@9�f�v�4[�J&�6�!1���j�r٠�� ��� �:�jĘ��q�c$Ju'@�۝h��l�k�t;c*��1B�:I��q)!�7qh9�4�٠r�������w��1�r,j@*�3@9%��"f�=��ݷZ�v���7�D���@>�Bw���MU_�� �C���r�h�����ȓ��$����������m�@>�@���jI'�(��s�h�� ����j��E֕Ħ&��<�m�gC��8��'hj��c,��Қ7&ye�&W�{*�cM�ڎI��4�[4]�@9�٠^�6�C�rD8�rh�%�V�h��4.Y�&b&���~BQ(E�L��4y�- �;f�b&b�m<�sy�.�
*�*�3*�4�H��s�h��@>�C��`� �����$��߻a��5 rh��@>�@��� ��f��fbf]���.0�,���*��ňH�-g��t�X�ؓ���8�.����w@m�'�����o���-}�@9�٠�4��K#S!$NA�U�h	ZU�D��D�}v	?�@>��@>�@���jD��2Š�VhIf���7�v�h
=}�ڥ�8�蚎I��4�[4]�C߱.��h��ɴ�7 �&9rh�%�V�h��4.Y�dϢeJ��E�-��I�	�m��nIM�^��;Jf���n'n���.L��d�w2�֤�,�pk�qe�`Ө6�%��vqv	�l�n���n܁p���i�Y�f7`g�<g� �ۆm�W;T��Ax��uYnyz���!�3��X�i:$��9�m�z^
¾8�ֽ��"+4ĤrO�8u��1l�]��Q��5"�����nS/J�5ٝ>{���u�Y�l�0�wۥ���-��s�װQ�,�z���y؉J��.1�W��N��� �,������@���bN%$�H�y$�@9�ٿ߿f~�H=��@=�怕��bj��t]E�U�� �mɠ����lӿ�%Wj��޺;�vA�(��?,���z���h9�4�٠��Pd�)�.*�3@J�V��fb�������-��>��Q�!ģ�&�I��;_�0����6����5ns�[��]ѓ7+�r�9���/�;���� ����~����3����hB����U��S�u�@-�3���[4�ڴ����߿$s�?&�Ĥ	1Ȝ�@9�zh�ՠ�l�{f��ct�8ʺ�(�����陉���V�$�� �٠r٠^;�q)$RF��$� ��f��"fi�������U�ߝ��I��ڂ�$����$6eJ��Nn� �G:]��N<���=dݪ2sC�@&�rh�� ����j�g��������%��q'�ɑ�I4�[4�*�{�hIf�1D�݇���Pd�)�'&�������s��O���Y10�"ff���h.y�rYcu�#��#�C�?%��M ���r٠Z�Z�>��t���&��� �Y�9��sy���{�h���}֔�g�i��q�c�K��3���,����C�	�Z��)pV��Erhܶh�V�s��� =�zh��<Ƣ�"jcIbrM�j���17`��� �y���k�������_���8��&��$Zo���[l��l�-v� �Z\k��8�i���⩶�@=�怕�Z3���}U<����y$���-39sndٓ#b�hܶh�V�s��@-�������{�JD�q<6q�A�6d��=����F02e��ջ�2�u�2�$��-v� �;f�[l�ϐ�4�L�jG'�G�s��@K4���+J�蘉���Ϣ���o�C�3��rM ������-�ffb^����w��@��:�S��	$Q;������h�u��,��f&&b*���w�JyD��1,�@�ڴ3M��� }��f�~�Y�)�fc��?��~|�}`�E	���.7,ȝs����#��t��=͵�N�s�\�s�ʝ��[R�wE�!�.��g���t���*��]�V�>d�qi����+�����:�Hv��k=�-�["�J�9�b�ų[��fy��mf�l���[�$��6�wkk>��ׯg/�ձ^hL.\��9�Ӥ���^ 9�`��uL>�m1[���,Y"Muvxt���k�ٶ�M��p��t�3GaӶ*�ĜQ�q��/�;���4�[?�A�?yhw�=�cq8�M6�hIf�1A�o4��{�h�j4k�� ���-��ՠ�l�m�yڒ�&H�n1�NM�j�s�h����zhޘ&'攎O��- �;f�[�4�[4_j�;�,�I���3�u3�s@�������!����m)��+���aن���m�!��9��z�hܶh������M��~Q���'7wn���I'����>E@�	533�1�=��@<�� K�o�G{�?!(��R6%��h�Z�v�?��bG�}4����z��JI#�&�$Z�v� ���-�ٟ���o�V�B��躋���������\�@�"+��~;N�����?�����"�Z'"��9���+��6[.t!�Z;����t$���ܟ#��
C&F���o���;_j�s�hol���(2d#��<Iɠv�վ�����O44�@?y,�9vAVU���O��@9�٠��N~�r��K�[)(J�$�
d�����H2��
�kJ@����Z�< 	�W�a��E���a����5B$��xFH���r�C`R$,�$$BF�$�� �3����	,*ŉ	0�*"Ĉŋ��H��$����dK�F,F, �1�ȁ
d �,!$
� @!=>��� Њ��b��b	�����+�0��@
<P�W�O�	3�{��{��Z�>��tD�E�9�C�3��īO4��h��h��4��YtfPa��VU�f�~�Y�}3�LDC�_�������4�q�QI#c�O!�wM�pV��x�+/�:�Lfz��J�"˵1���nHؖI�v�ՠ�Vh.X�f"P��@j�
�ʬ���pr- �;f�v�� �������ٟ�f$�x�5���j4ۓ@;��r٠w�S@9�٠^[�c�o*��*�4�D�W���<f�'����y��"�� ����@>�j��&5J1�NM����r� ����f���P��Y�W����JA)zT]2�Nt��kps�����]5۴S���f~��֔�O�9�{�����@>�@�,��s��&�U���^e�f�yr�s5A�o4���l��bG-��4�����%�h4�@�,F�DEP���i��Tt��D�X�C�3?~��}�4sy�\�C航�h[aUyU�$�!���w���33�bﯧ�i��X� s3.d����0��"�oa�)��#�Fn�-�]�H��YQ����f��Y,t�#��Oj�6���!r;����	CWF��4t��aȑk3	��+J���T;�b�탲��svl5�`����3=q(b�q ��<��ys��� X�d6�%N�9�GnSۮ�fթ��7���C]W�0C[&Yul���61/mHM�{��V�uA:�vx�֟˗E��q�	v'��YTh�HWu��KS�55�D��M6������^٠w�S�?|�������ؖ6k�����\�@�,F�w�� ���c�l?���d���<�@���ƀw�� ����4{0O�)��`^a��b�sy��� ��ye4gpM�(�����I����LEsO? ��Z�K4O�
���9��is�ۥ�nֳ��.T(��(�[�\@-�%����_6����f��ҭ �%�~�o4n����T���j[n�����WAp ��&2fbc��x�����{�f�x��J8�%#r- �-��Vh�"*���@Nۭ �r��Wy&�mɠ�� �-�k�h{?g�K�����}�Ǎl#P��$�q,�>�O����rK4�9�����-�]�Б
Q����&Q��;��v�μׯ5��YcWhn���iV�{�f�rK>����sy�&��~iH��28���hm�@9�f���[��ى:�	�����rM ����s��9����r� �-���uF����ĢnM~���[�;n��K4>�������qx�Y!"hXܓ@�v� �-��l�r٠{3�fy��r	bs�):F^4�דf�/[$�z;c����Pƥ8Z?���H�A'�H8�R. [��4�٠�@�v� �v��i9(�ܚ�l�r٠v�V�s���fbb�|�UE���XFav^fhss@�v� �-��l���&�q�I2dx��@�v� �-��l����D��"	�
�@����y���1?4�r~�Z�[4�٠�@�v�߿/QV{���eM̝��,��j;jy:��Kz-���IȎy��6�P�C��> ����s���ڽ��>@w���9��i���E��4��h�ՠ�@;m����z5����Jޞ�����{4��h��Iģ��8��@/-��l��٠v�V�e�+8�n~rhm�@/{f���Zyl�?n~�3�N�EB-�*mV�se�皹�G��	�	A���-ɹ�!%�K;��^�uc�дavZU�%m�U!�����:�\F�v��@��\�q�u֪��l˴ӱ��j]�I��`�݄��ּj�7=c�'09�!��mU��p1N]�� �y!�G+�-�sVq�XG�J�j���.�z{�ϝ�܍�Ӷ��pF�V���n�zs�d~w�w==���Iؗ�)-��j�$B��،\\�v#�nV��s����@���89ƶ�d�c�p��h�ՠ�� �h��L����y6��9ZU��f�rK4w,�3T&���ҊI�3qh��M �i���33=o��|��s.$ۢ�)������?L�]���4�������٠}��\i���$Q(��@r���Z ��h$�@��m:őPMe��a�Af��z�{Ոw[� ��0����O�{�"m[���33�?��@�� �h�Y�/;A'n(���JE��͹����~ȋ�x�h4�@�iV�Gr��I��Q��4�٠��@�v� �-��n%��F���ɡ�����������4���@;�f�r����<���Ebr[�}�����X�/☘�k����h�,�XA�J͞zq.N^�����L.�8��CX욷*ku��Y�tdӛ��8d ��s1����٠��@9{f���V��\�&ۢ/�*�/34�,ߢb"*��y�'k�@;�f��Z���6�D�rM$����$�w>���� �Z)�,"?E��C������hi����xd�#�I4�ڴ��hol�^٠Z�cN(�sq)�w���b"'舉�?����h���m��{��?M��i��$-qF�[7B����m�'^�d�c��'�i�2#u����� ��4˖h��9���@.��@�o�,f��2A��4��h��hy,�\�~�����AWV8��̚�ȫ��;N���i�D�P�}4���of	�֔JE���@;�f�r���4:"b"6""����30^��\V�m����'#�h.Y�\�@�|�@;�f���h�n��)4��-��ݒr��k�)uiW��Ȅ�sKT+2%˶��3@<�f���V�w��3��M<�;�F�(/�A�X�@�}�@;�f�v�� ���ٙ�����$��71G�h�4��h/l�-}�@3��b��B<mɡ���?$�y�'�Wʴ>����|�hI�X�R'd�crh�l�-}�@=�z�������� J�wP��h�����1�3�PJ�aZ��A2H�8�q��j�S�x��x�`Z/��C�I��8���S�������@�����k���t�wO�����~~�_�-� ����`-���K(:mjnͶUV��mu\kc�M+eAy�U#��+('�D�m�U�㍭���-�V0;cjͅ��Cql[�%���UM���A`
�U�mx1�h!�n5�J��4rsu�u��햎��Bj�0'��ϋHv��(��W�nZP8��(]��j2j6��;��H���۩ÃGR�:�r������Ɵ9Z�"�Y�ɧu����;� S�٪V�}�Q�U���Ԭ�r� �l\�UU*��p/kd ��)%�Pu,vΊ�M��:FZ��H��ϋe���kǕ�9Ρݝ��n�kui����vZ4��s��%�4���`�ɤ��-�l�NR/nX��@J�s��	���v^]n�W*�O+�F�	��\uy�lU�Nt��P�m�gt4�tM�9���!��i�N:F�l�Ʃ������9��հ���v�S����7�a��j��рٝ�m����8�۔�nŻa��S� l���6���gc)2Ha��qp�9q���Y�k���g�9�Hv�hlX�f�q��YnZP9w6Df ������5�r��=t�,����˵�]�"^��!R�[���`���Uڐ�q�Ű�eU�Vڤ)�6��U3a@���u֕�耡wX�<�J����Yq�Q�U����Z��nz

]�.�ki[W-��y5�l�$j�.0�� ]I�GUFN�@��֑jU�V�QN:B�۹�i�ꖶ����G�.�k�&��Hp��v����ڭ ��/��,Om���q��'d1��[zC�ce�"g��w5�\����.��@��ɑ��P@�K��$��ɸ]��;qUX��m�n�˱�m���tT jH�3��Լ�Pu�Mm�	��lCu�+�mq��q�r��U�*�]tӄ�pC�+i�v0�V��{q��V��Ej�����#JۄT�)k�vKfy\�=	����6L%�<��<�\"�~b
|��| ������x�4O@�Y��|8���7A�Uւ	�:�3>�Bԗn4r�n9{N7����fy�+i��vi�5e]�<���=v;#u����06�f����`.�EY��n�Ô�m�n����8�D���5� YÉvYw]�F�� aŅ��#�څ�]����c����KWF�);]v�ֳr<��H�<N�͕���2���nk��al36̰∗�7am�+dڸe1E���gt	�_e�nOi99u���I.g��v�ѱl#�*מ�V�vߕ� ^K4.X�&b#� �y�'f	����dc#�@/-�ol�ܳ@J�V�����:+�wL������rM ����^���ڴ�٠}�]q��h		�h~��?%�h�u��f��13M��7��P_�"�`�I&�k�Z��}���}4��h�v�c�"�D�Ly\�wM�.1�u��F�F�x8nu�{�4v�5_�����=���#Y1I�������@���>�����u���eE��7f͸ff�$�����* E[�TU�os@~��@;�f�315G�qk�D��lnM ﯦ�k�Z�[4�٠�A4ˉȧ��nM+�Z�K4.Y��"fb��y�_Y�Ɵ�Q)F28���h�Y�\�@J�V��LCdc.�W�m���Y�&�nh��<�v3r�F�<�6�G��łU�������)�t��5~�����h�,��U�1����`�hq�A����4_j��Y�	r��&b*�o.�XT�FV]]���7iրw��6�f=DAI1��~�o�@;�٠^�T&F�&e�efV�w�� K�h�,��b&b>������h��T^��YWw��	r� ��Wʴ��h��].�6xyM�I��XeD�{��6K���A���笚�G��5���Q]n��k��y�%|�@;�f�%�4�ঙr9"2dx��@��� �-�ol�^٠w�bXӱ(��#Z�K4.Y��TsO4�:�=��6���?19�@-���4_jп�fo���+�4�M��$HԂi�4��h�ՠ�@-�������o�x�B��Ig�l+<�]�`l�h#)��s��
�2R��B0X�s��HrI�Z�Z�[4�f�r���¡26�(�8�hyl�~��6�h4�@Jҭs3T����Ff^U���hm�.�9���m��@=�zhw�f���lrMM'�v�h�Y�	%��p&�Q"�c��&�k�h������I�����$��wy$�P��AE"�/v����W,��m��(���]�SBX���8�g�Z�0/O��X�=����E�d�y.{%Jڲj�U��ƺ� �:����S��y�Y#�m�E:nv��<�+%�̆�Z4�8�.&E�ē����me(��d'm�ɭ��Jk�mi�qS�a���
e����9M��Ib���;��l�v��@Pv�0���z���\�^gk�ww��`��__o{��LJ^�L�Ӓs�t�`z�m;>=F��h���[7�C���I�Ͷ�����m�@/{f�k�h�z	�b����rM ��h�l�-}�@/-����ɴ9�r9Mɠ��@�ڴ�٠�������	"I&�k�Zyl�{f�^���Ubdo�R- �K4M���O4��h<�?ՐV�b2�&�㫬[��ˢ1��xH��T.��֦���� �V�sfئ�V�6�i�.�Wʴy,�?w ��]��Ei!%���ځfb��$��b3��h\�@��pUՊ��kG��4_j��f�[�4��h�LN��'&LMG�^[4�٠��@�����pM�8��'#�h��@/{f�k�Zyl���&%�#�#c�8d��V�g1Y��lRY�iŊ��Շ9܉
f��q�$��٠Z�V�^[4�٠r��2!�đ$�@��q@����� ]�4�R����bR!��@/-�ol��#�ӈ=������Z������<mɠ�� ����h�@����5I�b��ɠ��@��� ��h��@2��r�"Dkam���H�-d���}�X�nARN]�5ۙx��K[�WQ�O+_6�~��h�i4�٠��@�,Ę�mdNL���- ��&�����٠}����f,�Χ�!��Z�\���L��� ]�4��h�#4��51�	������Ľo�����גI�~��I�z��RuD �H�E���3�o$�w��vf$ƣD�M�ڴ�ol��٠{�~�o�m��4�6��"EKT�<u�{:���n�{Q;)�V�(�\�������ș����qp����ol��٠Z�V�e�+89�9#x��4.Y��f��� ^�f�����a�I2�ܚ�}4_j���h��@9΂i���E�W��%|�@��	r�31U޾��Loͬ�ɓ�8���&�[�4��h�ՠw��LI��ٶl�X)X�3�[=�F^�Z���=�k�9/mn�%J�fŢ-3�U�XJ�^B�˙��2�p�[�cg�'|n>ujњ4ۣ���5�b�zÞݵn*1�gs�Z��I]�����t'f�Jc�{N��e��K��G+��T���	B�����v�.Y�;��4L��р�h:��K�#��f�Wb�Um�ܚ�wl{��߽�ή���~=E�6��lm; ��D�cm��u�&�ti1��9����oڑ29�	��&�{޳@/{f����舉�����|�W�wWY�q9�h/l�-}�@;��h��@�u:��Lj1$9$�-|�@;܌��bbf"����h����V�dL�JD8�h�i4�٠q^נZ�V�gm�ŎcrF�.���f���G�11�_������i4����9#ciL��,<�
P� �����v��!�s�,¸3@f�&5�b���$�8�k�-v� �;I��� �:	�Q�Y �8�$�s��AT��6��0� �@��PC��/�A@��=�M�w��� ��7���߱"�D�ߛX��'qhM��	%�9���ͼ���@�~�.e�ܛ�칻��y'�?�Es?������@Jҭ �H�{��]ը�ۉț�@>���j���h������ĠA'"�d�b�<M�������D� N�^�;���{���bz��Lj1$)$�����hyi4�f�}{f�k�m&D��Hڎ'�w��@-�h׶h�V�3�~H��=�LIȤƤ&�{���I<���M<�� #MlKBZv$d�;R	��� D���D��x��
_|.&�<F	�S	qBBzD���!@H��H���]�@#�I�Фe%=G�˔��x�m�)
��B(s��(�D�F�� �T�}O����#~ADP�|�w����}S=���;�{y$�^ܚ��L68�%���I�v٠%iV�{�Fh9������
ʶ�Ә�A�MɠZ�Z����m��{f������`^��O##J"㱫���/����۾wT�.�p��\�e��Fv��*Ln6�)&,N4��}��m�@?w,����@ݷZ�l*�U��a	�$ɠ�4����j��ۓ@��U6��sdNDܚ�{f���Z8����8� |�h	,�UX]�Ln1$(���g����_- �ɠ����;�����[I�20R1��fV�~�Q������h����m����\zG+(U��z*sh��(�n�n6�vv�m�\r���M�M��ٜ'"�s&�^[4������ ���4�ۍ�n<�d��ܚ;^��Dݟ;V�r��� ^K7虚��)A�
'1d��G�z��rܚyl�8���rĘ�mbRLX�i�h}3^��4�y�z����ʴ�ڱ�r(bq�2h�@���|���N��������鈙����+�T�_�n�ɗl36�&�ʷl���[���u��z�<��t��m�5�:�FѺNԜ��� �!A��~ٽ�H�m�ɥ/j�DK�j��(#�̱�1�`#f�<o]�ۦ��sm�s<]�����욆î�}�DӠ�+��e��&���j
m.���½f��ZQ�s��LQQS��q�Γ�an��f��瀹1���7��	��gtk�m�w�^������������\��9�:y��qa��i�:�D��e�*�I��dNE$����@�}�@>�?߳��wޚ�蟒�`L�&������hܷ&�^[4.v����L�����N- �����f����%���z���r�c�S�E172h�@��k�/_j��nM���X�Mɑ,���@��k�=���Y|� �}�yl�9ޘ���EE9%�R��=X���:Lx�/�A��E�걞Xl�,LI�!D�,�A���ڴ�[�@/-��uv���Lo���#�]ܹ��O��ww��T��P9�?]��<��=������6�Lr(by�h�@��k���fb^��hv�M�T�j1�M�9�h~��&��;���@��,� ^K4�UԘ�LRE�R=������h�@��k�>�cx�8!8�!��黥�6.�;/7 ��C�au�^��dث����s[I��S#j8�_Wo���f������� �w�@;۞b��2Dԃ�M ��o�3?~��]�z��ZW��k���fbn�o躋6��#2���˼��?�@]|�E?�g陕EDLM���~�� ��总���Ee^EFd^�zfbi�N�\��^[4�;^��X���x�8��#W��u{�f��L�M>o?���@]|�����3� �3�?�^n�(�!�nh��Ej;a��ͺ�D�;��1Ώa1"ݸ.��P��8������˝�@�}�@��l�ܱ�j1�I�8Ԓh�r��f?�"f.ϝ��@t�ٚ ��o߳�~H���PX�%"Q#�=]��:��&�^[4.v����X�YYf]�^U�h9�ff"�'�f�|��4'�߻����D5Y#���b_b{��k����5)���i334y,�>��N� էZW�fhm�����N���,<��%�tX������H��Ս��������v~\��Mb��ܟ���^�ՠus�M ��h���:���1�H��ڴ�vɠ�� ���@�,M�u�X�N��z�}�t����ŉbQ���������\]�&Չ�EO#����f�~�Y�.�U����;m�h��j1�I�8Ԓh�٠DDCX�~�o3@���W�3��$!�$������d�*�n��P	V�ۃsӬ�0�k���νmrV�^�w1�7&������Ų KǙH��8]K;k�!��:ns[t�琭�@����G/��"v���|�o�ae6��l��8ب�����4��f���[F�aT�����5��va�=b�h9vNe���.��YVQ���A������k���Gb� N�	�nk9�=��5Aq���U�7<��f�!|�l/G:�ʋ�%*2��n
�&��u��Um�@/-���h��Ŏ5�`�mG�@��&��~����M �����/_j���b�A2E�rM ��h�٠^�ՠUm�@����3R��k6�����@�}�@��&���}�w�&�����1�rM�����&�^[4��4��t����wrk�'"n,��-ۭ����lZ�_)��6��S�^Yx��'�yz�M ��h׶f|���-د�M���G��I��͹N٠^>ՠUz���$uwǜi�1�JLN5$��_M���?�%���4��������D��hB�3C阦�:�5o4.Y�⫚y�{���X�X�)&5N-��f�[�4��h�ՠs�n�h�)+ЮMCŮ��n��#�k�Ds0�ͱbnM�Z$Jdb�A!�$rh��@9{f�k�]ϐU�\�v�x�Q��,X��@9θz�ՠu^�4�ٿؑm�6����!1�rM�w�d���;��>PH��@�����o��}�t���RzDԖ!�$��*�ɠ�� ��4?�?c���-���M��4�H�<��4�٠[f�k�ZV�4��e�]!a��>ͺ^ʡv3��9\�m�XJ�덮�9���.n
ᑫ��}m���h[d�{f���u&,�	�4�(��-}�}�^���z�h�٠Z�X�X�)&8�ZV�4�٠[f�k�Z�nT,q�����I����/z�h=�Wʴ>�&	�""&!EN=��4��5��y"ō�94�l�-}�@��&�[�4��ܮ8aI:<[�b�i�c��lPlv�7݂�̧@1�6�B��P��&�k�Z�����c��f=`w�}�_e]���qQw�r4����&�[�4�l�-}�@��pM�F�6��L�ol��,��LDU7iր$�f�{Ȳ��SĜ�9&�}m���h{ۓ@-�+�Ԙ�A��G&��� ���	r� ��� ���`E�T�`Bā�$Na.R�ۇ�dyk�%�%Ms�f��%���	v$�k�ۉR21Hp�@��q! �\ >(�꿈�0��0,����=4��,
@�cĐ�`�������^<�da��FI$*�d��	
����cZ�DZZ�0��0D�  �"Ń"E A �cbE�@���OE�@`N� �U/~��?<�m� � -*�j�v�q�,Ǖ��:r%sM�V06B۶�[m�{��{�K�:�d�XK��^xHs�;E�s��kn.5h�Ob�ã1;p�UwV,+rڶٶ�"bKoNٮH�M��v�y�nw!\�WAWd]�y����.f���T ��Y��x'z۫����<�x�JǇ��:�D�͘��q��n���s r��m\�jJ�;�<�];9�j3����m%1��]���X
R��A���Z��T�* ��ki3FMj���5+�+*\�#*�@��[@�5Sc�[M6�v�]װ��v�N�S����(�V;SYT�l�r=ܐ<�-���ZZ�jڕ\@8��J�Of�R�įl�4���'���l�m���׬3���C�RZ�1<z{ny-���@���b)^�A�Sa��n���s*n 0��nj燄�S�N���<�gp��İȃ��^6�
>�R��0&Ų�r�1�����(�=<�)�<tb�f%�)�����y4�O]���6����|��p�n4�X�bj[;���ǩ�Њ�gPU����xz�\˲�v�%rڶ�ھϝ�*\��p�-�Ͷ�M�N۹��i
$ݱɊ��vV�H�d�AZ͋m�D��j��P7X�2�q�I��$�t���l �x�ml�cq*k�q��ʨ�r�9-Ur�k���ah����(����5y5m�e�u�)AmBF�R�걎	@�ݫ@�%�Sg^��i6p�qh�c�e��W�PnR�P�\�ӷ ��&Wiv㎧i� �3��j0��0+qgF^:&�v�ڥ��7b �uD�6�Km�6uTN��$�4 �Pڊb�ex	��sD�5<�F+�jÇ����"�z�[�'iX8��$6���5mSШūc�L��V�&�\���u�Wڔ���r!%ͺ�:�ۂ���73��E��׶��`G�n����{������S���C�� x��/�5�" CO9���	G\a�s�y��O�>+�RH�n�����T��jV��Z;/.qZ�f�r��@�Ni�S"��ɷC;�\�64=M�K=�����Gv[-�8�ȴj�d��l�o7�zy��<ON����?~6�M�-A��G!��q�c�{.� .`y�q�q��L���]V�v`ʙluM�كƑ��Ʈ�@��9w���lTߟ�ww{��?��aF���3.mOO�y=u�:�%c��e=��Y�n�٘�+�^��cN�-RY]�����yl���@�}�@���K�a!�m̚yl��A�{�@�w�@>��+�ŋbl��F����5$$��6�@]|�O�&"�I8� m<�9�ěN�D�,�'$�-}�@;ܣ4.Y��L�D�W�y�.yWqN�*.���̺�� ���}1M���<ߦ�k�Z�t]epI�Q�Q�Ni1�'B������ꕀΰum.8y�<�Տ#�R
4)6�p�ol���@��� �m&�s�cn�M�I�8Ӓi$����r�!��<�۟�^I'￿����������d�4�(��-}�@;�I��� ��4]U���Q�LR8�Z��3?bV���4�@?$�C�o��;tT^]T�D܄�{f�}m���h{n�m�������˄.�\�D�D)B�s�F�n��4FLvG�ZSa#�NtJ�X��'&�}m���h{i?�f~���_M��&�=�'1d��9&�U��*�&���� �������U16��9qh{i4�٤�߱%䳪�視_]ݟy�yG���wX^]�艋��f�w�}���h{i4��m��717q�34�K4��N� $��%�4}���N�3�H���j��z�OU&����9ED�`��`t䤿����|>�R),Q���Z�ܳ@-��l�-uV&F�E#��qH���f�~����|�h6�@]|�@U�j*��%��	�I��� �i����w�@-�zhw��j��D��7&��Uͼ���@;�,Щ���ʱr٠s��6�r4�,s'$�/_j�>��<� ���$�@J��yxX.����p����D���j�Tskku��Y�FR]�^"��4�|�o�߽��yl�[f�z�V�Wn	�Ei��y&�^[7� ��z����4���n�M�MĜjI4�,�_*���EP��� ��Ӣ��1w�8y�@���;-x���L��w�����Kı/׽��Ȗ%�b^���Ȗ%�b^��ڜ�bX��}���Pt8�n��>{�7���x�/o{7�,K��9��߷��Kı/���Ȗ%�bw�����K���s�9�P���,�FJ�i�ͳ���'��Y3��^�\��Y_��A]��*�[X,��hDD�\t%�]T�0�J�9�6S���]]�W>���$%$�e�F)�s��*5�*gb6�\�w>���v:-grs.Q����Lm\me����=pg�����cs3�����?���.l�\��k��<�j9�8ۘ����1O�\*Yĺ�Լ�}������w~~w_��?:�,KM��ͣK.d�m�m����q�&��a�͜��kKpsAڵ�ɗvn'bX�%�{���Ȗ%�b^��ڜ�bX�'~߻x�D�,Jb~~�f-1313��E�v*d$�qp��L��O�OW�E��(%����׉�Kı/����ND�,K���x�D�,K�ۙrtܹ�3L.n�ND�,K�oݼO"X�%�~�;���bX�%���<�bX�%��ݩȖ%�b{�ys�ɻ�f�\���%�bX��ӻ�Ȗ%�b^���Ȗ%�b_��ڜ�bX�ȟ����O"X�%��g����]�(2Y�����������\11,K�����Kı;�����%�bX��ӻ�Ȗ%�b|{�2�ٻ�54g�����4	�s�l<�)�㱇��]J�rY�ͥ�*�acL�_=ߙ,KĿw;�9ı,N��v�<�bX�%����r%�bX��������L��]��p�V�]`Ӳ׋�,K����o�T?��L�Ȗ%��sq9ı,K����O"X�%�~�wjr%�bX��{��rm���K$�W��bf&bf'�����Kı/}�w��Kı/���ND�,K�oݼO"X�%������n�m۳.�t���K��?}���<�bX�%����9ı,N��v�<�bX�%����r%�bX�����vQ��[��bf&bf'���ND�,K�?����ObX�%�{~��Ȗ%�b^���Ȗ%�bw��G�P7Ob]إ�ۛh40F���;+&⍹���\��4p������s�n�ND�,K�oݼO"X�%�~���ND�,K���x�D�,K�����131}���;al��<���%�bX������Kı/}�w��Kı/���ND�,K�_��L��L��y7'�v1�B�l�ND�,K���x�D�,K�����K ~�B��[�8�&�������%�bX�����ND�L��O��I$���V��wLK?�dL��~ڜ�bX�'��^'�,KĿ^�n'"X�%�{�{�O#���ow��������h�|�bX�'~߻x�D�,K���q9ı,K�{��yı,K߳�S�&bf&b��=qz�5%m��,�6uwE��V�p����+n�Xy���9^�!�*�eC��ıG�w���oq�����>9ı,K�{��yı,K߳�C�y"X�'��^'�,K��w�ii���v�˦]ٸ��bX�%���<��9"X��s���Kı?w{��<�bX�%��f�r%�bX�}��jt�Q��[��bf&bf'߳�S�,K��=����%����/����ND�,K������%�bX�}v�˓��f��0��ڜ�bY��02'��gȖ%�b_��鸜�bX�%���x�D�,����$��hƢAhA!(��xD����jr%�bX�~��.awrn�f�ss��Kı/o{7�,Kľ{��Ȗ%�b^��ڜ�bX�'����'�,K���~�?\�aO���q"):p�DI!�"A��ͺ�<������l5��~p/ǉ0��e���w�ı,K�����O"X�%�{�wjr%�bX��w8�D�,K���q9�L��O����yIam-��w�,K�����Kı=�~�q<�bX�%��f�r%�bX��{��y����ow���r��#c���Ȗ%�b{����yı,K�����Kı/�����%�bX��gv��{��7��￷ߪ�U�����%�bX���w�,Kľ{��Ȗ%�b^�;�9ı,Os߻�O"X�%��}���7m6�ٗL�n�r%�bX��{��yı,K��v�"X�%��{�s��Kı/oN�'"X�%�P���T���A=���䛲a�,3a6JsGN;F���ŹQn:;�gˬe�<�m�v��������2 m�Wi�f�(�j�=�'5�OP-�(���<�=t6�sqt]Z��&�l�n��`eJ���@���Ͱu�s�.͍��;�j nv�P��8�>��]��sFyN�]��u�5�[�|��#�xolh.NL�풌��rK]�Zt�� �[u�OF���{����������B�^����-�"$[�m�g�[ƚ��<o:�c]]��^Nv�q�L��'bX�%������Kı=�����%�bX���w��DȖ%�}�����%�bX�v�'�s3Hn�.n�ND�,K�~�O"X�%�~�;���bX�%�wx�D�,K����i��(bf/���r'l-�"�����%�bX����q9ı,K�~��<�bX�%��ݩȖ%�b}����ቘ����O&��N�2��,��'"X�)"g���x�D�,K��~ڜ�bX�'���8�D�,�#2&v�?n'"X�%�{�L���K��n훹swx�D�,K�����Kİ�������Kı/o���r%�bX�����yı,H���{�Y�r�e�ەu�`��W�e��մ3���3Ց�gK����r��'c��� �'���NA${~>�D$}�ڜ�ؖ%�~�wjr%�bX�����+���i%v]��131?�N�'!T| =�&>����K����'�,Kľ��ڜ�bX�'����'�?S"X����l�nZm۳.�t���Kı/���x�D�,K�����Kı>�~�q<�bX�%����r%�bX���2�'���Ғ�7x�D�,K�����Kı>�~�q<�bX�%����r%�bX�����yı,O~�s2gl���n7v�"X�%��{�s��Kİ��;�Ȗ%�b_w��<�bX�%��ݩȖ%�bzg������_-��tXmbݽz�Z����eϷ�Ŝk�:ڍ�VF������?����X�%�{��,Kľ{��Ȗ%�b_��ڜ�bX�'����'�L��L��y7'�v1��	dV�Z%�bX��{��yı,K�s�S�,K��=����%�bX��ӻ����wy=���}��ʯ����jJ���Kı/���jr%�bX��w8�D��zQ�#(EN/�zL ��W>�e ��{T�X+!Qx����M��B��1<ֆ�M�c�����X�&�%�<B`��<@$}	��<|8�	��x�Q$D!�H"�AB��0�>u�P�dH� 7P�B��"��a�C"	z*n�Qb���H$X�A�H�	ea`H��E�� XԁY�BH�J$�(����$��d�01b$��Be I(�����ҩ`Dlx�jE��� �B�?*�0����.��������:����	��Q��A@��v'�/�ӛ�Ȗ%�b_�����%�bY��vE�I+c��"n[1i����1!"}�w�q<�bX�%��?n'"X�%�|���'�,KĿ_����w���{���~�:ET��~ou�bX��ӻ�Ȗ%�a����߷��Kı/on'"X�%��{�sqp��L�ş/zi�S��"�GR�k���.��1��$GBp=x�1prJ��07c�v�vf�t˦�'"X�%�|���'�,KĿ_����bX�'����'�,Kľޝ�ND�,K���R,�4�	-�\1313���0�Kı=�~�q<�bX�%����r%�bX��{��y��7bX��$'�IP��[1i�����w;��8�D�,K�zwq9ı,K���<�bX�%�����Kĳ{�r'<B�RqPr���130�ޝ�ND�,K��{�O"X�%�~�wq9İ>�"H�ߔ����b{����yı,z]���م۲���7q9ı,K���<�bX�ȩ�����%�bX�g���O"X�%�}�;���bX�%�������X�&v�N� ��F�;E<:��P=�ݴ�u���+hA�V�-%Z����Kı/���'"X�%��{�s��Kı/��w�,Kľw����131wθy�J��u����ND�,K�����~�L�b_����r%�bX�����O"X�%�~�wq9ı,N��;��ې��������'�,Kľޝ�ND�,K�߻�O"X�%�~�wq9ı,O�ﻜO"X�%����i�3m�e�w�,Kľ}��Ȗ%�b_���ND�,K����Ȗ%���
]�����q9ı,O����N֚n��.��������0�Kı=Ͼ�q<�bX�%���q9ı,K����<�bX�'�*AD��F����&c�mݕ˖g\s��vv���z�]��v�V�t�y�bn��gk0��Z^݆3�d���^9�+i�m� �u&�z�#:�5n&ؙ��h��*Jl�fʝ��V�7�RqV���4]v����
ݧ�%��79�3N�k@f��d�n��K�S��l���:�\��
�;-�/GgR�q��z�b�*�Z�Y�I��� A+�tv8�1Rw{��/�xqp�P�*�#r� ����8����u��lP �����k�rS��V!��77q?D�,K����q<�bX�%���q9ı,K����<�bX�%�����Kı=������7sB�fnq<�bX�%���q9�F9"X�����O"X�%��;���"X�%��}�s��Kı>�&�wH�Q�Yj���������z�.	bX�'s��T�K�A!�2'����'�,KĿ��Ȗ%�b_�����YJ�%W�w���oq��s��T�Kı=Ͼ�q<�bX�%����r%�`	2&{�߷��KǍ���뿥�1H��{�oq��K����Ȗ%�b^ߺn'"X�%�|���'�,K��}�ʜ�b]�7����ϣ��N��Q2ꎚ���'�xSu�J�j6����瀉M<�R��C�\���ۻ���%�bX��Ȗ%�b_>�w��Kı;�gr�"X�%��}�s��Kı>���p��Mٛe�34�ND�,K��{�O!�*I���B�tW������L�b{��S�,K��}����%�bX��Ȗ%�b}ޝ2��َQ
�[��bf&bf/O��Ŧ&%�b{�}��yı,K��M��Kı/�w���%�bX�O�fd��n]!�fK��9ı,OsﻜO"X�%�{{ٸ��bX�%���x�D�,K��w*r%�bX���\��r��hf�&f�Ȗ%�b^��n'"X�%���{�߷��Kı?gs�T�Kı=Ͼ�q<�bX�'�|~�s���Oh�uv�ƥ�����vζ#��l�����]<�k���Y���Ȗ%�b_{���<�bX�'s��T�Kı=Ͼ�q<�bX�%��f����oq�����*�xZ�R���Kı;�gr�"X�%��}�s��Kı/o{7�,Kľ}��=ߛ��Os���}������ܩȖ%�b}����yı,K�����K�0S�?`#⡢�D�%��>�'�,K���g�Ȗ%�f.��z�VJ[evٸ�bf&%�{{ٸ��bX�%���x�D�,K��w*r%�bX���w8�D�.����nh:��kO����bX�ϻ��yı,N��ܩȖ%�b{�}��yı,K�����K7�����c���=�h.�\�ڎ�(ɚG@#!�֞�ɇxÚ��tc5�skë́6�7x�D�,K��w*r%�bX�g�w8�D�,K���q9ı,K�{��yı,O��32gi7.��3%�ʜ�bX�'����'�,KĽ�t�ND�,K���x�D�,K��n�"X�%�����.w.[��I����%�bX����'"X�%�|�{�O"X�%����S�,K��>����%�bX�N�s3�e���n����ND�,K���x�D�,K��n�"X�%��}�s��K��C� ���ǂ� �=�w���7���{��??���{MQ(��<�bX�s��ND�,K���������%�bX�����ND�,K����\1313��ߎk,�W%v��T���<M�է�'�y�ՔTI���y�@��i��c�]Yy�ߛ�oq���w;����%�bX����'"X�%�|�{�O"X�%����S�,K�����p��R�+����131^߻���bX�%���<�bX�s��ND�,K����Ȗ%�b|�>ܼ�u�8�Z}�7���{��<�{�O"X�%����S�,2&D�w����Kı/��ۉȖ%�f/��jp�vી廋�&bf&'��n�"X�%��}�s��Kı/o��ND�,�L�����x�D�,x�����ҷn�hb�|��{����>����%�bXG?^��O"X�%�}����<�bX�s��ND�,K�'@	�-�n_)���m�.۴���l��w�9;����sm��n�;^crp���,��O����v|���Tl�5m;��ᖴ/��(�;�gc����M�Y��<��W3�W9kq�jڞ�������Y7D�u�B�Y���em��[*i�k��\������.�k��gn ��C�v�n�X�mͮ��tg��W����6H=�nw-������¢| ��!�ɻ�n��r�ݓOO<v��~��x����YtG �d�#�fγv�\(�2#G���=�w���{�K����r%�bX�����yı,�ݺ�)<��,K��gȖ{��7�������̖�����oq�X�%�wx�D�,K��n�"X�%��{�s��Kı/o��ND��7����ȯ���TJU|�~oq�X�s��ND�,K����Ȗ?�a�2%�{�q9ı,K�߿oȖ%�`����.l�ɦ��2��ND�,K����Ȗ%�b^߻���bX�%���x�D�,K��n�LL��L��W�BB�"�Kl�[5<�bX�%����Ȗ%�a�G=����{ı,���S�,K��=����bf&bfg~^�JK#�X��^���3�箹�m�
�{vV�쏞]�N�Ł�Lݴݙ�]33w�,Kľ{��Ȗ%�`�>���Kı=�~�q<�bX�%����Ȗ%�b{ޝ&L�Keȫ�%���&bf&b�zLZ!��� $�H��Mv���K����<�bX�%����Ȗ%�b_~����%�bX?}��L�734���7719ı,K����<�bX�%����Ȗ%�b_�����%�bX���s�,K��߹s��e���\��'�,KĽ���r%�bX����<�bX�'r���Ȗ%�b{�����%�bX�N�s3�f��a�3s7q9ı,K���<�bX�'r���Ȗ%�b{����yı,K���'"X�%�����?]ɻ�k��MHU�y�N����n��-�Yv���+�����Z�鬊��K4ĥW�����%�be���ND�,K����Ȗ%�b^��q9ı,K���<�oq���{�<0a�VT}�7�ı,Os߻�O"X�%�{{���Kı/�����%�bX����'"313}}<�WkCR���ٸ�abX�%��w�,Kľ{��Ȗ>& �Mz �"�y��}�19ı,Os���q<�bX�߯����VcNZ�w��7��,K���<�bX�'r���Ȗ%�b{����yİ?��3���q9�f&b����78R�r*�In�ቘ�K�{���Kı=�~�q<�bX�%��w�,Kľ{��Ȗ%��{����g��x�;;uv��]»6]I�����蹰���Eas�H��771<�bX�'����'�,KĽ�wjr%�bX�ϻ��yĦ&b�~�����L��]�Ȥ��6���Ȗ%�b^�;�9�#�2%�}����yı,O��?eND�,K����Ȗ%�b}:M���Zꢴ��^-1313�}븹ı,N�s�S�,2&D�>���yı,K��~ڜ�bX�%�ߌ���.fm���̻��O"X�~X����S�,K��>���yı,K��v�"X��5?����D����x�D�,K�?ٸYZnJI�<Zbf&bf.��鸹ı,N���9ı,K���<�bX�'s�ܩȖ%�bx{>�^��c&j������+��l]v+�1WO���u�¥���/K� ����"X�%����"X�%�|���'�,K��w;�?�?��6%�bw;�������{��7��������]3�jS�,Kľ{��Ȗ%�bw;�ʜ�bX�'����'�,K���y��131{�/s�-�"���/"X�%�ܽ�br%�bX��w8�D�,K���'"X�%�|���'�&bf&,��n(y�:���ɋD�,�?�lN󿿳��Kı?���19ı,K���<�bX�"~���LZbf&bf/���E'�k�q@r�'�,K���y�Ȗ%�a ����x$�H���M�H'��~�	 �'�(*���(*���E�TEh��+������
���E�DO�� B
�0����"(
�1� �"("�0* �� �"�0V"�0��b(� ���D
�1Q��@"(  �@��Q_��Q_�E

��PU�E�PU��ATW��Q_�E�PU��PU�PU�ъ
�2����I� �������9�>�=�                  @S�I()  �p ��@ B��� �*� � !B� �HP DUQT� B��"�`  �A@  )@�@>�'v�6�f���ٽ��W� T�4֘��15@g�ס� ��@uLC� {��8��` =N�T����t�j � �� g`�ץS�iN�Mt    �
(QT � :    �     �       T��hU �g�&T��T���RΔ3���Y���3Je��� Δ��K�nyj�j�Wp y�$ɥ9cٻ��SvqU�  w� �)!,�@�Žj�&Ebj��5.��R��+6�jwq*ť� c�g�����׀�w.mJ�i.����罕�4��u�ڥ���Hd�3i�,��6U8�   AA (C@�U�2ʦl��j�����sVm+��eX J���6�ɮ�.�Y����O=*��e9e֮&�gJ�� w
d±ڹ����R�    =
Q  2 �fݱ9e�\l�dа �7��qg�����x���ӆ���K&� .,:�X�s�)Nz�'��,���WNAՀFꕉݓ��z��vַ�����a4��M0?I�6Ԥ�A�� <z�T���A�F=��J{(�G�  E?Е6�%)P  !HI��"�@Fjz	��/������������MBR�r���=��m�g�����L�_�� ���@AS��"�������QEaU;������ '#�������a�a��e�q�F$6�
_���	?#�,R �pN�� ��b'�<R��.	��`X�H1�F:#F&�1Г	N:����i�1��0�����Kd~'n�TB�7of�4�a�sNЌA8Y�[,�m�+a�+y�v�N Fs���m	O���/ٯc�l���[����Z��C��D��Q���������z�J~�����sXi��kEa���TG9k���;X32�q�x��/1#_��N���A�2�df�����.V���U�0� �4m�����k�c�E�9�1TK�Bc�����di]�<�3 "�#<�1���Rl8������6h�ӧfy��fh���f���8���F�|<����Ѿb� @Kx
\R�4�e׋��N��|M��0�1�)%�Z�Y�����(<����'8�c��6(g	�ӯ4h�)��Z��4,�@�K?����Bc��A���nMh��k���B4���Y��,�f�5zF�0�,cp6Cj�1��&�3[wZ��<ќ����0�#0�V�3L���z�l�х��x���c	��I��t]?��uD8�8�L!.����Ft������0bhL�!��X��.�a��%�FV��A�A��X��_�ӿ�u񃆝�32�N$gM���,�~�0�Zփ���k���'pd�H���k���ߵ�ލ��k�~�y�Q����FFO5�\0ňЃm3O��B[,=���^yg��4�&�`Z�3�bXi��xqߏ��~6`0c&0,mo�kџ]$&:CHFa����	H"k�2}ۆ��zx0b�v�ņ���I����I����0��c	<��q4���۳F��[0�sQ��f�L)+�H�ߗ4~�Á�!��������0�rK�������bH�[��s�k��FC�0C���z�cx������^���ր�R�w��y��9��M�$���4/��S򮗨�4@ˁ�g5ae����$0tmc@`N����6$�	�N���A��4n��A��i�L4m���<s��k��CS�:N&���6 A��&�U����+͖����e����,�`�i�4b��)n�uT#��+t7���/�嘆�*l�*��ϭ:+(>ˢ��>/�c�]W�V��8G�r�e��s\��Z��� �6:YG �}A�� �4l�������gxDE��d�i�0#Ae�ý��dp�&4�<'5��?�~�F4���=<,��y8j�Cf���Di3�#��PN/�ck���8ɮjc�јLlN��
hv�@��Hik �& J�iP�H�)�CbI2� T��!ЎՅ%��
B�XP�]�F\*�`����+� ��% �	R�FsSF����R�]��$0Hɬ�г'Q�2��$�pѰ��Î���kU����I��k����14�j3v�|lCF�$i��F��ڟ�' Ѱ��$�d�[����i�d`�ٶ����	 ?RF:9��ӕ��8���>8ߏ�w��A$ᠳY����Ka�{�0Ŝ`�-n��v�a8�����bFF�X�n�I�j8��Z�Ũgg�A��W�m'�ךբ�f�|M\˘1�Vh6S	�LR�+\9�qݨ������1a-o\��$k�*3Fx������D��	��ͧg�Բ����5�l���x�u��i�qᎫMAoY���D��xkÆ�\����$I�~j�Y~6ΰ�L�É�6x�-j��<c6����Da�f��Ѥ�Ʃ��J����%����2� �@�a8���0�m#S���GS2"ދ�9��A�L'P4�{(X6:d�
 ����ˉ@�N<0� �OWc�,����Isz8��c��6k2w�,f�r5i�戍�D�h#Fݬf�3[ۄSY������X#A3�����0���3�X���=ƧIA
lM�hd�Jc8����}����ONy���N�~r��Z�ekp��Qy{<3���xI�X��%F��Fa�<�r���9�|8x��ddae�����no������*����2x�|��c����:6s(	H*̠����2�0l�,�
�� ��� rLӓ�$$��p��6)xm����˙�ц�2$��9��i����<7���5�t���3���X~%$����ߗ��0yh���s\6x9�^%�e������}R��(04ƍ���S���$�Ն��\��|0�'���a�����A����oM�����Fa�$��̳ �4Z1m^W9���k��e���Q8������S��f��k��g_}��?AI$!&�< 1t��H�����0I0@B���w��y���o^{�g�N���~ʳ3�Y��XH�����O�a����<󆹾z��uh'!�bG���\��$�z:7<��9��2-���y~#D4𘖁1�	d0'��	�H���Q�󑆙M�8QigKQDi�3�kXo+���F3leM�9�L��2�l��2L�f�N+���iv�˃��a8�c����b�O�t8eXa�	1�y:ՆԐ�*�r����S4�գ�d���U�0v	k�	..������wf�h`�PkV��k7j�@B�j��BGA:�t��~����ػ����o���s���_c�bu���U}��>��뵔�}��e�_/�U���\��,�U��zs~��L*V7�e.}���G����o
��ܾ�A<)]Њ�����}�N���>�fP��
�ee�0���e��,E]'��~����˿f:3*���՝��Y�U���?y�fkMd[��������y9�x��>��|/���˾,(���e�8��L����w]�Q/�T
�(�UA�pv3O���>Ŧ���w�n>|��r��1|��tyU�m���qU�t/���.��2��N�窓�Q�+��J�e��f�������o�[����UR����0�Y����R勗k�J�S���ym�Б��y��Ee+�����6$����o��� ���˖�{���x����aY�l�Öh�Ѳ76��f&�|±�R8�>�B�Z�._p�����pUE/�t�}���A���w�tX�ʾ�UoF�ב�-F�,�dFg5������w�۫�vهn��+��UWϴs2��w��2��e1����|���v�}��߬\�{T<�Z��B�>����e,Ͼǆ;�_.輤RUu�]"��s�'}��N��Β���5Z��I�؄�}�>|O�q���5�7���vxs�ro7�7�Y�/��������uϾ�)u��LϺ��w�]S����w)�_՝�Ms*�|`�k̸Y�[��FQ����\�:G3���7��������K8a$��Y�+�f��-�Xh#,L�cj�����0ՙ�����/��[����c�Nj�i<O�..��ߎ��xlh|XMZ��d��ia��d��Hf�^o)'�ČXi7̌�`�ٴ����|L�z���RY���9���afZ��DN����6᭾Ta�g���$�t&ݶRY;QS���݉x͕��,���7��o���4l�_�[�h<ӆ��)��$c�$��~��Jl8l<a���C=?�ɡ�n	������N������o�  ۶� ��  l �� p     H  Fz�9zi:���t]v�H[-Qd�&��m���VA;8��Uq���\��W��0/�.̓�'���6�63��N�D���w����!f19��8;d;�f�}S����n�S�ѵ,uD�G;Qu�<���m)>W)n֮Z��z�I�I����_��J���� �<t�$�H�.��[��U��ux�3�g�S�����v�p=���q�D󴝪�\��\v��๪���h��c�jl�5��Tb�"�$���,����+Ì��D��yr��UEm�U���;��.%�j�tIŔd��R�9�	˦�.���ic3y'������y�n=��k�f����4������m����ݵ��$q�s��=.nҬ27:4�5;Kog�,Y�[�\�!˃X�k��q�*��b4Kb1q�۬��H�l�χqE�|��P�nX������!y�6�{iXM=��Ӡ@���l�nY�Qv����f3�l����Euvv�Y,��� -�Mn[\ �-� � m�p[C�[E)�86�    @p-���bD�� t�vճ����[��`$|H n� @  -���!�m&�}v� m �il��  �   ��h��  �l��� ��   ݰ6�g   9 �� �m&m�� u�I���$[Kh<�n�-��kvݜ� :BN��t�iz�U2��p�]�]x���3��hl��(.�-UUm*�d�v����W��ݴ� �,�N.B5f�n&�G6�@<�2�6�ۉ`6�Pm.+mՒ��d��4�����h �
@j�N
�4��������j��]Um���UUԻ,\aَ��y�ɒtu�+���6����;�c�
t��@U� ]5�p8��u"CR�;���W.ݵ��ږ�3̨+v�%�-�酴v�	6�W�̰Ͷ�[RH8�9V���Hj�]�V��rm��l�� �[�Ā7m��@-�@��r H  ��l�ְ��]� �[%�mHkX  6�e� l8 [R7m�/P��mj��K�g@�J�-����@pm�Xn$6�^Ԛ5�!����8��Wf�Ci�V���  H��6��[e�-�i0��  �-��U�[F�ۀ 5�6�m��m ��m���mrI6�` b�4�6���6�m��  �q�mK**���_@_.�L�Bmp h��h���e��n�ćvZ��Pm�8�J�*��
�c�%��9��i��	��vSmKR��ڪ�����V�j�r,�1�Z�S� ���_��c�#�ҙA�tUUʠQѦ��F԰K�GD�Z*٪A�Ilb���T���s�J��m�AhܭV� 8[x!&�6��6ؽ� ���k#m��F��P	6�m*t� -�4�MY�"�ku2�v� �m ��ٰ�� 5�<�UUW)l�&��@A�R���&@*��ZtHR�P �jj�q����Wf�j�%�@�mH�^/��)a��d�5�I�  �[p$�m&��=`$�d���[��]2�UA@r�� ���d��5��j@��6�6ٶm�Ͷ	�@� %� k6��`�H[Jݨ%��� 2f�I�P>��h�@Z��� @�_���l #�[@��6�j��G@��ë'g��:�m �[��m[pn�yV�^vN��Z����5h�v���U+/l N�F�e�`���A�cUlYd����e�m��,�濟}����pIT�{;l��pb���=f����ӷm�V^][UVʽ�d0�C�`�6�a��������*smE�鱐�� [M��}�|�kP"!�UUQԷ	�l+;��(cp,��v����ֶ�At��Ț>8�8����  �<`m�u�-7m��l��6�[q�6��d�]��mm #E�]z���V��k�ٴ� ��:�`m�]ͺ� ��6Z�.�dٶZt�Հ�`8 �8 mI��u\z ��H d �mXkI6p h  մ��C�UR�*0"ƶ�ݬ-� m����*֠-�e{�i]#C�m���p@ֱ�i�#]� 8m�` m  $[@p 6�@ � ��ٶp�  [m�m��v� �`  m�E� m���7�Z�$ [@m� gEm��kz��xm�6�gl���%�Q���C��l� [F۷d �8 6� �-� 6�[�&հ��m��h               6� ��Hm�$J��7U!�0�V� (	c���&�Z���UM��`  [&���l 
��t��K{jÜ[%��m�mp -�8� -����ki����t�5P[@ �m� p� ��mm�@ �  gۻl  o*����>�1���W� �Vh  �6ۀom�ݶ��@	 -� ��)m6��v�[y���4ڀ   s���n�L�!����  �� [@;6�i�m   	l�[@  �p 8�l ��ċh -�l��ې  �m٬CT�i0  l$��  �`�   H �� �`  �          H��6��4���8�  ���)lHŵ:�
l5�VhH����U��4͝�[$Yr�M�n m���l�I����˵@*���eZ:�nݚ�`m�j@$q,� �d�ݶp    �v�m 6ٲ��i�� -���ݴ�6 m@�  mf\���!   �    �M�pl@m�H�ܫ�T�]T�+���%`1����'"�Z �`�  �Yyol ��lݰ�� [�� z��iF� 6���\����*d�<r��*�Tv��  ��i66�`q��᪵��D��i�\I ��Lm�$H-�  �  l�`��    [@�  ���   6�    �m$    ?}�����        �  `�  �  8�H�*��vGr�UJ�Ύ��`*�y��-����: ��ҏlΐi`��I]�v�8 ��p �  m��� �`�@ $[UGQY �j��@;Al���$	K� r�n�@UQ.-��g�{ kX��ֵ� ��R�l��JK[uv�,Ɂ�� "ޠ����m�( ��m��m H@@J��[�Yw`9��U�`�b@ ���t�Kp%x����c@�WQh��e�D��3X`�k��p ���     [@�   � �  [@ lH�m�[W�M�A�v��m� �/��_Uۄ@���;Q]k���i��@�����Zж� m|   m�6��e�    9{�݀%�6Ͱ��S[���,��` *���T�d�i��p.ݰoӀ�L�,��~>�}�� H$4n� @[A߉g�|�{d�ɶ�M���Mn�� h       �`       �     hM��ٶicHm�n�������4�kXR��n�2ӱ!u��l8-H��n-���&�� �I��`�0	�QQ89bZ��n�m�i�[% m�^��k���AKI3 6�T����UHS4(�j����M�td�N�j��}q9vȫ�V��\�֚օ� ��� �&���@W�I�+�*Ԗ��9:$�$�6��T�W�u�'n����-�-U[� kn�m�v�ʥ�V�Q]��*���C���*+e�`X�6�Ie$nAmv�M^�Bh�j\�.�U�)<���$Ia��f��M�m �l��6Ͱ���k�����Tp@J�������$�@m�9��*�r��[F�V��!�&�$���d��l^�{&�N�e6z��x�Dp��ut�t��6�m���    $H/�a��;m�8mԘ  k�  $�c��m�m� %�`iX 6�H 7Z�h �X��  �ۜC�J�2�^�D�S�*[#]��Q��v*�j�ӽ��m[�M' ��'!V�^�5��E�&�Uz�z�����ݹ��vZ��{��(*qQ�U���<u�?�..�*����� p qFTF>�(��x��@���'!4".��R:h� �� z��<�?����'QM?�%����F$@�N����pJ
/�z0��< P��a!0����V0�(�`{�����CC��t�� pҠ����OEQ=@ �leBnM tC�)���x��?�w���Sc�D0dT�W�ߑ@��6�#��7�����C��v�"!�M.�<�`��|v�����Q}�Y����!ꎄ䜪��ʊ(j&�&X��[,�h
J"J� �a��#,��%��êy�����D��80���v�J�����U"UA�<@ځ�"�����P
H`&�*�,�$~�߳V���Y��-�I�[�4�H��8�Ls��]s�C��i��ca�]��rO������	�/8�x�q�F��nd�z͵�-�s8Z��ճ�61Xŝ.U݇'\vӴ[��#t�gKp���rfe��ͧKm��PR�4Z�����݇�#Aԁ�5Jy�R�*�K+�R�8[��4eunm�J[���p�["4�2f�ۗgl�����'m���\��OLמm�]�m �Z.,�F3��me�@N5�ŕ^u[�5=g��w���u0p�!V�5l�������V�Ҕ�c�;a'vq�m��)�iy@Uͭ���Om�s�Lyk�v6,���um���	6ȼԼgI֓�e��6lӪ^��2M����ڎɶLqMQ�Cq�N��j�PE�Dk������ur�&�2sźSѢ��X۶P��m���Zv*�Xx�v��AY6�N��jF#����vN�vpT��g�
�w<��P)Y^'FN�ヵ�CZ��rһp7m���@ !���;�ʅ t3֋�������i��{]�  
�zA`��a�C��;I��'6���m]��m��e�<`�
K)M�t�[-I��n��HM\�+u�v�V6��um�VԫJ�@UTp����Q�k]�gu!�vn��$M] ��J�;It���+UVU�$K�Q|�rԷ	Ym�yv�w�IӆT��];��R�Skj���m�� �U �
�
���9j�jU�`�b@"Xΐ�4�i�VM�ʜ(
\�����u*Qv�{c���I IU�띰�t�b��m�7sfv��J��&5�'�/hu���B$ӖJ�n�m1�H{�%-�Oe� ��B8��nz� �rg��S\�E��ɷ8�r��Ͱ���I�!�2v�AE�CB�����ɜM/�<m�Y�,$���c�;�3���n.]m���HHrd5mĝ�&�=�ۡ��[�WZ�{��s��D�#,���� �
"6�"�|C^�Q�M� 	��wV��7��sY�v�m&8�(Η�lY�+�cR ��	l�մ�A;����۴�<��f|����#f{td�9��	��晹�q��w�MB�[/�T�gN(+L�e��TO
�-5�ڸFܙ�=l)��wl�mM�1�]����MuI����ûX���.q7`�	�M�m�rp��a��J�W[u�z���oq��iT�:��{�}� }�<8�ð�ϲ8<dݗ&d9�Gy۞PcX��7����B,�9^��� ߷_�r�ʪ��5�{ҟ���v�[m�v��we��r���Us�����<��ՠU�W�~������Qae���o��	�2�-�x[���IBh��Ct݌�o �و�"ݗ�E�/��N����(l��mU�e�� �d�)��l� �\������pw�\�=^�p�	�)���[:���t��{sn��V��U&s-���6� $��	�e`k�`l���F�j�Zb��Hv�6L�����"����*�����|�mzo,�9�d�F@�y.�u�Nܔ��K�	�6L��$$d�i��91hr׿ff$��@��w4��o2U$mH6�n= ����4��W-z}�U(�25���Hx�v3s�\kl����81u��`��=��@6����*Ӥ�&�������	ے����٠��c�0�$d�@�rR�"�/ &�x6G��n�$8�i"B'1hrנ��E��*��� H��3
�J�+4I��/Nq��R��e`��E�Di%��c��؛w��<l�X�ڋ ��� 紱271Ȱ�	I�^[��M����e�� �U]�^�Ry��0��i������[nz��w�X�T���mؚT���4t�N^�;�!�~�,-��l� �&V;�$��б���W-{��<� ��f����h��Z��Td����(ۏ@/-�廚��W-z��w���S)�&29?���h���Ws��\�!�&�(�(��>Us�^�r����c�	岄բ���I[�m�K �d� �#�&ɕ�T��5r(ہ�@nG�dH�T\�mۂ��t������lv��G6i)�����XcV�`l��dx�2�UUʯ�v����S�nx��c�RG���l�Xے��x� ݄j���5��H�M�����ŠU�^�^[4i���LƤm"!�&�6䥀E�/ &��vG�}�ꍱ�!�92'�*�+��f�}����ޘ<�� {z{hן�'<d<���m��>�����Ƹ���9	�ظ>�H�C�^�<:�n�F ��ȩ�Ӻ���*mun����M�E�v6�m�n��R70��ڶݺ�b�	8V��\q�5�T;aeS�9Ł�T���[����Rٗ�zH�2%$�˅�.jgٛtu�c�z�%� ���!�v�}{s�<�lqz�لwq���_g����q�v���@ڜcr[����}��`ۜ�=>��6�ɶ(Qݺ�WQ:���H�?�{���n�������{ݥ.��w�)JN����R��~��┥'����սY�l�f�l�z���JR������'}�N��R��~�u�)J��v<��/{�fo-j��l޷nַ�)JRw���%)N���\R�����c�JR��|R���n�.���X;����9QvK┥w�JR�}��┥'wl���9A�TF�]�&4!1ݫ�yĥ({����R��}�)JRw�u���)����)?�}����j�k6*ƺ�^p�糮�^�Tn��&��71g���7%%/���ɪ��̥)}�~��);�{����s��\R����ǒ����w5�f�xlټ�e��{┥'}�{`�4"���!�L���qJR����J9D�s��+��ݗc�����z��JR����qJR����JR�{�w�)JN�<��=��}�:���H�?{ݷ���n�w�?n��JS���k�R����w0y)J{���(9�W�v+�ˤ��ۮ|)Jw>��qJR�����ك�)����)J���y)Jy�s�3y�f�s����"3�(�b���Iƌ���=��AC݊�Z�� \V�^!������'}�]�JR����\R����ǒ������)?W�����kf�z��o0y)J{����9)C�~�c�JS�}ߵ�)JN�<��r�Iv����4ݤ��9A�PW&��y)Jy�����z6�!�U�lI��\�JR���{�s��+M��c��tӵt��\Ü)O3��\R���빃�JS���u�)J���y)Jw�滬ٸ͛33Y�޷�)JRw�u���)�{�u�)J���y)Jy��u�)J���~R�Y�����UWN��ml��͵�pZ{=�nwkS�	K��w渵�C�JS����R�=����R��;��R�����������o��M��M��Wv��9A�PW&��s���w���);{�m%)Os�{�)�+�w��;ۦ�tm�>9�p��}���)I��{hy)J{���┥}�v<��/;�t��k5��l޴f�[���@�$��~�<��;���qJR����JPp_D	[�K��#�;��R�����ov��Uou����R��=�u�)J���y)J~���┥'g�և�������ߝ���f��z�k\��7X�8z˄��:�\��GU��f�u���^$��z���)JP���c�JS��{�)JRw�{�hy)J{��u�)JOo{V���(�Mɞi�y�V׹��FrR���~և���s����7c�a�Ps�'/U��2��Е���\R����u��)�w���({���R��;��R��w�7kZ՛3fQ�[ݛ޴<��=���┥}��JR��{�qJR��������{���7�~��*����m�v��}�ǒ���_}���)I�s�kC�JS��{�)JRx����;���q�������A�S���S/q��@j�3 ����mڌ�\Ƭ�EӲ�T&"�� ��j�9�T�c�k�@(v�K�����9y�4�m�^G.�N���Q�c���۩ �m�ʅA���:]�����9N6�U�!�a:bU��#�b5Lu���ݬ�6ݺ�

C
��HӴ`�ɗc�����\�]��ݽ�HAL~���{�����_s������t并"�Jz�:2�`������IY����6l�k6[�oek[��)J������);��w0y)J{��u�)J��v<��/;�fo5�Y��7�����)JN��]�JR��{�qJR����JR��{�qJR����Y���f�+{��o0y)J{��u�)J���y!���N��}�)JR}�����s��j�M�6ݶ�9�r��6M�%)Os�)I�}�s����m{�y��{N4�[Lq��m����%)Os�)G�?w�C�)����)J���y)J~����	A���N�=�������0[$P���v{c�%�[��x��������	����)I�}�s������\R����ǒ���{��JR��{�v��Y�v��ѭ�Y��%)Os���	F�D�ԥw��y)J]���R����w0y)Jt��}�j޷�[�����ַ�)JP���c�JR�����)I��{hy)J{��u�)JO۾~bt��6��V�s㜠�(���)JRv���JR��{�qJR�l���9A�Q�۔�Wv6ӥwNշ�JR������R��Oa1����┥���%)K���┥'������r�.s��yݺ��
��lVpfۭ�W�\�Ad��ff�q�ݐ��{ݡ�)�w���({�{��){��|R���ｴ<��=�Xw�����F������)JP���c�JR����)I��{hy)Jw=�u��<��=�b��5<i6�rg�y��}�w�)JN���C�OCa��M2��DM�<S�`��������v� ~�W��[߮�[@��NStT$BA@S0CU`K�98��c��x�P��&Q⚿�"z���*���8A@�CT~��Ѱ;�%��+�1!�@����g��
�u�0px ��Q�=E������ :�����Os���)C߻�ǒx,9)�]w5�f�5������R��I���f����s���������_2F\��}�)JR{߾7fkY�s7kf���v%)Os��\R������c�){��o�R���{���`y�}������c뉲bNa��E���m�ֻ'`÷F�@�Jܩ%���R����~��淫zݛ��ַ��R�?����JR�}�w�)JN�;����s��\R��������6f��5�foek{��)J_w��?�g%)>�>���)�w��)J����R��;�t��5�ַ��ݻ5��JR������)��{�)JP���ǒ�����┥'�v���n��ؓt��s��E$�R���{ݏ%)K��w�(IFN�x �US�I��4<��<��k���Z�ovk[┥{�v<��$'��v��������ߜ�z�����D��F'�ص�i�Dٻm֜��f��Sh�\`�8��;�T޷��)w��|R���ｴ<��;�{�)JP���c�JS���5���5Z�fk-o[��);��`�R���8�)C�}�ǒ���{��JyA��vJ�&�]�NշJ��9A�����({���R����|R���&ܢ��9A�Wa��tջ�w��R�=�{��)w����)I��]!�)���┥'�����f�kV�oY��Z��>JR�����JR���C�JS���┥{��y)��������?������C��j��M�O.��.{C[���:u�.�v�3��;k��s��9|�r�w+�')t��a{"!�����S�פG9�V�ecl����������#�c��4��i�Wkm����g���g(={r-+�m�p���3��,��P[y�sʡ�; �Cם����GZ�mY�b7n]���և&?O��n��oC�}N:�=��-ʌ�ڞ[2�:헙�	�Ѹ ��Ѻo:+v�9���!e�e�����m�v��߾��<��;���┥{��y)J]����)?^罬م�6e��o7����s��\R����ǒ���{��JR��罰y)Jw=ý�m�l�խ���y�)J���y)J]����);�u�JR��]�qH����q�*�ӌ����L�O<����{��JR���]!�)��{�)JP���c�JS�{�k7��h��5�ַ��JR������)��{�)JP���c�JR�{��JR��sܿ1$��������s��:��nn�vyۛc�v9�^	|n�Z�.4c[!bm%)N�)C�{ݏ%)K�����'�����R���忳tջ�m[Y�Ps�ɲ:���**�jR����)JRy߾�%���س���(9]��~�:��J�I�-o{%)K�{���)I�{���C�x��>��p┥�{�ǒ���j���i�I���m�9A�Pr�˄<��;����)J���y)Jv<�(9�WM[:T+�HCcV����{�xqJR����JR�{��R���;����Ȩ|{���ū�G�]hj���;��f�ۃ	��Wv��u(v+�]Wc�oj1��Y[���JP�߾��R���{�)JRw�u���)���R�����u��ֳY�o"�k5��{%)K����)I�}�s���{��qJR����JR���5��[uke�֭f��)JRw�u���)����R�W� �K<Dp���ǒ�����������wi1 v�S��sr��;�wۊR�=����R���{�)O(9Sv�U�9�r��Ӊ�V�Lm�Z��)J���y)@|��}߷�)JO��}�<��;����)J=�����]�Er��l�!��g@�0���L��"�1!{v5to����\��#QZ��>JR����┥'}�]�JR����)J���y)Jy��tN�ۢ�4�HM��(9�Tݸ�sp�;�{�┥}�v<��.���R���s��l���������<��;���┥}�v<��.���R����w0y)Jw;��5����Zֶe�oz┥}�v<��.��w�)JN�<���v.o�w\\<��9J�+hI���M�&y��`)w�{�)JRw�u���)����R�=����R��?wV�5�wf��[�y`ڻZv���.�8�k{<���&k]�֮Tp�AM��n��vZ���(9Sw]�JR���)C�{ݏ%)�v<�(9�Ww`�wj����T�W�`�R��~�u�)J���y)J]���R�����!�)�oM�6o5��4j޷��o\R����ǒ�����|R���빃�JS����R��{���vlֵ�5o-�o{%)K�{���)I�}�s���s����?�����JR���όݭk{��fkv����)JN��]�%)N��{�)JP���c�JR��{�)JRz~����@�ш�=kn�v��ygه��ݢ�2N�9�L�LA�״��Y�@����X�7����GO�x������[����][`�^���mD�<:=�?d��>�v死u��Km�Kp�a�U�+$'���nS�,�8�UZ��75vи�+��g�ř(��;���u��M����̛3�s���=�F�A�t��ӡi���<q:	n�nŲ���m<ȭ��vMu���dm��I;%��l�+b�Eo�I��o{������~�y)J���y)J]��w���%);���y��`y�w�^�<$Ć�LCn=R����ǒ�����|R����u�`�R��~��┥'��{�j޵���ef�Y��c�JR��{�)JRw���y)Jw����)J���y)Jw�^泻�[ӭ���Y��R�'{�����{�{�R����ǒ������JR����5�a�37��7�5�`�R��u�s�R�=����R���{�)JRw��ޡ�)~�3�����V� �ܖ�q8��2��fM1��D�x�\���B�a\ƧH�e��)J���y)J]���);���P�R��u�s�R������ݼ���zٛ�̵��|��/�����	HU�UN>JRk}�z�����׽�)JP���c�JS��s�nֵ��ћսe����)I���z����{�{�R����ǒ������JR������U�F����޷�y)Jw����)J���y)J]���?�l��{��%)O��w���{��ֵl�{��R�=����R���{�)JRw��ޡ�)�����)?~�V��.�`���1xÛ�N�ji�`�e��]�9᳖.t�1rD��Ҙ�J�ǒ�'�Y���|R������C�JS�׽�)JP���c�JS����`�l�1��NM��<��/�����	���w�┥���%)JM�9�r��&�i���!:�*v&�JR���qJR����Hb���ʇ��������JR��{��'��}�'�m��-۷v�s��r{��y)J]���);���P�R*�s��Y�Ps��ퟟ�N�.�6ݖ���������|R����{�C�JS�׽�)JP���c�JS��{�"����ܑ�YIZ2�Nœ�mc� m8(Ĳ��9ӬL��t�#ad�o�R����w�y)Jw����)J���y)J]���({{��嬳[+[޳Y��JR�������}�ǒ����}�)JRw��ޡ����s��Z�M�7i+�!�k9�(~��ly)J]�{�)O�"������<��?����qJR��{k���BN�Ҷ�6�sr��TW){��9�%)>��oP�R��u���1B@���ף��?C��ly(y���'�q<j14�ӓ|��0<����P�R������┥���%)K���┥��FY�Y�[�n��{6�V�y���8䍫���.��
�#���w���┵*vM:�w������߳�R�=�{��)w��|�O�R�����ޡ�)�o���<���1��-��<��-�g�g�fb8��/�￷�)JO��oP�R���,�+�\�R\�+����Y�+m+t�vZ��>JR�����┥'w��<���Jk��┥����ǒ���{��oV��ލ����o{┿*�'ﯾ��R���}�qJR���ݏ%(>DR\����(}�߫7��-n�oy�[�ג��{��8�)GȨA���c�)}��o�R��v�v�����$`��ܢ�4��(��z��1��9�u��ŕY		aXR8AĴ)�V#��b2�SL��QqF�qeL%qd6�����R�0�$0�	@I2P�8F&�,D�(HA�0b�X��aWt�2������Cˑ�:It��?f�ɋ�BMx���'1L	�L%�(`!��BHL��b�=�����@<Pݽ��n��{�w�o���&mmJ�fjU����$e'۶�/\����RNԮy�Ql�d�<����<�9�9�z�ֲV��PV�D���N�����T��)�0m�9�e��q�@���a�V�c�,�o[��S��;pp@ 5UNRV��������VӻmT����|�&�Yj��1͜M�yD�2r%����pV��#m	Ų�ɝ��+8w��ù@��mq�Z��F�YG���0��h���ΐB�A�oX��X����&�+�3�\Y��k\�I��FG2qZ�j��}��eHIı6j�s�M;"\��]����-���ve�I�.Z6 d��F�S�iԼ[�;,��Q�r���xu�nr�ֱ.�0��M��� l�U����Y��-+�UN���9�-
b��^�O+��=k��AM����%Fp�@��J��;vM�N��d^��Ľ��jK[�V���J�u��A+r�H2�����m�C�x�ʀ�@ q�k���.ͺHz�6��$�+Y˳^�m�6� [v�;;H+��!�h$ܻPfe,Ѳ� x.���ž� ����l��m�n �g�Zs�0�a�\�Bڠ��]�&�շ@P��b�����K5i�\%x��6	0;�;R��k�PQm����61�Y�ӴR2�U��l���3��m��ԙ-m۞�H�*)����WbeiVmmUV��   �I�J��@�&73Hm�9\���6�̩�) ���nܸ���m�N9We*���Ү��\��Q�]�XK�knU��ͣ�eZ�]��ի��\�,HLP��{E�a�s�٢�j�^�&ۖ�]��kh�V���+��m�2W�s�" �p�l睳�X9�0A��g�t����
���v����p��\��d)�V.{�֗I����V@u�x7Mp*�[�u@VٵrK��ۉ�w-.�����~)�M�1t/�@}v�Aj<� �{����֭oYY���n�͓�n`n��j:�1"��]�� a���kkg0j9'[@4�h�b���휹�Km;�;1��)׎u��Df�c�kv[��M����W(���IhX��&ю	�&�{g�CZ�qOM��7՞P�������ms���ܺ�l Mm������ͱ�s��K��=n�\��+�sq��g��l��;k<���&�O���w��G�qƨ�箎��;J[:q���	
�ɍ���k�����r�]�w{��>�����Zvn�����)I���<��.����)<��v?*�y)J}���8�)C��>�_oYfo+[��Z�ly)J]�{�������R�����%)O��g�);���y'��J{������v�Ҳշ��9A����rR��u���hL���F��"��(J3�(J����ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�}����(J��"��(J3�(J��J��(L���(J�}����kv�5���Voo�(J��0J��(H��(J�����(J!(J��>�}�x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B}�~��(J��<���(J!(J��30J��(H��(J�Ͼ�����%	BP�	BP�%	��P�%	BD%	BP�	��P�%	B~���x%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP����}�5�z�kxo[޷��<�J��(H��(J���(J��"��(J3�(J����ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	J�%	Bg�}���J��(H��(J���(J��"��(J3�(J���߸�J��(O3�(J��J��(L���(J!(J��>�}�x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B{���Z�[�5����g+����tPC�tF�����m� ��6b���s`h��f�ݷ{��%	�`�%	BP�	BP�%	��P�%	BD%	BP�&}��o��(J��J��(L���(J!(J��30J��(O�]���(J��0J��(H��(J���(J��"��(J����P�%#BD%	BP�&f	BP�%	�%	BP��%	BP�'�����(J��(J��"��(J3�(J��J��(L����h��6o{�Y����(J��J��(L���(J!(J��30J��(O�]���(J��0Jx�~1��!�
�my	BP�	BP�%	�`�%	BP�	BP�%	�����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&}��o��(J��J��(?��Z�(J��"��(J3�(J�������VB��{��m��ݷ{��f	BP�%	�%	BP��%	BP�$BP�%	Bo��<�J��(H��(J���(J��"��(J3�(J����ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�}����(J��"��(J3�(J��J��(L���(J��~��(J��<���(J!(J��30J��(H��(J����~���ц�lս�y�P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'�����(J��(J��"��(J3�(J��J��(L��ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP����	BP�%	�`�%	BP�	BP�%	��P�%���$BP�%	Bs��<�J��(H��(J���(J��"��(J3�(J��9�L�LH�b���3s��<���0J��(H��(J���(J��"��(J>���P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'��ǂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	������(J��"��(J3�(J��J��(L���(J�{�	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�{�����vv�T�e)MHuA=�l[:yi��u���l4������/�Yg���լ���P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'��ǂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	������(J��"��(J3�(J��J��(L���(J�����(J��(J��"��(J3�(J��J��(L��ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP�w����Y��oFf[5k{x%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP�}���<��(J!(J��30J��(H��(J���(J��>�~��(J��<���(J!(J��30J��(H��(J�Ͼ�����%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	����J��(O3�(J��R!(J��5�%	BP�$BP�%	B{��9��5�{�oxk5�o{�y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	����8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP����~x%	BP�$BP�%	Bf`�%$���J��(J��`�%	BP������(J��0J��(J��(J3�(J��(J��>�}�x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'}�ݚ޳z�f��޷�(J��<���(J��(J���(J��(J��(L��ߞ	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	���pJ��(O3�(J��(J��30J��(J��(J�߳��(J��(J��30J��(J��(	T r~�~؃�(o�g��Z3f�����k{� � Ѓ�n�b A�@���>�}�<�J��(J��(J3�(J��(J��30J��(O�߹�(J��<���(J��(J���(J��(J��(L����<��(J��(J���(J��(J��(L���(J�]����]1ԗ9�/�N�v�����5�p[v��.¬���w<����e��7�z��(J��<���(J��(J���(J���~�	BR}����%	w��|���{��%	��=�o7���fj٫{��P�����9	B]���)<���y	Bw����>�����Ω�
3I��3L�<ý���%'��ݏ >X�O��~�	BW��{<�3��/<�M���<i�!�'������ly	B}���pJ���ݧ!(8��V��{�o�R���v�Mڶ�LT�����9�r���qJR��~�~��)J_}߷�)@�}	9�9A�Q�v]"����&����v�Wle��a�(t��GGf�l�v*K�.���9�>��o{��~��{�������JR����ג��{��9�r����*ح�m��wV��0�R�{�w�>D'%)?}߷�y)J}���qJR����JR�����ouoV�[���)JN��vJR���qJR����JR�{�w�)�s��!:Vn�SiZ�W0�(9ʓ^�8�)I�{ݏ%)K���┤r�˅sr���-lM4RuhV:coy�)JN���y)J]���);�u�y)Jw����)JM���R��/�tt�������UYl��EY��Y��n٭���u��-�"ծn�g����.�l������t7�53uvGwa��ݶ��.�kހ�n��I0�����G����6�FT�[����DF�M��ʹ.#�v\���4u�n�Q�tݷ=k���m�i]�h��s�����%ٮ�anEܖ�!��5�� �	:z���ZI �|�vK�s�oz{����V@�F���Gk��=lOK�F��kmų��]������pk��޳z�l{)J^w���JR���]����{�{��f.�)>��ly)�{��]��.�b��E�o9�r��6\+�s��I{W(	$� �c�;�֢j�Mp�j�l�$�� �L�yf�m��?S�*�q8�F㍵�I&`�$p�$�� �c�����nH��4�Y�[e4_*�-�t���,Q��71���8�H�5�[����:��n��9������dn��J@��94l��k�Z��[�4�qT)��q��$7Kز�&ɘ$� �3ԑ��<�4RuhV:cm���� �c�&�M�ʴ�\L��g���;#�&�m�X�3 ��j�[�Ġ�bM94�)�Z�V�yn���@��9�!Ha�D�M��6ܷVH{{$���b]ݗnE&<��GOK�t�-i�U̴�X��G�ʴ�w@-���?{E+�s�G$�@��wܮU$���=<�`^ŀ}�ʶ+N��j��x&ǀM�]r���8�o�h�w@��nx��<�#o �0	/b�&ɘ&ǀjݺ�10N1$7�ʴ�w@-���./x,tjH�� �L�PS{t.nXxZ��}v����[op������������B��m`d� �c�&��ʴ�G��`8��fǀI0	/b�$�3ܪ�G�#W}� dLLI�&���t�-|�@��0M� �ֵ�m���t�6ف�W���{ـlx¹\RGzk��ڴƒM'n�X�3 $��	�� ��,��s���{Νڻ)�W.+�/�+�ͻ;z����Suu�ƭC9�$�M�pLS$�9�s�{{4�)�Umz廠z�nx��R�;o �r,)��	�f I�繞g�bG��S�"M����� �&a�${���=/�XQlV�)6$�28��]�m��ڴ]�@=�8ՌI%<c�M� �٠N܋ ��Xݙ�]s��s��#�����n��t�[O3�p��͹���-S`^)ԛ期Y���h���vܧ.9v��6�h�ys�e{=����ѐ�s���n�HΕ1�m2�yV�SLr�G|u\6�"�cl��䖼+�bع'�8����j#`g�Ӣ^��ma,w].�L�n1�x�zy��g�����<���C8�`8�����s6�:�'Vzx����Sq�����w�}9s���^٭�۶%㗙,�aښ'Y�nylk��Lޝkur��<y���:�Dk�����>ؒ�,n��	6<�kQڶة�Wm:i��I{6L��s��<�Wޭ�rW24�8��#�E�{m� �c�7nE�I{�c�tՖ�8�x��yf��;V�k�Z���?+U���<L�M�v�����w@-�s3���;�3�ݙn�nŲS���
�6$��k��7L��'`��fm���Bcan5���~����l��lxۑ`E�Z�S�@��wı��@�v�����#�X�D�6��9��<mȰ���&ɘ�kWq��&Oliɠ^;V�U�z廠���Ecm��x��L�ŠUy^�6L�	6<mȰ�M�t�.��ⴸ�nP�V������泰]c<�ͮD�&5�E1���L�I1((��;{��	�6�_���A��z��By$q�`�m�@�v��k�/-��KB'�4,�,h�M��r��{�r�j�)Q��� ��JPC	����uXr0!�6��z᠃zWh~&@�$�����;F �v��`�0D hۚb<@�&�l̈���Ja��CQ�+�@�c� ڀ= #�Q�E��~�S������C�D^��fî�*���pW�����*�~���=\�S�)$i��k�	�< �G�M�QH���%c�-�x6G�lx�ᇩ//O?m����ߠ��-A]�b񗛞Λ�i+�`�m���y}W��Zy��k8�S���N7&�q.��h��Z^���٠[�"n�")��94�j�"엀dx7c�>�Z�����(�p�*�נ�4�y���@�{:h�>+��H�!�'#�mx7c�$�er��D��x��;��Cf���~ ��h{k��f���V�d��#"��3�\	�jp&^�ꗶ���McU��0��t�F�Fڃ��KG&�x�Z^��l� &�xV��'J�I��v��.�x6G�v<mȰ	-lQ�M2c���@/-��hrנ�j�!Li6�q��l� �r,-��l� ���v8�a `,jI�^;V�U��}�wʮ���*|�\�P��oύ��mѷ%�Z2'n�-�����wg��K��{ N,���ӝB�.Jb��SŪ,����Ț�z86��!N����mI�v�:�:nQ]���ݫ���{t�ՔV�$�ر�4�
n�*j��uT��2vYgz7j�9�U]ine��u��c�vWu�F���3d�:�m���t��{���!���ZϮ���˴����|s�͹��74�q$Ҫ�穀���O`���\8�4��5�	F��f��N/@��:��٠�4�j�?z>+��D?���� I#�$�RK�7���n	$� )$����@��h[^�[l�?*Z6Lhp�I&�$p�"�^��Iջq
ba�F��4
��@����f�m��-�m�b�I��Ʉֻ'h4N;r�X��:�Ć�<�kCt&-W)DLJcM�c��[^�^[4l��W-z�#�X�)�M8�nNUw��|��+�$��^r��o�x�z��f�o���D������� �d� �G�dx�kQ�܂1Ĥ&��|� [l�{� �98h�>+��E77#�	$x6G�I0�K�;ڎ��}���E�s�M�/;\:^�ΝDf�Xг@=���&��2�������9�=lT��~��	#�� �G�|��#mLrA�AI4l��W9^�[l��@�s��LNo$cp�]�}�U����4 �X��(�������w����/�r���bOLcr= �ǀ�<H�E�/ $�m��Q�7&�_m��S@�䦀I#�r��9׬�j����m�+Jj�V�N��z%L7����
��^����#~8���x��~�)�[�M �٠����"��#���R�f&�`�< �c��|����[���x9��`�Hh�� �c�$���o��z��U�-Һ`�o�������=���7\0��%s�������t�bn�&�%Ȱ�e��< ���i8��~]��u%�k�/�����E��Se;&NԵ���Ɇ�H�h��ܮm�[��I�6_�\��{�~0֯TD�LxL�r= �٠��@��h�)�H�q����4,dP�ɠ��@��h�S@-�hy�\n�;@����	#�;4�f�^r���"���)pT�ـN� �G�v<H�m�k l�@<=��]ݪ�kdIP��L�\6q���1ąش��[N�х�S�sv�k&�A���j��qΎ@1�Iy��<����um�9j���\�ý���v�֥��mn��cǷO8�ŭk�,C^9���Mcb�PnW`��gT��
��j��!�b�D��Q���'al�$�����`,ڶ҇)]gvv��v���׉��qgՋ�����L�>���nU/ft��ݭp�,Aӣk$��M:L����TB",n�s�n���SY����4��< ���\� ���}���Ut�t��&����h�V�}�s@-�h��Qjcx܆&7&�k�h�w4�Y�v< �uD&���WN�b��	�2�I M��	.E�I{tLx�" 㙠�4�h�V�}���9���bN��M�A�'GV�I����ɄL�$��wI�h�XL�̎�#U\�x�cRM ����j�/��h���,N�I�ɉ"'&�k�X�8u���X;���ǀokZ��#~9���@��W��4��4]�@��%R48� 89#�	$x7c�$�d��}�����SI? v���j�*�נ�433���D���RcM4g���i�킥�m�N�i y����<k���&7��bcrh�M�mz�e`ݏ ;��L`�I�lV�d�I2�nǀI0��bN��$�4RM� �G�v<8�?�*B&���o�~���r�ޝ�u��ț�ԓ@/9f�m��*�ס�33�{٠v���(�<y	�d�o �8`vK�	$x7c�>_����n�40,l��7\]n��.�'^�t�ȹ.GT�lp	��ƛE/-�'��� ��^ I#�͏ �8`��T�#1b$��m�o,�-�����>���&,~)ǐr7_ {�� �8`k�$�X��M��$X�ܚ�S@����e`>o*����\��s1fǀE��Pɑ�'�[�M�w4�f�m��.qѶVE"��90s$E7m�z��1E������bK'W��id���R�4�a$����4m��m��S���;�ΚεZ�&&�7mI�$�=ʪ��{���y�éH�#IM�O�v&�[�S���$��ı$��!���UU˻����I{��������s�Px�bn%�/�������Iw�،I$����K�9\�r���%�$�%g���8��9��$�l�ԒJ�g�$��ı$��!��%�qr�����U�L�HFVa�:o�<D?���$���`4��~�L�4��Ƒ�}�~ h cG�����i%�0	��� �0D���|҃��8��X��,(���F �%b����q���#-�CZ� ��R��1,�����h4�3I�f1M���Ӛ���d�imjB���� ԈL�x�b�l�b���0$I��8&�1�1��0�-(�J�[ܙ�q}����9.��K�^!(�QJ0,�L�$,����0�3,��p��,2��3�lU4xѠ��b�8C��$���؎e56��ؓ���M�\�>~���yoz޵��{�ҋo�E��n��M��h�KiW�n�5���j{+맇�-�l��l��=��wa�kq����j5�ܻqy�8��G�M�
Lb,�WLW%�Gw��k����+�n�We���*��G��ۨ�	M��	۪�j��A�ݒ���y�V0��]v�G&�.|6�[SۦS�W�C;[u�m�	�V�8���(m�VgIdva-�{�+TurXuIl���`���n�B�6J�9v�ee�ݮ
�᫡��f�\���m5P�Qbƭ�nƞ+�g�fё�s��S��E����mn�<��@���V�1Қ�1���죳��p��;�mA#��":��H���I$����H���V�
@�t�vܱmqvӅ�@G4k�i���.5�I�������.�t��Τ�l�86�J��5� 2��rv 9��B�����9mZ(Z�m����]l6*�0�*��֡Ֆ\-ˊ6ۂ[(�t:+�%�\�qmp�P�GD��B-˵·�ko]-��� �m�cX������6�������P��UU^[����(u��&��ָ�ܽF��\�+W$.Z�us`2��
�gK��[q����ж��a.�l���&�I�=��r��؃�i�\��͞U��q��j���m��:���uO5�+\����1� 	uWKR���-���m��m��0 ��ޱI�KcN���79����fuV�إM�\T���6��r��蝓��+�1���a���+t�v�$-�T^$�݌^�(��I��+Ŏ��U����h��;\�y�i����R��)l��[@$ rA�|�i��*��1�a�O@wX2-؃�y�oE��G`v6v5��׎pTivA�\prr�W]���l؋��w4J��Y��������H�i�[���N�H$h�d^�v��ݣ���\��<n����pE���N����Ҩ~y��A���g���Y�۽�[�ݶ�z�����w:F�]2v#� V57Y뫝�Z��x�h��lV;%��6t�jw.��3�B�.�n�)�{]rc�{bg��,���s�4����a�*cU�< ��� T6�
��'��\H=u��kt�%g&s�m�������Ɂ88튶�ڇ��6yHh�Z��'Nw/k۷g�XЪ����LWa�T�ژ�\W�PF�u[��\/n"�[(�P�q��v�ǋ;������~���}�ۊQ��}I$�����$�s�Il܇�W+�]�{;�����B69�bR�NOߒJK��Kf�>�$��5�B[$}���i+WQ�<���ũ$�{�>�	8�$�[6?�BR9�Ē[sc�'Bt	]�RvϾI{�ʫ^�xx�Io���$��b1%�UU��}��IJ�:�Qd�cc�$�5$����ߒJ�u�Kf�>�$�$���k�Q�������,9�:}�m�s=9��R��wGNs2wiʸ��e��S�tGN*��������Kvd>�$�$�]��$��H�m��#<R@Ԓ\��~����2R$E���2���o����w�o�䒶�����Jۛ� �<��#HV��H����$���$��b1$��k��$����ɚ��#m�I	�$�����$��b1$�ܒ��$�$���Ѝ�`ĦA��?~I+e�jI+��H���I%$��JR�Wn�t��-ضV{i��37k�}V[<m��<U�b�݅7F�G�#J�ӵe�F� ���"��$px�II#�]���F$����v$�N���eZ���$�{��+���{��ߒK���jI*���\�]n&��1)	�$���ߐ���-Jꪻ\9�p�T���c�;/�Iv8�$��|7t.;*ݫT���/r��W�?}KIz��_�$��Ʊ$��G��%�W�6FycǉɋRIW�_��$���I$����	.b��U]
�$QP��g%�t#���3���d��Y�F�h�wS�(����;QY�1/1
��m�?o���$� ݽ� ��X����,�Yn��> ����{%�X�8h�9B69�4L�Drh��Z�"��W+�Iw�~0��� M[�r46H'�huv��h����{m��3b"���nU�~�w�3e���۫m`H�$x�`���o��{�������F.[Q7H�O^p�{s�$�rv�U��b:ڎ�\b���-���3�f4�X�����h��Z�����-�Aׂ�La�@�8��s��$E�z�����}�� '��{�:�i�⃋	���8��@�l� l����M��8�Չ��m�ۼ�0d� ��T�x���ɚ��=i"��/of��>Uʽ���r�;���X���%QDn�ߛ����YI�X6�;�gN��-��L.�qm�k�^�p�ՙ�j;�ێbò���Tvm;u�8�i�ݳK]ݢ�P�;;^Ri�ح6AƵX���qJ���O�`�q�l�$ 	���t�d5��`Ɲ�C0��u���-�����y��]��.+��Yv���s���z����0��G�qx�{=G���l���dJ�rFyK�8.���=���( �C'b�b G5s���)�J''�9�JhW��H�6< ����cv;V�l�5M���ʮ$w�~0zy���q{lbS��	Ǡ~�S@6lx}�%�p`n܋ ;ZjV��	Z���r����~0�ذ�p�/�H:�Y�F�9$�9�Jh��y|}�� >�<)���V�d�������T瞸z卸�i#�a8+0vMқ��M8�r���$4/y^��G �l����?r��{��~�_��(�I�8���j��٠su� ջ/=��==���ˢ������π7��� ݽ� �ݗ�}#��KB6a�L�Q94>�31[/V��� �G ��հ����4�V��5l��z���{<|����{&��Ԧ>&�ui]:�@�Ԇ�]�r��4�Is:yqn�U.-l,�f��m�
��H�6<v�/W*� ���@.t�[�y�Mŉ8h͏ ݽ� �$��3���_��g�����Lm����h���@ⶽ/�<��1�e���@��u:�nc"�	<NE���W�������r�4q��ń�N'�8�ָ`�[�y��<�[%�jl�����h��i]��Cqˮ��[��;v��b*�ݳ��4�⑓�n��x0��	$= ��~x��X����\�}�� '��;���4շ�n�ş㜪�Q\�"~����� �竜�����U�~����L�	2%"r-��|���h�٠s��h�����b���r�}���y���`Ns��+�Y��r�z)���D׉��ۆ�{$x�R9��Oz��#�;��e�����(�����]4�6 ܷ�;�`�hr"s���(y�g�v��5_�{��/ >�?W>@w�� ݫ�}cNd"rbO�h^� �m��dx��Y��\�s�I�\G�X�M�n��x�{� ;��*����z�.w�@���b�x0{�7���W)/���Is� ��^�r��K��� w��v褝1!6��ذU~�U~s߯������Pr��WԸ�#�{�]k_i��f�Z�F���v���v�v.=�8�(�� F��u����F��Le�;��AM�:��s��n�k9�Xm�tp]qm1)��Yy%DOn���n�=c#v�N���Ǌ���ɸ�A���Ƶ\ӡ�m�5g�h�o)J���p6#�R(H*ۉ{x�8zd��8p)
S�nb��[�6];p�N�n�����e�EFM��O'o�{�3��#n^7�^h�Z7n�]J�� 랉\�<	���Sv˧��ڶց��׀I N��s�U�	.y`[<�'WN�V�@�� �H��UWo��	.y`wk߼�3ҝj"`�bn,mǠ���7ob�"ݗ�I%h����+�c���{� �H�;��]���-�:�m)y��NE�E�/ >�< ����ذ�����2�خ��:Z�]�K��wnō<d�9Ͷݷ�mӞN��Z�}ޮ�gӧ4�q�K���{� 'dx��_�A�'� �����Te�J�6�M���<�ꪮW�ʔP�.��	�]��9W���k�^[f�y�$�w���)�HRM�<�����\H����v��-�Nյm�.� �H�nǡ�y��f>�{��8�ߠ�1�y�$;w�I N�x��X]�x�{��߻���錷YXU.jݮl <�Ru��^��s��/n�$
gh��~�>O�ڬt�msl�o���<v�,.� �H�	��#�C�$]7lv��7ob�$yr����gߐ���-�:�m)yӤն�����#ü��9R���� iIX4�w?y��b�� x����䓆"*h��}�?y��&ҡ���P�����̊��V��-���ō�XN&YdN9����2�K
0#2�Z��ZӚ�2j��,1���̰�#,�����lq���`��ce��YdFfA��`�~[!���x��C����=X8��C� �'_��7ʿq��p�o$$L�q��c�	ݏ ݽ� ��/ ���}J��R��WlI�� ��<�s�9��[<���h�s
 �o"��")R��V��귡�g�B��P����vWdm��ӥI:bBm���`vK���@/9f�^q�F��L�8��@��^�^ M���ذ�ꔅ1� �G�~Vנq[^��>U�q[^��W
�FLS�7#�@�^�{�l��s9G8}Ew��fKvh�R`�x�<q�$�@�*�5M��I�l���w���[�C�s�Jf뗴��,��wQ!�㞹��b��q�8��j��2�nz������[�^ }$xT�x��X�!��HH��ӏ@?[f�꼯@�ŀj엀M��}J�e�^U��	��W�� ݽ� ��/ >�?� ;�<��1)�M�����[/V�Wo^�~���<U���V��92y!24ڶ��l��UW;~���"������U�(��)��>��5;3{њ�y��^�%U�	ɣv��uK��]�����S���6;O^��6�5���R�&�\tj:�u��W=��ON�q{dK���t�Z�DU�5[��
D�D�I�1�N�k���g��l���Ϸ��z�՘8{v̯m��P¸k���\��[u�捵�.]`� F����q�c��L׍��:�;���������n�ts�ڑr�gN[��w&�t�;D�.Gk�t�2�u���=��>76g��ͻ��~�x�l�v�/�\���,�e;FLS�7&6��8�+�9�ʴ+k�?+k����ΐ�`�x�<q�$�@�_~Z��g����]�^��xJ�m)�x���RCC�_{נ���RK�7ob�7t���j�;LlM� �H�I�{#�h��-{�p��Rcb��1'� �Ѭ�m7�U<i:^¦&9k������q����wV�o�{�x��X�"��� �"���BIӰv��{}�WCD�D��_�\��~�9U���|��٠U�*��'�Q�I��Z�ՀI�=�y�\���HN���M�v�X�����r,x�gz��F^�Lh�ܘۏ@/6<�G�/���z��%�.��۞��m�0ر��Ų�2ss�G+l^����ښ�L�x�Z�=x6y�S_m���j�*�@�[_ߐ��@���q��A�Ȝ�@��U�~Vנ���v��K�025$�H��@�^ M����`l��O�{�U��	ǒI��/���@���@�����{נ�w��Q`������`l��|���dx�����߿���[����f�-����sKB�mݮ޺읶�n^�#��"���}GmV:i��^����=� ��h��Z�8�!LN�b�@���@.���ذ�K�ܪ�H=�W��v%01�1��v��@�*�亯z�W{נ^gXF	<��4q�ʻ����^g{�r�/��P���|��}�h�I���dy!�hI/ �I/ $����`B�U��qP�:���T�w���~�Y��z�&(��nt��5����9�����������@/���v���?�a������߱�`*ut�n� ����r,-���k�y��6qt�4$�X�m�-�y`���������"�QՃNx�n&��*�@�[^�{�f�|��V��h{z�)��4��	ǠuI/ ;�<v�XV�xr�k����/�
���N��g�;�u���%S{�қϚ�O�\�g����Ͷ����9��zcq��W�q���ۮ���������9�]�<���˱8ݡ���:���b�2�
��.�Z� ��Ӯw�P�6b;s�<��\���h��Pt{a����ɝ�v�tm�ZL�4�WI�l����v ��]��賯P�y�}���{�����Ι8��}S�vR�6f�͈͗l,�l[�=��v]�#��4�v2c��rcn?@/of��r,�IxT��	��#��$<q�RM�v��mz���vG��*�"l��-:`��Ӷ�^�� ;$xr��$I�<K���ܺ�!�M� ����y���g����呂}��M�v��k�/�oc��1��I'����8�ZVנ�f���f^t]���AI�)0p)2k���6z��VS({�͕�ng�[u��1\�����}�B1��!$$�����*�@�[^�[l�*���Hc���k �Iy+�ʯr�\l�=����<x�Z�r�
dy<�#�@�[^�[l�8��@���ږr�s8��Ɋ8�>�3>�33�ﾚW���[^��3o����ɍ$<q�'&��y^��fy�}��y�O���W�������S�$1�S�1ƌN7.jhf���/]� °�]QI��e�q����G�MP�.��x[%�fǀv<��^����U�I0N&4�n= �����WI�O<.�x����]*���Bm��<�wc�?U����r�#��4'����Us�u=�x����>P��'�V�&��x���vK��� '9f�WP�0i�$m(�^���\�~����~��~��< ����~n���i��Z��ZD�9�Pd�̥˙J�[��0ۜs3s���ūus��)%�ݏ 7v?s� ��z�Q՝�ɋIc$�zy�4��^������3�;ܤ;	����6��o $�x]���ʪK�������=�N����a$$�@��^��;��]���+�C� a������b�$��<�x7�궽 ���� �� }Se�g�yn�˂����t�<pZ���ڳ���dC����6$d���x�r	)�)#�����;r/ꪯ�u{޼���'b|un�l���U)'��{o�X����,߼�<H��F�4�6�rM�~���� &�x����T�)��"b��h}��{��ho{4wc��\����`�ʽ�J���m��x6G��;�+ >�<GW8���!�ws(4S��
O�SÆ��l�w0���s�@���J�Eb:e1w�� �6�C�0p�FlsZ��1���25�\��p����1��1����+1�ȳ�0�I�(,���LĊ,ɉ�+#,��Ȍ%������-�[֢�i�-ڐ\���,�+�{5!�ѻɸ�̣���.6�un���,�4JX���u�#�*�qe �݌�'Y2T�;#�[App��ax�Vۭ԰E�B��vF�n:J*��U�!��MU#3���:6z���5���v��i�r�ܔ(�zS���R�1��y�du�nζ���l 5�kO�4�clBx9��n{�p`�(P�n�L]��c�F#�Я<�u��2�WT�m��ymt�T��ó�ؙ�a�܎M^�\�P(�i�m�T�Q\�6ٻ:���rpu��-��P�3h�� R�G	�+�ӥdOAq�r�he��C�M��˹�s�I�6��ʓ��x7�7n�]��
h'�&��+���M�&��m�Mv �m����R�u�v�v ���W��P;�������X���n��9�Y݀�v�;h�g�p)ԛ1��z�kh�Q�U1�n��=�&����ګ��H9�qb��	��a��nJ�� 	RF�� �G[��$KdF,m��/d.ێ;mnƚ��l @O6�ܬ�j�"�'>ڞf�M�ù�v�9z���L���@�b�����P�&����eU�+Tn�i��ui�Izۄ����6�-�[mЂ�hے^m��j��:�{T��j��6v �)[`;�VV�C]���3�t���ͮzV�w�K3<v�n�\��3�uh�U��L.�� 9�X`mp֎�d��i3qYsl��������{vi:R�jXyv�痓�"s�#ngR���g��v�vVڥ��ml�Kc\�8%l�p�G6{K���̪���jy��WD�8��Q;���#���U�	` $ I[5Љ�Z��A%ڸ��v��nv��8�xKv2'��)���� ���8�&Ud�:۱�C�����d�͋Zz����;��tF��q  %{-UP�m����,B���яH=u�y�4�1փ[�!⎁��qBm�wR�Pt,� l�ʫ��_ ]�=5Y�4oEj�Vf�9u8�4��G�Wuuzٝ��EN���mƖ���˩�{HT�j��,p"']��-��c������ˬ�fse4WL��mz�A-��[�T�Z�c�SuMvw	�Mզ,�JU��f��^�6�8*�a�X[�������v��q����*ݰ���Y��{5��5�pnH�q�G�X�ێ^.۩A�+�˴��{�'\�FS�j�#�ˢv�OhcR�����; z7��Ymq;h��˻1�V n��	�2��#�UUW�l��9�}O�3&<NBA�4���ǀv< ���ܮURF�F�aC���t�t�� ���x&ǀ�&�`g����Y�I���w�W+�K���of�o%47<���3����"���N�[����ݏ �^�ޟ��w�zo,�;_�jGdmș�nU��q�Hu귌�<7cu�����D�<v�z�AS����6lz���2FҎI�}��|���l�\�|��y��z��wV�ݔ��f�^w��UW3���L��wc�&���r��J�ӥJ�\��;w����ݏ �0����j�(�5�0Y(��s�`c��^��R^���7j���C�Lhq������٠�f�s��@�.;q��y#NbNOd�i�kyD��pX�l"E��ۦ6�%$썒/�����2G1�&<Q��}��@-�����s���{���==���U�$��Zm��=���&�`�G���GN�b��)�4�٠I{�r�II }6< ���X4�6�rM�ʴ��h�٠� wuJBt�uj�be�x����< ������mB��>*�^d"aݮl u+μ���XIn��El�j��Rd��&<Q%�ɠ�� ������>RK�>�E�M:�`��M��������Kf���u�L�521�4
��@�I/��G��< �<��Z԰��lm���&���/ $��wc��U�r�������7���UҬ��ۦ�m��������G�^ 7�����7:+e��+<RULnw��B;��l�*v��B�bqqt�Av� wv<K�`-��I Mۈv���t�X�m�H៹�W9ă��x�{� ;�{�Ăl^�'M7Che�v��{׀H��8��zh�gM �UkqB1Ȉ���)/{�x�y�G �dx�52ƢI��D��@=�,�;���z~+�w�ʮ���*��%A�{�̽u�Ft�3F�e�ռ�Fut'LngZ5,�s�^�h��<۷N��g��]�E��bڛ#��mnK�m��*�Ơ�Z{���M7,Ӥ�{V/��9c �v�x�N�ΐ�S��$�]�n���ֺL���j��-�nΆ;e�[RFԆҵ�3	��K����������k���T.��k]�'kp�q��b��t�v=���F}wf*�7q�e(��t��.J�G�M����!s����0'l7)���K͂'JU��~�o��-��I wv<wjbj�N�[M;n�m`-��I wv<Wj�9���Ǌ�9!�#���� ;�%Ȱ��xؤ�ӫt�m����ǀIr,�^ [l��:��0nci�)$�-v��^ I#��ǀJ�uj��-�[��[7��4�Dy<��iͪ�NGf�G^�c[�+��+�ř(�m�?����m��9f�k�h«[�y����7��]��4�����@p9w�@�_j�?.Z��x�TQ��WE�e�o ;�&�`-���Y�{�:�cS��#RM�ʰ��� wv<n����av��-�i��l� $������S@��,J���$��BpCě&Z�jz���6��P춥�v�V��rv١?��x�}an�B�� ��� wv<Mp��G��@N�;4ն�m�vG����<�)�^ N��b�� ���$��@�|�@���7y��+�W�_�� }=���!:wmZbe�M�-��M� &�x��h��^LPi$��o,�vG�I{ղ^��'N�˦�X�f�rƁ�NkZٌH��^ɣ�.ة��"�1��Q(�,x8�ӓ@=�,�$�� �l��lx�.+R����5qI4_*۟͜]����}�y�fbE���Q`��NI"qhg�< �c��ǀI{�?��Z��m��I�>�3���o������i]��r�*#�FT 	D_\����2Gwf�{U��52F�p�� ��x��`�#�	6<�s�����������ضT�^s�'St��x���n��6G��+�{eZYG��|_m+b�n�$�}����l� $������HN��V��n�k >� I��wc�$��=T�z�z�hv5i܌nM �of�s��@�� �m��8B���$�c�94����`�G���R^���7j���k�6�D�$�@�� �m�o,�ݏ �*����%��]�j��lWFK;]���H�6M#�v�k\��Z�7\�k���7S�3�t�Q�k�8)�1�WdnX
�7@_���{Q~=�f�c����u���y�s�*��k2�vg��đq�����'ݻ5s�H=s��cǂ
�8۱c�^Wm[J��N�m�հ��]�$E�mc�v�֊���vCC��E9�58�۪�zĸ!��ww~�����ۮ���.0ɒupW*��7�>��Z������Դn�t�`sU��BF�l$�vրM���� n��U\�z�V����~ŋ���IG$��w� 7v<m�X���b��N�V�+o 7v<Kذ�\�r�;��h{{4�r�i����(���`�G�lx����HSq��AƤZ��4���3>��������z���Uy^�ˀ�u��9»k�"�������I�7fx�c��E.6���s]���H�A�����yf�n�xSe��G�N֌���#Ff����o|���{�c���8z�ew��Ҙ �*�#LF(�`�i�~(!�n{�������|���o�y�G9�����yo#p$�@��y`�G��I�y��� �Mj��$y#M�27�s<�3�<����= ���4����h����bf-�v��� ��� &�x�ذ	ەh�	f,#PRcI�p6��en�`b�{�Eb� �rb�-��[�@0������#�N7�r~ ���Z�ڴ��4.�n7���5�@��� �� N�x7c�r��d^�)�8�x��R-�}���,�s�����$0Pـ>8�l� �#a�m>���i4�0x�ȯ�(���� .�!�AI#����0�K!��(�H��% E	L�D�Y4C̉O 9���Q�`(�!�~T4>��?������~����^���9U�U%��whj�`�X;��ݏ �����/k���3ɤ�J��[�]��nǀN�ŀN܋ 'v?������?�뛎}L��V
a�Q5�[f�ֶ��b��N5rv\x#���#)��M��m���;r, ���s����h�������2'�}v� ���nǀN�ŀO��}J��m�#�~ �/f�^r�>Ļ�z����� �Wz�9�q�I&����^�� ����'nE��IN�x�9B4�x䍬j9&�}|�@���'z� ��< ���V�L��8�ա�F�֢���qX����X���ۢq��]L̍LB���Ǌ5"�/�ՠ�W�v<v�, �*��v'`�6�I�_yf���a���}_~Z��W�fy�bGy��TK&<���x��X�v^ N�xt���F&�,� 7&�ػ�z�U�zy�4�9f�����G��ܘۋ@�n��?qzO?�;'�;r,ySk�2B�� �b�ۑ�vBrn�W��NS��-����j�+���L.�I��M4����V�wn��͹����Qs��S�;�<�gp�9���
ܑ�.�{�Q��Q�e��g�:���FKKn�5��왻n<�u�\�N�\n�Cu�qm/j�]�v�TK���m�5�Zh�c���	���p\9�<�݆W��w	c��y㋵�\�E���.h���=��q�6�}��h�s��m�n��i�ۄ�n6�9[�&�&���>x���~��A�@Q�(㏀�~��yf�}v��? �v��:��1'0�9"LnM ��x[%�)��nǀE	6�F�q�II&�U�z�y^��Ď���y{4W�u�(�q⃃����x6G�ݏ �Ix"T���Y	&)#�m�|W���^�� �M��}ݡ8���6��6���'vnܶ�c4K���݁6{d��m�8�q�Ƞ���@9�,�*�@��+��f��u5�cO#����]�{�s������5{=x��x�fV�5�v�m�lnLMǠ~W���,���<J��s@��z��w���c�i�8������=����X]�x�v^�"�1'�#�A�4����*�נ~\�z}����$����m�A�F8#Y:�9.S���.]��D�X�%��������B9Ic�F���\�z��, ����ϐg��%��&[��j�m����=��r� ��� &�<�r��<��<H;Ժv"27�!$���_}���W����BH�)��Cuw��z�V���!TC���6���r���<�-���{ N�����"�x�rh{�����s��_ {g���+ �R�e�^dn����Va�w��h�S���{�E�-�K�����B���f�x\��6���� 'v<wfV;{�=�}W�˺i�Ujݶ� ���?�ʮU$zOe`��h�j��<H��WTbN,�����{+ �{�q/m�� =�� �U��"��(�hw<ϳ��3�y��r������Ww��x(� C��ID�p	ECP�j�Us�*��>�Wv�):L�mR�ݦ�;{����y��x��Xm����s�q1a踈j��9�r��	z3n�u3�F�e��pnX�o������4�y2�l�k�o��nǀM�� ���@�N��0LrH&���,�&�ŀEݗ��<����TR�I�1+o �{v^�_�U\�U��ߦ�}{��-�uF���67#v�v^ N��	ݙX����3��~����^7�E������w�@����~��xyW����Ws���*��hO�0��'��6�z-�VZ�j�Y�ĂhM94pj����� 5��3]�.�:mq�Oa*��[ ��"�ˋk=uFx�0r��4���֭�BӢ]H1���3�nMB�a�(�qK�T� �T���W��fj����=*���c���g�6[�$E��{��񞊶8�Yx����6�oQw��}���n�A�}l%����N�Z�&���߽�nn~�Y�\�јu�q���kkz*
�r���R�-��]\�:�i���L���e`���_�׀lx�UDcpqDB73@���ٞg������w�_yw7��8��Q�b��țq��W��@-�}���h*�h�&��$���_lx;��n���+�K׳׀M������Ӓ`��}�\�z^� ��4W*̮F�c�N3-]3s������Jl�$h�z^�y���Bv�1�Xbm)��\�z^� ��;���y{��w���i�H�1��x]�y)�*�/�<n̬-�x���}O���BiP�ۿ�=���'vea����׀yl��U�]�\k��v���W){g���O^v^ [�4+UDci�F�$RI�Uv^v^ I���ǀDD���Pn�pUrt���!N�y��l��g<s.������W��qqf{Y[4�6�[=x&ǀ���e�E	hv�ݱ۴���m��wr����"���W8�6��\.���m������U���/�*5�G�d�sk��@���u�X1���۬-�x]�x&ǁ��9\��߻����ԑH�1�n=�y^�N��	ݙX[���5K�wm�����l�]-Z��[l釢�Tfv�<�ް"�&7�77b��F�5�;��h�2��e�we�v��$�񧑥�@���o�g��[נus�z}�hT��18(�pm��*�%�vK�	�7fVջq�O	F��C��g�.�w�@;��h���+�]���] k7���U}_{�i�ۂ$q��_m��.�W9^�W�����"`d�� ��b�c�K���o$��b��y̛��P8/	h�;�B��؝��Mٕ�E�/ ��?��33���y��}y5��LQ%m�n��"엀�< ������q��x�mƣ�@��^�_m�z��r�I�� �׀M���(�Iڢ����o��nǀE�/ ������
bN$�c#�@/9f��.�x;#�;]�Ur�;�+�I�T='hXF_��&��<p����a<	�`D~1� ���K�>L xf�-�$��I�f̟OƓ�C���,���ΖVNe�3XFaa�9fe~߇��M1�8��e��?���%X`hњ�ю�Ϸ��v��=v7���z]/N����=���������R���UmW8]E��FWz�eu�{n+r�moa:M�;Tۋ��h�x:"v,����k�Ѱuv�v�c%�3�uk�����v��m)�M�v�������F�ZKP:+]:޹�.���tj�n7&�&�-�)M;����6:�KP<A�?�|�o��Ҭ�5)��f��tf��W$��^7j��h�z�\��u��k�0����[q�Ηnmɱ�mb�3u�J,��8m���ֲ����mg��)Y�Pv̱���u�j��ۙ�v:f�eڸV�*
Mvum��T�Pz�u�"Yy9�9m���0u�Fz0;���v|� �5Vݱ��:.�W]�'[W.'��,���p+�:�ͭ��J��t��hn��h�(-�UĴ��WdݖӮ����³�E�V�$2���I0��6i#[\-��خ�0t�Mtiۭ�eऊ8��tҡ�������A�cnk����ő���Z��wiP�V�y�ʶ^�i��a�Sg�x�Um�ݶZ�U�ʽ�l�qU��6�BLΩ���5��l���m�m�m<����n^�cmNے帠�/n�d=�^�55[mD�lN�������%6Q�d3�77GFR{e�⸓[bG�%}���9�j�ڕiV�
���
h�8ٺ-f��; ��=���M�9p���F�~R��e#ZB�U*eR� xl�m!�W�yy�!��vYӄ2��
@��s�Ѷm� �� k�kj��d�[Zh烑���@q1�2�[4�Nn����:6P��TL�ks��.GR���ۃ��ݖ�,�[T�.��O4Q�Ki+j��c�ʭJWR�*;�,���5y����q6;r��UUmUUR�KV��I�'�f�.����F��;=�D�ZGz,�z����/K����#���v���x^f�&�ݮ���YCH�q�+m��Vѫ��@-��*K#�����`mҫf���=�PV�f�{��Et�|���HW�&�:��~��Dڡ�o��w�e�N
 p��	��R�������y;Q�d�p�h�C�����:ڶhCg�j���#[�T����=�!s�n�v%�:�]6�%�{!�d�y�U�"�����@ ��bh�1Ű���NZU4���lu�f���gwi�󧪑�Ƚ����+ؿ7n�w��uư��[e�nF���0c��S�ܙ8Ԝ�P�E&�8�M;V��*����iv�t)ݶnح�d�a�9�N�5oD�=d��vɒ����Ϋ�[#�{���{����r�AX����忽x]��vG�v<�v�*16�0��9�U�{��y�� 吏��\�r�ʤ���/Z�v�)�v�� {}�N���"ݗ�Eݗ�}SS"e:T]X�'m�ve`n��"엁�s���W��� �N?+wN�Z�t�6� �v^���z�z� ��� 'v< �M�v���X�ذɒ�� ��������5�m��P�F�aM�N3(�r96�rdn/�ur���٠�6�,I�}������![{ו_{������ >�� ���hu��Uy^���>�b���d���x�x�ذ���vG�j�����իWm�~�9��9����׀�< ���[��I�0JjE�U�@/�� ��4�ʴ����h�"��y(N���ѭ�t�7mm�!��%�죮ׯWZ��L�bnDB9�@/�� ��4�ʻ�9U�U|��O^��L<�>*�1��;o 'dx�ذ�e�� پJ�y1���/*�*��M�};�x*AH[ƃͨ�Y���*/��@���T���N<�š��g�y�f?�����呂[�4�ʴ��ﲁS/�h�շ {}�r����������h^W�s�:�XF��fȎ���Z�]bU���]�F����(���w{޾��/V�Κ�m�=��E�/ �l� ���P�C�<� ����\�zW���٠[˹��#�H�	#�*�/ 'dxz���R^��V�'� %��������l�-���"ݗ���ʭ��T�9��ojE�ڧ��(H�M�]���fy�w�������f��9
���q���S�Yt�͛�˹�\�[�-/�u�W�[Mی�<'������Z�
�+��f�o.���"��$$LM��=)��l� �fV�y��9T��_����l$F&��>��M�]�?���K���@������X�&�y!2�M�]��k�*��@-�h�r��&E$N��VנW+��O_����	6e`�Uv�%t��z��9�2�8���s�\% ���um��f�.��vn�6��+s5n�`M�mv��^�]��W�����+vx�MBy��B�9&3ۧ:�K��{h�\)�Ӕun��lM�}�@���)tu �қ���VP����ݎ6�<nI�l��c�����Hn66�A��8�zvm��7O� �9۴�]pl6�m)��Y�{��w��'ֽ;�iq��u�ʹ�+V��l�%�Z8rhq����4�Da)�~W�zm�@��s@�ڴ�k��H�$q��I#��H����/{׀E�^݄0T���cwCm�d��$�9^�[l�?s)*��F<m'	��X�"�"ݗ�H�<���Հv.��G��,RE�U�+�m���s@�ڴ��P�ݚ��s\/KOE:�p0lN1�ye�9]�m�a�Q�I� {1��M��}��@/-��ՠU�^�~�u�bn,�)�drh�f�y|���7O���|���@-�h�-�L�F�q�"rM�k�"�/ $��� wvZL�j�"����w1u���{�� ��Vנ�Z#�#�8�����<�����we�[���c���VV,�k�.�3�{�	����>�gc�&�����͎���e���m�ݏ �\0���W�zy���RF���#�x�ؔ�㙠w�t�*�����@���h�r*�NFH؜
n�]���\��}��iO@�X�JFe$i��Q٘��Q������ʼ�^������~��E�%R?���_}��@�/w4]�@��W��]b����	��m��e`\� �d� �G�j��~SJͺ[�bz0�GS���'�/ .���Y�'M��T���u��z��E�^ I#�&ɕ��V��O��@��� �٠^[��Z�ZjT�4�0i�$�@-�h۹�|Ļ�ޭ����=�LV$�6[I�������9�^���e_}���U��{�UŐ�����T# ���%�pO�ٰQ|k�>�|���;�7��F�f�&h�V�U�����w4����~s�����n�n������v�n�ŷ,�]ېiR�ۓkn6w�\��{����$���Ф��>_}��m���h�V�����)��ܑ���;��h۹�Z�ZVנ�]b���y 2ɠ[n�k�i�y�uv��{���NPSjA�7��K�`M��H�	6e`we�Ɔ�Dp�p�*��@-������{���`'�EdM�n����d#���C�<�;���wh���������m�1��il��BF�#8ǘ3ю�[ ��6/��}[�H�;���Hމ�zm&�N���V;��K�j�v��d��5�ns�F@PV% T�Ӣ��I�v�m����������įl�Z���i+��B����cT��vtίl���]�&�{m\��i&�e�UU�����c����7V�z."�����מ�k%��eܕ�մ	�L�j�H�ԊbII�1�#�����@-��S@���yK��H�m��o	$��f�x���t�:�z��f��Gy㫱�F<hh����;�Κ[��I N�x�Z�m[m�М	��h}����@;��h��hw�1w�ޚ�;�߄�I��rD��;�y�����y��"���*�������H�Td�:�E�UY[���ꦚͦ� B�&�H�`����uvKL�lt��צ������:����V�wl�n�	#�_+����/��\���� }6<wfVz��l��4МR<Q7���@-�h�]��)�_GU�bII�1��@$���2�	#�v^݄�bMժi�����N���=\�{���:�z��f��z,+ĝD��	8u��j.3Ҹ:���gfr�Jp3�zU7����)Ǎ�7JL�-��\�zm�@/����*�NE�1�6�-�x$� 'dx�"�r��ϻ�߅���Rc�Ȝ���}���w|�x"o�`FL�b��bɁc9R@IPx�x�*�CHkdi����0��D?1��FXHZ�����Br)0��	�c�&SH�@�2 Q���`�&e8�`����!DC�&AN-�	THK$2Y��b�@C!��_��!��{��C~b�x?�1j"4����s��~87"_QD� H;� �Oô���������lz ��mA+��sܮ%��ڿ�A�߿^ M���һb��H�rhu.�٠w��Z^���f�{U��,NdmĤJI�Z�X�r���z� ���Mٕ�D�t=��]��v&yz�SҠ���m�%���B:M%܆y�>��ܔ����}���^ I#�'ve`\� �.(�ĉ �I��@-�h�]��j�*����y��fy����ؘ�s�H�i�M�߷4]�@��W��4Ǒ�؛���h�V�s�����W�}��_�" �fc��#����勮D8I��$Z^��ꪮU/{����$� v���h�M8��c�7j.)C6�d�Ġ=�`�8������Q��tR�����{���	ݏ ��X]�x���&�I51(G&�}��߼�3<H�_z��^� �ٿ�:��S'26�Pm��;�ޭ�r� ��h�w4��bjһC�V�� �d�-�����y�c����@�����b	 ��9�@-�����)�U�{�U��Q� ���|赯�Vf�l8v�r�b��۝iC\��W9�.�B�vy�n���G��&�[Z���J��K,��v�2������ӑ�8����@������m���.�\���˷l��ۨ[e$�m3�fe4��i6z�Ւ�8�N⚷��$��-��5���;:�J�%��rt�ɺL��-�Eu:�m����Z���óN����N�<m��	�s{�ߧ{���wߍ]%ݢd�X�+����a�֖��2�r`�M9�3W$v�.b�	#M<RI�/?��4l��W9^�[l�/�>+O<x�Q���Hឮr�<�����<vL�wZ�Ĝ$��&)�9�\�zo,���U��^�{+ ������Wcm:�i4�Wn� ���6L�I2�?��/]�z���)���,�1294yw4yw4
��@-�=��[��nغ4e�c�\�Nx�N7Z0p<;��Z�[�+�i�mH��#��F�LI��-�s@�� �٠^[���&�i=�n��[�ʻ���qA J��T�Љ�����_�����}��)�r���b�A�G#�m�����w4
�k�-�D��ŏ$�&�(��/����S@��W��4���U��4,�ڎg�=�?�z�z� ���N���ԩ��f���.dV@M���p}�0�6ٶ�mZl�W�M����Q�p�CG�yl���<wfV$�X��gTa!�F�nG���f�_yf�m��^�癉�K��X�L���o|���{�U��}�z!(����y�<���נ�{4ڭ�c�(�N(��-��^� �٠�Y�z�r�I�q�'p�*���^�����e`Gh*^R�Hh�G���`ss�b�� \�Q\������<u�n�6x��D�9�$BNB9�[l�&ɕ�M�[%�kZ�]�Ut�q6�G&�y˹�[e4
������c�d�6,�ڎf�}��hvK�	�7fV$q5m+cjcpJ	�h{k�yf�yn怊�&��(`�G}���ʿ�������$Ndc��ۏ�{���<�;{�����hrנw<�3�n67�NcI�u�m��J���@*H�м���3��Y��!��ɓ$�����yn�@��� ��h��6�q�i������Z��f�yn��9˄��D�~'$��\����@��s@��Y�^�9�$ yv��	$x�2�	�2�s�^�޽��3��L$�6�8��/-��'d�0�e��<�_s��UV���8�;T��6��1��v�䭺Λ�(��G��t�A����sv1�X,a�:���+gi�������"פn���=v݌�3�Ӯ�v�1�:N�۲��/Gkm�ʘ'8$���".U����:���{ On۵Q�s��ݱm�t�Խ�<��x+����ڶ��m��kp��U�"�@�Ȥ5糎C�q�"&zwiܗ;�њ�7��Y�g�(?¨� ���{�������gm��<�C��
⫎I��5���k�;qhu�.ݎ�ܷK�)מ�lc�o�7~�0�e��?�s����{4�Ψ�����IA��-�x$� 'dx�f�=3ɲH�ɉ�$NG���f�}�sO���Ur��{}� �׀on��v�J�:Lv�;&V;&Y�E�/ $�h�[�mD�J27�9���f�� �G�Nɕ�w��&��賫E�z܋��I��=v��݃n���c��.YB�3��yY�7j�:w4�߇����6G�Nɕ�|��=�`���I��][m7n�l�;VUeU�����qF��3�����*����\����*=�encxIM�������-`n��	�<{Pq7c�t�cM��'u�X[��l� ��+ ���$�8ǎ�hs���@�۹�_y+Z���)�G��p7Ar�-5t���m���jѪ��BЍ��r*2���_~?v�c���ߤ�~���<w\��E�/ �n��Zj�t:,v� N��	�r�� ��h�[�i��$��9�����U���뗊(�"���+"r�.�}�{{��z�r� ��ny$n5�E6^ M��l������Y�yygz��"I$�F8���f�_m���Y�U�W�{���H�x���OB,�X	�.�s.�&�ks粼aN���{��mq�L������M4G'���h���)��nǀoj&�aWH�[7���U�}�5s�EQ숺��}���Wm���@��9�$Ln),�"ݗ�v<=��W=���='������$n@nH�r?����y�7����o�_����*���V�EC�S�����3�z�_N�cME�L�x�X�r�� �����ߟ��<M�[�bhؕm����2Y9��RZ�t�B�؍���ظm����h����r� ��y��z���ۚ�����2AƢ�*�+�*���'d��&�Q`Iv�6����x]�x�X�j,-��/iZdncy$kq�wy����5�E�/ ��/ ��M�V��t�o ��E�?��Uy���������}�*�EQ_��EQ_�ATW�aTWEQ_�E�*���"*����((� �)
�2� �Ƞ�� �* ̈�"�4
��(��?�E�QE�*��"*����+�"*���DU��TW��"���EQ_�QE؈�+�DU���d�Mf�cp�f�A@��̟\��>  
�          ��RL  P��@ �D"���PP    D* "U)J�	JJ
 
 ��D��
����  
�P
�   �PP�1� ��zj����\Y��gӽ�����>@�zS'�g��k���{q���������qe;����׻�����]�[���3���+ӓ�X }]��O'ݪ���i���0h� 炀
 (�  ̀���n.�;� �Р �  �biII���&������4�FSM))���g'@Tbi�����M�;�������s)GM"h�4��)Ft�R��vR��&Ri�&��HJi��� 
� @ �Gr�SK,Ѧ�ggI)K���)u��� �%9�>�}�=������8= s�������=| _v���ϥ}�˺����r�{��x�K �ӓ��X�|�������f���¨��P   h$��cn{�^����zw�An�=/� >O�S�{�yO&���z��;�ϥ��+'ݥ��u��[�+�{ދ��>�O���N
�i{{�ϩ��@ ����������[��w�ҏ ��PP�� 
R�� �!�E,�﫟}��ms���xƓ@����Ӑ�t����:u�  �<�Y�\�x  N^���iS ۪��w�Ο!Ӹ������>_l���q���/v���}����> OI�L�*h  O�5T�SM�ɐ�O��Oʀ�ت�m(�j��T�Д{T�)   !HI��)�L��x��R�w��k��K�����,׻.�v�o�I%UT�z�� U� �
�� E� *����*+ �����Ǻ�@���c8E�pޱ�98���iذ�C����Q�&,�0�:i&��`0Lb������Y�������h%��UL�Bɡ ��J��b��6��M#f;�aŲp�q0c$d�c&`#F�Df;�a;�FZX4�`�&$oy�4d�X�A:6�g)����X���f�f0����t���k3�mĤ1��\a  .FF�����3F�FAc���a��cF��k2��5��[#G71N�����a�A�EDX�M����d�$e;�E<�Ӱ�Fr��it��Eo�dV�G�@e��\��f*"�DE�8r9184���v�eR�ř�"�����3
Ih�kZm8c&��1�$���^6�;S2��"#3{���V�X��51i`�#*r0,�%�ă�['���Lqׇ��F��\�1&y9�,-$O,��q��E�W��
4��)1XFB]8� i`	RU0PЄ,�I���bT�L0��Cqet��*p]4�HhȨ� ��p�qdLM$2M��f�����0�#���t����@��BC�&"����
04�D&�ޓ$�30Б�Lt��GI�"� �%�\5��$�,��l6�&�"E�16���� ��30��8F�Q,�m8�S�q⦷��k1�5&Z5!�8���p�k&�ٳ�RIVkol��Zvx�N&��jIa'���;I�0ѩ ��8�������%c��q��M�ZCkf����f��uPb0bBBK&�(,�Q���1�X����Ddda���(�%�,8$�6�P�Yp�EÃ�7瓘bY&\�������#3,�� ��s̢�l/#-�I�1O�8�6��BL��Npg癎��BY��9��#&:p�Êi�f�Fy�<����Y�3U� �գ2��	��3yEX��a�����6q`��y��6սq6����1������3�7���*q4���*����8�4H�hH04���P�PI43�%BԘ��DK��g
 ��:_lѷ��l�bcq&�Htm��%�d�,�,�"\"r
@�(Ƃ��Ym#	���@���$�NZ��ap�$�B��J��se�$�T�l�4�(h��3�9v�)RN��k�&��[�1����1@X�q4Qʈ�*�bS 2c�`�24ld�&�Ih|	�HN&���60b�8D(N'����i��#5	xBx��@��0��O�bpt�EY��@�#�����j����N�q�A�(م��ih"�O֚�k�~EV%t�H�s�.�+M�͘�ke�P���e�n��k���9��ʌ�� �#[�Y[�y�¥���u�8g��-o�p3�T��<���qbq2/o���ZB1��0������b�m��~Iǆ<(��Y@h���Jf_�&���6n��Y��X���+�I�&ߚ�6`THa�J$�����D�7������� ���C&gc��a6�$0Mf��mF&��0�n@��A;i ����q�8Uj\4HZ��{�kG���<�ߛ�v�ǰS��z ���>�.&"J� ��,���\$�BC���8T�vi���a4U@@��5�pe�S5S���2����Y�PeQ��\"����G �D&j�E���sTl��� �4QdKa�Yd���ZMNffd��`d�c��� �IA�)�Af�24�8$��٘�H)�6&b�C+�|��J¼ShB�~OD=w�ә�ѱ� Û=�Ѱ8�0��������<6�1�XhHd�!���v�� ��xs�'������x:I�F�Hb��[��	0���7���2ѱ�_�u�B�.	�qԲ�����ھ�@�0��\5��<e�k	��\t�N.'���H8ˡ���.6��Z�kV�&���`A�8�q�p!4�lw�E�%�Di۵�1��h�5���IӢ"�h	 �h���������Dh�DᥜA������9s�Rl�i,Ѥ�֘�h���saĎlѸ�ݸ����������A�xܮ�[��C`h�3Z哢޴��t'e ���S��s<Hbw?~)�@�1U$���w���[Ôw��jz�X�/߇�˹�w)�����}����E[��w�[���k��W{�Y��ej+�?��A����ׯ�dB�)A��	V�;}���(�w�����đ�ߟ���@�X~w���~�?!�ԃ3��<��^/?~���I/�����_�V���[�*���u��n�[~W�w+��Y�u���[��Ù��*)�3R��.r�����_�S�ݨ������/�~��y<�?x]�G��qx�g���1����q�e$�:���9��Q�����s�{���q�jlx�@�m�;�#`F!HtI���f�f�5p��v����x��L<=���h��\��zD�#����B#2ѿ9]Pޭ��%��`�ֵ?�1���̳*�aA����8ٻW�H�~<
^�;_6h�4:(����h�͎��Y &��3���I�3A��vp�qc�gChK��!���k���lۧ.����h�l�ddY��tZ-���ĒM� ����N @ä,��+~�\����#i�Z�FBaq�~���Cf���5)�a�ˇ����գ�cm5�ښ�p�Q��!>���⟪&���Lu��+[Ӌ��Ӏh��n��1�i"�<��-<K��E~,U��Cr.�D�h��0� &��Z~�^�>~ �dxΉ��Ĕ�ө&�p�X �;6s&��9Ġ֭qH�1�,���բ��јe�<��[j���
���xy_�Lw��iR��x����7�;�{��'ǥw#iӬ��?)KI5f��Ѕ$��Fh-61���I��jq������8D�8&��}?>�����1��8��K�2Ag�����y~y��9�$'v�.�2&�)	O)��:0I\���LM���gA��>?�<#;8��,�:a��<<���h�����|g)Ѵx�����ѳ��x~<<K$#�7�K��=<߾	���p�Cg���PBBrd�8�9�hه�t���x��b�IŇĜ]1C�=��k{���$/����?��Tf�]��!��w͞���0l%19����pќ81w',��ߓ��5���f�ى�r
��aa� ���?k�j:mV\Q�ȫ@mq9j9ß��NV��4d�>[6p,4m��# 6�vfZ�VS:5Y��#4l���9�i��#a�d�#��(�U�Il6���W���7�   l �      �    [@        ��� �  �H�[j�    �pm�� sl�Ŗm q�#��]5�m[6�d��(�4*�X��T�UKʄŠ+�-�m�8�@ H �� �M�l���`p�h ��p ��^Kl���UPUVҒ��-UYI�em��=��a�mW�����mmm���	 [@ �l)A�g����  p 8[@   -� u�m���E��@4�vi%��m�uR��y�,��-MV�mI6�^�H�k p�-�i��V��  m�$��Am 8�f�j�!mH�VV��Xr���UYV�����	��c��j���'j�]��R�U^Xy���l$�U�����K��UT�U|_��O�1<��1�8४�=k��6,�l�G�Y%�X뜁PU�D@[N8D^dZ+Zi �[D��[R-���+Ŵ�|
��)��y��]F�m�^���^�m��0
�ZE{tʨ�WJ�]��<n\�	�ZU��U71��!���F�B�nݹ�ړ�h$ � ۫m�i  8[E�H��i m��Xր� �cEpɶյWJ�ʽU[/7��5�Kp �UR�@E� I"���[u�v-�  �a��    IÀH��	���ݭ� Q\P�/*��;ll�[v�����@l �i$�m�� �o���    �[[`-��&�\� ��X%����\&��[v�m�H���m� <T�0�ڶ�WF�7J�E�)��Pd�*��g��|zmU�\�vuJ�&Fڬ��UT�Ҳ�Fs+n-�2hٲS�i[v�[�6��S�h�P�6��ɺd�ڐ  Ѡ݉��L�PRp UuT�JAm�h�     m� �-�  m  
ksm�i��[@H ��*ꫫ��f��V�-�h  p �� 	�R@Y��msl�l  �p8    @ �` p�� [@  	��     -��]    kn��Am-� ŵ,� �`�� �	�6���i.k��  � H   ��@$�    k��H6� $@    -�  �� [@��m� �  �6崶��im  �mm���p�\�6�m�  �h  ml]���U*Ԥ������I��`s%̕On�K�e_7[�[<e��y��s��F7]8�26����s����,�΍ˉ""�9Z��PO�#�ga������hN�P����/kY}=V�J4��rC	M<�yہ*�C�G67;1��V���A�|!��]����v�[sY.�d6=���u�] �.�P�j Mİ�I�CNu���A�z0�.՚��U.6���-�+R\ݱ6� H mm��g ��6��r��-6�a�ȗ([d�c�X>O�����qje]YQ�)&V���3vN%UU�i����
��j�C���A�6� p  �`�
v�m�J� ][Qm   $[V� $ �hh�V�sm& Hm۶-�m� m�m�9��f���` �> �aͳ���[m��   $ �� [@m���$�I��		-�m���� m� 9���mmŴ$�bY@ � ݶ ��I4��:�����V�X.vUz�(
�.��u
�P�+��p++�1$����oQmm�M��l��`�rgXj�6I�ϾH|�cm�vu�ā 	�M���ӣ�� [V��`-�$d��`�m�.t��-$�m��ʽ�@7���cLUU�[@m�����h�5頊�T�D��l� 6���,�n�0 ��z�j�@�Z��V ��+AmcY7Rj�p��L���Nri[�D���9F��n4���I����}�n��O$������ �7W&�3��j��T�*�խ�t��  [I$RȐt�Amsm�j�W�8:�5\��^�%$[x��m�6ͳk���+g\J�U�v��� �l��M+U�sZm� b�-�ymp��,���v���n���@m�m �:݁�Hq 6�ޗ��H���  l����I�H떨 m�m&mf���V$ċo	 �u�:��*�ٺ�eNRT&���6M���x������ ��շ��u�=$\Զ��I2�pm�kMUUR���6%XH�	�ٷd�Ip�6V��p#ku<��HMJ�(9��ʩ-ʵ@UAg����a�l��@!���H�Y0 m�1�� *��UUYF��m�ݦ	-� Id��M� m�4݃ZŴ�U]0 �����}�m��̳:\� ��  &�*ڂ��RviW�sJ�ր:���m�� H $��Kn�����~6ϭ-� �i�ݬ�m� jm%��` �lmU�f�Kn��� �.�8[C�  6���[F�9�lm��� ��   �}�}��5�m&��    [@Бa� kd��Ў3t4�p�` �@6�P�^�
(�4UT��m���n�[@ $ �P  ��M��k�-� l �H$6���r��À�9�@  �\  m��t��^�f�Y}k(�;m�J ���lp�j��9m�`��4���yU�q��m�m�� 6�  m�u��$�� ��,6-�  5V�8m���a��6�m�n�d������ZU^f8��[pb�U���ǎ H���V�I����eW��u��i��u�Q�n���UC�*�Y�V��$�7naxk���ln5S�v��(7d��h+i��.�C�S���n�s�@<A���zS$ m�~/m���[D�o8[:S�Uu*��HMm@Q�r�l�u����X���HM� ���� 6C8    �^�X��U+ϥZ���+�l�����mm���ed%V��Gt:��.hn���Pn^��  �WG*n����m�� $���v��s�;v��ko[KM�u�0�m ��kZ��v�ҫ��;];H &Mk� mUdl�ʁ��WʩS�1q����j�`h���mG�[E����v���B��T�Sd^{&�9�Z.]ٔg`kT�G!�;&,b�H��6a�8��t���zJq\&��(6�5W�@���$,֭`UZ���[�SR[��vV�ٓ�,v-� m����s��n��"��` �  � �� I����`	���H[�t�d��n 	Lի�ّ$� ��Ӏ��qĉ "]n@Ԁpm�i6�@  �D�6۵kl�J�+*���U&z j�A��[�i}Z�i ��ta&۴�������F�ۃ��v p[m�d��H$}>���� ���Sl��/ivJVV�U��WJ�����/Z�@ H◠�T
��\M�KUyVt�m�� 4�nհ���j�i   6�[p8[@�m��]jg5��۶�t�p��
� ��mm6�m�m�>��ؐ �` �m� �����[�@   i�wL, ��Ӎ�����oRD�޷�.ۘ6�[p���b&�V|6Z��m��m�5�'��� -�6�r�m�h 8 6Zh���� m����
]��I�L䁶ŴR.��$�u�����F�  6�����	�{]5�o   �d�k]zf 	�kwM��\̷El�� "��3�&e�w��lcku[ ���_]�  m� ���^���h    ��\դ�HHj�8A�Ί��
�&�dsr��[,�
ZL�V��  l�YT)\�mAq�үm��@I��ڜa�`m:�U{g=R�T�T�n��kmٶ�[sm��Z� ��T6 �]�����	+�A�m�-��a�� �-� � �k���Cv݅���@ڶ     ����sK����Y4W<-�ll6�  H�6� | �� imP����.�;q�J�P\ @ -�  ���oZ�oP6u��[I�������۳�� H���\�������U���m�gn��m����Zַ��{ٽ�o_�����QO�X_��� ?�����< �*+"�LQ���!D1 ���O? ��`Q4���x�	�� �	+�=�~C�H#�E��&�S��'���G��)�O� x*�V�(�Ut�Ș*#�qx�������"z�A0ECG�
���P:�#�G� C��z�~ �!� �� �`�H��D
�Gi�� =DE��PM���<ބt��t�6����P@!���QU 4 �A���V	 �&$Y*M"�Pb��"��_V|A�pv��}E����� p pL4�)�x"z�P*�~G�<qu��v�iD��)TA,)�� �W��=q��� '� �]����a�CNfRVfUFA�qMx uT�;��M� �	�Q�A?!���U���EG�/�+��_S�G�O��� E��Q %����w������V���������� ���6��V�����m�4�m<��܁i�IJ�3j2�F�]�1W 5R��x%�^݊�
���azsN��m]rfjWQh-�粫W`0Ɍ3,i�@=���������˭��;-�����.P .�)�L��ĬK+r�UL�km�p��	a�s<�\�,ʧ�tJf��x��b�xt��W\�s�֫��j�5���-Sڗ'4N�b�k��2/,9�rl ��� ����v�� �un,4�^+m�e��eLR�q�m��v�F�:P�]�2�&w$�R��Jvmf�������:q��n�Cp�S֎���-�$��"�2U	��[uR���Gr-�K��n�m]��;:a��8p�(�8��Y��c9n���dޜ��I��-�$��Ô�5�+������-���+�Y�ء�a`.+���Kd�z+q2���:��
̛%ʵ�(�۶S-��d�2�!�q͙xZۃa\�3����m��C�}� �<;i�v�t�#q�:��Xm8;i�I�n�u݈m�I�N��mز�ɰ]�)nyV��yܼ���F½<�P�&����Wk�8����6�*^@f�u��@⭪U�TÎ$��EȘ��'$�C���^�%��tkl�@8�θ��=�vl&�9]M�.br�g[�k�
 �]YUWuԪ�'f�!M�ۙy����Uv��YAɞ1��;s�X�m��F�s�֡�'�n��#Z��H��ʁ	nM�*�G�+�9FΟ ����:��'����T��L�,��lBmgF-���2��m�;r�%�U��UOF<yjGSskv �;q��c`�Xv�r��kv �WM�˶An�ҵ�∗��v�j��<u{e^������m��a�*U����'[5	r�*�GfӲ�VQ���#c�R��7A�z�V��]&�z;NY��Y�ff��LC�A}�F�.
�H�O�}_�@8"p�Q� �IM�J�J� � Y�'.@w-\J Z'j�P8Z r�]����M���ܝ���i�k!�(�]�1H�<m�2q��U���Z��B���y؎a����u�\Tx���{zT�ns>6�MS6NK5ȸ8�=��KR��6^�m�z�Q�:5n��j�#O	��t0���O�>Ԯ֮5�ޜV�kV�_;BfP73k�o=�ٙ�oB��Tq�#�V�U�AL{p숯l��<vp�!��9�<��ȁ�Xt��h�Ih絠w���s��v���w��ȜBpN4ۋ@�f��J���*���vN0ޜ`��uh�K�HF4�LI�hwJh����>�@�e4���<�9���L��� :��@G6=��+?b����w��Rd�q9����-� :��� =�l2���ֺ��6'�V�]�v{65���r�S�+��R��ɶ�c���a��h������׎Z�s��oU�f�kY��ʼ������U:��?Q^��
	�W;���W{�{�����:���I��E�G!�^���r�͂ �sP�&ݘm'�Ĝ49�Z�)�wY�^�����"q	ĜI��z� =UU�U_�M@G6�r���.��u�s�A��^�V����b*ڃ��8�;�	�ہ���r7@����#�R��s`���d��i̊'&��/[��yϪ�/YM ��y��~��z��&I 6l����ʿ{�{�����r؀�Q��B�2�#,�((~莑s�/{�7ʻ�{Õu[��@L��dx!8�l��y�f�m������z�"��s� �5$��x�$������)ś6��q0�][3�̃4�v6�ms[��P9(��;�yr�o{����ת�F���I�}�ۚ����)�wY�uvĆE"K#s0rf��>�yU6wt� <��n���<�e�����N$܋@��h��h�?fbV۹�{Ϫ�xK�&5NAD�njI :��Au���U���&�E�G΀~�o��W���v�-i̊'&��-�s@�U�[e4��4̥s$r'�Ĥ	Ȝa�mBS�l�h�&�%\�q��h�����9�US�s�I�H	������Z�S@<�ݟRI/�;��`����Q\�KE��h	&� u��	$T���-�vdX�0BNcbp�<��h۹�yϪ�-��[�I?�����A�ʹ$� <��@I6�r�]�!�B##s0rf��>�@��8��{� ��ŀyI%�"j��J�ֲ<kgb��8��j5ͺ����
��E��h�C([���z��f�bTxa��8��-Ͷ�r�n-7F�W�t�v��`}L�+��֥�#vN~��k�_}ʂ^t��R"��[��'��H�C��݌�;-��÷^]7� �p<n�6����k$��k��\MÞ���n.��/8H-O�:z��=w(�v��}��|7_9��j՛6W/l=�4����Ƶ�v��ӹ:[��ܓ7+5�C�C�7"�;�~Z����n翳��h���9�D��Dp�<�r�ȩ=6��/�!v�'2(�I��z���e4�S@����v�b�sɃ�I��� #�x�ʪ��� $u{�2dq�0#n�����:���e4�߫����46ڙ0���L7�CrL�vG�X��d3�]��-�%���0����H����@���/�S@�e4{�3/�'�5ۏ�w���9���u	"t�T�R�.�OL�_k�5��y*�?{{��ȜB�����[e4�S@��^�z����`��N$���4>�r��/����ȩ� 	=m�ڸ����(�x�7o 䲕W���@��4�S@=�mQ���'0`��֚�'72�Y��lu�^��5�8,�Ż5A�0��,GQD�B�����/t��z�h{k�;=v�b�sȉrE�o��3�*I6v�� ��u����/�ʀ�$S6�^��r����\�*+��>��k�T_DS����*����ʿw]�1�bX���N^����h�S@�e4{�e�$�F��ʹr*@F���=�Z��>��fҸ�<Z��q�tf{g��&�^��X�[S[
�����{���>_>!��������M���/�ՠ^�s@��&D��8�7���7��x��� ���3�&ø�+�dMě���~Z�w4/Jh�����tK�)M8�R-�~��J������t� �vi���Z�W��8!*(����ʼ;���3{5�l�#�f���M���;��h�ߝ�m�?�Cc��\uə�x*�u��p���v=��GE��x���'�B��6����Э��� ��@G"�gJh�]��0�KsI�@�_U�T���U]��ذ{����L}�!������cn-�����4�S@�{k�=]�!�c�dr��4y�͂��1�*�q��@vtv	�2bq'��z�h/mz��� ��f�U*T��51�}NM���n8܅#�9lm��u�]��ְ���-��8���A��ݐ��9;F�F��3�x���Vͳ˽�nV�\y�W��)A�;Wmx�+�����}���kZ;^�U�8�ݫd�y�v�#lH.E�x�V�/m[��v��+%-���1S��H���#y��B��Ⓩaf��Gz�������N�Klڝ;��ӆ�vu*�^"�pÙ��[ݣ3f����p�{*ҝ6 ��
�u)�S�^�,BU�E�����5ndj8z^�=�������z�h��D�y"��ӈ7wȩ�=�9�@v�&%�W;=v�b���#�f��e4��0���~?{� ��ŀ~z��Z�\827���<^����h�Қ���aX�$�<i8h/m��\�}�k�77�� d�m��Ӫ�&�����nj�Q�Wa�a��D�Ʃ]١sW{��:�W���Z~`�EHy�͂��x�c�9�G!�rf���M���d'YM�}V�z����`�&'�ff��� ��Z6��9 =&�U\�w1��r�z�������4�S@��:%���&�n��o���T���������}�6�����c��v��]�F���4���ΛNU�`C��ɫ-�y��Y9k�D'G$��Jh���ץ�Az����J%��L�,7�� {r*@8�7�^KM�Wm�0w�ŀo����JUU\*��XY��`�!�S��0* Ɗ�$���]�4����h	�Q����&��},pK/�1��x�pD7��E�?vQ΅x�_҆�߀8k����*	'� x-��~Q_�L_�;P�%^�Q�o�{��((y��~��<E�;v"��Q	(R�,ʪ���{�,{g�UI~a�ӌ?*�J�����v�u�+��5.AuR�Hs1~{g�RI��og��UM�ob�;{�r���Ԓ_pp��]�e�ww.�,��7E�Ka��a�%Y�u�Yt�d�n??}�佢��]�e�<�I���|`�]�ߗ�;{�}T�?�����U?���W�Yr�܅��wobϩ/����ϻ�a���$���oN9R���}V���_1��.E��U*�w�~X꤫�s��v���T�v�,W��6���F;�:�,���ݳ��;zq�~��ϯ+G��!���|#�4��� ,����O�Xr�4m�q�h%�� �l�M�9 =絠?7���!�B]������å��V�WQ<�EJfs�Zp�k��r9�`�nPa �Ih�T���͂�E�Y2E?(�0iǠ^�sO���v�����<ʟl��p�&��H�۳��M��8�?Uw�����rI6z�U�g8D�7wWw�Iv�q����IS}�ذݜrI~aϞ�_U�.�Yd�`~���������̯���r�>����_� {���{ݿ������\��De�3r��#�;n�K�y�lavM�:������S�bj�Z܇��v�^vx��h:�ܽ�2��<�α�ڌ�Q�/�([������qF��cv���eޞ+#�NvξI�[�e�h���be�qv���q��V's����B��<��M���W��>��K����.�Y��[��2c&��z�#%��btݹ�F�A�܀��^R�ʩR������I(L��Ml��1=L�1�,[�ё�m�7a�����7���m��S6����?~�I*��?,�g��R��;zq��*T��{;���p�r+����.G"�I%I��goN9%_�ol� ��Šr�n��8$��r9���:���z���JhqeƘ� �R��u�M���^��/YM��,�����8h���:���z�hzS@�:��p�O+f��D�r\M5v�ml.ct�@�o'<-�G��!�2b�����4�)�^٦��4�U~a�݋ 纭�9�'!�oN��ܫ��}���&��Q֫������ץ4
��c��b�n1��@�Қ�w4�3?%~��@��>4뮉��6��p�/[��q�͂ǰ@:�H]���c�'G$��Jh���ץ4�wʕWi�y�wj9`�Q�we���aIn���vH�ջm�֎ʌ��/�W%�]����7��C�>�O��Jh���:����W���JA�I�@q�ȩ �� #����,�����f4�^�s@�ҚO~��i*�uK�%Uy3f���L��2ʙ1dr��4=]n�^��^��<�w4
���eP�����ۆ���W9�߾����R7�@vaN[K��9�quֆ����b*ځ����;��;�������E��o�'�K@vH�� {�L��&H�q5��@�۹��٦��Қ�ڴs�h�)1�D8��J@F���=�Z�EH	~��K�rb�#��;�S@��V��{����z"z ���oϮU���ici}��x��_]�@���o���M��M�{�T�&I$I���g(����f�'�lޤĈ�ɪ9������Y1�~nLcMŠyz�h�S@�zS@��V����Xʙ1dnfAI��� ��	���*@z۬Xʡ1H���4��4�i?b^^���S@�ʣ��i�G�Ih� #{UU���?����&�I)��빠^�D�� '�K@NW(�2�]�F��V2q���4���;�8���9��-��:�m����{i� �N�\��r��h����d�	�m�����d�cbu]v�I6���m��\�:F\*U��pb��r�*���gqh�<��cd�6�O�5��!��=`�9sE�k�a#��m�1�u���;+S�l.{��ɷnƛ���|���:)��\y���z\��O�����_D8e�.HHB.��]3���r���nxٺL^�:q���ϑ$�2[�����s8~�{Қ�ڿ�U����ŀw��6Ӹ;�9h.I!�?=�{$�����{)�m)�sI�@��V��۹�^�M�Қ�n�K"O�Ɍi��9$����`�8�<�f��I�׀z��2�sQ��'�Jhl��}v������W		�D��.Jg��b���xp�5�Rr:�n��h��8�K��5���q~m�@�e4�hm��/t��˗#��5nA�[�Wk��|���j
�v�hD�T�>I%KԒR���� �͜`��o����j�&H�q4�IH��q`�L9Ro{���� �Ǻ7�Lm�!�f���M���=�4��{�ߖ��sm9������� �� =� 䊐�`�����}�VÒ�]�'he�n��g�<:Ŧc�!�ev�0����=��k��NP� ݙw�tG�@9"��� ��n�K"O��?H�4��o߳?bE�Ɓ~�|hޔ�=��,dX���c�`��L�٦RT�)*[Mfci�����h��Xȡ1I���3DUUm��� =&� �6.\�w��I�G�Қ[)�w�S@�e4����L�;^�W-B���#��U��^-���3=��-٫%'�~��kQ�!Q��p����@�l����hޔ��Z%�Lm�jI�6i���Uvot� �o��l���#犯$�I�8
 ��N0��^UWԮ����t��?x{5[Wm�6�����S�gs�7�\����ܮ(���
T�	��Q�B`�B	�!Xa(H!_�!��pYt�����N�#������*���F�Ӓ�Ȭ�w��� �Z��.��o��@��V�紨�"q��'fۉz�q]	=��z�	�W���.��m�۱lT�uŠj�j��c�~�g��� �/u���_UW���� ���欎9ܻ�`��L�RT�ʩ+��x����7�f�ʕ&�z����+q��;� �o������U�R_����i�w�����ZY!��N$܏�*O}���ݜ`m����U*��>��s�ӑ]�q�����٦ʕW�7��;��x�n��1]RI�IF�B!	fR�=]Ê��2 I*MH�	*��P��P��Ғ2E�+ �C)!K,���"��P"$pH	Haa��TĈc	���&	
���B��d�XI�1tI$IK�!"���C) -n_;���*'�"h�� �	d ���d��XP�M3*~Op�b<݀�)8X$���)�I����C5�6Jl ��77�Ÿi�D�h֍i,�b�EfF��tPf��[���l8{b���H`�l6a��J�>t� 	HfH %Y�	�O�=�㧺{�ӧ{���>N6�H���B��l�٩m��P�ԛiű��ې�f`-�������)M��r2�������Pj�\n9ݟ\��ڞY��5T�ks=3�Z�n.��iv3H�B�v�T4Z�u�fᤜ�J�;\��̫��]��Wm$��m ��P2��kg�m`�`+�:�mGGN�Fy��s]U]9��M����*���ٵ`1�v�.�vlŻvP��h���̿>OG;�L8C�v8����e��j55˃	=,]M���jU���@�']4:8�����Y2]d��m�s���UWn�e8*��ء=�D�;S�7m�n�tk�Z��d6J��;j�d;�g�^f����"W���Z�)�u�+��6�-<dڻ�C���kW%2�DQ#��Hީ�S��۞��[kЯnݺ����r�x+�mv�qtïe�q���ݏj��u=��6�v�ք����m�V|�Y��2����m<�����d�kvn���v��"Fϻcc7h-�p�;���M4�a�N]f6�^5��Q8{p�u:��Q�؞F�����)��Y��K�ۢKl���˥����bt��H�;+������3�!a����v@g�u�mq ]R҂�����+F�Y��$�5sr;̀dN���m��%��6�U��b��w�nqsє�K�ŵlm�ݳd�Z�U��5�� �dtQ.��[�y��6��:m�`~EpQ.[���'Wm�w8k�ǰ��m�2�n� 賟hR٤$V|L�/E����!�"8��ݷ'�K�*�N`6�A��뙞T-�S�Ղ����ZظM��S�(�$
�K<5T���ef:[��Pl!���Ŕm &��L�e݀[`��#�v�� �+�vn�y��|��_!y��&zU�R�e��.��Zy��;�r�<�+�:�k�.�UeL�<kd ne,�k;�� s��{m����*ͦ�'.��"��A��'��#�
"¼@�=Q8�=�]��,�u�t���2�s�������v����9�9�^���v.6%��z��n̪�ěd�(n�Ca�;\�s���ym=�d��ӌqֺ���;UMp��[f�ܺ5�m��hޏ$;r�pI�Xt]�\۴���m��:p,��훱V#/e���g���Eۗ�FC�&ք6��p�U�{m�-�7l������zs�hݝh�M����T�,W<�";T1Z�����<�����u\]W(�m��nlU�U����H��K��$�����o���|��ʪ���8�<���5m���-;�����*�U��$��UR�}� ���~��T�����WNJw�wq��v,}�i�U*M�׿-�|�jH�Y b�f6����T�n��{� �}�`rI�ߖ�w�&)1�����g�r��*)/z��w�ذ|٦ ~���Mv���Z�㛐�M��͇H8��]uY�+�-��`��S~��>'�s���Q��@M�@OH� �6��@?M�m�.8˹wwp�7��Y�I:��[H�UU~�K��ϧ����<��i�*U��}ϾNEwde�\���;~��ߺ���T�U]��s�<��X�h�b�dlMI4��hޔ�<�q`}UO}�� �N�cVېm��������*@?M����sפֿfZ�'v��4��nj�IU�X1̜��Ǧ*�j��XnAۊ���|�EH���_j����	�%�:ԑ
�@���NL�/t���>� �/u���ŝIU&�z��j�Ԉ��,m�@���@��V�>����7_�}��}z|h�UF9�cQ'$Q8�	��r*@F�=W&�@~��,��(�q$�Zs��f~�톁��h�j�<^�X�cQ�s�՘*���ԋ�\�ۗ8ٶ�+��b��[��q�NEwde�\�C�~I&*J�w>� �999?w�}pA�rrr~�}�A|������>� �998*J����\NH�nIp�IW�RNBBB���\|�S!!!�w����A�A�A�A��}���A�A�A�A����$�A�A�A���}�V�fk[ݙ���|�������g!!!!����!$!!���\|������>� �999=��xk3Tf���ֵ��!!%�$SP������������������� �999?w�}pA�rr6����A�|����� � � � ��3-_a�ћ������� � � � �������������B���\BBBB�w���|�������|�������.k����HBE��/2PT��j6fBB2-c���r���>�����{l�w������������~��!!!!�w����A�A�A�A��}���A�A�A�A����!!!!���}��ƶk-淭�[��>BBBB��ﳂ�?ʂH��P��������!!!!���pA�rrr~������!LT�1RT�IV���1H+��n�m�y��A�A�A�Aϻ��8 �999?w����� � � � �߹���A�A�A�A����pA�rrrs����C�Yq�#�X�*�*J��*��A����!!!!��Ϯ>BBBB��ﳂ�����+���~�ǂ��������߮�>�{3{�oY���z���A�A�A�A��s��������}���8 �9999�~�g!!!!���\|�����Q{���"k���ʳY�oY�Y�s�m�זWc�-��3�ܭ�ۣ��h�9W(`�rr�犭ݹӥݣk�܄[�),������l����uq����M�wmt�4F��nw`�Zx�;bf��}�h�s�ZP�gJ�ژ&�����W-���:�ڮ6ݹڵ]��nI��1�����I��єDƥ�����㰻!��"�N_3Z�h�ѳs"u`��c6�n-(�� ��x��Z���e����kv.
ݧWm)u]�&\7"���숕Is�5���~�HfL��m�7r�wT�|*J� � � ��o����A�A�A�A��}���A�A�A�A���� � �:���￹�pA�rrrs￿�k5����[ۭk[�>BBBB���>H�H��P�������� � ���`�%	BP����(JY�P�%	Bg�?�pJ��(O3�(J��`�%	BP����(JY�P�%	B}�>�<�J��(OقP�%	H����(JY�P�%	Bk0J��(N�s2����l5f��8%	BP�'��P�%	Bk0J��(Mf	BP�%	��(J��>�|���(J��?f	BP�%	��(J��5�%	BP�&��(J��>�ָ%	BP�'��P�%	Bk0J�(JY�P�%	Bk0J��(O��~מ	BP�%	�0J��(Mf	BP�%	��(J��5�%	BP�'�k���(╔�I���܈Y�Yq�ַq<�$�����}i9&I�d�{���'�d�&I��x�rL� �YK�q���I��K����\V�\r�\.��I��K|��)~)2��#�'��O$�2L����\O$�2L��w�I�2L�$�����ں�Vsd3g�%���a{!6[�m7j}/]������J��ݏ��i�!6���2d�&I����q9&I�d���v�y&I�d������MI�d���������L��L���"�c��%�brL�$�<��v�y!�Τԙ'����rL�$�>��}q<�$�2Sݽ���Ҳ�)oM��E��Ǽ������y&I�d�_o�I�2L�$����2L�$��]ى�2L�2���i���I��K�Mȭ�����m���)2�)o��e/�&Rbd���19&I�d���v�y&I�\����],)2�)2�����؝�;��w����L��Ov�'K
Y&I�w�yۉ�&I�v��i9&I�d���v�y&I�d���{]ݯe�"VY�e��ÉĳOm�6��kWkH9��8�tZ��շ����I�d���v�y&I�d����NI�d�'w���I�d�&w���NT�I��K͛�����%���e/�d�&Iۻ��|�N�ԙ'��Ϯ'�d�&I�}��brL�$�;﹦R�Re&Re-���Wq[	q˹��NI�d�'���'�d�&I��d�]�ԎI�;�9ۉ�&I�v�}���$�2O{�5��kur��ww"�_�L��L��obt��$�2Ow���I�d�'nﶓ�d�&I���É�&I�e�;�0��5r�mے�N��I��K�74�_��2L��w�I�2L�$����2L�$��]ى�2L�$���s�Խ��@voJ��5��❋9���حh�qK��y7S�C=�[j�b����L�$�;w}���$�2N��;q<�$�2L�uݘ��$�2N��;e/�&Re&R��o-�m���,n��&I�w�yۉ�&I�g{����&I�w�yۉ�&I�v��],)rT�Ҳ�)?y�n�N�N��W���'�d�&I�}��brL�$�;����L�$�}׽ͧ$�2L��ni���I��K}���ڐ�5o[ى�2L��R}�����L�$�{���NI�d�'w���I�d ~׊�WE�7���f'$�2L����ȅ��%���e/�&Re&R�gm'$�2L��}��2L�$��]ى�2L�$��yۉ�&I�|�ߝ�~�.V�ma棒�.�f)�t;�y٥�)6O\s�p��ŦƖ76c.�ַ��O$�2L��~���2L�$��]ى�2L�$���2L�/�K(�f��������2O�B6��ַ���&I�g{����&I�w�yۉ�&I�v��i9&I�d���|8�I�MI�e�}��f�XIn[v仃��&Re&R�{8�_�LL�!�^�6��'�cRjO~��O$�2L�=�Z���&I�~��5�3��b*m�����{��7{���^�d�&I���É�&I�g��]�9&I�d���;q<�$�2O���5��� ۸���r��I��K��,��&I�g��]�9&I�d���;q<�$�2u�si�2L�$�SG�ws�v��۾��<�%^���8�5Ԫ�IxH�a��[v��[W�'8�e���G;�R�4i5P��;|�ѕ�pq�^�\�f�\x��Cn�8��M���H:�JtG ���hO�lnu�xg
��ԙ�pq�z9H���i�9�@2��u����t��v�����ֵ�H���/�9z[Xۛ����!uN�Om�<�t Nm�T���������%�S��y�QZ��O-�39@��+�fٙG����ޤ%A�g�+qqɑ'i��m���|�}��&I�}��c�d�&I�}�n'�d�&C��m9&I�d���v�y&^�{�����5�ۊ�W�w��7��$���2L�$����y��2L��~���2L�$���щ�0��L����B�Ԉ�ˍ]�2�ⓓ$�;w}���$�2N��;q<�$�2N�;��d�&I�}�n'�f��ow���76���bY����ę&I���n'�d�&I��x�rL�$�;����L�$�;w}���7���{�>ߋ��^kJ0o����2L������&I�w�yۉ�&I�v��i9&I�d���v�y&^�{�������o���O9tdh-�ͦE⶞���:8匧�������n�7���m�Cfӑ\��\��:^�I��K����y&I�d����NI�d�'���'�d�&I��x�rL�$�?{w9���N\de�%�)~)2�)2��6�rMI�2O��|8�I�d�&w��lNI�d�'����O$�2L���ϧ�ÌVn ���oq���?w��q<�$�2L�uݘ��$�2Ow���I�d�'nﶓ�d�&�����v�Ԓ��_�L��LL�u�؜�$�2Ow���I�d�'nﶓ�d�&I���É�&I�/tz6�j��4K�:XRe&R�=��v�y&I�d����NI�d�'���'�d�&I��d�<oq����７El�(.��kش����S��vsmK���f�U�5�a�4^:kxkZ���L�$�;w}���$�2O���O$�2L�;�wf�y&�L��[�gK�I��I���_1\�l%�.���aI��I���w��_�NL�$��]ى�2L�$��yۉ�&I�v��i9'�kRd��}־˫�iF����oq����~����I�d�'����O$ɐ����2H��)� �� � ��!����z"y��u��k1����z��!�SXFI����|�v-!��� �Oј��$mj`:TC�_ w�J��mګ�
"m�E�%@=} p0�*?�x z{��=�߶��d�)��n�唿�I��I�=Ѵ�CW,�ݹ.D�aI��I���sL����NL��w�I�2L�$����2L)2�ݽ��)2�){��5����o+f�{޷q<�$�2N��m'$�2L�����O$�2L�;�wf'$�2L�����O$�2L��e�un����X��fp�$7$�-�=6�t%I�] �vul��r��*�Y�|��$�;�����L�$�;��NI�d�'}����I�d�'nﶓ�2�)2��_���;�7n]]��R�Rrd�'{���2L�$���2L�$����rL�$�;�����L��{�������5ƚ���{�L�$���2L�$����rL��Ԛ��~���2L�$Ͼ��10��L��^l�Q�#WF\i��)y&I�d����NI�d�'w���I�d�'{���2L��ړ���K�I��I��߷�Wq[	q˹{���$�2N��;q<�$�2N�;��d�&I�}�n'�d�&Iۻ��aI��I���鵰��vG�[S�S�{O�e�z�Gc"%�g��4檩cuy�+A6���oq����}��v'$�2L�����O$�2L��w�I�2L�$����2L�$��u�8��RH%-�w��7���{��~|���L�$�;w}���$�2N��;q<�$�2L�uݘ��$�2O{z�[iȜ��+rK�R�Re&Re-;��NI�d�'w���I�d�'{���2L�$���2L�$�~}�@�+
� V}�7���~��ۻR}��}q<�$�2O�ϸ�rL�$�;����L�$�;w}���$�I����؝蛷.���)~)2�)9;��NI�d�'}����I�d�'nﶓ�d�&I���n'�d�&I���n+ R�X�7M�{}=�麝�+�m��󲛚ȵ�AZ�iL�R�q�x��:���|>|WfY�"JK$T�[��Y)���㤺݂o'd�\=�{,��Gk*f��s	ʶqwn���X�i�
dt�3V��F@��I���t�<�mr�pgn͠�v���4f;y�jD�ljx=ͧ�P���rlYf��w��j|�ʱ�@uܶ���ݛ��������|ڥg� m�m�Zݸ��^�Bcf�s����ٯ7g��Ҕ��.&�J�Jt���L��_����2L�$����rL�$�;�����L�$�;��NI�d�'��6Ց��#.4�ᔿ�I��KM�ZrL�$�;�����L�$�;��NI�d�'}����I�d�'u��pWq[	q˹p�XRe&Re-�sLO$�2L������&I�y�yۉ�&I�v��i9&I�d��ߺ�ë�iZ	��w�{��7������ǎI�d�'�����I�d�'nﶓ�d�&I��yۉ�&I�~�۹���2	Mq������ow���ϻ��&I�v��i9&I�d������I�d�'{���2L�$�_���[MQb�WU;R�t���k�g��W�B�ؒ���k�����!Mq<�$�2N��m'$�2L�����2L�$�s�q9&I�d�w�t�_�L��L���rF��;���nKI�2L�$������0�¢2�+��'���<�$���'$�2L���Ϯ'�d�&Iۻ��Re&R~nޖ�D�.�ܙK�I��FI��x�rL�$�<����L�$�;w}���$�2O{�8�I�d����-�S�
��K
L��%I�}�Ӑ�'n분�)?y�ݧ!);'{���2L�$�����ݶ���,��R�Re&Re-6it��$�2O{�8�I�d�'{���2L�$���2L�$��w���I	-u؆�����I�8Z�'Tv�'�2�P�����b�Zm�ɴĳg��x�2L�����'�d�&I��d�&I�}�n'�d�&Iۻ����������uz�V������2L�;�wf'$�2L�����O$�2L��w�I�2L�$�����{��7�����7#@���ݒd�'�����I�d�'nﶓ�d�1��T1PH0=ѹ7&�{��O$�2L�?w]ى�2L��^��Ӹ���+nK�R�Re&&Iۻ��&I�{��v�y&I�d���19&I�d�w�v�y&I��ow����A+
� V}�7���L�����2L�$��]ى�2L�$���2L�$����rL���{�>����[��X���uLinj�I-`����[��pP����M�ټ��kw�2L�$��]ى�2L�$���2L�$����rL��L���K�I��I����A�Jse�{5o[ى�2L�$���2L�$����rL�$�=��;q<�$�2L�uݘ��$�2O��zo[�P$v�e�2��)2�)i�K��&&I�{��v�y&I�d���19&I�d�w�v�y&I�d��w��ռ5��%����&Re&R��sL�����2L�uݘ��$�2O;�;q<�$�8�箹'my�I�2L�$����TJ�M�{���oq���~�c�d�&I�}�n'�d�&Iۻ��&I�{��v�y&I�d�����ߎ�9�V��ȳ=L.�s��v{<sl�z�Q�.�ť
�U�7#@��19&I�d�w�v�y&I�d����NI�d�'���n�~�Rd�#�)2�)okyʹ�'.0�Y�޷q<�$�2N��m'$�2L�����2L�$��]ى�2L�
_���)~)2�)1W��Hݷn���fff�i9&I�d������I�d�&w���NI�d�'�����I�d����.��I��I��om���3v�����L�$�3��vbrL�$�<����L�$�;w}���$�0���K�I��I��V�zJr"�[��brL�$�<����L�$�;w}���$�2O{��O$�2L�;�wf'$�2L����!�}������#\�N�PȸpT�I����-���a.�f��Ux��ӧj�Љ�m�aۙ�<K��x��98��cRnt�q7Uf��s[�鎋F�7Xƹ�7>v�Go<��5qi��gMںŽ�vL��ۭ8�OC��������i)�}�FV��OOD�u�
8�P�pԼKEg�dvҸ��;n����M�H�NJ�7���H�^�zН����1��ᵒ'Rp�"��B�VlK���6YŲ-`J�a�A�tM�Ύm�K9m������2N�����&I�y�}�q<�$�2L�uݘ��$�2O߽�n'�d����}O��:9�=�%�>��oq&I��yۉ�3�5&I�}��brL�$�?}�}q<�$�2N��m'$��7�����������o�����I�g{����&I�y�yۉ�&I�v��i9&I�d������I����{������tWS\{�ovI�d�w�v�y&I�d����NI�d�'���n'�d�&I�����ow���_�p�L@:�|�2d�&Iۻ��&I�y�~�8�I�d�&w���NI�d�'���n'��oq���~��N�C���[���k�iK��uڇ��WQ<�L��k��Q��론�۹c����rK�I��I���w<O$�2L�;�wf'$�2L���yۉ�&I�v��i9&I�d���u�ݱ;��A�G���I��I��ŉ��ؘ��rd���;q<�$�2N��m'$�2L�����2L�*^�~��%9rX��D�aI��I��}�n'�d�&Iۻ��?jMI����q<�$�2L��}��d�Re/|��5dj�\wpN�K�I���'nﶓ�d�&I�����L�$�3��vbrL�$�<��v�y&Hoq��S��Ύ���J՟w��7�$�<�~�8�I�d�&w���NI�d�'����O$�2L��w�I�2x��{��۷߻p��#���ψ���5�i.%s�z�rS����V�
�5�Z����w�2L�$��]ى�2L�$���2L�$����rL�*L��ni���I��K����wr'r7nK�:XRe&Re-���)~)2�I�v��i9&I�d�{��8�I�2�)n��t���L��[���������F\�!���I��KM�],)2��$����2v|�J+��M����NI�d�'߻Ϯ'�d�&^��߿( Fp�q�V}�7���{�<�~�8�I�d�'{���2L�$��yۉ�&I�v��i9&I�aI����n؝Ӗ�1���)2������&I�y����L�$�;w}���$�2O=߽�'�d�&^�l���1���e���i��WhXPᛉ�:y:-z-�צ�g�[q9&I�d�{�;q<�$�2N��m'$�2L�����O$�2L���)�)2�)y{��P�\��Fk[��I�d�'nﶓ�d�&I���n'�d�&I��x�rL�$�[﹦R�Re&Re-����5 Z%ɭk{ݤ�&I�w�yۉ�&I�w��8��$�2N��;q<�$�2V�4�XRe&Re/o����w#Y�n�y&I�d��w�'$�2L�����O$�2L��w�I�2L�� z�r=z����k���3{��7{��}�������ę&I�}�n'�d�&G����>��I�d�'��Ϯ'�d�&I��x�s{��7���������+lIT��11��z�R��Ͷ�j�M�(t�c2i��`8�*$k|�7���{�����r��$�2N��;q<�$�2N�;�弓Rd�'��>��I�d��}�g
� V}�7���{�������O#�gRjL���8��$�2O��}q<�$�2N��m'$�2L�?W�{m�t�d.��)~)2�)2��;��d�&I�}�n'�d��R}}��'$�2L��w߳��&oq�ߎ?6���,��=�7���� ԟ��>��I�d�'����rL�$�<�~�8�I�d�%�5���fR)2�)m�ܣP�\��	���2L�$����rL�$�<�~�8�I�d�&w���NI�d�'����O$�2L�ـ�*̉J'�aYdBIX	!�V	-�:,�@0B�#x(�+HL�b"mRIHT�CA�-��&���������0�c�H@�� ��o�!��ļ]��vp���ohmJPgh�Q=L���? xЃ�~3Vjp6���@�{Z !0��!���R���S�<����#m��[@-�p⁌*Wn-ʨ��v��A��.�6�5@I=:4lbZ�,c��T�՞ �U*�:��6@kn%�^j�� ��l	^��sq�y�L����6�ܻ����'�jQ��:/ �gr��������P�N��W�N�լ;�����j�n�NWh۲�WR
ٶ溪���  �]
˶�]:��������Ů1�"ۤ!Ҋ��,طev�]{Q��d��5�vE���k�Fv�eh
G.���GF��RF���p���̺%��d�EqimkX %�a�\��l1<��u�$q۶�MJj�Α9'Z�w]y^�691׊`BzƜs&����"FAZ��#����u�k	�a���^�]���kT#�42-S�V��:�E��l ������u��[c]v��7N�u������/g����nkmPݸt;+������ ��l �QF���:wt 1.�tv����;l؊����W�v��k<���M ;�R�W w=��ܥ�[�  [�D <�¯'8���
�S�#S��uvJ�qNk����"�댫���C3�=L�n�]�i�u���e6��pͶ�qu9:��rd�F�[=]R�j�A�ݩ���6n3��MM.[d��V��)�'���X$�o&�Q��;"k�ݱ���0�7���lDmb�l'RR���t�C��y����K�ía�����d����*�=K@[7���vuԱЊ�[��lgV���q��p��N�4qcj{���;P=��1ƭ�W\��n��+Fh<�N�G\��O]��@��N��Î+��:��� ��m�i�C�r:���	�0����9iY v�+`h�Ɠ�	[V�N@��I��-�m:GKt�C��&I���+�:��%kQ1��%O$�g�li�-�T	k��t�N�l�URfͰ�̧m���T��Z��Ohf�kF��ޭffk+7��DLS� |q<Q1�6'�S�P;<�^kv_���k7�؄�3�B�ntu�X���� Z:��x���-c�yNzI���NtB�릵� �[ �]��jm�8w<Q<��gK�n��:ѫ<�5�Ӯ�]V����]��sm��CnX�؊��,��Ԯ9�qs��px{ n��ygl�uCrsvNucr�.t9본�z�6���E� C[p��RH�$��f�Z4��$���{�q5�XP��p�[��΢J���͝�.��۷h�n8�ی�E�f��{���?djDZr仹!t�)2�)2��7�Q�&I�g{����&I�y����Eo�jL�$��ZNI�d�+o׼ڒ�B]���.K�I��I����vbrL�$�;����L�$�;w}���$�2N��;q<��u�;�n���@����j�=�7��2L����\O$�2L��w�I�2L�$����2L�$�s�q9&O�ow���_�q\T�V���oq�/��R}}ϭ'$�2L��~���2L�$�s�q9&I�|"��]�������L��^�d���ܱ���,�{���$�2N��;q<�$�2N�;��d�&I�}�n'�d�&�٥�)2�){k�V�!$m;�ֹiT�HH�ٶfV�������
Zf��xrK:��9�ym�%�CV�v��xRe,�$����'$�2L�����O$�2L��w�I�2L�$����2C{������u�nVOKx�|��{�2N��;q<��LC��SB�*ϲ{&I�o�I�2L�$��y�q<�$�2N�;��"kRd�����2�ԁr���K�I��I���ŧ$�2L�����O$��D�I�>�>��2L�$�����2L�$�}~��ճ�iZ�������ow���n'�d�&I��x�rL�$�;����L� ��'����rL�$ʖ߯y�%\��wN\2��)2�(�s�q9&I�d}?w�}q?I�d�'����rL�$�;�����L�$����'�v��c\�lA:cM�.��ۗ\�WY�d�����Vr\Nr�/ާ)���ۉ�2L�$���2L�$����rL�$�;�����S�=�rd�R}D�aI��I�������r'&��5��7���&I�v��i9�$�MI�}����y&I�d����f'
L��L����e/�/�Ҳ�){ݒ7�q[�rc��XRe&Re.�����2L�$��]ى�2dC�EB���Mɮ��\O$�2L����n��I��I��ݒ۶Kr�jn�y&I���׿k혜�$�2O��}q<�$�2u�si�2L�$�74�_�L��L��m�����wn5�z��NI�d�'}����I�d�'nﶓ�d�&I���n'�d9&J{��5XRb�*e'舘F���;óA�>ç���4�:���A�p�7Kq��j�A�[2��m�����{��0��{�I��w���C�d9&~��9&C�w�yۃ�I����?X΋\=+rT�w��7��쓿���$�rL�?w]�Rr�!�;����L�$�}׽ޤ�Z��L����Ԋ�Iwv�iˆ*�Rb��$�~���NC�d9'}���>I��ơԟ_o�C�2�!�߹��w�w��7x����~�⺫%a��I��9'}���>I�����Ԝ�$�rN��;p|�!�8/ˊs�E�$�ߵ���I���Z�fp�U�墷�w�w��7x����7�C�d�w���C��&w����&C�}�n'��I�)���ﮭ�]E�k��S8�$e���K�dի�&�u;s[���7"5e�ov��2�!�߹����$�3��w���!�2��;q<�$ȦR�f��
LT�LT�{��m��r�ѻZ�n��&C�d����NG�"0jMC�}����I�}}���r�!�;�����L�$�=׺-+	6��G"٦~G�F~G��n�d9&Iۻ�NC�d9'w��>I��&w����I���"d��nۆ��،��؏�N��9I����v��&C�d����NI��}����C�d9=��O�3��6)�������n{������!�3��v`�L�$�{�����!�;w}�I�rL�$�ꪽ�,�jז��E�v���5�V6��F���ڸq#�W��m֑m�h{9�C�ӭ2��$�k�(Mյ�K�L^��tq���d�nդAtti��n��
�q�kv˗/Zڸ��J�c:\��q.y8���U�9g[�Dq�;%E���@f����Ȗ8틄]�s�6F���fy��,�E���]h�|��-��Ϟj�:����z]�n��յ�w�\ur�vz�b�h�������YV��mȘ����.-�TN�:�ڴ�����d9&I��nNI��}����C�d9'nﶇ�d9&Eo��e/¦Rb�R�f�ӑI!n�k[޷�C�d9'}���>Gʌ�I�}}���r�!�>��}p|�!e&R{��)`�������۽m�"rE.˹�*�Rb�Re-6m��
��I���n�d�'{��r�T��f��R
_��챻cm�c�P�@�D���3�m��I����sOߚJ�+Z�Iy�ȒF��<�i��H�RjI+ݴ�Ē��֤��ݧ�$��ӏ�6��1�sr%���<��
�ӓv�Ɯ-�ۛm�a�x��Q��)��jI+ݴ�Ē��֤��ݧٙ���=�����RIs��D"���27<I%Ϭz�fbI_n��H���$�v��>���!����q�D<�H5$�?O��@?M�h��.9�	~�nԕjB]���p��~�gG�v�� ��z��h��X��"�s��x��� �T��z���� �vlI?�'.�H��˖��8����Ր{8[\���]Z�A��+�*筺xj`8�*�<NG!��Y�_l����b�?fx��gƁ�}�Ĉ�q���!
G�_n��6m�#{��/�\�U~�s0=��m�8�jn�o�O��7�f�|�Y_�V��W�+�ϻ/ ��g�w�D�,m���C��/�ߍ�����)�{l�h�lH�Y 8ۆ6�Uz���w�������)�y�e	g䆇'm'�d���J����']P^�øu�M� �ֲ3�,�KSȜ�7�}�����{�>�|��=��}�?<���Q�@��cϩRM��8�9�����3�IU/��W�6�'#�r��$� ��|`�W�_]�@��b�*��D�9�I��w%�`rO��� �o��n͏��*K��MW$�RC��`�vF�ww ���c��o����W�����gW��/��2s�7LO�u�F�è�]�,�f���..]���uVV��QO�8bmŠ{l�h�S@��g�}����"E6�X�����㘀~�-�6m��\�U/�]����e����wpe�0�����~��䒦���l� �/ݍ��A'�In=�����-��}��}�`}J�*���׀k�z6��RGwwnG�y�6<��{�~�������~��>�T�/`�QS;�EYxƞ�G[,�u�mT���g�ѳ[̉[l=F�:V�(��n�-��#K�M�{�mV��kSl�t$��dQ��1�k���<t� Yzm.Λu{sPbI�a[��F��vg9���k�r� �[�ݷm��X-�5��ٛ���1Y�v9�X�=s�u�'�6�N��4�n�T3�@\8�рz�\�ڲ�4UVӺ23���K��~uH����ejz�]�����m�`s�r��c�ͳ�� ;7K0�E�_l��*�^�޾��?g�w�O��>]�$�9�I�D�$��U�o>T�U6o���{�G�~�f��J�;�ؑndM9!H����m�-�ҚW��:�Q
)�n�qh�,Z��4
�W�����z_������)"�j&G"�<�)�Uz��}V��ŠZD�W��k$\�M������t�-."�{��5g^'EF���{���R۫d���>޼�/�x��c�RT��v�0�ߢC"�I�RD��@�_U���߱`�8����V��o9W�w\�����$U��I��6�I)��}�m�;��\�#�j<�Z͐��f)� �#�h^��*�^��ߺ�>T�ԕ��~�<���N��/j�����ϯ�G�����{M������/�o&5"ndx��E�+u]�tn�ns��Y�q�k+Y���G뼿}�H�ndM9ҎO@�������b�<�)��Y�u�4�(��cmŠ{�͏>�K������L�/�x��	:�X�Q<#�h^����w���]��J��3*2�)(J�ԁ0�I�)K�C,@ �32HCT��OA �Eog񠉃jb.�1����0��<�V����5�Z321�F�����k5�#1��
)K��!,��h��h!�Yi��$�؆� ڠ��(@�o��
b/�&
��=>Y=����y��ޖ-�m���&�pDp���U�s�@G��@?M�hǰ@Oc��dr6�Gr��_���*����E����4��4+�*%�D�6�̒��f|@����n�xڧ=aS�
��,|p��JRRD�O�$���IH����/Jh{�x��- �|����ɑ���E�yzS�H/_��yߖ���b�*��RX��$�d����z����ŠyzS@=��m̉��&�rh+����O��<�)��_���5��������}PS�$��qh��<�)�r�^���נg�
��1��ɎcR�ݝF鵍3t�����=dM�V��zI��o�OaMD�,i����-���4�����/z���'pCp@;rb��1�6y�c��ȤI<�ȓq�/mz���>K�ύ�~�����?<r4ڈ$��W*��������1�\{>��||%���J8�I����M�?U%K�����{� ���^�U*����m���iSa�][�v��h��=�o%�[��FQ�
A�9S��7mٝN�vF��7C�P��v�y�³ɣ��]n"��,����n��40ͫ��#;��..N0E:��lv���n��՝F���gc��'�4����cn�un�ڮ��][Y��V�t��m�;6'�bU��q��kv�c\�lu��vX�c���/b�mR^�#�l��{�M1"��֖�B�%$�Q�צ��mƭd�A�{U��sd�ֵ%��q�8&I!����zy~��<����/�<�`�� q���䘛nG�w���=��h^��<]k�����id��I?4�ZW~Z��4�K�~����h��"D8�4�n9���M�ֽ�}V��>�@�^�D"q	��4Z��v�|�z��~�f�������Lm��y�8���Z�ݱ���y�'�hmcnۄ�X&`��g��Y�������x�;��rb ~s.�w�RK��nG�y���5Jh
)Ҫ�*��UU$n���s��;~���L�M$Ӌ@������^�bW��h]�h.���9�Ȅ�$�ʟ��׀o���=�u�|���4�� �S��16܏@�_U�}UU����;g����5歖9.�Uծ�r��pۧE�2�[��[c�D	�m���C�9t�d:�/i�"�ͷ����hǰ@vܘ�~�-��7l�dq�ۏ@�����^�޾�@���$r���R!5�#����� ��A��& ;���viH"r$�zb�/�@����^����\��=��D�O��6�IH�~��`���1 ��Z�s�U�}�o��N�<�\���v�f�c/Wܒ��y�^��%3=9[^��_|��}�|�oM�]��$Ӌ������ֽ�}V��>�@�qh�'1��C$��<]k߳1"�-��-�қ�ff$o��ԎI���z�~Z���?�~K߬��=Wyָ�LQO�y��@��-��ۓ>qs�U����9U�*WJ����x�;��ˌ�([�wrM�c� ?W+�>�:y>��9h���o�K!V�$;4��Wk��m�m	 Չ��{V�-A�vs��$�4�����9h<r�r����d�����!�B!�ND��@��V��>�@����ֽ��$��獤�/@��-��_���Ihߡ�9���i4��/>�@�u�@��V��>�@8���2I��G���1=�Z��x�7j���c�۾��QzN���(�j��7,s��cu�vzq΁۬Y�i�����sԘ�@Ғ��X�dӺxy�r-^h����L�0nt�N��`- <F#�����L�{�v����@eD�r�+�:%NgX�*���];W\#�����K�Jvnu�d.�<�k\�klY�m��e:�Ʃc��dOQ�ݷ=`��+�r9�?ix��Y����X;rt̭L�5�m�(��dc�����mE�+c������()�H䘛nG@����<��@G�Z�����nm^��� �qh��Ϫ�<]k�/�տ~�H��A'�!!����$Z�ߖ���x}UJ�o���{���6��5dr1ۗpQ�xJ��J���׀}����=��h�U�y_X�ȡ��i7�}v��}V�y�Z��zv�>����V{]q�z�B�Jt�zB�YQ�u�\�3g�^�'��/���ψuy��F$���:���/>�@�u�@��V�{�YQ��� �M8�Ϫ۟�9$��_g^��s�<��׀~~���\��C�$�hs�h�j�=��h�U��X	ALjG$��r-ꤕW�U���� ޾����� ��� ��q���f�n-�}V����|��ݝ��z����� �����OUL��r@'Q۪�e�m͕ct�ᛮW'
�c��ű3@��ƵnVF������@u䖀��-�Z�6��Bq�iŠy�տ~��s��uw�^}V��}bC"�C�q��[Wk��U��{���� z#�*x�=��`N������ʻ���Z}���~x�FӉ%"�=��h�U�y�ՠ_]�@=����LY �m۸���׀}U�$���|��Z������)1�Lsx�#"V�Z�Y�"Z���R!1�0��H�:Ɋ��P���Cp�E�y�ՠ_]�@��U�f~�}]�h[���5#�cl{����-�Z<r�y%�ܻ~�8�Ɋ)�� �qh]�h�U�ԕ&���x{}� �wq��E�rH�Ϫ�<�j�/�ա��3�`�p��*���}��������7E"��cN-�v���Z�������
Hhj!���˪r;RSr�k������W�*�{PW�n��$P�pMDӋ@��V��>�@��}UU_�y������RU��]���%�<��@G�Z�$�y%��UʫA�|��LP��66��>��;V�yڴy�Z��RX9�L��E�.<�'���v�� ���^�_�~���[~��ƤrLm�E�G�Z��y%�:�K@*�eW	!���W���&$c4{*+�Ci�pG�`��HC�	Dv�(�'�a�����5��'�<q1�LB��Ԡ�,1�?�ѽ��p�L�rB&j"	_$��ￏ��� m���Ё��m�e'l%q;��+c{Lu�:�������4�7F�\.���e�eE_5P^z/Z�'�K]:l-� �#M+�YM60�=F�3Y�6e1Ŷ�)�bΒ���k �{V���2�ˮr��+�=��v�6V����"�Ps��j���N5#���;Z�V�z��tF��tt���f�.��Zɤ�^�Y�f�cl�%���$�m%�Ex�K&k5���-�vYUm.�l����"��1{!��m�� i�X���� �^�i�eZ�j��Z��vT%ٹ�7�G�uq�0�d���`�jˣvἷ�!��,nK�,�r[�K�H
.-1e��Ҏ�v��/\���a�{k�a�R!a�UV�m=�:�J� 8�1(�7m���[��q���-[��mt7i݆1�b�y躮y5!��$U�P�Z�4���t�[�L��y�2��i�+`�d.g�\���7�`^G�;iكkOB\�Vʵ��ΒG\�WzӏP��p�����n��KV����L�"���kh���k���Ի��lV�� �,�ri�e�Vq��"X�e��Ɖ.��rr�J-�;Q��	p��&�� ��,�$T��t��F�Kd�0A5V��;M[]�ʘysU�^��6���h��u;���o��\�L\��ٞ"�VBj�gg��Sq˰쀪��-�mu�n� ��c@(G�9sn�V���m�L��QM�%V��G>�ܝ]I�:�vj��B�b(8]ٷY�` ����Nծ8(0�m�$�g��Of�y{���t�,��VٮH4;cR��+�W[AK]�R�z�N�\�p��+�)^�iYݪ5¥j����eg-8����R�F�Ptf���I�GhR�+m�(��y\�t]i��^4�(\U��d����UU*����Cc�Y�:�2��6���*��HV����绻�wI�0P8�M��t�0�������*�w��C���A6�P;��e����ͣ�ۖd^(6[ǜ�g��Yd��2��m��B���P�Sup���L����<�r�۱FI�-�3@���d���(�������;C*�gT���s����z�6��-�ƱծD���i�Fۇ�j.8�5r�[� ٹM��m�d]�6ǚdda�Mkr���un��3�E0���m�h�J�-�Omǧ�:Z�����w�����/k�I��j�<�X+�\M�D�0>9��..]����S�S"Y1~Q�Nk��ՠy׺������8�;���d.U��y��h�K@u䖀�lx寪�3�G/��E	���1���|��S@��U�^}V��}H�"�C�q��Z��3���ߍ��-��>J�S�gs�;��md��(��i�p@y㖀�\�l���}��:��@u��т���U�ہ.�J��n]A=GMaPs�r4�t��kL�{��������h�cn/ ����<�j�/�S�33�]�h�}�K1ɓ�9$�@�מyԪ�U:�Գ�?��o��������[~��ƤrLm�E�}�o���x�:�K@���w[H��P�)��>�@�U�y�աԕR~^�^�݈�#!r��[�$x^9h����� <��@~�s����luj�� �a�G�r�.���fl�%l�^�Q�yD�N�����{����M�����~�_�<��ݼ�o�R������@���i2(D8'mŠ{��=�u���׀~��^|��a��[jO͓"i�Ǡuw�{Ϫ�2~���/9ڴW�^�z{^Ta&(D�ʹ^9h���x���nl���/�,�&L�brI��;V��>�@��U�yϪ�=��
ı��Af�RtcJ�g�nJky�p��Dv]usdě��z4�fk��"$X���=���<r�x�:�K@v�I���Zo�4�4y�Z��hs�h���m��s�n4�h��@�O����Y�uw�u}B�$�F8����;V�oJh��/��?{��?dweZ���I�B!�8�nZG�@y㖀��^Ih�*�t$f��KI`�>!]en�Ӎ��o+�zTw�Y����+[f���A�-�����$�-גZG�@z�2��I�8��iŠZ�����=���|h���Ԗ�&)0d���?{{� ���^��߻{� �y�wX	��I��ȴ��Z�����Z��Z��� ����d�x�ߺ�IU%�N��6�����ʴ !� � �T{�o�c��p���Q:vGv;\n`.v�P��ֱh������Sz�M[۫�Ͳmm�Xvٛ-ĺ�{��h�S)�0�{s+�M.#m�+eS:c�Ѥі��.��R�k���G[d{��{X�m��ۤ�t�j�A�d�++�i�iܽ����bN�L*ˣ\Btb�Q��Í�\<n͝�Zx�v�D�<ҳ]p�>��\��4�Vu�����{��ĝPt�֫I���gQ�mcL��]u�5�1U��]'O'3:m��f�5G������>`��- �9h<r���i��n�#Xԋ@�@�}V��>�@�V�W�D�"��8�n-��Z|�̒��9h9r���n��i��h{Қ�ڴ=}V�m��=^וI����iŠZ�Zԕ%������x�ߺ��e��w`z���U�J��v(�v�:�ὂ�=6�i*��K��-���8s��@_�:�K@I6<r�d��<��Z��rEwe��ݚg*�J�R�Ī�]r�2d���ր��-�=&n��$FX)��>�@�V��;V�m��-����?6�NI�&Ih���M�����i�Y&1ōH�9ڴl���>�@�ڴ�#�X51@s �6��N3ʗU�U�[�^g�O��@�N�,Ki�E��q��Z�S@��U�Z�Z��Zz����(�q(�4^9h	2K@u䖀�l�L�eb�n14�qh�V��;V��g�ߗ�� ��<��s\�����ʼ�KRX9�H
L�Šy�ՠ[e4y�Z�ՠrꀡ2bj8��f�$��9h	2K@u䖀g�?;�ڲ݅i.�r�Eq[�E�2�[g��[�3�Glgr�K��]F�:엚 <��@I�Z�$��`�v݂$C�ۍ9$Z�վg���}��ӌ�o�|�J�=��Tn���I�ǍH����h�M�}V�k�x�ͽ-ˍH����:��_*���|`��<v�^�UR�$�J�ED�q�#�w�y����;�l��J&�X�p�=��h��@�@�_U�~����}�a"R71���n�d����V<�*r�qu��+:ܶa;��/���W�I$��k��.�۷q��/���<�j�;���������K�I G12H��<�j�-�M�}V�k��3?~�H�ߘ&LR9&6�"@}�߄�9h	1�@u䖀��M�,��X&L�4y�Z�ՠy���IU>��0��$e�*��$�@�ڴ9ڴl���>�Co���7�lF�dH��c�U�]�x�h�ۜ�9�\GY:tMe�9�T�lt�y��rE]�=F��:kZ'��m����iv��h���j��FY,EY)��ܺ�v��k��v���mO86;�nKv3bR{9��]�;���c��I��.�0�ȳn�O�|��*+km�sl�&;��M� k8v�<4���`�^�ʴ򢵲�C'{͋/4�JIC8vh;C�.��S�Yz�:R�#1lNp�3m��l-KUts��j�J?�o����������o�*�J�����{_�ǒ�q	��z�h���ՠy�ՠ^��6~r%N,J8h��^�������T�U]���� ������	1B7�M8��ՠy�ՠ^v���M ��,N��\���?{{� �R�$����|x���@��Z/jB��JD�2��I1V�L���d��1�D�֍:l�V0��ڀ�nLi�E�^���Қ�j�<�j�=W��,��X7�����k��4�`!���P����%�+U\�RJ�xw���:����� �n�!�~nF9$Z�j�<���RM��� �oy�m�Ց��"�����:�}J�%~�}��>���>�@��Z���H!�&�H���Z<��y%����r\v�+=]����:S���iC���흗g�t=���S��{����/4�u�f�̟Z<��y%�#����	1AG�M8��ՠy���7ݚ`{~�ΥI6w�|�HLX�-���h���=ه��`N �A[N&	 ����0J�@C$�5,�}#W5���̦+���������	�a&h��%�X�↭�I3��B�fxF������#��W�0TG��	 ���A��z��c@x@�x�� �;�y�r�;��@�z\��1�c�h�����}�ׁʕ?6w<���,jc��`�p�=��h��@�@�e4�W�_AD��$�G�!�@�Qۙ�i�m͉I�y��C),p�@�u+P!�~mƜ�/ ���Z��Z�4����=��x�}Ѳ�ԁ"���ʹ^Ih���Z<�����,�$C�6��/YM�}V�R��o��m�< �u��r7.����0>~��xm�<����<I(��\�hy�TK�G�ۋ@��x|�/{>���|�=�u����z"����ԅe+I�d�g��׊��q��՚��nI����m靄��a�����䖀��-Ih���`�nLi�E�^v�����/���}��� ����R�����8j`�qh]�h��@�@��Zs�b���f9$Zٙ���女�|��ՠr�נ{]�2&DH���06�׀}I$�gs��{�ʮ���~U��dM���w_��|�ߵxmus�s�e�E�՜C��ݖ�;oV��4s�ܵ��T��ݰ����]�<Y�Ʒ;Y�J}���~"���v�l�,�#c8�"���[q5�Ƨ�[Y�m�g�!�N1s�	[����j�.�&�m�9;[gI�m��x�m���et��гf�� P�j6�.�ntm�P��Fw;D@s�u�޷��������d]A@�u�n����g��nG/=u���;tsÜ[m��(q˛�Cl�k ՓV^$,���=�u�{~���vU~a��|���f��D�iŉ'��>�@/[49ڴ�ՠ�Z���<Q�&�N- �l�<�j���������:���9�,�$�,#�hs��䖀��- G&�7���6`�nLi�E�z���>���Y~^ {~�hs�h�V�͆L�
H1�L�˘��긆ݢt���W9���ڞV<�Ӕ0p@�L�z��� ���Z�����H�s�r3�-
���|�r[��������ל�{�x�ߺ�|���dj@���@�@�wW������uw�߾����J(�@�$ۋC�r���O� �O� uɨ����5�?I��	8�y�Z�l�<�j�=�ՠy�6W$R6�H�Mw2T�0;r��z;)��W�k��m�j�5������ŢX8dyB�n/ -��y�ՠ{]����:���=���$�s�$����ou�R��l������< ��ٝ_*�I]�����!�w",��x�|�=�u��T���TeR�*�UVa߳���k�<�w%��]�[���U'����� ���Z�j�-�X��nF9$Z�{� �U*�6w?�v�s�<��׀|����M���%=,�՛e�G�r�.�c�L�S�΋�Tc���v
��΋F�8���{_�-���=��h��@�{]iE9��q&�Z�)�g�Ԫ�޾��u���?{{�>�l��-���E�x�p�:���/;V�%�|����@==V��p�&(��Z%_RUJ����{��� �vi��RJ��fW�0W:�-�ۋ�K1�I�7"�<�j�?W+�O��@s'ր�$����n���H�m#N3gU�8tu�qÒw��;.��q)8�r����w_���l:Sc��n�@�g�Z��s`���-���,� ��n-�}V�yڴ9ڴ�ՠu�`��?7#�<}�׀~��^|��Wu���7��z��"2FCqhs�h��x�ߺ�>��}����ϭ�q���ۀ��x�{� �$�ݛ���ݜ��u��*Ԑ�B��ʥ�{�|�S�����F�v6�W%��w:�L�Na.�dB�����i�'�֖�Ɂ6M�6yg��Ui9�Q�`�n+	�B���]�kl�ۍۦb��s؉OV�{:�]�\���n��OX�u�eWV�e��B��tۓ��[(�\��[s��Zi��������@��D*���?�|wo��>9�e~Pv����[&.��-e��ו�:������=�{���%�5sT�mM%����a��#t��]Z�zF��;�_=o��;	^�d��tB0�o���?���ՠy�ՠ^v� ��R�28������7��y�UJ�g�}� ��{Ϫ��V��s$�#��r-�$�y%�<��@G�Z 첋��
G$��c�h��@��U�^w^%I������K� 0���w����-Ih���䖀�߿k��M�䈘Y'\3Ù.c1���g2μ.���!QqOy��3X�g7��UZ<��y%�#�/�W+�d�����ȡ�2��@�{&g��^ՠyϪ�/;V��V���1H���qh��@��U���?%�|�k���fI�H�m8�n���~����v�s�?{{��RO��� ^�}�H2H(��Z�ՠy�ՠ[e4y�Z"�MU1'�4��Y���b�pQ��!Gc���fNzh◦�%��"�[�,�$�(܋�=�m��=��vx��H�@ �Q�IW�a���o�w��h&�ג^��3;���,��������ߖ���}�ti*0$� ^)����q�\�rgU�;� �K7l�C��I�m��<�j�-���K�^�w� ��e��1\������-$� <��@I6Ы���l�լl)y���D���*��am;t�t�m6�N�j��":�am�c�M����`���-�Z�RF�۸ӻ�`{~�ΥT�;�q�{_�-�)���R@��Q�����ly%�$��9h��u����$L�.T�'���}����_�׽�W�
'������ύ �P>�Q�I���"�-��<r�M��$��6p����]uZAԍ�zt\3+ͳ� ���g�&�m�������Ő$��4y�Z��0���ꯪ�R^X}��� ���K$C��RH�l���^�m��;��h]�!�B!��bn�^��7vi�URI&���xwN0}���Dɉ��Ӌ@��h��h�M�v� �h�I��(�q&�4k�l��޻V�m�кz��""���$�2�B1,!$�,�H� İ�$�D��Bz��qfa�1"��T�@ZV� -���&�Q<D4����	$Ē	a`���Ia��0L1��9oV�:�F�eI31n����'|��}�^Ǟ]����~Q=��&���&ȍ(I�&h�&�F�6��D`��1����`w��s{�������p񢥤��nk	�2��nm$�Eƭ���i҂M��dn������-��TUԓ8��<b��9���Uc'E�w<ɂ���a8`ȵe2���3t�]m��2��ô����v]��0����A +� ,�BY�&b�5mU�9\ܺ݉s�2�k(p��UΨ�`�AU��-�R����YMۇ�j��Fu�:	,؈�r��4L��ԩ��eP�'M�mVi������=�Y)�r��m�ж��IjY�`u/lU���K���� uT�	&�P�Z�u��uFv9Z%6ҎN�.�N^�!-��g��v9]A�5�<6���^�i���cst9#rfn#Yv�
6�m�74c�f�Ы���2�9k����0�{m�����7Q��يÞ�Gm����bͮ^� ��8N�:N8�6S5�\�@=I�f)���v���h�T�j�(��m�j�(@F2�汐��o�8Oa�뉶��׵s@Aq�w[��Ͳ7]�J�a�0^��G�t�X�R#b�d\�x�m�;2E�	�N����8��#�ΐ^"f����+gE-�q�8�:}��ܡ����Y^��I88��%7!�ٶ�@����edWa��t].dm�����̏$h�E�i��em���{!ݛ���s����뭭��+�F憜���c��j�H��`���'*�"�hv ��w9����y狎��tJ����4��Ѹ �!d�3�ŧ�]�mj\�v;L�s�I��Sm�6V:t'#2;P�Q�%٫�ˮNJ�z)�)�̻�sF�R���t�ڨ��T�g�����f�jRZwm�K����L$5*�5�nY{n��shU�m�������U�N<W�4���<��f�ث�=�
�Q<q5���X�;L�V�� +��K��UU�-��V���j�(�U}�`�@�����Vz
w@��jd#D}�=����ww>���U8��8�/��ΗJ�_��E s��3==sy�lOwUƫ��M���ɦM�n�ၶ؇r&̻�p�m��#K�۵��v��C���:�Okb;u��;u�ܵ�qxK�����.�,k�;bFrsl��7v�v�5q�L���)���|-�ݙ�]n�*�nup<�i�њ�;K���;T���j�٦ġ�9�C�+��N�ꕒ�2�&3P�նn��W�����������V��4�nK%�m<�3�A�λ�ӱ��s/i�����Vź�=���D�1�.',q�w�}>0}v��)�{_U�{��I`�I K���� ����U$��;�q�{���ݚgʩR���X;�.D�ˑ��8�<��ׇɾ�`m�<��c@�I��{Ϫ�-���ou�|���S��� ���mX2�H�rH�ݚ`%�����`��=�P����̉�LL#��C�.��S�X�^�F��;1�5i�$-��-Ut�Ic�Cp�<�j�;�U�{Ϫ�<�S@�ګKTL��M�M8�{����� �� 
~�k����U��>0���ϕSgoqmd��r��i�f�2}h	&�גZI�@��m��K��n�ǁ�R��*�U~������Z�r�x���2II�p�<�j�;�U�{Ϫ�<�S@��*ܙiF%"S�m��T�Y�l�È��Nvf]������g�-[ck"�LX�ۑh�M�}V�m�}_%J������7��"��KFay����`���-$� -�ZX���$�@��hs���\�\�W8r���&�@u㖀s$�e���W-�;�`uRO͝� ����>�@��h�k�(�q	ĜI�ǀn�� >J��{���8�?{{���7��P��Ë��`9���)t�M��2J�P��9����F�Z�w�Rk�=��iŉ� ���@��hs�h�M��$���8h�L������ӌ}�ŀy�F�qI ' �8h��@��i���便O�ﾟQ���B9��6�Z�`��lM��]��W��䪮o�{5h���,�  �!��@�f��]ݜ~�����L�6^�ȯCcnH9F8�nZy^�p�r��=Cȵn����J����c6�wo�kl��yڴl��z�h]�!�H���&�^v��)�^���S~������"�C�8�n-����L>UM�t� ��o��Y��(�qbm�@�e4l��yڴl����Z���$��Q�wf�ݳ������L�T����US�c�
�Zt�m�.A�mʶE�YD��W��G� �U��x���A������;�j�/Q�\��*P�ΰ/��vH�����"�Ɖ=;E��]���1c�2κ�b��]^y��ۙ�g�s�Rɗ�r��`�q�X��M�m�Ͳ���4b�BI��#1��K�۫�lX���l�f�Vplc&" 7]\����Ǩض�k����T��rt�����{�������J�]\9���Y��Jp��N�N� U9��i]��-j�����M�ch�ϟ��@��h���m��:�.X�#����"�-����_�Ɓ��O��h޻0d��N����)�y�ՠ[e4m֖0C�9&1I"�-����Z�S@��U�uvĆD�8�17�v��)�{Ϫ�-������~n/��st[/V`GI7hv^�j9�q� �nӺ2t�3X�:�q&�Z�)�{Ϫ�/YM�v� �h�I�����I�h���߲���$�%JA�N0|��o�4�=^�RX8d��$Ӌ@�e49ڴ�S@��U�v{e�L�LM��� :�K@G6<r�͂�� �cP�bǉ�"�/YM�ߺ������@�@�kif�&E��XV
+:�!붧b�,�̛"�Y�v�F�<��#r`��		�'��M���<�j�/YM�tk1����h����;V�z�h��k�$2)X�P��49ڶ������2$�uHp`,,T�"��~����}�)�{��B,sq&�Z�(���-� :�K@�e��36���I�h�Jh����;V�z�hs��ۍ�%$�HH���J-L܌��������k��F"�4ܪ�;6�M8�n�)�y�ՠ^���Қz�Ia&E&&�"p�<�m�#��� #��XJ���,hmȴ�S@��U�^����Z�۳@�I�p��32��f��;zq�~��^��bP�*�դ�T���w�~��-�$��+��:��גZ9�@y㖀������߿�.����%1ujȔ�N*;$պq�*�%���]=�R��gE�5M��=�z�h���S@��]��Y2c�8�n-�}V�����4�?{{�:�6�ŵ%;��i7��-���<�j�=��h�k�X8c���iŠy�AגZ���9h������&�"p�<�j�=��h�괯=��r�M":�
�L������[�Z��<{e2ac0%�W�3�l��`0i7�n�[����F�^��'-�]6au/�v��"��se� ��o73vk�Ju�c=�����k��Gk;� �V2�Ռ�<wk��rq�lF�M�٩�m�g�k�{ls%e��J����:E��dm�vUN�[�����n?����FN-Ϛ^����������s��~{�����>l�C���'ZR��n����+&���gi��џLs�]OE9�ck�-7�Z>�����<r�sa����րo�Ѧ��Xn�{����-�6���o��-�C��I��1�I��YM�v��}V��>�@�]�!�8��It]��I?6w<ݽ�y�������{8�=�����������<���9h��@u䖀�����M��Vm�-��n%X�zd:�]Q��g����o��e�6�l�^FF�Q��.}z�� ;mށ�g��z�|]�
�#�p������5RT��U$��RT�U%I�fm�� ���� ���^>�|%�������@���Z����}V��YM��H.H�#�u��{����-�Z�ly"�=�ݙ@��"�=��hs`���-�ZXz�ں����m��d��N��k���i���v'SÖ89$��9?)&1I"�<�)�y�ՠ{Ϫ�=��h�$2)Y$��3D^Ih<r�x�:��}h��?�&E�`��i��k�-�~�9~�-�C�px�F	���@������HF.AFc I DT����,C��LɄ�� 4�`�� :6���8�S@L�B�BY$X��CBMB��d��`JC��bF$���A@��AD�)KR� D�̤BL4@TI$,AC)%!A C$�AD:S�� �ef�����$L�EB$��x�C�&BXF�%��t��#>
�h�	�\���ҦiM������,	I?�4�{�f&`%fFm���<���^.�����q�Y,[�r1�.!c�PN� tU���1!Dx���ӂ�	ݯQ�^��S�]���}���� ��%�~n"cNF��C���nE����o��$��`�<z�X82B(�qh�M�33�>�x�}>4{�4��\Ƙ�! ��a�Z��4nC�ca����MU��e�t��"�q�8hs�h�M�}�}��wN0zލ�)�ȅyy�h	&���	&�גZ����I]��}xGKq;����$� :�K@I6�Aeg7w�$�(�4l���;V�m����ݿ�g�؛�����D�G27������]ݜ~ݽ�n��6���??w{w�jM6:��	�(���R+�̔WZX�n���ݹ�J�,ܬ����6����|h��l���;V�{m�?)2!�"m�@��U�ԕSgwN06����L�6����(�������O��v��)�{Ϫ�=��%�������@���wf��ߺ�:����%}���|��A��%&�r-�)�y��wf�����>J�����BI����������uj:-[iݧ)�M��<���n�|��ٴӚ�^6$oh�7�E۳ 6�N^M2f%�;
n���ۑ�g��m��Q=n82��V�Dg+y���'[��|��tuĩn24O;�u[on�P�-�8�Y��3��-��\3����[uv����\+zN��6��&x����c[����ۅŮ��\�\R�Bg-l�ͦ�o{����������9yU.�cFu#pޛ$ȷdxu�°�|��6�N]��B�-�v07.~���}M��$��`���YS���IbjK� �٦&�v���ӌ�v���$2)Y�`�4y�x��0�RT�~��<���6^��I��q��Z�S@���@�f�R~��x�w�)ȣ-܎�����-$� <�K@I6ӟx.�A��SLvq`����,�f2+뺽s��TO'������&t�[zdʪ�6/�}������-$� <�K@{�#m(�N�0�� ���y�W���E
z"�&���Ux�)/��g�O��{� �٦���R%&�r-�)�{�ՠ[e4yڴ}��H����М4{$��`���-$� #����~$��#�@��hu�|�ﾟ��Z��X���6�I��Ǌ��3љ�.���M֩N��� �3v'%����3�D�G27�v��)�{�ՠ[e4/Gq�E�`��m��z�h�h����;V�� ��K$��Ȇ��7���^��<���2�HUE$�SIU�v�^�l� <<��,QE�r-���=�j�/YM�v��v�)2'�I'"p@y䖀�����g�Z9�@;p�5��e	�@Z7*X鬫tuW6�v3�
]��q�ali,�86���q�v�͂�$�s`���-�uzD�#&�4����;V�z�h�h���o@F\���#X�L�@G6<��͂�$��[�,�d0n��Z�)�y䖁er��+�9UʤL�orV�"�0pn6ۋ@�e4�?g�����}�O��ou�RO�z�:+q]�'mh��)l��Jt�zA�N�G����:��$7S��D�X��&D4�D���u|��S ���}I/�;zq�����-K�Q87"�/YM�v����=�j��߳:��RdRbn r'��x�ߺ��&���x�ӌ_��F�䄊)��Z�)�{�ՠ^��~��}��;��H��`��ƒp�<��^�%Iv�q�v�����{�������9nm�1�+*�t.��ֻqX�T���t�=lo/`�7mb��˸.�rZ�T�3��(v[�Ark�ϖ��D�(Hc����2j#\�V1�t�l\r�;M�kh���ۀq��q9mh)����h.�˵�m�i۷�X��sϑT�4��WA-�4�,Ig����e���.�I�i�FͶm�疒�ܐ���l��7���ц���h�P�Q~�N�w{������m�\N��B��g�fsW-z��\,r5s�uG�B���n����5�$qx���@���@�e?���u|����HdR$�9���h���͂�$�s`�«�ʻ<���"d���m���ߖ��;V�ʪ�U7��� �o������.)e��0jE�{�ՠy�S@���@�e4�UtH&D�#����z�hR�^����oy�{�� ���ږ@k[�)��꥝�fg/nD�v-������mR�!u��Y�����챚+|�?2K@y㖀�{\� %��e�j�#��� ���^U*N�)Rk)W+�\�Us���� �^IhzG�P�0Bnc"�=��<�)�ԕ*o;�{���w�-P��%����s`���-� <���vĆE�Rd0N��Z�)�{�)�^���}C�w��pL� ��]t�\Ue�7��7R���m�Z-��-W��{�����a��,���m�~��� <��� :�K@H˺��ͭcNL�4{�4�S@�@�e4���#r��ӆ�z�r�=�{��6ĲCD'� HQ��U_� 7�|�߷*�����Q���$��$��C@�@�f���4����q�s���)#QIEY{���lo`��ly%�/\���H�L�BA7 ۃ�=u\K�ڜL���*$$�^��.���{���wϜ��0BncI8x[>4�S@�@�e4��I?F �C@�e3�UT��;�v�� ��f��{���H���C�y�ՠ^��}�3����}~����"q	����ǁ�UI/�%I_���{����ە�ʲ��!���YϾ�Q��K%��Ɯɉ7��M���<�j�/YM�y��#di(�q�BI����C-�iG3�r��<��]\�1v�`Z�Cn	`�4�E�N�)�y�u���9R�_*J���{�� v�Ѵ��$��ND�y�ՠ^���Қ�)�Uؖr�&I�!H�������גZ�qmGb%��V۸`uRJ����`�8�?{{��T���q�olT��n4)r��L�K������߷�ʿ�TW� ��� ��J�(��� �+�TW�@Q_�UEE� *��� ���"Ƞ(H��"�2 H�H�Ƞ
�4��H��� ʒ( B�,"�2�()*��(
������
�������� 
�� *������𪊊�������
��𪊊�ʪ*+��Q_�����(+$�k/��/�ă+0
 ?��d��,�� @         �@   �   �� ��$%������TQAE"(@ J    @ HBAP (
�J�  �@ 
�Q"�� >�����95�^�5^������ �{�,ov[�}׷��;�v��{� s����e�� 7{��& >�.�1������9:WpҞ�iq�w��L�n[���p+�  =�    )@�� �_[rz=9{���{������    '���&'p �nR�zt�ݼ C��ӓ�y���Jd����ɸ��9n�}��烛}엛+ӓ����� ��(   ID��e� ������._f��:���zo� +�> P)ي  �P {( �@�c   �� 1 4 , @ "  �� �:)� 0 �@@4M  ;�   �QH�
0 �t�M Q�@ҌA�A� 
 �ɻ>�MŻ^��a����O.{�7ϓw��񻱫���U� ��쫽��5<�v������l�m������n������.]�x��xϩ@ @)$J V N|�g�޳�u�y:�����@�>ӓ�=s˻{��Yǻy�]�����)����cx ޼�"�ӎ ۵�z���[nN�n3�g� +�{��������s�oy���<�q i�
��)UC#����I�f�)P  "x�T�M52����F"{J�ePd21����j�*Pd ѡ�DHjJ�D `������?����������G;���Ez�*��(�
��*��� �+�肨�EAS������0���9�x���$׏�$>���x��A<"��\8y� ��q�|̙���4�R�N<?Țb_ W�7w��Xn��L�o)
0�BD������#RdJ0I"$�F��	"-��!���<`R208p��f[H����ӄ����o	�c<KZ�D������-���BZ�������J��BHSZuC�ԍ�5�ݐ�
1�%� ����ar'c�Ms=<�0s��y5�1���.$�0)��
E��������.+��D��A�T�Ѓ}$b�Āz��4x��F��B�J^H��i`���+�~��/�H@Ȕ��<3O08~q#P�P D��8��6�
�6$�!}h�!�=>�:����}�̀`Ʀ(H�7^�0ϵㅓ
�5�Ѝ��4����9l�FS4�5r��!@�1<`f�HS��(c�<v�ɡ3-'&�p�hc��ᓏ��i��!���x�SG����l孱̀i�J`���&^@����T���T��O��?�H��a� '��٭��܉�����✩�h�_��u�BQ��A:�!*0B� �X�@"�h�`$����R� `,H������R �*. �v2T�58�(
$�A�1�"D E����
A�0� ���"QĜ�b��p^#,jDb!�Ĩb�������	(� ��A
��@ bq�F%D��b9�I
`jo-i(���WS������@�E��(�X8:�ĭ�J;�.�)��(�*(�H�	�� �B����[d�#dF@`1-4�XLb0M��+���/ՍL4��1C@�@����ƊB�����l���`::�� �A
�SS��e���20�H1��cD�d� �+��Q"E4H��R��
q4=ZK��;O��S����^�K�H�A��E*�`�"�X�*8� B��q<<���6ْO ���%�ad������$a����A�嘰���CY��bF��A�"�����n��|���&	��b�@�z,B���B,,�Đ$����.OMh¿LӔ��4�t��;�Sx�@��'%��0�@ N0ܳ7r�!! �HP�au���l*me	YRH$S��^0���+�aLC!�dXp�7$@�0ܩ\!$�H�$�sM��L4�p�~�|$7w�C9����ԍ
i��			Mԉ�0*�
�n���XaW����̹l��H���݉8���N��@����<��S����X�"Q�M8>0c,���N��sNn�#�(���ٚ�4�5x�/)]�tqÇ� �c����I� ��2�0c���07��K�#S�L��qw�~��~�/��J,�C��OU�ӂr$�G���r&��jĈŁ��)��0�9��2����O����Yn05�)��F1!7�y�:�B�nxd�����y��a���p��8��c2K^���_o3m�3�a���x��B]98d.2��p�4���.k)����R9�	��xs�I��a
D���jGLt!p��n�e�aM�Xݓ\ ė	���g�o��_<!qӇ�̞�$t�<9������
���76.Y�d��=������~�Iyu%�J�jK�bO0F,f6!bx7�-���E�[B�,�2�IrДiBR�(����
a-�z���L��w+6����3Yv�d��0��	ZF�RRB[Z��P����%)YjE�ah�V�F�R��������
�
B����*�ZF����+�!������Bo��������L� �͛����ϳ5���y�/�!��/���&��@Ä'z�K)�s�|���S�@�F��M<�Eq�@��.o<�6�~/������2Ji��Uz��Ha!20�a���12I1�XL%V4�'m�SH�V0�Wr! V��@ӎ��n�
JX�8�0.lreS�I��p:�ZL7��ݷ.����
�c�y!$<3y�-�G0�SJY��5�aXCx��:������!b����d�"��e��GD�r��I�.8Z�2	�l �B���+&B0��Q�cFT�_�yMxC�	�#,�h�c�2�Ŭ��K1�d�ԒRbF����J� �'`"@'���Ƥ28!"zaz���K�x2�0a-�\��FぢŀJ��D$�� ȗ�1�1u:�&�񱐴ƺp�4���p����Y.�!$)��<�F%����I�	OP�p�g3���*:���B旜�F��r�J�hCŊ���48D��p�F\��%�e��0ԅ�� �J0�cLaLe0!rIL0~�|	!L5Ӽ��愎Hk!���!&K��I,�.��&sy�%�NA��`��:��MߘB�N�Z�J��D��������FF@�U_�<��Y�2�A $Ԡ�b�W��b�	�ϐ��Ȯ!�L��b����A0�L���%0�!aY���ʑ�e�[I��h�3&s�x�,J�K!!V&��W�7�HIFՅ0׏�<����<�!sT�H��4eaq!3$�e��(x������<�txJ�(y���ӏ��n����K�!vLHp+����pX�$d�SLx�h�X!�fo�y˚��Қo�q�$��sN)�rB��y�9Lhdjdd���8�K���0��IJ��	��
�i��鰸D$�w8�a>>B#�������4�z�������L��S=!YN2�J�xK�+
�����j0(qa����NKIn�+����Xn�p)���0o�T�<�.�<��=� i�)���o<ЗF,缙[������s���NaC|�~���CY9��=��.^��y�/���n2�s���ut�����
ě�y�O�{�4� ��� L�hA���=�7d����߾=.���w�"oŌ�NXO<����=9��)��p��{���za癞m�}秾}�P��������p�/�ϏHS�㐹��ˆ<4�|ee%����ϳxxu�cL7�xro3�l�}���9�St�x��F���y�aa�<��8qt�9�<�<|%ͼ��y�<8'�)�hř�V{�|8l$x�='����xg��)�'9��7T�,��X���r�S����t�a.��E���>H��4	�ސ�O����LXpO7�D�qaa�|���L��xg��20�9�<��4�XS��n��a��B�6�>����F�`K��	��X�x`¸:l/�X��u�"�_D��
dJFB�)�.o8x˧q�HCz�!']=ad5�#L4�:����cL3�THq2��b�&�����       -�       h    ��H   ����[kXg[x l�܀�['Qa�i���O�>����W�S�	e�=���� fU��um|UT��]�y�H�Z�kK6��m,V�6 �m���nW/�M�� ��oIx��(H���` .� Ams��]��� �lm  V�m�\ ;m����$$$�jP��l  m   �H  ��h�--������m�ٶ` ��  m&  [d�88 &ٵ�l��qlױ؍t�z���j�t����'����}��pv�us�[����*�l   Z-�� J�cv�.�ڢ���Bj��ȁ���S�� H	���l]x���	 6��t����4m�5ͪ7L����U���@ H�I�z�Dn��9�I�ZڨXvp%IC��UR�P]$�8�t�]:�]$�|�[W���m"�a��g�ћ	�ԇ#AU <��UX�rk6�z ��h����nh�㊛��\ [%[!��WW]��յ)u��)E�M�$�8k���mgUT� p�WM*����U\P��A�Ζ��'^�!�Ю���g�Ft�@|�(�_Qrkq*���n��v���泀bJ���U�T�U�ڵ�-���+q^�m� m�i{K=���m׶�$GH� d���v��H�[楒��I�0p�[V۱�O;'ƺ�mom��l��+�yA�Vڪ�)`��k���28@��eٮ����l��� ̫P	�M�m��gS���	 ��M��5�m��Rַ[&� ���mb�H%�Kd�m�Ӣ�E�f�u�J���m�<����6�	v�l�Ҥ����Z] ��i�!e'b��]�m��ݶ �q�� 9W�1�{�tUV�m�TWDk�R�vZ�� �6�\�]�[[mP\�&�n�*W���\��ˆ]\�[�����%mR��ږWj�ej
X�uK�0��h8����yK�p�n��Im�Md��8 �b@ �[RHX��-��l��S(�p*-�i^`#�f@�,5�5U���v������&���E,���8��m�P e c�Hx��$�K$��m�r� Z�IY����0t��[E��]V� *+KUe;f��묧t��+�i!m9�v��┎�v����ck7����� s��8��k�����:Z��v����eiT+-T��4�U[T���U[J��Bu�h�n�}&I�Bmv� �m:j����n�myp�ڤIV+��[��a� �-�!�k�j�28���٫iI@U�yZ��I��)\*ޮ�RC�J���J�*���5��vCb�V�kL�U��m��v�[@  �ŵgQ�� �$[I�mm�:qi�N�<ݶ���M����ܩ$�� p   ��T�*���;K�UUG  k�-���Z��[[H�����I@�H6�Ջ(pl�A]om���U/<�@lcIu�4��Y@��k� �mI9����&�Rl�qsz��B7<X�aj�A.i�lm�ڬ�UUU<�r�R�<!*��lդ�6^׀N j��-��6�ܣ�gn� s�$��*����%�t��g�� �Ѵ��Ƞp���uT��sUT4��f�H 6�-�[Aa�Nm��.�@�hR��m��bCck� �����8N5�,��  �     ��j۶��`<�}��}�UTp*�ʀ��kX;m���6�S!+�g��e�z���� �9���  �h��]l��iY�� �q"�Q����Į� "�ݛ]	 ���f����í� 8  �2ս@-�$�B��   R�8Ӕ 8H��,�	l������]U[=�Ԫ����@-�[���05U�۴�  p6ؐ�6��H u��<�������]Ҷ,�Ė�	I[  [^
ۀ4��]�j�$����� �@�E�jͰn���lp �	.յ�RUE�`���p6۔�9������|��k�x��kR@��,��(	c�-�������Ndݝ�[mm��`�f-�V�TjG/`�F�[7I]e��.�M�<���Y'If�n����a  ���L$ic[H�y��7c�� 4�N�Z��J��  [I>o۶Ŵ��5�m���e��n�5T�Msa�	�%�I�W֟  ۫�z�	�����@k�m&�n� l�.כ6͵�`�l6ݎV��[F��� ,��lٳ�Z����[l   �emlUT��t�T$-��`�j��n�� kY!&�m�P [xu�`��n�-�k;d��|o�������зt��  p�i��[S#Gn���m��h hp9�  $i��l����m�H�`��gm�X��K,�����JY.�a��;\[@ ����m�m  H�  �i     D�@  ��-� [Cm������ �g mݰ-�        m Hm�ڕ�  �@��� �ӆձ5T�m�pTcT�TK�l��  m�m��5]im� �+mn�m�ne[X.��������Y4B�hʹ@*�a�j���m�m� p �	h@^������]@��*ԫlsu*�,�$6�t���on�0z� �    �}� H  H �8   	m��  ���l  �             � !m        � 8 �H�  l��@m�f�`�m��` [� p � [R  6��� �Glim���    ^�I/Z ��m�	 z��\Hm�mf� m[ r�^�m����M�p�pm�� �Ӥ���o���lGj��h������E��6��	 mm�B۶ÀZ���[A����	H�$;vv�ض�   G  �Ԁ 8 �` �� 8 $ �    � �e�  m�  �@      $���   �`�8�h>�@   m�  ��HA��m�f�6� [@��~�m[ H �M�� ��l �*Ps�Uj���[��L���
��Um+�@�s�[�kZLr�6�� ���Ӕ��[T�����k�&��i[�Iͥ�]&]6� �oY m�H  �����  ��   m�    ��H  � [@  @  :�X` G�� ��]n8t�� �	 '@�m�m�v�Lp� 6���K:�_�N�e��p�%y�.�4j낹T���U!4�eD�n�qͶ	ԅ�m�m    �M�Z��݀�� ,��V��m��U��
��*��UUU�ZĽ�7*ӲJv�׶��	��T�v�d+��` ��sW).�7ki���� i6��:$���WU����Z��Z��D�om�N��[�R�+f�[gU���Z^��ə��v^Tۧ���n��&./9�g�]UW���Hr�/c	�j�6�c;-�t�@M��̖PI5IUYy�j�*�@ ��V�R�� m�   ��2`����	8�$� ��$n��m���I�� -� ���kNt��  �` ۶�   f� ej������@UV�[@m!��Yu�qm 5��pm�8f��[��` �  �vͶ-�m���[x�cmv�$Ͷ  �I�$   �  M����n� p �V�f��m�   �j�KVӀ	v���cm�m�@�klF�X��Ճm��� $�Z���`%UR�wih$�6�t� ݫ�  �q�[I��X�������mf��җ�gZn�� ���B����-7F��@[Ri6����km$k�Yۯi�J�{a�IMMU6�*��vy�=nl ��6���J�UUJ�n�F�
�+�.Nfm
�V�����j�h �nr� ����mm��`��d	5� m�t��ݤWB��@T�\�p� �j�Ym5�p[Ik�i�4P����&�V��Э*�-=��!���I,����m/
"��(��
E�0��$�H�?�
������
��"L4j���z
�^��C� �
�`�@��'�)���� �P��� � P`z��!���EoA4 �;�>�'���h�Ġw� ��O��a�T�V�,G��A��Q��$� �H��B+T��!�j*�UC�S�
P|tQ@0�@� ��N�5S���	� b�PC�D�Q�Z=<8�P�� �7��_�LUuZ�,_5@�P�C�����%=O|�� k�� �TS��O@�QC�����j"z����@�POT������x��;�`	�>1z�$P/�@*�'� ��O��!��z E8
Q�d�z!AT8!��=À��C�(����t@A=~0��~�(i�@�� �+��?�Ղ�����o�@m��dP����1�ZĎ<V2��@��N�[JK��څ�2+�b�ZNґ���HM!)�F�&�Ѹ莻c��+j�Eօƍ1��7X�ҌI����nNL�\vn"ۃ�����R�j�۝ m�ͭ�u ��Fȋ;�=pma��p��n��Omn�;1=�I��5X-���V�xL$����J�n3�V�����A�]e#�;v\=tT���e�9�evM8�b�;L�q_\���Yu��7&Y�t�tgmԚ�0��t�	�W
H�Z�k��f���r%Q4Yq��='�LH��*B�p�r�lV0�iZh�`x�u�L�-��\8T�۱Iϡ��X�уm�˶-������ڒ�B��vv��`����MA[��&Fg/C��=T�J�E&�@��֧��<���L�<1J�P2�Q�r�����3����:�&�mígv��v���<�#r�ݷn�淳��ˮT�Щ���{k�g��6�7F(g�d�Vu�e,�!��H����&�,y!jr*9W��W�6�R�V5�9��&�0�na:yJ�(	��.g�[s*<Y#,R���R�eL�yr�PWUUXv��T�3v"�	⧇��8T�v�gn�<uT�ێ6���K��j�ҝ��sn�� ���T���t&�v�6[���vzcb[=��.1Z�k=�g..,�뭭��ݖ}�Ϋ�P8ky���)�llA�l$p	9���Yl5A�7['E��ق���j�`5��l$7$E:-%�m�
U���#���\��ș9�by�lu���9��:YZ���q%��!�zTЄ>��q��.{��l,u:Lo;BmY��v�D[�unګ.�,S�:�z�cA�r$p�Ql�� ���B�Q*��9s/%F��
�|)Se6�ۍ�������h��@���w`��*�1�n�Г��o2cj�+sNh�[,X�.H{D���;T��d�mب?§� j��D����b��P�O�X(b'tA=�	����#�?���4Ơk��4��������W���2����蝈�ո��Gn�
5N�հ���h;E���S���Vې5j.8p��3��_kq�ҙ�ץ�<��s#�u��Ƴ66�^ ��S�����T����9���#���]�=lM�<�\��;u)���X4&���\���
�<XRB���,u;���Y�w{�w��w���� ʣ��S����>s�'(gv{<'��e~0X6�6��Ő�^�@�{�����/�U�r=kjc���(őJ���u���B�!%
d��`fN�*�@�a�j�C��9�}#�e�L�e�;�"`��g��N��h��
���>W���DD=ͫV�Jk6�QN[���S�"ݖ��\��2GL�ؘ��W��]�*�%���fh1{u���<�(�y��6��.x�\��^S�,1����̹d����0"ݖ����Yfdۚ\��nrI�{��<X�0^�N��Vonu0"ݖ���-��)K�"�Q���{Ϫ�*����^�m����Bz�)H�#qhI-�Ւ[I03/b`��w|�#�yBȤz�ֽٟ��w4y�ZVנr���45�"�$4�Zv���uC��nT;=b;m7lmʖ[���фI���S"�&�z��h��
��@�zנ�Y�	D$I��9w�`f^���Il���H���Y�sŝdƠ��dr-���^����]cN+` �h!lQZ�(<
�m�nh�ՠ_<Tn� ��$��r�Y%�$��2�&RK`uj��G��LLq�۹�w�U�k�ٰ?=͛�B�N@�WT��)�4�)9��,Q˷�vr,�������n�h9���ۿg�@��8�!9#�8�π����*���z�޻���*��<QGRL�;^���M�}�6v��==V��wV���yBȤz��z�m�:"a$�w'y��:l�o[N�)�L�=޻�y�Z]��� 	�D��xW����=�`����t�ʠ�j�Ұ3/b`E6[�$��01�s��R�fڢ��ۉ�\훞P��v�m��8�r�mh	2]����}�}�ڥ��/]��"�-�ܹM��_}U��<�����1Hd��qǠ}�j�-빠{Ϫ�*�^�����mH�a�_M����0"�-�ܹxj�\Y1'r'$���?b��U�Uz��;V�o]��v
�=O�ƪ���`k�ٰ:!{+���zՁ�gݼ�x��@�A[�KhD�Y��!!`4�㵿9��]p�1d������ۣr0ݱ��N.pz�!m��hU�.�:�C[d���-��`��n71�.�X���gF�(�+���G��s��q���ې��t�ۃ]d���nմ�7�mɹ��'nJw)�	��������ٷT��[%�ݮ��c�����,[U*bR�w`�ڮ5zom��?��Rĸ���ָ�W�bv��T�;���+���jۓ��B������AkA��w7!Zu�)�n�9.&7s�&H�HjG�}���h�t�̽��UUuS��TbR�\G		��#�-빠{Ϫ�*�^��^�w������@QdNf����@��z��Z�w4��βcQb�j8�
�W�{�U�[�sAf/�Z��+�DB
I����=Ϫ`I���d�Se�?}_UK�.�gY��w=vX�>��{u�`�9�iH���.Q����<��gÑ�+ͷ����ݠ|�נUz�����j�\Dœwwv����'���9C�&'U��E�y�e�&�5_RGshQ
�<D��jG�Uz����޻�˭z��9�G8H���R�������0:�K`E6[��\�K�酹�y$�~�I? �"�V�O��ݳ`{'5���;�HA3Ci��6ʳ��:�Ɯi���X�t6	��V+*	��f:������^�@�>�@����4d�*�j�u56�͛�I�6w��ݽj��u�@��R�A(dN?����}��'{�xr~TĈ��G���A���~�6>Λ�Xk��䙒��w���c�V�l��`f�����W12E&E#��|�נUz�����w4Eĭ��F�I�@���Xzs�wi^��.�ݧ�]U�]�yy�m�{���&���)1�ԏ�*�^��}V�m��˭z�u�s�,p��5#�=Ϫ�-�s@��U�Umw�!���L��SN�R���;���2�&RK`w.D�4����&U�U3Jâ""*P�Ne�;�gg$�{���!H� ��{�sAl��̂nE�Umz�{+����Ձ�Nk�=��L�n�J�魷����l���.��n��s%�����-�c��n���c�M���g�3�������m�m��=��h[^�����1�Rji�����"��S&d�;�g��>�h�W
�L�HG��f^���l�r�L	6:`w6����H�����
�W�}�j�-빠�f~^���ֱ�8�G�CO���\��&�L�ؘM��߫���H�U���3��nˆlۭ7ɪ	V�t�\�3�۬�]N9�˜�)��]���J�x�u��Z�[�cs���\i�e=gv���=���Hv,獛ո��#�on�xsź��mX5��'j1m�B\L���Ӈ^�ZE;h�J�;)����-�/;FY��xp�ە#n�
�M�GO�6�a�-0]���5�y�X�:ۛC�e�Q���w}���_�vW#qҬ�{B�n�xxݺ���&�3庙݂�-n:�g���1HLxӑp����h��
�W�}�j�;9X5IH,���=��0"�-�ܹM���_$wm�p�6�t'3T�{�6�N���}��4���|�R��K$��RG�w.D��c�e�L��`uj�GZƘ�����o]��������/�����ZqqW�c�I����Nݙ7' �T�i����5�`����g���v��@�GԒB8���}V�U����Z�w4w	T'��R)ə�y$����(b!<�T"AS����"`I#�e�L��]�ZPY����z�v�޻�<������h[^����T�.5�̘�"`I��2�&Se�;�"`mc�D�,��:j�iX���I.���{'�����IBK�ro�:m��͡��m\���b-����Unt]��ɗ\��7�M���u�����??m�ܹM�����ؘn�%�茑)'棏@��ՠ[�s@��U�Uz���9:�4p�qh�xrI��o'�l`G�$H�"��c$�X�WSc%�=�K	��IbP�!a�ĈFI�H:����)C�
�	$FD,V�_E�'hf_��'��I	�!HL!D����G~�"�OσĊ���,�R!ġ�F_�҄(U��E��8'����tS�V�1���+�<j*���| ��q ��I(��7�����/�;gy�興l�'���t�%UU5SJ��Jeo;�oO%�d�;?BI7ݽj��Ѿc�r�U*��P�:���}�7ВM���v~J}�֬��|�/�>P��B���Ԍ���2ೞ�R��,�ڡ���z�T����2gق�UҼ��?�ww�?|��ww~_�̝�g(M����
!?J1�r�Q2�ҥ*\�;�z��舉�v{�g�P����ld�>P�~a��<D����eUU+�D'�[���	GOwO�=����P�wu��,7����
RQСL����wM�l�O�גO����$����CU�~�����?��q��鑨9&5z�v�T��l����7(�[o�,0�`eUz�d���7�V^�e�un�Y�l$n�)����k�I`�@�s@�'7���zl脛�Os�7	�+���K��c�I+��_�=��g(�o�oM��;ϒ_�woZ���<��9��2G�m5$�?���z��Z�w4�h{��,���yxۏ@�>�@���}�����Xr\��r<���R��s������]��>ޛ�����HP�po71�$�EIM#J4bR�fQ6�hd���g��q+���}�c����Np�ݬ�_kl-���u��\h�	7Q������i�h
�����TӶn��]n��ڎ�y�a��y�G X�7Sp�ݔ�av�K��n:9�d���X|
d;\8��.)�\,G
���A*�j��s��N�޴�g�j��i�F�LY;:x�I�n��%k/n�����wa7��e����+��\�^�-ۍʜ�Lu\�;Ӽ��K��N1ٰj�m�ʪ�X�&��������/�3gy�~Q	>�������`�*�J
�����9������(_�woZ���{����}J�U4MUD����3gy��ֹ~`{{������1�s��jf�T�54�gv�� ��U��sf��Nm�;p�R�U	��Tꕇ&���`s����3gy��ֹ/�����ߏ~�9y�=�W��K����]ռ�;��.�9�J�.pP�S�.�b��OYE�U���{zl��vro�zՀ{{������K$2<��m�n=��/���1�R&d����ÒO����Ϸ��B]&4k{2�QSE:�)sT���V�7jϔ(Q���3z��<�\�ƢIy���f�U��w]�޻���u���NF���M�����h�����_m�{����;����U��&i ƀ5�c����t��es�f{�g&��rkp�{���,I��JI��#���-޻��[4
�k�<�
�hn)���7c�,�l�K`w.D��R���E�p�$Rf���@��^�~�ٙ�`D(�@0�	B�P�Lקu���V��z�t�F(AA7����ʾ��yڴ��� ��T���I��ԏ@���vB�IGf���y�6�f́����<;���]�[�l�Ő�nz�{M�x�n�-�l�n��ե�n�\�f�LY��f�`w.D���rw�H��$���^�3*v��;V�z���h:��I�#PĤ�@�ֽ�;V�{����@�x��ɃR(�����yڴٶ�?f͇%��W__M���s��I���o]��~��W�wW�}�j�9w�9�&A)�MF���6Q�a6�l��Ѝ�l��1�\4MǛn���<V�pk$Rf���@�ֽ�;V�{������&�(AA7�Il�Șv:`b͖�$ߢ�H(�)m�#�>�h�w4/uz^���xU���F�<iȴ	�01f�`E�-��f��`E����(��0�<�L�>��
���{+K}�j�BKpz�D�Թ��U�JW3KRp'U=�s����sG�|�6�o��sU��^κCf�9K�d���]!,Fq� �؏\�neg�m���V�i�lu�!ء˹;;U� ��8�z�vs�Ξi�n�WZ�^0+�*�;���Z�q��ga.�p�w\
Y�7[4Ҝ�K,���G�C�.(m;s&t3]�L.��:�v+k�n�=�{�I�}��M�4�±���vY���.5��6�n8� MY\��ť5̙z�Rt8�ʹw�&��[���f�_��۞Vd��M*CuN�����?{+K}�s@�Ϫ�*�W�|�����K���	�0;��0"͖��o ����`D�cy!�)3@�Ϫ�*�W�{��/���>���'�y.Z��`E�-�w6q�2GL��L��v�;�����㑩�0&�C�st)�l��	���k�s��ʥؼ�.ԼQ-�R= ��f�}n���U�U�^����T$q�Ŏ9&�}n��{����U�`� A��T@��{U�W�W��������`͜`j�K�����T�UU+��5��6l�	&�f�X�֬���j��r:���+�-�l�e�&H釪��^�Nvl��M*c*��TK���5�6l�w4��hwW�y{���F���mŵ�}c3�ɻ���@�m/�.3�"�)�K�y� �`9$�~Q���w4��hzנU�@�q����X9sSJ��Nk�P���wM��7���͵͝���wNd��C�s4�{�6o�w9<<R	�0E���xrI��]�fF=*��:�S2��M�C���;;�X��v	����k�/��Z��Ja�����VDvV��<ޛ�uzpc�L�4�Q�����7u;�u8�uk�St�Y�#�z�;R�~�o��e�D�b�0�<�L��w�hwW�W����;7�X�^��S)�T�T�0"͖��vyl��==�L	��?${e>:iSUS�jly�6�v՟%���=�>}�M�����e������SU6�gw�`vN�5�l�}	ŉ~ �r�@?�?���g$����3̦�9�MM+}9���ul�������w4#�s�1(܀LkT�l�w=uI��"M�*�ns/EZ�3�5ْ���@[�<�J6�_���=�v́�͵�$�K�������T�7U53*j�l~͛�D$�IL�w}j�ϧ�v�n��&�5���U-UK�0�jl��V��g��#W�~�l{�M����gU9M5T��*��XtB~��v<��f������+����X�	"fȴ
�k�?�2����;w�X�s]�ԯȸ�"=BBP(C�k!�c��G�C��*BE�	I�b`���X�
���� b�`�� ���
`1���,���Q��F��@�# ��- �+�ˆ���HK��)����^X� 4�X	�EH-D�!�b��0|�X�C�
p�V1	eZRT��B�
N�bB1`HL�B*b� �|2cF1�!��.S�,���0�A��,�$`D(WT�L	L�S�q��$bI$O5�cH2H1d����$�"��
���L2��2����B�H�j�B�!<��� `z+�G�%*,
�.I� �Fa�pO5cP�g�z,uN�AŔ�I�����!P�M Pr,���&�������GP5>��3�7ww33t	$ �jk�[�$^������0%nP�'N�uղ]�۷�}WR� ��Y`(�]:��ب
ړ$F#7J��k�4��e.�!l�M��I���{woe�.�e�9�\�ݻfU�|�V�v��]���Sƻ"3��dqE�P�q��HGu�j1Ÿi��)�K�N���eF�:F�cg��f����P�m���9tj�S�'	�:�:6�j�<$bQɝ��v����W)�]�Z�s��gb����۶��"+������:�T�/A��S�;mkv-�r�,��:�̀�-ڶ��&�h^�H9�V��ág`�)-���nT+�3��L��$ ���;�eu�9�\��ەv$GV�i@��-Ȕ��n9�������Z�iV���qj� �=�-E���taD+�:���iIJ�&t���F����*���ct�7R mco'\���Ȁ�GY �N������H��]��s��g'm:悮m^u�Uժ�(�^h;=h�<�U>@&A���q�m���u�y��ᜲ��l���U-���� =�x
���8
��UUl��-2��Im��.΀X����O���/'3;x54Y<��gqvM�k�U����N��w��B�p $
�5U*������
�y@�{e�İm\���%m�3F�����qrJmm��@8k[�-��a�m�3m��I�N�u����v����k�\�����)�������EF�@��2�m��	&F	 d-�fY%��6t���@\L�v���v;`��A��xt�?Lk}�Ӽ�w"e��S U�h��f���⃊ܛ]qx��`�.4� �]
c�0��x���J��S�V�����9yek��+��F�r�(���+�1��`;	�S����m��A��2r[q�KI�s�n�ju�����IGA�ƻi�y_e���,���.Ŋ~AJ����QE�_�u�&���~ȇ�w��!��4�f�et��
�vY�Py.�Gjx!{5�u��(^�i5��q��"3hI��9����#6�&u��kC.��ٹ������]���糶�x�N������۝�|�$�*z���gnL�I�Ӟٲm;;8�
�4.�a���H�8��Ȥ��i��s�\���mK��8U ���X��6���7W�yf���������w�OWMo�m}�v6��.��� v��c2�vX۶�##�y��R���;.��0�&�%���9�}l	�0;/b�Uu�����J��
j���MT�����D%)/����}6�>�l~͛��|�L�R�5E]��L��&Y%�Ԕ[=lI�L�Įb��"&�Z^���e�&�釩g�<�~��u|�\��̩sS`c�l����}�~�;����z�ܲ;!�6F)��28�i�m��<�����,A���݋q�c��N%G��-�2F�?�8�z�hW�hz���]��U+O�"�I���rf��ϻy��H	� � |���$*�^���^�o]���բ	DHH��E�Uz����>�߳�]�����⥐� �Q�i��Y��lt�콉���������1���d��?$��޻���ZW��;�w4��d�jA�MYkrr���nL�n���rN��d��U��]���"Q'�`�1�&hW�h^�@�f��
!~a�[j��boP�&UQ��w|L��`nlt��c�e�O�I�r5��ML�J���S3S`noZ�7smY���(H���;������8�&5�51�Rf�o]�������}���@<��Ȧ,L��<�L�>�����Ϻ=׮�o]��\Jꘖ,l�12%��J#�w[�7 tV�vv��9ݹ��d�Y��v
MJC�ZVנw��h۹�}_U�_<T�0H$�n=��s@�������k�>\�.���G�|��:`v^���(�%�76:`r�qؔI����MI���ZW��I>�����$D��H���{ÀweW�Ld���Cqh[^��{o��wwZ�?l�V���.�Ҫ���K;$���O5�RwF�Ԗ`��a�sm���A��LSl���7#�>�h۹�{Ϫ�g�*�^��<���	���r-޻�����k�>�h/redS'�L�L�=��h^�@��ՠ[�s@�a�V�Dۍ���E�U�^�����m�����׊�BbHJ@�8��>���<�^ڰ=��v�ݛb:�8P�	3���v��}����9��u�q22�HL�z���N�ػa�7Z���63t�<9v㱬n�wh��>wf'5j�`8��d;!;s�xbS���V�j���:�ZS�p��ݢ��ۅ�{i�;�tnsHp�,:��'[e���ɘU�]���T@r�V2�*��&�@��]-rZ��Cn�1Y�rl�(���x��	��TL���Esw�L�f��6�˔D�".+���ݾ�~��2݁�\ꭓ��S{r�[��nO`�x�iγ��uM�[%�7N<K�4��Z�=��v�͟�D~a��`y��=N�*G35B���`{Ӛ����Ϳy0$�遛Z�
��˙�47�U����Zy+n�h����|�����{Kᛙ&]���2�� �`�`�`��������lll~��Â�A�A�A�A������ � � � ��߿g �`�`�`��t�����n�7r�sv�A�666?�~���� � � � �������lllg�߳��A�A�A�A�����A�6667�����8;.�ܛP	p�אc��
�	�gs��t0!����]:GL<1�5�w���lll~�{��A�666?������ � � � ����x |A`��A�A�A����8 �p�����vۻ7iw7o �`�`�`��?~��|��& �A� � �����|��������� �`�`�`����ׂ��D��A� � �iO�ٰ�n�f\���>A����������lll~��Â�A�A�A�A������ � � � ��߿g �`�`�`��t��~�$����fnm���lll~��Â�A�A�A�A������ � � � ��߿g �`�`�`��������lll}��L��e̍�ܥۺpA�666?}��x �?����g`�`�`�`��w���A�666?�~���� � � � �d��p��)�a�Ssq�7R�v�]Ӻ'��<gy�O����!�����{�r\.�nܹ��� � � � ��߿g �`�`�`��������lll~��Â�A�A�A�A�>�����lll}�;����.����.�pA�666>���^>D���A �`�������� � � � �;��8 ��������lll}��~���7r��t˹wo �`�`�`�����|������g �b��^�R<A�>��?��pA�666?���ׂ�A�A�A�A�w�'��t̙�.�ə�pA�666?g���|��������pA�666>���^>A��C�A����ӂ�A�A�A�A�	�~��ɻmݛ��ws��A�A�A�A���~�>A���߷���� � � � ����� �`�`�`��}���� � � �������n�k��&�H1�{SɎ���NU������{vy��k+�p�\j�v����|�����o�ׂ�A�A�A�A����>AJ�x�zl}�6牧��@���OÎ-�w5�G������yڴ���b��H����y{��"�[�r&�:`f֩B��e�D��˚��B�!O���M��?|���V�\%��BK��e����o7rF��G#x�@��ՠu��h^����@�q["x����&۟��a��I�K�.y��0��M���ݪ�M@���{��}+�#XI�jE����s@��W���� �?��r�3��F5#JD����ٳ|���=�����W�d���L*�uESM�T��}�X�;�ϡ(�������V���ݔ�֩��k�1}�j�-빠y{��m�˱g7S��H��8��-��l�$�`w.D�������U}����~~���c�i����qM��]�ճ�c�G`L���+�{7I��f�F�m����;�I�r���</S�'�r��ާk&I�r����r=�z���?︃����b6w[m����[^�pR�P���^��U�S�Iٰu�Rs,k%\�q�v��-]U,m���M���Gc&��n�.f���Lm�]��噛vnC.:fm�g�?���y��ǿɎ`��h�����3a�6˹���Y�u��v�Nk�ln^A�,�S\%ʀu~���q�ܜ�I03kU�=Q��&�zm�^$}�)�[�s@��W�}ߎ�'��j�����v:g��l��{��=і6�F�Yp�-�s@��W�����s@�{�; �iI�Yw�S�l�7g�0&H����;�ۿk��3��9���ۉa��l�ќ#�[pt<
j���m��\�[��;|}���
BE�I�?����빠_[��|�W�Z�p�P��G!��&��빽	%P�d��`c���ڰ?<Mcu<	$�O�73@��s@�^�@/u�{���r�A�$rbjLп�nl�Y���0&H�ܨ�b�'�$�M8�
���;�w4�w4���,;�L��$q%�tM�k�P��݊xdq�	���ٶ�	���2\^�$�3�r7�H��]����平п0��`c�rsu5�74���Sl��Se�"�-�����H��c�	��I��4���
����j�F� A���z���ѲB!(1����$����$�OC��W��a&�H�HL�<zB
�(a���M �q��@<�	$A����H@Y��N	��B��.�D�x	W@4*_�T�A= ����?#��� @�0O3���9$�[��|�K�� HH�)#�*���YM޻����׊��܊8�mH��e4�w4/uzW��<��W�1D�X�E���3�r�s��i|�q��+���n{\�t����_���&�LY��M�����9��c�A���18�h^��
�W�}�)�[�s@�p+�أm��((��*�^�����o]���^���u{�ơ��=�YM�m��ٳ`�D%J�Em�l����R�~K'0J8h���<���^�@��S@�0�l�`ӎ8Lc����s���grn�q����tۚ�4�/Z��X���I��I��4/uzW��>���-빠}���b�$$X���d�����7c�T�l	.������q���-빠|�W�U�@�rn��'R~$qh6:`b͖�&I�r�L�R��b���<����Y�}��o$������ �T�ŉP
�T�Q;�&��f��vvV����^�"/n�f��x�<�;�t���t�J��c6���X̮7<���l�Y������v�9����Y�Cr>�cp\Ҫpn�"F7�Nv�t{	��݊�Y�l�l���VΩ� f�ű*�vL��[��ی욘��/��VL/=��t��tv��
�������h�a�eD��ծRL��ܧ��@�n�����n�w�o�_����J#f�1a���m[.�Ļ����c��	�3[1��0�(�m�IAG�[�4��Z������I=����=�;Sn�LY��d���Z�J_>K�LJE�^빠y{��*��@��ՠy{�7bM�JH�K�4/t�Y%�;�"`M���ۥ����F9�,JH�
�k�>�h��h^���\U��G�H�?�77�Ý�[�[!���X5�6��<�칺�5m�,�k7"C���|��-�]���^�W�zːsu<�OÎ-�]͵�/�B<�(\��Ž��M���ՠ|��!�	!)���^�L���Șv:`f�(	�]��P ��B�^��>�h�L�|��=���I=��H�drhyڴ�w4/uz}l�>�rȬ�(����yT������܆�r�[��:��uɤ���$Ҏ~K�0R-�]���^�_[4��Z�{�l��"K�"��`b͖�7$��r&M��p��1a1G�Ĝ�@;���g{yZ��`� �AH 1V �PK�~�I=������h�Y"nD�15$�>�h�w4/uz޶h.A���#�)?8�6:`b͖�7$��r&r�G��cs��]�<\�r9n��ۓ+����hQ�퀳�&�u��:�(y�x��,�ld�`w.D����7APOSLmQǠ���;V�{����@�~�D���H�%��Șv:`b͖�&I�*Ե��hC�
C�v
ow�`c���ڰ��q�
'η]�潓3����H%�$���^�^�hyڴ��h���X��dM�8��e=�u��[���`��]�"%a����q���1�JH���@��ՠ^�s�?0Ǜ�`wJzL�UNf��br���\��6GL�ؘ�q�ը5\�9"��#�@����}V�^�hyڴ�˖B$<�"�Rf��9 �N03.D��GL�B����Yȴ�f��;V�m����Zf{3����`�?'2H�� [m4;���oW������ ��ֱts��0�w�r��s[�E��q���k[n�N�������ہw]�];aB������l��nҞ�]�\۶��@��s�Qb�[��q�n�Eg�mT����٠�nֆ���!c�.{�,���g�ݹ�m���m��Վ�<3m�VW�S�t�f2�!sk���Zy���������oNhvi�-��)"�^��;��e�Ԓ�V$ث�ۏ������n��K�.s�v����GLˑ0	$��k��P��RL�`n�ڿ�(��=������̭,k2fv���D�93@��V�[�h�)�u빠^h:�A"8�A6������4��hWj�:�Tn��NHưrI�wt��m���ڴ�f���݇�/����ǒ5#y*�t�s��.^��f|\i�`��l��cw]ŞP�>�Ҫ��uT~��Ձ�gu��vlΔ�<�vY�2GF����[ C�O�F�b��e���[�� �ٱ��@V���ڮ#�h��@���@�n��;V���ʉ=�OH�ƤzwJhmt��T�����.|�+��K�L�:`f\���Ilˑ0�b�Lx�5 ،x�B���1[��=�q�q���8�2��ф��c��į7\u��s��e�LRK`w.D�ٱ���`�#��i����z��Z^�������F���k-r�l�Ș6:g�-۞L��[�س���G2I?����h���{�6	BO�]���O)]4��&^F�9���������:۹�\G��,���R8�o�3�i��l]�L�-�u�[����a��ܾ���Vנw�S@�n��}V����{���)�H���Z[03/b`j�[)h�|�+�1)�����}V�����Jh����r �Ln$�&hWj�9w��I>���䐤�<8���g�~��*�`A�"r&�Z+k�;�S@�n��v����왶Q5%���cA�y,�����n.8�1۵�&���,�Ն�Y�������:`v\���Il[J�\/�$#��rC@�n��v�����Z_&���+��L����UMM+�sɁ�l����:`w �B���P2���r�	���7v��-빠}]�@�~��'���I�Ԗ���A�&�Lˑ0"�-��}��p�5 ���W�����P>~��cP��	�b9��"F]`(�@�����B�B�HD�T8���Ed�A$����  @�0B��X� ���%Uی��$�d�,D���<H�-K�+��bAbCtc�拨���$YEB��)p##����J�*@��V���B<cp�	F Pv̥`��V	�~E?:����Ʊ�Ka}j<����H�!)
��H,��P��C2�D�dJg�_~���{�ݽo�~ݾ��	8�Iiլ��IF��[50��=��W��5&�R�nIm�*��&&��L�ԥ�.v@�
��� ��f����b�6+kҸ�/O���\�il���ۢ�n7��r<�E�8��ݗ^�%��Џ$
�z�B��2�&1���b����s�����6	3T��$Z4q
�ނ.t򍓓�`Ȟ]m���9�J�=&�1�YJ�[F�Z���1�k��m�5R �$�$�Q���E
����[��x�<li8�0���.6éG�Fw\	�иwZ9덊W]D��R�y=Y	^:��<邴u�nxyx�x�L�S۶�T��e�����f�7l�N:��r�9z�T�k ���հn�n��j)H�:��n�� �:FP("�8�#̅]Lv��V�ݸ��J���meT-,�
����Y�]\�i�U��3�����X)X���ZL��lY�q퇩�+�OI;fs���S�6��+�{4����pj8i�X==Z�����ʭS���n
�ڪy�\��0��#����.��r�M��8M��<@�ٺ�*�Ma�);#U�.��2��p[@��f���{l6[K��%�%9�k��|�jZ�ng��#t!�mj�`-�����v	$-� Am��`�Y����7�q�:�핌pմv�&��:��iN�]D�E�5l��$,=�m&�i��4����\ޠ^��FB�ڥ�uȉm�թ�b�޸�n�v���s��89�f�%^���^j����sn� �J��dm�e��-�WL�2�hg�Gl��T��8�t�m[c���ᗔ9���XÌ���*n�qd,&6��I��%���e)Ikڍ@GWS8��8�ڨ-��R�A�՞�y	�ی��d�P��&u��$����WU)��=���ư�lv�����׫���Ѯ��npv�*���r����u�s���j�p��@W�S�����LNy⨧z��ʎ�P�����뿈>�����v��B���ч:u���M4��y�<n��4�䇞Ԧ�N���v4�����]�mHf�����r�b��VL����`srY����y7b�	v��8��09�M�ٍ63صcp�l�G(t�0�23g�@�qM���68ت�[�I�5�q�G[���łr�]
v�a�R�6+�L�W9�gx�إ� �&N��;��&ЗS��q�L��F���+�z1S�xcI�b9�n�u�q��r&Se�ﺂI����z��5�X���}]�@�����-�s@�����I�9n-����)�[n��v�֎MՒ	�K�=��4z�hW�h^�@�v,���8�O��޶��;��7sj������P�6v�~�s���;=GnR�g/tv��2�l�q*��]0`�<=V�L�T3w�z� �g��0$��܂Qm�nZ�d�3N�7sj�$��]
/�".!BK�$��_U�om���뾈P�3c���MKUT�GUV���0;.D�$��iV�!ϒ(C�M�@����v� ���;�S@�sr0�$���4��h�f��Қ�w4�m� m#p6����ކ<�g�.l�zg)G�x�Hp��"@�5�@-�4̭,��\�DG���vt���5T9���Ӛ��3+K��ݽj��;��޳@�v,���5#��#�I����y������WH+U���"I+IAgv�X�\X�ꕵEJ�L�uT榕�$�BO�[��;����t��[�hz�T'��M8���L��`w.D�$��eȘZ.;�ǺZ�k��qڝmj9ۘ��;"e��\;=�C�f��^�a�fN��)`f\��I��ˑ0"�-��U�����D$��z��v�����o��H�X���b�@uU`fOs�5�l��	7�=��;{���%�,a&H�qhu�@�����N���$�PtP�{|�o$��G'HH)$m,n8��������5���
"#ӈ]+�GLv��Z7:}�7�����5r�n��X7nt��\����T���S4*��? v�U��g*�*�^���M�w;�Cq)(nj��9��DDBM���lͮ,��@�9T'��)i��ŠU��sy6N0;/b`w>���.5�E1����M �l�>���*�^��Yպ�����h�e��g5��6l�V��5�v���k�eSc�PZ���t;nՃ�+wlפ����뛱[a��b��fz�;��^ϛ`p�̓�����}��3�v��z�)�(+A�.�q�Jn�
�<��ܢ���!au���M�Z�˃��j�q����r=�3z��M��y\8m�dۘ9���뱃��Z�V 7Nx������,��x�|�"ڞ����;s�ջ#4]Q� ���2����k8�ɬ��rF护����HJ��ٜH��"G�8_�Z]�����f�W%�	a�$	#Qȴy�7��76����?l����բ��b�"�����z��@/��_ߒ��wW�|����cm&bo&���;߻�O"X�%����֧"X�%�����'�,K��}����bX�'��L3�n̳3m��s7x�D�,K��v��Kİ�������Kı;;��'"X�%�{߻�O"X�%��J_���f�%�v\�X��7Q���l(�tSm�8�\ِ�7\뭮�����˔�ݵ9ı,N�~�q<�bX�'�����Kı/{�w�����~��,K����'"X�%�����Is����7wL����%�bX�O����r&D�/{�w��Kı>�{�'"X�%�����'�?y=���w��Vo�f�!��w�3*dLʙ����O}��3*dO�{�*r&eL��S����'��ș�2%�w��r&eL��S�I��,�M�4��e����ڙ2�U lN�?mʜ��S"fT�����{�L��S"Y�xn�"fTș�3����{�L��S"S?�v�j�hOw�ܧ���=��~��=��D̩������MO"fTș�3�~��O}��3*dO�{�*rB�p��2�f-Od�)�R���%�4��5q.�uc�ݐ7p�vcvv�]����-�1��M֗v�n�����dLʙ���592�D̩�{���jdLʙ������Mڙ2�}�����2&e�;��w���碒�Cm{���=�Lʙ����=��D̩�>�����Lʙ2�{߻�O=��3*d��&�"�?ʯ9�ș�>�?�3�mܶ�m��2���jdLʙ��fbr&eL��S=���'����*8���t8{�NA��jr&eL��S<���'�ם�S��w����)Q:i_w�3*d���ݩ�~���{�L��S ��𚜉�S"fT�>�w��2&eL���w3�3*dLʞ|ϻe�B�k���.n�=��D�S ��rMND̩�.S�G}������2�D���̩ș�2&eL�ﻼO=��3*d�o6��DN.�p����]�eA���V����u�����J��J��݌ݭ��592�D̩�}���jdLʙ���ʜ��S"fT�~������lLʙ���592�D̩�I�rY���]۳37x��S"fTȟf�nT�?���ؙ�3����=��D̩�{���S�3*dLʙ����=���E �9��Tȗ'��۲��nɻ�w7nT�Lʙ2�w����{�L��S ��rMND̩�3*g�w���ڙ2�D�7�r�"fTș�=���gf�ww3wm.n��=��D̿����<�S�3*dLʙ�~�'��ș�2'ٽە92�@���S� s����?o�jdLʙ0�s?arͻ�vnl����S"fT�>�w��2&eL���P��y��*{2�D̩����x��S"fT�?w��S�3*dLʞ�~�C1���5!&$���ɕ�Z��D�䆊�d,�3f�乧�h$0٭�3w��2&eL��ov�ND̩�3*g�}��{�L��S ��rM�<��S"fT�{���=��D̩�/��L?lI�(Ow�ܧ���=�����'��ș�2��$��Lʙ2�}�{�O}��3*dO�{�*r'�'�)�jr&eO����˞��˻n�˛�O}��3*d��䚜��S"fTϽ�w��2?ʐݩ�;��nT�K�2%ʟo���'��ș�2'�os75����.fɩș�2(�ݩ�����y�L��S"ww��T�Lʙ2��߻�O}��.P�I�{��$��Lʙ2�M>�˓�L�4��e���{�L��S"}�ݹS�3*dL�~ O�J�������jdK������bX�%���x�D�,K��	ޝ������[~�E�:�vh��s4+q�f�v�mY�;���n�3���*)ybI���^��K�P��J�gd��f�$P����E����l�D8�Ӝ��c��Dg��h���ˠGlv�GU���}�*����4e��Yh棶]���gؘ��r�u3XV^6�g�i���,;��)�9։�<V���%���Ͷ�a���t��&D��qۅ��{��ϝ_�r�]�3�N��7�؋�6곷��q���T$�e��U�;=[T�N�}��K��?w�q<�bX���ND�,K��{��g�2%�bw;�r'"X�%��t���n��ٷm.n��<�bX���ND�,K��{�O"X�%��}�Ȝ�bX�%�ﻼO"~@ʙ���g����.��S�,Kľ����yı,O���D�Kı/�}��yı,{���bX�'��L/t��˛3wd���yı,O���D�Kı/�}��yı,{���bX��=��������oq���~���@
n�Ȝ�bX�%�ﻼO"X�%��{�S�,Kľ}��Ȗ%�b}�wr'"X�%���6}{�nL�7e�얶��<�;Pz�,�@I:�Ca�#��c`;N�dq�t��s&��nl����%�bX>��59ı,K�{��yı,O���@�A	�L�bX�����yı,N���75����.f���bX�%���<�E�@X�`A@�S�0 �a�Dؖ's��"r%�bX���x�D�,K����"&TȖ'L>�e���ݺ]۳.n�<�bX�'s��"r%�bX����yı,{���bX�%����<�bX�%�v^��Ra�mݷsw"r%�bX����<�bX���ND�,K���x�D�,�?�b~��HVBd&Bd.�O����UNf�Nkwx�D�,K����"X�%��1�~��ObX�%����Ȝ�bX�)�f���Bd&Bd.�-:��D����<��[���C�s/M�쮗7q�C�vu�����8���z�:_�̵��[�w�����D�oȖ%�b{�wr'"X�%��}�s��Kİ}��59ı,O=ޘ^�7.e77fKww��Kı=ϻ���_�k�6%����gȖ%�`���ND�,K���x�D�,K���;�r\�ܘ��Ȝ�bX�'s��8�D�,K߻�S�,j�/�m��hF"A�Ph��8+��$dH$����#KH�0� ) xcxB��y��� 1���5H�D�-�1b�OS_�#!5[��|����0?@�)�O,0q+�Z�D�B&)�`�A=N"5<Oz�b�衈�ʕ�	�~A�!������/����yı,N�{��,K��׷�\�-�r�n�ws��K��`d���S�,KĿ~��x�D�,K����9ı,O���8�D�,K�>���m��k6KsMND�,K���x�D�,K�@�k�~�܉�Kı?����q<�bX��w��"X�%��m���s��Yq�xn��]m��Z�S �lfdR�d��7���맷J��u1��sw��Kı=ϻ��,K��>�s��Kİ}��4?$�&D�,S����L��ONo�SB�sHsnf�D�Kı>ϻ��yı,~�ND�,K���x�D�,KӛRB�)p���]���(�US������'�,K����jr%�bX��w���%�bX���܉Ȗ%�bw>�s��Kİ~fvᶛ�n��f���bY�?w���yı,O���"r%�bX�ϻ��yİ1�؉�OA�DAd����"X�%������n\�nn̖��Ȗ%�b{�wp�Ȗ%�bw>�s��Kİ}��59ı,K߻��yı,O���a�nZe0�p�'�ys=�=ѻd9�MA�m��[�շ.έ��=��ݞH��E�|�����oq���g����yı,~�ND�,K����<�bX�'��w��bX�'�=���s70��2��Ȗ%�`��xjr��DȖ%�����yı,O�����bX�'s��q<�bX�'�}ٛ��L�l�暜�bX�%�{��yı,Os��9��0ș�~��8�D�,K���Ȗ%�b|a��&N�f�v왛�O"X�*@ȟon9ı,O�����yı,~�ND�,��3��߷��Kı/g�i��幦�Y���ND�,K���8�D�,K�߿xjyı,O߿s��yı,O���9ı,O���EC��������ϡ�C8���1fH\�,)j�e8��cQ�\J��SH	� &�d��Z��*��[���n�\��Ų�:w2��j�<ט��q�4v���q�#��9q7�\,��L���W3�U]��3dRm�R�R���a�D��#n�0�@��8��l����T1k(�s2���g]N��[t�rt!����5v�D�l�J���#v�&1�m����i�&��۞�r`������Ӳl��UNf�S559HL��LQ�p��Kı;���Kı>ϻ�@��DȖ%��?~��O"X�%��)۟�i�6�.��S�,K��{��'�,K��>���,KĽ�{�O"X�%��{�S�? ț��,N��/��r�Jn�.l�yı,O���p�Ȗ%�b^���Ȗ%�`�����Kı;߹���%�bX��nYs��	�v\r���,K? 2&~����<�bX�߿p��Kı;���Kı>ϻ�D�Kı<���<���3tۻ�O"X�%��{�S�,K��G��y�q=�bX�'s����bX�'���8�D�,K�v���e6ɻ��5�L�k8��y�m��/T�������75����e��S�,K��{��'�,K��>���,K��w��'�,K����Ȗ%�b|a��&N�f�v陛8�D�,K����NB
��A�R�����ؖ'3�����%�bX?w�ND�,K����O"X�%�}���M�ܷ4��37p�Ȗ%�b}��s��Kİ}�xjr%��!�2'~����%�bX����"r%�bX�wo�;6m��s6�3ss��Kİ}�xjr%�bX�w���yı,O���9İ?
	2'w�����%�bX=�'n~�m�웴�sMND�,K����O"X�%��}��'"X�%��w��'�,K����Ȗ{��7���}�����:�b#0�;%j�^�����m	t
h��a�.Y�<�<Wi��칗6q<�bX�'��w��bX�'���8�D�,K�����D'�2%�bw��~�O"X�%��Ys��ͷ��D�Kı>�����%�bX>��59ı,O��vq<�bX�'��w�����,O?��.xٛ��7tۻ�O"X�%����59ı,O��vq<�bX�'��w��bX�'���8�D�,K�>���m��k6KsMND�,��������yı,O�����bX�'���8�D�,�@������Kı:a�ܙ?7f�v�e͜O"X�%��}��'"X�%��w��'�,K������Kı>����yı,Oʿt�7��%�.k�3I�#�q���D�'��OL�|��N�v�,�����/,��6Cr��s,���'�,K��gȖ%�`��xjr%�bX�}�vq<�bX�'��w��bX�'��}��2�ݹ�i�����%�bX>������DȖ'{���Ȗ%�b}���D�Kı=�����'�2%�ܲv��ۻnf��f���bX�'{���Ȗ%�b{�wp�Ȗ?� �"dO������%�bX9�j�Y	��	�������ʒ��33gȖ%�b{�wp�Ȗ%�b{��s��Kİ}��59İ"� W��J�h �D������%�bX�>ܲ�L�3f칐�w��bX�'��|�yı,?(������%�bX���~�O"X�%��}��'"X�%��vR��p3336Mv��Kc�e-۶����p��h�(�_&7Y��b�;5�f�L��yı,~�ND�,K���'�,K��>���U��bX�'����yı,O�����61����B�!2!fw��O"X�%��}��'"X�%��{�8�D�,K߻�S�"��0PBզ��NG*f[sP�P�BǽR�$D����D�߻�S�,K�����Kı/�v�I����r���"r%�bX�����Kİ}��59ı,O��;8�D�,ȁ2'��ۄND�,K��N��%��ܴ͹�O"X�%����Ȗ%�b{�y���%�bX����"r%�bX������%�bX�A�Ϲn?�g��`+��\�)�3+�[e�pm�&9r�\na�6��ڳ��!�V�:zxv�vX�rB`	m�ZƧd&��6-�e��������u��2��|t��������c�m��Xj�vԖԆ��\�v׃���˽���|�["�g9aŋ�+4٦yZXC�Ӌ�Z����Z�LLَJ�6oaYnZIs��]����ӛ�MyЎ��n�ɺ��[6<�\�q�m�����`ݸy5Z��~���x�͔����T:��P�Bd&Bd-ξ8�D�,K����ND�,K����'�,K������Kı=���;�]�2���L����%�bX����"r%�bX����q<�bX��w��"X�%����gȟ�r�D�?ܲ��Y��p�!.�9ı,O���gȖ%�`��xjr%��ș������%�bX�gn9ı,O>~��<�I���f�w8�D�,����	C`�����"X�%������O"X�%��}��'"X�%��}��Ȗ%�b|gݙ����n�2�sMND�,K߻��'�,K��>���,K��>�s��Kİ}��U
�L��L��
�j�L˪����Ԥ�@�Dl�nM�/[h�Uـ���b�Ϯ��^/�wrp�̜�K�7mٚe͞'�,K��;�p�Ȗ%�b{�w���%�bX>����bX�'�w��O"X�%�~���Le�i�2���"r%�bX����q<�������L�`�p��Kı>��~�O"X�%��}��'"X�%���O��f]ɺM�����yı,~�ND�,K߻��'�,K��>���,K��>�s��Kİ~��.vi&����nf���bY����Cbw���Ӊ�Kı;�����bX�'��{�O"X�%����Ȗ%�by�yl�if�2��)��8�D�,K����ND�,K��@�y���8�D�,K���jr%�bX��{���%�bX���sm�Vt��t�Jxz�܇c<c4��5V�sv(�,��#[]I�E	�û��r%�bX�g��q<�bX��w��"X�%��w��O"X�%��}��'"X�%��ײg�	377L�6��Ȗ%�`��xjr�X�L�b}�~�O"X�%��w���,K��3vn�!2!b��u5�jh	c���"X�%��w��O"X�%��}��'"X����� ��@�<,O�g�gȖ%�`�p��Kı>0����.�ɹ�fi.m�yı,Os��9ı,O���8�D�,K߻�S�,K�����'�,KĿI��2�ne�ve���D�Kı>ϻ��yı,?�O��zj{ı,N�o���yı,Os��9ı,N��{��4�-M��Mr�}{����6���bKj�ɜժ�&ol�6�BL�g�w�{��7�����Ȗ%�b{��oȖ%�b{�wp��Ry"X�'s��gȖ%�`��s��Mݙ������"X�%��w��O!��"dK�;�r'"X�%�������%�bX>�����ʙ�������.[s0�Җ��'�,K���܉Ȗ%�b}�w���%���2&A���jr%�bX�~��p��	��VT��˙n��r ���,K��>�s��Kİ}��59ı,O{���yİ?�<T����D��ۑ9ı,O����͛$���7r����yı,~�ND�,K�o{x�D�,K�>��ND�,K��{�O"X�%�����-�����[s.ۛ�S���P�t����u�N��T��I7sm�4��Kı;�����Kı=���D�Kı;�w����ؙĢ�޵P���L��[+^��:�.��S6K�x�D�,K�>��ND�,K��{�O"X�%����Ȗ%�bw��oȟ�2�D�/d�i�s.��-�7r'"X�%��;��q<�bX��w��"X�%�߷��O"X�%��wr'"X�%�߶�gf廙w6�fnnq<�bY� �����bX�'��^'�,K����S�,K��?o߿gȖ%�`��s��L���6]��S�,K����oȖ%�b{��ܩȖ%�bw=�s��Kİ}��59ı,M4"qRh��UK#Q6A�CY�
ЕX�W~j����:��C�Y�c��'�x�Q)M�H�RG�� IAM�<6�h�^$�>��O�T��b�	 S��}�n������n߉�'V�0[�qlj���66���`��ui*:��g�w<�ha֩X)iV7c��]�v�j�ZU�Lƶeq2ʪ)�[��.��E�.N#-��y�s��{C��U�3N�-u ��Eb�'m�6�fO\���hu��.�u�Z2=m%�ǳ��"WX� 7I �i�eΫV<,A��=F�;tM0sg�T�:�<ӷY��oa�+5��2Y��hs�;�p˞+�7b|��[bSd7��Ҍ�劕ʆ͉�����"O�a$!gZr�CI�;lbb݅z�n������j��5��u�_^h�cqȬ�Uu�/S����92���	��.�ҫ�R\��pkm��rdƸ�ϡ���Ԛڍ��R��O�+R�i��I7M���U���hZ쌣�i�Um�����P��=���m�)9�Q�A��6�`g��8��۱8�gU�ۈ9�[��,x.�q���{l��=�6q<n�עq`���n�M�R�""$�h޶��CnUuS�.��s����Ѫ�F�r\�ݶ����p�rp��mn��+��N�:O�`c��M2�I�AD�� .����� -�]!�u+���X�s�$v�k+���w$�����b��ڐ�`6ݪ�P9��j� ���h�!ٲ���)���PE=��v�t�l bU$1�׫�8�Zu4��YM�<4Y�l���4������ޤ�2I��q����<6�[6ݣq���ng9вI����n��l�"�ݰ��m<K����9#uWH;T���n"���u,�UW;h���n��w)�@v�f2�;�{Wh�Dk�0�Y�;�\ny�%����� ��6 +A��D�+-�����sY(��_mu.Y��J�[7n5Q�H�[��Y��Ob�Z��@Q����;h����Qm�ĄŽ6-ݓ�r��n�[%��.3nݘaL�̤�w!��	���>@��� �NEUSU^�>`��
�p�S�w���������Օn��t괫R%G���x5��v/��V6S�A@�a���;��g��y'N]Q�ٶM�7kkcpH�n����\m�#�:��N;�=m��np��[.���Y�v�y�l�ܕΫL���G�UW�s�!����U��vn���6�;������;F!쵧֦zsϷ�v<�EJ�Ն��L���&d�k��d�2n�*�৞��չN^��N�[f���/i��	��8Ir^�j���6 ��=W(�>�bX�'�w;�9ı,N��q<�bX��w���'�2%�b~�ޛ����L��\���z\�u4��ʜ�bX�'s��8�D�,K߻�S�,K��{�s��Kı=œ��Y�B�
HL�����E5S4n四���%�bX?wMND�,K��{�O"X�%��gr�"X�%�����Ȗ%�b|g�˹�����f�n���K����?o߿gȖ%�b}�s�T�Kı;����yİ?�������Kı>�v����dۥ�f˻���%�bX���w*r%�bX��w�q=�bX����S�,K��{�s��Kı?&����rrn맏�.�d��ob-�e2��砯k��b0��n�ﻵ�}�&�.T0�ܩ�Kı?������Kİ}ϻu9ı,N�w8��ؙ�2J��p���L��]�ç���f�7,3.�q<�bX���n�!��	�2->T��"y���~�8�D�,K�~��ND�,K����'�?�ʙ���3�ݖn˸l���S�,K���w�q<�bX�'�}�ʜ�bX�'s߻�O"X�%��}۩Ȗ%�b}��%�iv��0�&���'�,K����S�,K��{�s��Kİ}ϻu9İ? �!un��/�&Bd&B�,s��[��-�B��ND�,K��{�O"X�%��}۩Ȗ%�bw�����Kı=���D�Kı?����?ofn�ۖ�n\��ڃղ�1��ڒL쌎K���^$��׳m���Kk���=�ܖ%�`�?]ND�,K�oݼO"X�%��gr��<��,K�}��q����oq�ߜ�~��`�`4bbND�,K�oݼO"X�%��wr'"X�%�����'�,K��>���Kı=�}~/K�fM�I�37oȖ%�b{��܉Ȗ%�bw=�s��K� �FA�Y�D#AxSbls��ND�,JB����_�L��L������
�t�2�3w"r%�bX��{��yı,~��ND�,K����'�,K�$����HVBd&Bd.�a��Ku3W72�w8�D�,K߷�S�,K��s���Kı=���D�Kı;����yı,N�4�gwI���Z�l��t�:�h�ݍ`3�=Ɛ3�r;����+�p��4��k^ﷸ��{�N��v�<�bX�'�}�Ȝ�bX�'s��8�D�,K߷�S�,K���ӗ�K&�3�nf��yı,Os��9ı,N��q<�bX��of�"X�%�����Ȗ%��Z���vG!S@ܴ:�D+!2 �/}�w��Kİ}�{59�� C"dO��gȖ%�b}���D�Kı=�g{'�m�7s6i�����%�bX>�����bX�'s߻�O"X�%�}�wr'"X�E�	�bg~���%�bX��r�ie���ٶ[�59ı,N�w8�D�,K�>��ND�,K�߻�O"X�%����Ȗ%�bw݅����w��-�x�m뜧Z]S�aq)pɲ��P�8.��=tG,ٱS������,K����9ı,K�~��<�bX��w��"X�%�����Ȗ%�b^���٥s2陗2f�D�Kı/}�����E#�2%��p��Kı?g���O"X�%�}�wr*�\�J\)!2m0�┺n��Ȧn�q<�bX����S�,K���oȖ?�!�2%�w��ND�,FB���_�L��LQ��:�M9���nfi�Ȗ%��@��?}�?N'�,K��;�p�Ȗ%�bw=����%�bX>����bX�'�Μ��]�0̙�n���yı,Os��9ı,?��gؖ%�`���59ı,N�w8�D�,K��{������κg�DY�k T���mb��Х:o/�Ϝ�;��1����ɻ9���ui�b�*vq�gk�x�lFC����A����,p;+�u!�q�d����v�zB�&�n^8'V��C�k�P�v;c��XtmR����sC�C.��Ԩ�:r��[O�k�M\L�k�.�n�eg=������q��\���x�ڎ�l�t�]ٸf\�LٷUP�����C��̩\��x��F�i�Q�]�훬��F:�汽�	�AR�ث�yı,O��߳��Kİ}��59ı,N�w8�D�,K��wH��bX�'~g{'�m�7s�n�nq<�bX��w��"X�%�����Ȗ%�b_~���,K��{��Ȗ%�b|g�˹��sm�,�4��Kı;�}��yı,K���"r%�bX��{��yı,~�ND�,K�>��ݦf�t����q<�bX�%���9ı,N��q<�bX��w��"X�%����{���oq�������n�EEkH��bX�'s��8�D�,K��xjyı,O����'�,K�^�&�O؏،���evL������-�SɎ�S���c���Ǐh��/T�#H�"��ڑ�{��Wuz����*��@��.�c�Ȥ��oNI;�}���D E��I'�w�X�l�͵`g�T��t���rC@>�Y�^��{��y�Zg�EqcM&≀䙠U�^����h�S@>�Y���CY9���q�{��y�Z����*��@�.%l�OG��`�r(F�9o;i�N6ݼ��uA�j��n9:�B^�\�\cb��Е�ob`͜�Se�;�w4\�r(��)�����̾M��zlf��w+K �xު����˗5T�{�6�fڲWDBj!%�	/+���,w����)��Lk"Ȣf7z�빠[Қ����*�^��<\7f)�8bm��$�A�w6r�M���lt�տ�~Ls��wk��tvK��ۮPv�d�OB�W��M=��y�$F�F�j�l͜�Se�;�02NA�ݢ�+�hn(�I�.��bG�̀{v����U�!6fA������S��[7�t��9���`j�-��憩���Ա��aГ�����������{��E�T�R��&~�Ӯ��h�2�Q6&`�Y�遫d�sc�I�0=U����~��l�-��bC�G\v�wg�Nzb�;�������#b������>�ݱP�e�9u�y{��`w/b`d���6]09p��&4E1���>��[)�|���˭{�����SnE19"�;����^h�נ}��h�r*�"BcnF�|�իń�Ӛ�:"������y�1cbxԃ#��Z������h/uy�v\9+�P�<��������1�ӮW�V��{	zwGom�ð��yݹ���l]��s��c�$�KZ1�66d�)cpɵ�d[������]�D�3���ض�^^y$��1fx�d�&��j˓��'��Wn���|l�q'�Z�9��.!��K1��5OB������^6��۔�sf�g��li31�������ܖ8��ګ������ܺK���nY�3kM���ԃ����]�1F�g������L]c4s]��g�y�ݭ,�ٲ���$��������_ʡ�URl�:�v�wS�6]05l���^��ՠ��\\s!J�4�4��ٲ�y�6}
!|�D)���O�; �xު�:��r��y�r�^���U�z�V���W�.s���HD�n8������B�!(��_|�=��V?ń�1^���D]�Y��3�����v8٣[\���V� m�v#�G=/T�]�!��_�2^����.��K`f\���J�l�ٙn����'���b�`�� bA�U<W1@44�D��@�?
~��~�9$��w���9��IBl�D�:i��ʗTHLԫ_oM��N볡DD7�;��ǝҬ�c�;�2j���S556�Т"'v��0=���01d�LY%�5��D��h���<�k���z��Zpc�C�#rAB2(�	Ʈ��'G��v��61D�b��}t�
�~������k7"���0R/�����4^���h�����H`�$"i7|�`j�-��r&Kؘ�K����6nJkz�"AR�$S556d�;��ݼ��Ă�H��R �c>C��Q�������V�,Ȅ&cp�#4*��2З�x)F(|x�j�O_����&s�c�'=��-	��4��e(R�"�y00`A@)$�1��N2�7�����.��@`!��ؔ"@�A��Q=AC��9�T�)�%��T@�> �GP���'�(Ģ%(_�:��`k�ٰ=��:�Ln8b�Šz��@���4W����y���Õ>t���i�T�It��6[2�L��0?}�}�ߟ�������]��,m ������n4��C;S[Ac������#f�F��2�EMJ��ޛޝ�`c���""?0����4ߪ�B�b�d�8�yؘ��`b�.���`j2	J��uN��,uT�{�6��eYС$޾ޛ2{����MT�E*D�n�l>Q	By9�*����`{Ӻ�	�/߳4�z� �T�H`�$#hMŚ=͛�Q���������u���J�J0I�(����x8���ǩ�n�o;��ۜA��m��]0�sY��u�ΚNq4�9}v����{2�T��6[6S�g])��)�C��vl���IG�BP�dݟ�j���}6�;���ٸr�@���7��;�������yڴW��=�;���m)D�����'���`fOs�1�l��}��[�C�BLx��@���@�-���fOsV=ݛ�l$�`�I#�w�����{�����rl�e�@��h"��yk>�Z��o�^q���<��K�Ru��Kn�;\S] >�l>z�,�-�#\o���FpޞیD��:�J�L�p��
����{�cD�d�y;uB�Ut�glr+�+[S�IN�6N�{=�:��0�;N���祫��c��1�7�I���t���q?sԄ�{5�*�96����]	�/F
�o{���>�w����y�w������vd��V���/E�\m[���6���o�ۋ�zU3b�u�9Ic���k�vlzwZ�1�l�(�Q�w;��Tg�E�L�9�H��r*`j�-��{T�lujS�@�J��X�i��́�Nk��(Q�N�=��Ձ��Y��SEQ"�\�3.D�ٱ�2�T��6[�)�3�TMMU:34�ܭ,��*�y�*�zz��"`w(���p�(^�rv7Wj�Q�sۋ�t�eq����Bi�=H�8,��#y#dn��Y�r�^��;V�ץ4v�,�ۗ4�nm9$����0�'� �U,���`ouq`{ӺՁ�Ǭv�d�5UI���ޝ�`g����M�Or����z#�%f�`�I����:��3'���sf���u���\$�d��H�yڳ@�z��v����Q����,y�v���໭؋l糸v}���.���O=�{*u��Q:e���u%U9��5�}�6�;��ǻ��J?0̞�z5�J�Ȱ�f6�z��Zs�yڳ@��vo�	Cfl���4�2��DL�>I;{���'��{NN�"V�'�9����}_-�X%\F�n&�8�9$�+��ϻ����u��6l�wq~�xۘ��Y�|��@�g�ٝ����w����u��Y�]H����qs�{/kڃնr�3�^��v13���w�Y'�1&�2r,�b�������˺��v��/��@�z�Y��$əM;^f���g�{��;'����V�\$�d���z޹0&\���r&[���5N�L��s29�j��BS���;v{��'o�w9 (0�
��W�1ϳ7�������d˴��#w�&e�L�}��O_@ͿySeȴ���vL�4�&�'	�|\��9'��!�e��cFwp�cv�k��+��z�,�8��
���@����\��.D�̾�@�,�#�7`�z�v��/;V��>�@����;���1�9�暰7gu���>���IL����3g<��X�*�U'$�&eȘM��̹0$����Ω��@�m�H$�@��z��߳�w5�y�6�;����p��Q�G��m�Ϸ�S�F�F���Q����ψ�U�m�Xv�Y�ϝl����ڰ�c]������M�Ӟ;6���Y2,�����}�Y��I`�R|eӹ;\:����Gk�nm�65��r�n ��J������A=B����r��jĵC��V�6+�:��n�Q��;�&��-!�j�%��dmY��\ݬ��/S�=[s6̎���������B��ܐ]����<Vqל�B��y�=���VWa;M�!�t��]v�=��0S����b�����"`b�-�n#T�XT˪��[���~ݛ�IBl̞�`r���@=�j�9xY�d��#_��[2�LRK`f\���K`f�.��!�#qhVנ{�՚<ݛ�I<��va�7�I�̺sM��=�v��9wW�{�ՠ|�׻m���^����U��s/9)�K��i��fv�;d.e��1Aͻf�����N]��*����d�e�L[%�������h3����`�@��U���y*J"�}ޛ6s��1�vlg�SS ���o��<��@>�i�����t�����䚊B�E!�uSa�J~���y�6�9���ޯ@;���a�I6�N-��ze�LSe��0
�9��m��3MD`��\��XP�^{67l{`M�%ySv��&�1����ٯE��&&��Q����&KؘqH�]A�E�3n��qR�Hd�Z�� 7�ܴ+k�=��w�Cfa���I�LԹ�*jl~�ߩ�'���9"�PW�r����uh+���wqdHK�j���ٰ=��v�s]��	B��Nm��V%��ЙUES�	���3/b`~�=���3o�T�՛-�JG��zz�ۂ��[K����vew�-�F��L5�.]���!/FhK�v����Ɂ�{�r*`j͖�̽���`%�p�Y&��yڳ��*�������}V�w#��țrD�һ���l�ؘ��0;�"��3iR%��]UM�%	�V�'����$�{��9'��@�#DB�ġ���z��͔���C��jB�L���rNSVl�e�L7��=�����8[���>4vK�]s���!��g+��+Ů;)��v�y�(��M��rGLY����~������&�O'�N)�2�A3T�~͛�ٯ@�[^�����=��P����j�lY���"g������0"��@;;���,$s�dN=�e4�n�˺�˺���K�� �L&
�@����9wW�ywW�}n�rI���&�B1.+$1~�� `�a�
�"A+�&)�y�Q�\c N+���w%�'���P��
 A*���T�*M8pdVmR@��Pؼ�F+�F)	ak	"FJ���1�*E��:t��曻&�l$�ݖ���uT���:MR*��	�k�K�� &FIسe؊!��m��MٳD]'U�J��r����n����c�5�i��-�c)�Y�Q�,�M���y֬��+`�m�S��`�5k2�8n@:6��K����q�}���2��H�56�i�h�}���'�kL�\d�3ú9���v����:-� ��!�u�;O]V���M\�Ӟ��S���ny��^�l�3�/.\H�[��u��=0�$�pu�Q�GbM���I�n�j�
۞�荣W3\D�ҷ�>�m�T�J�U���uŭ�;䂕k���}��5�J|��R��'����=]T���e�#c���q�u��S��p�=X�ӷe��z�9���.9��N���i�`+�"x�M�M��������Y�M�7PA�q�l�m�%�2�`�^.{Lp���p�h�!i��v����da�m�ˠD�U,Ơ�g��Fz��ۤ1V;n�ۇ�2m[*�5I��^���$�d�k��燀&���p7q=T��O���wQ�?��v�JUA�jx�e�v�]���X
q����Ҡn����Š�v����n�fL��������]BQN���m�M�ΐ��\�z�6� �)�kn�:A�� $-�$ mHv���ȹh� �*4Z6�S]�C��[n�(��n<�mmlh�gYu��nl9zG�6������#�H�\����J]����i)m��l�'L�e� f�e5n�m�i��Qm�*7m��\��4�4��s;��ۃb[e,��5Ҭ��UK�q7k���m��A�Ə-Ю7;�W��FW��J�e���^�vFh5�� ԡ�K�vT U!�C����%xLF8&Ө�S�R��-X�lT�d��VLa��8�D0���t�c/\�l��F틓�����j�Y�i0����b�/Jq�ͻm�rn��s-�A\D�G�ȁLp�qS�@�D
����!�/�x�_L�̓0ۛ4�������RC�MEhɬ�صZ2���Ϸd.R�x�7�^wmY��v���kv��]I��z�1�F@�n�*;l[��wkn�<4�C�6f�tc/n�v�i��ƭl���=��H�,Ef9��֐ݴfvS4q�.\�!��U��������6�]i$�N��w3���&Й�+wB�l�0�P�Om�C���ӝ����盤��ٷ	������C�3�f�<���-���Ϛ�֎���$G����w��6��Y17J4���?����]��u��>�w4sA�d��J?�I�癳ВP����`{{�X�6o�JI�6S�g�t�T�US`y�u�;�:g�����'���{����*��1H�h#�@�[��r�@��ٰ�%	'���=�<�M8���)�R�1�l�(�����>ޛٻ�}��?͎��ܭSd犡��=yn{v��d8೷9��벛�x���my��颙&4��<��@�^�@�s@��@;;���,$s�d�=��^����A=�0_�E 培��ÒN����@�^��`%�r(�I��D�z䎘[����`un�`��8KT��L�R۪V(_(IBP�+��"��������ܑ��h6r�V��G��#�<�W�}Ϫ�;��h.������`�L�F`A��ĲLrkk���ݸ��&v�/%���]�8	���>�X�5 ����s]��ݵ`~y�<�D(I~a�����M��r��jh%74��[����`wob�#`_�z�:SH&j����`y�l��Q	qz�@"8��,TJU
%G��G�v�g$�����'��6K�rIUJ��J�U6DDD(S��},��[rGL����JW�ਧT������<��6��;�/�y�s�<�W�wT�;!�l��8�F�"z�6��g@���N�03��t�]mӠG�������	L܊%"JbQI�^����>^���h^����Vd@�-%�S�$����7o�L[=l�h/$u�1��y棏@���@��l��BP�y�֬��v�S�Ή�eS��&f��С�s�l��V�9��@?�������{���$�i��K�C��U�f����mX(J+w�ˠn߼�Y%�7	J[�
��[u�I�������p�s3/�h;h���Q�&(���j`G&h��ˑ0:�K`fH�ܭ���\��$�Z��Z�v�޷s@��k��
㹓J��̕B*���s�2GL�ؘ��`L�ڙJD�Ĥ��n��>�@������M �#��Y'ƒ�4�����:��v���j��ȧ��~���2�l�m����͹.�fWm6"�>ݲrc�m�=����;�id��M�G��_�#�ػVqR(u�e�Z���.!��t�VKLm֛]��^p���=<���Ny�s�m�1&�}�����[R�/�a��s:Ya�PMݹ��£�DSv�#�w�d��,�+%�,��رu�I�^(Ы�n+jn[pҘv^ܴ����.����������������;f�-K�����ɯm���K�'��k��;�6z�v3�P[�s�쁦�'j�W�9w���9ၓyd���"`{%<�&*�n	sE����ICf��6���̜�0�D�˻E��hJ���:`n\���9Kڴ�wq~��`G&h�j�=�,l���3��=�G�\�md�$��h���<�W�{�S@�wW�{=��ŘdcdƠ!
9ۍt�/mJ��m��N��c��O4�H�e+s�7X,�����@������@�����9.M\��&%0qI��]��@� BE
���T�N�~�&���Ւ[ �4S�ˤ��˴��`b͖�̜�?U}Ib�z��\X���Ҕ��%Tĺ���P�|�05o�l��01d��ͺZ)Ϧ�6�	8h^�����<�k�=�j�>�.*�C��&!�!��\\S����5WR���.�\GeK��tV�ֹ����l�$��������z��_ߢ���wM�����@�˦�*j���$�eȘ�K`fH���k���47#�=�j�<�k�"��AHA�@���B�;��Z�9�l�x�ve��ԡ�T�>J""���3;�X~ݝ�v��\�w"i8%1Ƥzd���K`flt��6[ �����s�<l�b닗ػ��km�r�m�n�`�������p�z����������` +��s��"�z��01d���H遙h9�`�y棏@��S@���@���h^��s�³���I�RC@���v�nڳ�$�ǝ�`fmq`{��4��3-�4����!�;�+wM��ei`�%@�P�(B�H��
p�o��rI��gK��HK��i��)��$�f�Y%�;�:`r��N�[+�&�QI���T����Mz7fV�*.W�3��lG؍ă����l�>��#qH�������;V�����<�k�<�+��$xE$Q�'��[2rY%�1d���F��w �n4�8��@�����ֽ?��b\�l�,1�{T6�T����K`b�-���&d����&	��j8�/Z�u��=�,<ݛ�	E%�Qyf��UEfU��4p�T^�v0��W<r�[��0]�n�s���b"�y�R�.���_���.��vm��c��2q�6���t';]�݋��Cg���u\����2&)�c��y�t�Y̦i�`*n��	j��{eUm���l��i�����55�J��7&Y�������v����kvرL�p�p�Ron�kŧ�W�ϳ^$+q�p�S}����t�.[nnM�mEv�c�z[�d�{�p'�l`��\��^S�?F��?	������z�e4]k�<�k�=��QƛƣpG�{�Z_�Q	6k��1�t�~ݛ�7y>�h(�M�.f�wM���נyzנ{�S@�v�Oq$n)S.�l>J��NwM��7����������1���U5*��n�t���^���[�~:-����$�*g
S��{Y��;R���K��s��qٱ���;g˵r9��V�
+p�!sMvr�]ݶV���sF5h��e���f�6rI���� �B*� ��(	wg���9$�ﷳ�O{kK���<R%�U8�SS`c���3w�`fNA�ղ[%���.}�$��$z��4z�h.��^����(�k�Hp�=�)`r^���c��=�ZX~�d��\�Zh+'!v�oF���Z�v��|��b��oiblHĤ0J��p�>]k�<�k�=Ϫ�=�)�}�¬Oq�H&�z�����^���������B�ُ�uL��ST:��GN�l����'��{9>�{��L ���x�SH��c[Jc��[a@8'�8��*��E�t�R	 L"�(h@0)R)��HB!Z!c$�F#D @�bFb��@�����@���#�Uؑ� Fu��M�+�W~��!��^�'�8��1<		 6@�O!�¨H�w��2t�3�\I
V�ʰbL"I�fB i�Ca�Zx�{��tb�x@ /�`�Q@����u� O�
���S�O��>g�=;���'o��rI�'�&fv�C�RRuU4�>J���wN���@���@;˅dI���`b�-����������}�`w'!�r3�� mHDG�H�Q���r!�G8�m� 1��೧k�2���mvv�2/�G���@���@��S@���@�x�n���E�RG�{�ՠ{�ZX~ݛ�۳(��I)�t���4񦣐"�-�O�yzנyzנ{�)�w��J������������~ݛ������!&�D!���		j�s���`n���ͦM,��9�v��f��%��������=��h��]dě��X�X�v��'-�{m;�1�i�3!�s�;/o&kVK�sJڐ�I�q�z�h���=��h^��,<�m��%�E1�$4��?W�_$n��`j�z���0�²$��81'�}V���^������YM�h9�`��y���~͛����=�,>I(�B����)�3�SS50:������=�,zs]���ٰB�B$Gw���?{��n�5����m8���Y8�)��A�+=��b��u��hz�nw���)]��a5F`���%�+r�g9��p�]�K&����m�sl�n�:����)6��[�[�nѥw`�%tq:�;����Yy�샦#t��=h�IU��s��gP(F�+!u.%�/��h,0�v{�,���_i�q�Dk,�m����gj\���<���#������}�羘�q�p��}�F�ɺ���wF�;fj�w�Z���<��OM�.Fߛo������{Il���r��(�UUTə����5��(I�oM����>���>�`��4H�$qh�e�;�3�_%��x`d���ͲN6ڐ�QD8�z޲�޲��9���O'7���F>���N�T�қ\�rr�ؘ�e�;�"`?���~Wm�mkM��HA�}�;�58�-�T���݀�ۋ@N�]RX�<�洕�`f^��ś-��6[�9�h9�a&%�܋@��W�ffL'�$LE^����=������'{��h��h狆��ێ/Ē=�l�rr�ؘ�e�&\�R�hM� 6$��>���;Ϫ�<���+���w��bx��
8h��0=��{=}���ܜ�)��rU�\U΁��u�F�)��k����\v���l�c<V:z�,}��6[�l�rr�ؘ�I˶�$C�C�Ǡ|�W�}�)�w�k�<��7���}33�:��)����=�\X��v5�i(�����>W���°�'�$�v^��ś-��6[�9r�l�(UI���D�S�<��6G����ί�@�>�@���^l�<�#��E�`uhw*t��l���&q�mg��w�5ϱŖ,dm��$�@�^�@��S@�>�@��W�_;�*q�m���Ĝz޼�r�&,��Se�$H�K�0�ǒD�4��-��^��^������v��	��<����/ń�g5�ܭ,.������µ�1ߝՠZ�cnGH��!�#�;/b`~����S����=/ߓVIl������]\΋
�'�N3m�N��+��7���1��5j���@��{��[��I��Қy�Z/Z�����V�`�4��^���s]�����!��,7���D�n��q0"�z���02o �ܽ����p�Q��G�8��>���=zR��Nk��"���;'�\�e�53JdӰ=�ZXB��t�^wM��gݼ�q}AʥU�oN�͘k��zk	�VA�Ve3���cn�,͹�m�sN����g�d�nY�c��q3�蔪�\em�v=id��x��v� Y�˹����o��r26q=l.��9v8���Omdȝ���3��y&=;��  YM���Qq4Nt�6$�&qn�U�� ��d��s7���v@v�7;�.QU����sv������x��2�w �W��a�����&K�6ff]͹cg+�3��|��Ɍ���VI-]�v9��9-t$9)'��F��Ww��9zנ{�5�(Q�gmq`{u�sC�UR�e��-��$�e�L��0:�K���-g��m�#���qH����땥�B��$ߞwM��;���F<��������=zS@�zנr��@��S@;��`�@Nl����-������}v�&�	���π��a[K����1���`��ON�����u����1Sq:Md��9��ٛ�y�6��������$�~a��`Z�Q��A����=��M��~�3�*; @�OA� �<�{9$���z/uz��<+�5�Q�H#��ټ��$�>��J-�����]Ĭ2b�m��h/Z�^��{�4�Jhw`��bO	���-��6[2�&f�����P���vK�.�Pj̡'=���i;6l��6Awv���1ӻHw�w�����J�QN�|W���<���0:�K`j͖��×6۸��dS$�@�������@��@��W�س�" (��������6~Q���HQIE%(���}���WŁ���6�	�22%����ֽ��^��Қ(Oӝ�`n�zL�uB�uT��MM��6[&�����K`wh���v�n��i��LI8�\Y��^شnҹ۞vt�î7�������޾���	�&��O@�Nx`ud��Ւ[l��\/si5��s2nf�I<������u�t��zlnV���3U�QT誢�i���6繳g(J��������9vW[S$��F(�z߿f%�INW����������6�D$�%�P�BQ�ǫ�l��L���N�)��E�z���>^���k�=��h���L$7!��lS0g�w[������j����<q��p箻<Z�h�m��.r���05d���/��_Uuv���)��)*�t�&j���ٳ�|�W�}z�h��h����5�I#�>W��>�w4��^������cr4��z��~�̉ϻ�+�{�`c�l�|�C�����<�M5LsD�U5J��Nk�/�%����1�:��j��J��Q��BQ���E�Eh �+� ����"
���E�A?�DEb����ATW��ATW�Q_����E|AQ_�DEo��
���*��� �+�(����Ex*���b��L���V���G� � ���fO� ��@   �         �  �� x>�*P R�� P��RJBB�E "�T  (  
 PU
�R�(� @!�  `  E  3`Oy�>�>�뗌x�wۇ��h_p ݍ��M{y��k�*[��ax�p;���ێ�| w���0�A�Mާ�#}k�8�, pV/#�}��<A�wr��  �@ (� (d� ﯶ9o��m���8�t��+�� ��|g3�{{�g��  d( }D� �q�F�ū�O����a��| ������/|���������
9�����������;���Uo �
R��� P �����m�}z^1��^m���#/\} /r��]][�k�N{�{���U��p��L� &�|�}纹�� 橎�n,�eݶ�<�/n@����'מ�9��y�vޞ}����|� P
�
�� {���wz�=ǣ����n�W� ��4��  ��N�M��A�N���(  " �<�E���<M�"h w{��s t��� 1=4��i�JoX�)��   :P 
8����Ku�@R PN��  	��|����g�/{��fo ������9�n  ݼn�o�g�7��|*��1vn}���Ͻ� )�}n�9F}��V��q� 4�Om)T��  ES���M�R� ��S��T�U<�h  =��FҊPa2 OД�)J@  �h�IJ�`�
��?���Qt�������j/��$�(�P����*+�
�*���*+�����UAS��S��e��O��4si)�6�J.�6R�ԥu���P��;|�T�u���̜�!��P+���1aw��$�H��5������tl��(р@�C��״�$)�#]l�]s��>����|���Yn+���P�#P�q���6m��0��to��]`��/f_��>�N}�+��CF����6q!WJl��F)�T���ϰ�D�8�(D�ibWO�jF�J����B1,)�x�> XS�ta����B���Q4��O�!u��!�{�`aI*��F���M�vq��4� �0�B��9F�!�H!�$ր�Fo�%��7YR[��yoĺ{
i�8��B%J��F]m���,:7�v6�`%޹.�}���)���Β�jm"��I����$��_����"fM�_gdu���|h����vk6˜s| ����D���i�w�ư�
�]1� ��IMd���tB���5�Bj�3R��l�ϻ��3{�f�k{>�4J�&���]M�^B�H�ЄH�� �.�����-���`�p�_gn���e#JԹ+&��� ՊE�"���U�Id;4J[ӆ�n-4B���4�2g%�$�5&�YB�F�
,��,�P)�U��E����)��
h��c���%�|��>����
L�.��y K�Ԑ���(JJO�h�"[4|oP7������G�� 4����%�֊D�)�h�͇3��#]1j@��Iu�Z��5���}�7�o5VX̿�|0}�.2,��P�]J�35��.��r� ��b�R!P��A���4kg	Nf�B�g�|Jk7˭m�H4�:˷���d;>�3;�}��Xƚ�.�%0�i0w\y�6ӆ�;q�I�fi�|��b�cp�4��58B��u:SZ��d�g8|L�M��9NR�{i%�4 Z���
 R�ĉ2�wz;.�SgA�̺�,�,�>�Gc��4��� A؇�ư�w�������,�`E*�#�bH�A�`44Mq���DJic@��4a��!B��A`A9 ���D�É#�BJ ��˭|b!�D�� ��MJ�+tj��A�$0c!V0L`hD(�"!d��3����]�6Mh%$R(|*q~H]d	.�%>�h�O�!$x$�	CSR�j�o|8+�S\H!R$M0+ ���\��ьHP���T����30Bl��5�O��C�J�`��Ņ�@�B�Y5���z@��W�b�nOI+�_h�.�D@�,BH0bX�H��A�D��)@�.�]��$.�\����n$�"�!�H�H�J�͈gIBNq�
ٝ��P��Sl9.��L`P~X���B�kB����1"�$!M"q"
d�(D�4c�k
:W��CX����XTѐ����H�H@u���A���#MXX@� F�l$�R�X�B��LSd)��ԁ蓬�#M$$0bń���� r��a�/�.MMu�țK��V�0 P�J�#]A�!
��J],����n�w�x�6s56l�N	$�x<�H�*!W@F�M8@�XkY��ɨo,�!]�
hb�S0�`F$ ��^$ XKi��X����r5�!!�ԗ��5��A�IP5P� E �$I��AZ�B��!`AB+"�P) �@B �`�X� `A"�E��"�` Ā�$X� $*��� c,@H������H� �D���RAVX�! b�@��B�"�4t�i�D.�$T�$H�k��$�X�)��K!�FB(@�F&�jŤBD�bDb$BI��0��D��
��"�+P 0"0"B%T�`ֵ�l��CYM`Bt���R��*���͚7�����MB�VȒ��c�T�!R���"$U4� @����#�Ӂ����Ra�SX� ����p�¤k)���.�����Xk
�$%�F;`�HIV44��k �qat�]� ���ÓDY�7C�8��h��tolB�A�A�a/�cM-$�M�M�0
顷|#WF(�
0�JQ#i�ke\tm�<8�0�ԁ
h6��
f�SN�rF4�Ue�Y�� ŉ
��b�!]%�ƴ�I���F�Ɛ�54�A��J�!�H���i"kD����zC�/چ��|Q��P>X	 ���FH�&�d�J�h@����.fA�ڭg�t��1?��Qe��'{�`�5��!�1a9o��{�pd�hJ� �a�V E"Ձ@�V2k�nԁ��E���H$BWC�"�
FB$$#
j��Yl�N\��y#�%4�0�.�HHr�ɭ[����B�%.Q��B�&�g#u�
�p�!M\�y$*Jhaf������ GZ���D�#$Jh�H���͙c�����&�BUb��Tk��]�$JL05@�R������	�6"aP���pbC|#\f���(¤(�(<�Y8�3Q$�0�k ��$�ZL�J6B����A��w�5��@ނ���2&�1ӽ��p���ѶC)�˄4��%�l�ѩ�p��h#t®�j��I8��	�E٣PӁ�d���a�L��"jp)u"ћa$HS�,����"D�V��H@&��
kO�,@���*:1�`S'SF4w��Rl(d�Dј�#�Q�`�F	�RF��%eR*��h�&�|a�{B�1��0�J�),�%Ve��*�DR��@�t�Z�X#
6^fwe�����k���80*An�wP��'�|&�,�$i�R,)��4�}���K�Ku���7���BT�*t���ᕑ�Q�y;�$�j&o�l%4I�}�٠40�O(�P�jSF��jic�E�Hh�Fl�fJk�ߙ�؛/0n�fs���_��}�o�	yϻ/s�4�
�`�_%��f�a8i�F�6��j;)N���fs��7���r:|�|�����n2���$!��ѐ�ɇ�>��.���zD��jFO�:�S\��I�|h!M,0 A�a�d#��1f��"�4ơ�>8F��#�*A���!XR%4�
�5�`a���`х�l��bC�$ i"T� 0�SP(�`� j,
E�D
@�R$J��wO����� h �� 6�   @h[x� ��[Ie8 ���ٶ�f��`:3K�It������l�ck�$�ت���$��0����p�v�%��r:t�m�I��C�U�t��b뒲�UP �p  3��UP<l�+0mPU �p�P�(������( 6ѭ�%�$��p-�(�s��[\��J$�I9��'Om��k^���[Kh&t8H���	&ð�^���B��y�U2�JCpu�Zۧ@��|�&�9 �m۶�����M� $H��`6�m8I �m[p6�-� m��V�K�Y�ۀ�`�a����  6�հm&���0۶ $ �  ( �bCm��� ������$m�6ɵ� M�8 m&�kn8���Kh$�V�q[*�q<(�ŵmUҭU��M��-�@��I��[y�m����������
�!�\peyY`X�$ݙ��;o�k�    Hpp
�n�.�����/i�u�L�m�K��AU��v�}����V�� iS���x�Wj�R��yV��������q���.�6x�5ur�J���-'竐ēK(����$�I8��k�yi����v��[Ge|����*�*�Օ��\8�1hz7+��=���	@Q�+W����@m���t�ր�NV��P��S�P��o%�� Ia��l6���I��' ��[d�:�V� �l �#gW6[�( m�!��S^�   6�6ۭ�޴;[��$H`h  $I#^צӀ�`iÙ8��(䂷5[V���i��� ]�c��	�����t���$���rA�mp� �A 6���`t�� ����A�U��V8*��8iV���Wd&��c�n�&�A�Z5�H��[p��u�mu����U��d9l &�rY;�3Ze��hHI��6NKx [G/Ie�` ���hsM� 
��`2].&�����;�*�:)zڭ�j��y%�RX
���Ғ�6�͖�f�6 ��oxq m��l;Tےt�Ce����[,�F����6��;�l㌀�$$��Lm��)������%�Iu��Ix[�#v)@��Wna��'k��A�v@�`��;�ʕ r��Mr�\�֦�(��`����ۗyy��Iͯi! ���k��*�5T�q�"`�1ۥ��һ+�wW!%�c X -���A�,��hÖ�	�J%\k�������ٺق9���lIնݵvʵ@C�&ق�Wi�!LC�
��Wf��O3Z4u���-�ۤ���5��N��N�B� [u&疪�C��.0�pU��`
(5�m�>F���&װ[@ 'N���cF�r�K�mv�mT ]��X�§,b]-��m��� $��o6�� m��-���� 	�>p��H�7�>�=m` n��ɲ�q���`���d�յVuђ�q�e�VϧNeE��î��dp� N.ٮ�BI -�m�� [@,�o [@ Ft�@ ��WM��T�˴ ԪZ $[KjĆۀZ ��+UAīWUJ�T a6Z�ꪭ�yr�5�E�� ��N>�@Imְ	4r�Ͷ   �	-��m�6���:�kj�e�� ��A��   �`� � m5�&���l6�H�J ��Ij,P5U� ͗��0����үPl++UJ�IE�  H	-9oV۷  �p�f� m�M� ԛulT���@@*ƦH� �`�p�wV �� m���ll  m�m&�h��6 �} iכ[@K��D. .�F���     � �BM����7�/^����kn�l�@��n�[d �����b�m�v�i���M� �8^m�� �T���&�M]���T��K�'���YD�KeN��̰qp�V��@�܆
{;-@@r��jU� �`�pҸ0[����H�K�Ʀ$<��*��N�5:ڝ�m� m�� �hIn��  m��*��U�Wi<J�\Jqv 6�Z�U�l$�z��@8�iM6�����U�Ij۠ؠ$�Y-��n$-����$p ��z�ZF̴  -�   [@��  H  -���      8  m���� [[l-�$�5�5�6��ޮ�Z�n���T��gi���F�z궔���e��������8�Z���A�l��V��q�2�P8 Z-� l[C��mm�   $�H	   �kh  m�  ���      p h      @    -��` [@8�`� @�A"@ h  �m �   �  �  m�  [@-���������aJ���r�l��A�H$ l�C4�6��Y�8�5\h��q Kҁ��  
^ ��m���   U�Q��۞@��ޠ���6�$lm���@   z�@l�Ĳ��6��� �      m�  $  h� � �x    �  $   ��   �   H    	 m�-� �x�  m�	0	     �m� ����8 �   ��k�x ��`�vͳIٶHjس�H  ۭ`m�mHu�   x< �[V��'^��H��N��T-�%�^��[f7 �X� H8�o��O<�i���Rӊ.̪�lʵT�o�ʪ�  �    �     -��   l�   6ض��  ��/�  �   �H8mp6ۀ��v�� [d  H �a�f��mn�`k�l�LN��V������Ur��-� �g  �I H�m�8�l��5ו��n�6��iq�lͮ[h �IGm��d��I/JC3�TF��������n���Ҳ@[@ �V�pTm*�t`�/J��j� m9��ݻl �H:@A&��鋆�O{�x�k$�c�����M��^��gdyt��Y��J�A  �m�@�� ,6����6j�nٶ	�kz� ����E�5�[p � �it��m�6�k[pv�ۭ�[@   X��H 5��V���������)� �k��ͦ���l��m�m    �-�Uu�U�v�삵)-*� -� ���֖�.˅���h $Hp��MkK&�]�pC�pZ�W��5� H��ٶ H��˶�ޠ8U<�u*��ض�Ė�    �[(ĥ@l��UH9v��@�m�p ��۵�]%���x�	  m����    8 	h ݰ ,H�m�pӢ��@�tr [=R��u� m#�l�! H$mٷإ8�H� �mm�@8H��-��`-�H�m&ͤۂ��ж��� ���p$[v��)ajZ���V��l�^Ϥ�Hmt��-��Ŵ ^�kh0� *UUWUp]6�6� ��Xl����̲���,�7m������)Z��܇  �\��m�v�`��$��'���ì��FM�Li-� �NSd 3��UU.�[T���[p�i���M� Kj@[�۶� oM���
P'�u���ki �˪� �c�m@��l�m$��5l@9  6����p��m� pu�8Cu�Àn�u׮�d��I��   ����M�m�m  r�,0 �]��l�2�o�6� $ 	-�� ۲B������$9�I�.m]c�-�R�V�A�Ʒ�m�kuT���m   M��e�	8���pe��А �"��dH�t]�u,��Pꪨ,론�*�I���8 �v���m�����6Ź-��l�	8|6�s�$i6��7$�5T���)RmqWR�i5� r�n�#K�*[���A� �8b۶��6�:���dB�3�"|�3�j��l�UJ��De�KkH��2r�R�eguG4��U���@�Sj(���^�e��f��U��5�a��krD�V=�7V���;nƺP��V�g�2�9z�g&�������n�8.��γ�]��� �{�����[F� %X�c��� 6�6�y}}��$� ���>���������w��*E !"X�~3H�(�!�������ڃt��p8"|���M���v� Ch���;Z��J��DT���4�� �v��|S��D�^��D�
_����pG�[A<g����C{��H�D 	�A"�#�BD`��E袇��>QGx��Q�����TN���)"@!P �D � ���EJ�P�lJ��E0>Ux�"�8��AڞҦ�"EQ|@8�.��"�G@/� �!��i@�#���� :/S����ʇ�NC� ��FO��xUN/���ŀ"�x�xS�Dc��@�D�b���!��ͪ��z�
*T�Q~E��>:�+��)�0TW���P� ��W�ߕR�GlpQ��h=ɷk�î+�E��9�g�gc�\��jyU=tj��Ӝ�Fw'-Nշq���r� �Q�kH�����tc-�PΞ̍cK�r�Ю�.m(��Qyv���*u˂�b�-&�ҳvt��i��n��f�rnb���r�3�;:QD�Ya6�	�G�la��0��|+�Ѱ��8mƸ�㔗�8�α��6Ƚuj�tcul<��jskh��Q=�n3"�.�-�v�<m-Z6t��<�>&�3I�	�v9q�������C�{�5�|��N��2���v��\��Si(^�t:�f��`�Ȯ6N�Ŵ�X��v��H��f4��lF㶌�s؍WN�tUeCm��FO<�2ZW��*��G��k�aX���,��M�(��	%ˤ�FvѸh;j����sD�L���!6G$�gny*.:P&vѸ��r�t�"6�,�T;mHi�����V��Ԇ)��8vvH�[���<
�@�Ut�9�VV�ڨ6�� 6��8m[���r���P��	n�1���YypUu]�Y�p]��� ��!m$-�W6 H$I%*�R��)r�R��Z�48�n��Bz�Bn���E�ḟ*����k�/G;i6�lHL��PlO�v��>�.�MU�F� T����xL�;n".&�dh{!��sɍ�:��]p൭n]�(�t�.(��ؚ�t�0.d��)2J�.��4BZ2Dd݇7P�c;.��8Z���R�K�*���������&$&S�6^�ӫ�Ʃk���8)tg�����	�f��[b���J�Ҩ�nȩuUӔ��s��T���V��9=�8����*S�nw9n�qy:S���м�l�Q<g�V�@,��v��� q�G�vѳ�v�+[���k6ù3�V8N�·sq)<a��������Nc��Z�Ѐ� z��F" ���ҜD�W��������~q/M�I:�9�x�Γ 4e1���/PCy*"����(l�bp��+�xz֒w]5���j%sv���k�b�Q�;Ta�.ݧN�ݹ��jۜ�� 6�[��W`�5���ٱ�id�-�	-���c)�/��(hڴ�M����׵����YѶ�<T�烶q�1�=��Y��-rs)A��L`�[U�:��.�@��QӽɽJHkR�Y�6�����x�y�d��L�+�Ϟ80�_�S���~��V���z�P�� {_^�@�GQ��7B�nI`w2i~�W9��$z��ŀw}�`����-�mA��@f'�&p=]8�k�%|�,���ԔĤ�*s��X�ݖd�����s�Ӏ��k���5�bI��|e�����rWN �ֽ$����?|���,��İ�V�v3���ٶ�Z�Y��Qm]�]�*q�m-&��M��t�.J��z��Z�	�샸f��_����grWN�S̐����$���CCJ$�BZ����?޼ ����m� ��-��)"���c��,��� z���gu�,��� ݩ5�d�O���&��_=/grWN ����	q�i���n�jM�����l��]��w�wS�l"�����u����a-���t�2p��Q�c�Z6��q�e,������m����������������\Z��n���O�$� ����W�OK��L�t�=��-{�ŃCi���wٹ'�w�71@��"	  H0�B0H�`1��� �f�]>�znI;�{6��Tn6�z��7��z^�g�� }�_ Y+�'��]�3[i��i�m<�.z�p޵���ޗ���*���E�� l�\�LJH�L]pu:�.��N\�x�M���~����殮_���u�T�%!��ߥ�nf��ͺ�.z�p-%њѩ�1���o�,������WN �־�\km%�7[m�����WN �־ �W�{6ڒbԛY���Sy�S�g�䓟{ٹ$�{�܊�(�Q*��bht"��O(���ٹ'��5[Ż��7�I3�>���,����V�vi`b�ԅ�ȁ�"��B�R#��r�]�Ip�U	ŉ����eZ�m�FνՉ��i4� Y+�=�{8��OUr��sޖV=^�RN��J���=�{8����Z��W�O�du��Z�֞7��3�Ӏ=�_ z��z��޻��Y�����سu��=�_ z��z��g���h�D�8�$�D��l�=Y�ߗ�޾0�n�P�J��%�B���G���ִ���bljݞ�)Cs�vm�8èm���c�7Z:8ȣ焞��N�˺�m��hŵ��4p���V�v�2uc;����2�8�kv�Ɍv������9�v����qV�p�2�Q>��W���󗕡�b|nW��%Ӏ� �GM���Ȟ,��}'=ku�U�d#wLӳSk5�-U��+3ۑ9g=�/&jp�ۉ1��+�SӞ�$gv��d�:0%�wu�"���dںa6��[56���vp=]8޵�����m�$ĵ��c�m���ٟD�n�^ ow^�7� �>֚��)!J��n��� ��������+���k�&j��V��o�=m|�og%t�z��{<���i��L�y��7�{��pWN ��� �n���K�]�T��L�� ��1F��s�q�Pw�3	r�c�N;\�	���6�)8��8�H������`�=m|�og}V5��֞�,ɫs&����q[�U<����|����Ӏ�ZK�5���cm��� z��z��J����`}�3j89"��H&��,���`[��8�Z����{6ڒb�v�����%>�����x��u`fMRF
*��&H�I(���1۶���)j�����5���k]��v�٠�$��z����ޗ����p�Mw�Hx��ZM7���tBJ&M�ذ����n�/V�J��pJR���{�u`w6if�9I)���"��w��� �������M���p�Ӏ�}j�K_���X�&����G� 5!`|�j�I_�K��}+�<�	b��8fk���<�<�Y9�\���s��1��]n.f�k����*)�5#?6���+�=�{8�t�>�Z��	q�$�
A9%����_�ʮ$w}<Xsޖ�͗�U$b����dS��GM�\���>���=e|�/g3d�Ԕ�G�ۅ��ʤ������p���fff\U'N�ɮ�����I���W�{��p�Ӏ>��7^����U��d��Hģ�R�[Y�.��Z��Vy�4�[�Ь��n��܊���qko�����'�� }�_ {se���a6�P�.9!$r���/�2����׀{��`t�J�M��ޘ��g }�_ z��z^�z�p-%њ�i���z�7���ޗ�������|��\i�S�1f�jm�����t��k�=w�d%�D6�W�WsU`M
��$�ٜ�-��� �d�6��v��`�i�=�5v��U�MbsayxN��]���7h܉�Ӄ�3�In�K��{F�/F����;t䞩��q�m��*늼w/"��`K5*��t6��"7gDRo�o�=����#��h�/G3*��L��Ƃ��(\�8z�s�iۓ6v2ɘ�Vd3��u]��^�/5�����{��������q��8�&��+��Fg��.<q9��U(FtFM4͒���9�M6�6�p�� �־ ������͒���kI�<I3�>���=e|����t�'�m�Lԇ��6����W�z[��OWN ����)�7cԞ�z[|����t�	-|�+�'��᚞��UՖU��7�ـ}�[��Ϯ����Xͭc��
Np�"P-�dI�� !�i�]��c@v�K�O8m�����ޘ��g Ik�Y_�og��A�����4o�$�9��Q9,�]�
=E6�`������Iq��O ���M����z�p�� ���mU��7�����M�=]8[_ z��	m��2�f�RSQ��1�Xn�=\�S�����X�v��Dm=�sS,A>u�qΡ���[Y�јi�솊��,ok�9�M,���l.���B���~}��,��Һp����v��n�n&���nm���ʤ��O��K �����a���B82IV��0^���Ԓ^V	
%BI"T�6D0��� ��X���4��kh!B4M���P�\�t�)-)*�H%��F$� v�8������"�,IZҐ��)�$�R*F�AHBK(A��d$�a��*A"���Ba$ �H�XDz���F"1���]��YY�Q8��h��T:�"�B�'|�qTX ���*�����H�)���L�G��'���=f���ך��cl[��,��=e|��p���>��]���f$޴��Y_,�Vu� �͖���zӦ�#m��n}u˜U��2X���j��q��˵�P-Yt\���*9C�RpNI��z��ιw�%���W�M�V�5��k��m�<�� ���Y_,��͒���k��@�-oxY_ }e|��p�Ӏ�e�����P<�����=w�k׋ �;f��	r���<EP9�[���x���f4�����	e��=�^� ���َ��,e�:��dP�F��M����prli�7L�ӝ�闄(n���qٞ�by�W��	�_ z��Y{8x��K5����g OZ����z���I]8yi.�ԓ�ى7�S|�k�=e��$��=k�'�͸��[0Y���|����Ӏ'�|�k�=���b���m�󀒺p���=m|��Xj��D�&$��)����W6b��4�D�#����¶M�f��ݻv���ϑ��u���npunG;Pi���gf�j4o����n�z0���c�N�J�k��=<����s��k��m�!�6rRg�,.��P*:��b�b��YvW������pۖy�Y:֚�̎$ۉ���K��q�ju<���Ɨ��A�1	\h�u�Vu�O���w��z[�̼�׫iD��*�n��p�`�I��@�K��^���ܕ��ٹ$���������������閮Bfkl�����Y_,�����,���yM���bZ�k�ŭ�Y{8	�{8Y_ z��g��7��by�Iog K+�[_,���.��f��ޣb�l�	e|�k�%�����po�����b��զZ���aӰs']�ݬ�����u�f�r��V�q��Y�z�N�suWx������7]�舏���`n5���j�)ܖnm՜���7]� 5� �n��t��j'$����͚Xnl���UW3���7��)fm7%:Q�A%6�������K/g%t�>�v�5���Տ[{�� ������I]8Y_6��Hz�z�^kLl�U��F��)���m�\�v]]p^�lt�i�k�,�M�-z��-M����I]8Y_ z��g��7�cby�I]8Y_ z��	e��>�u�n���j� �����`��gyD*5�@  DT�t
 Us�jn����vi`w��*I9
�޴��[_,���Ӏ%��ֱmE��JA�%���u`zB��8� ����w�tN��2~��[C�J�Xn�ѝ��/R��fK6�!5��CU�,\sU3��}U�]��}���-��=m|��p6K�7�5���$�������Kog%t�=2��k�ǭ��� z��	m��$��-���z:����ǫ^���,���Ӏ%��vﭯ��@�{L�m�c4m�%t�	m|�k�%����-M-N= �4��1%՗�-����A'�Ŵ������$^�k��5�SW:��o��}���6� ��,u�0z��7*wSf�57�6����Kog%t�	e|�ٷ�m��nkbI�[{8	+� Kk�[_6J޴jh��4�jo8	+� Kk�[_-��͒�M�Ѧ��$��Im� y�x��`�ـ$�4�D{o��*Ӓ�X��[Gf�����v�n��,@�7i���)	����8�ˌ���mc�蛛�TdK�8w[5خK0���F�����چ�ό��m�v@�mڳ�Wt�嶕�^z5��E�g`����u����F�,�+���6��5bặ ���X瞎!ݞu�p�)8��v���&� �F�s8�q���<���]�/�{�_���a��:�)^�
�שS�:b�@�.8������3	8����#��)�@7���%�����pl���z:����cK^���,���Ӏ�e\�k�>���f�li�lѷ��Ӏ�e\�k�%����=Gu,׭��!��[8Y_ z��	e��${�����*I9
NE��;����^�En��j�$�Z*�5p�sv�
��磉��ˡJ4N�n^��[mu�W�]�S�++_6���Ͽ;��[��-\�k�=�V����Y�e�.f�w���� �1*n	�	�)�E��{�ܒ}����}-��&l�o�m�x�=�=��������En��v�5��c�O^�����z[��I]8?�r�=�����<�N22�j i�`w-��$���Z����M�EǋjP���0U�fS]Q���tT%����3q�5h��M�μ#7�ޒ~J��{e��=m|�������b�G$�J�������~�W�zX��Ձ�{�����*I9
NJQ�`���=���vET�78�[��lۏX����kbI����Һp�j�K_��=m$�ǭ���V�햮 �����q���~�k+�j�ed�i��L��� {@�A�Z�6�1A�Q������Z5=�=���������[��]��fjCL�OV�����z[��z+w���W��uCF4��-M���p���=������]�3P�i�lѷ���xln����b��_�$B�""&u���&Z�ĳ^��f�n�p�j�K_�og�]8��%�kŹ�i�i.�p0<�nT�:�����Bb5��\MD�	t���ܔ���;��� ��g%	G���XmK�W6T��p�lI7�z[��zWN�-\�k�=�V�����ŭ������[�9%&���5�b�5N�UM��I�7BL�=��������Һp�v�5��c�O^�����z[��zWN�-\f�g��!�	����l��ɥCQ"�LML�8�� �FD�@�`c#���RΤ4�A��#	�#�"�0,�!� ]]����������U/HX#ke�GA,����$HB���hM2�!��]K�0%�e�Ji# E��kMZ�0Hŋ�"��b2XA����L�K�pŀA�p�_��1 ��.�E��}!�d�$H��b-1E�T�����GH0H���E����H�CH@��0�"�*1��R�+�F���� �(0E�Z�A`���(`���"M,F���CB� B�J�����C
�d5M0i�#P5	�X�+�M,1+�#SC Ħ�	MkL	"h#5("i�) T�	
��V�P�Fj)�QA�@ h#��`CK5��i��Z�(�U%V4"`E�K� �,$�i�R�"�*���&�M�h�D�7jm�ȴ#��uYߤ�33-����`[�֋\��ywcb���m��$�a����^tkx�qYd9wp=���Y�a��ތs� ��]�2�����3A ��m4U5�6'oK"�e�nin^�UF����� ��Z��1hH^͋�Ji�ϠκU�9��_�o���� �m�a�um9�˝�l8V�y�m�ոS���G]]*������SF��W�\�'8ocOmc��&oc5b��z�c`q�d�2�_<��C�+��g��H�wm�[�z��[�v�śh+n��gtbz�t�9����=��q�;m(�r�5۰�k��n�)�%�IZy)��������νp�N�J���I6�.���s��n�`馡5t�J$�v�K���<:�m�vVUV�v��ÖV��d#�K]��Bɽ�r�ַe�F5c	�<��V1vͧ�ا���tm�xUڞ��l��1;A1�U��Y�C����,�v2�`���U�Z��!�o(l�{-�����	�dL9��ۭa� -���	�T�Y]rU��n���h�L8�;��ӡ�Ζ귰Y]��mӉK�g��+j%j�U�-�^A�V�[m\���Ֆ=o�㜡�F�y%,��SWf�d�V�;��t�j�Rʡ����oR�N;m���'kj�;!J>��@uC� ���g����B�h�Ԅ�ݍ�,���(�z���؆ػ.�˔卲[WC�b�`:-���)��6�j��QҮaUq��[
��x*�a� �6۰gN�fj��Ux�\+QۍP����=B���̳Fխ��Z,R�=/���d�ݹ���@k9�<q�uTn6�nc�8-�ڪ�6.�aBk� d�lD �ǈ)݀j��2ͳ�]�6�(����cvt�l�/��&�P�lR��4��g�ۏ����Ţ{]�;�IF��V ��r�W�@�..T�񓞻 �Bl;Lֳ34qA�n�8�Wh�D� q_�T����MfM]f��Z̶�Tm��F�ْ^��݋3��R��^d7�u��{�vc~�,���wE�:SsS�ĕ�N.�S�����1�Ghݵ��iEKu�x�죭C�0�8	]m�jʻ@�,�vɻZ3^��Ѧ�6�v�F\�Hm�Y��p�];Z��GX���%�w&0��]�8woWY�sǁ
�t�c�K���둝;9�۝6*�k-�X8:�rsN	�x�mj\f&���i�����
uc�Y�6K��5�����g�]8l�p������{JT�Q�R�U��٥��W9�q#�π%�����pg���M6�4x��ـzu��kw�(P�u�b�5���;��:Q��7%(���=-��=+�햮�lۏX6��3[M���p�Ӏ��W zZ�L��Q�������1�Oc	+�:kL����Y�����]gMD�S-�����Һp�j�K_�oU���6���n&*q������w�k��T�`A#1`�F�D%$�������=�ٝ	)�6��lPM5%EN(�v��K����zWN�-\���,LZ���z5w�{[ŀ{]� ��u��
L�������+E*r$㨄I*��l����W zZ�K{8�ˉ	q�f�v�蝌�m�&#��a��֘��4��;"�77I��	R��XY����x��\�B�!��N�A�7Y�&��o5���k�=-��=�`uf�W)#����@N�*)H6��%��8E.��}��-�� ���[�"��jBTRR�U��\Y�|����������{6K�7�u'��M���L�#�=%��=��o�w߻BK�G��Wn5�p���́�����r��̗��*�rS�9Y�q=z����������K�=k�>��[N���(��%��ͺ�3��־ ���	��{L�6�k4M�"�xz��[_�og�z��,Ե1����	-|��x�x�]��Ӏn�wM�֓Oq�7�S|�����p)w�$��Ѭ[[I-Ǹ�u��H�@�M*���	�k5*��[��<��#9�X�p�lI7�z���H�� ���[_풷�&	�Pky���7k\�BQ2�^ {�� �o2w��ѹ)��LT�5"��zXۻ0�	L�wb��Ӏ{S��M�U5v�U]�Wx���w^�݋ ݭs�В�����͞c�"��QD9,��,菻��� w}������$�A�E �����ֵ�e-�\��M����˭H��L����m,K�l�F;X�������W����z��͋�ո֨�rMA�猩/�Y�z�Z�Eհ� 4�1X�5Dc������3Om$�\.�:ށ��U�ι��(ۍ�1���]\�cv�C.՝�=�Ŝn���и��p�bv�D��n���h66��A�n�&���>	$�JƖ�K�2�w�ﻻ�{���y������벋��'��ώWV٦{l��i<������ͭ��:�P�D���?��`���>���9��{޺�;����*lp:��+ ��y�&C��x��X�k�}@��-i4��z�7�[_�og"�x���H�T=`�7ssSē|����]�K_ }m|�J޴�8Dؤ��1���,�z|�{���n�X�em�rR���F�V�˭�d_-�94�#`�=4um��K��v�-)�[�4�ŭ� zZ��k�=m��$R�2�ڵ1$�x,M�7��w�Mm7� ݭs���r�I#��<�NE���rX�Ob�xK_ }m|�d��cLֵk�4�E.��� ���Z��}��,�Y�h�cѷ�%��>��ֺp)w������A�;L�9��ˮx9�ݳ�s+���u��ܺE�R�V���"B�V̼�q�$�?����Ӏ�K�%���l�{�{��5j���7lϢ��>� o���ݗ�s��}"Q�'Q�))G]>� �n�PG��rK,��w��v��nJi�Hr��X{�ķ}�`���<ݳ��"������}�Ud����hI� ���Z��H�� ���M���c�oX6���ckE�����Ƿ�{�b�v���vC��y2Q�놜�AGTӒ��l���y��s��+�\PA���ٱ�A�A�A�A�~��6 �666>:{�5i��sZ�ɖ]]d؃� � � � ����b �`�`�`�{�߳b �`�`�`�~���lA�lll{���M�<����ݟ���Z)��.�4e��v �6667���6 �6667�߿f�A��������A�A�A�A��߮�A�����~�k.�YMj�2��3b �`�b�	MA]���͈<���������A�lll}����A�A�P��@� �{��؃� � � � ��}�S)��-�.�ֵ���A�A�A�A�����A�lll}����A�A�A�A���ٱ�A�A�A�A�~��6 �666?������u��k2f��kZʝk҃�k��Kԥ�9�a��dݸm���c�.y���Y&��j\����� � � � ������A����߿f�A�������؃� � � � ��~�v �6w�����������Z2�aK����� � � � �{��؃� � � � ߿~��y��߮�A�����~�y�~�ֲ\���Jk55�͈<�������ٱ�A�A�A�A�����A�lA�QH�� �?�g���A�A�A�A��f�A����O~�jh�e��5�)��͈<����g��b �`�`�`��g�]�<������~͈<�������ٱ�A�A�A�A��߹�L�[���2�.��A�lll}����A�A�A�A���ٱ�A�A�A�A�~��6 �666=���]�<���� 8"	 ;����ړ,t���untHF&��I3��݉��{�7˴����k�kT75��cyz�N�S���s���V#�VWK��;_��ʅ��W,9x��-��X�`ݧWWR��l�E�EdeL�QԫUsm��L��r���ۃ!�Sc�=��p�6R�]��J�F;fx�4��˶�GDl�u<�2N�8:16��X�����{�=�+�?�zq�T�,�a��V^��Hsٻ11/,.����:���z��\����Z)�ZɪMff_=��������؃� � � � ߿~��y��߮�A�����~�y�=�!������e��f�A�������؃� � � � ��~�v �666>�{�؃� � � � �{��؃� � � � ��}�S)��-�.�ֵ���A�A�A�A�����A�lll}����A�A�A�A���ٱ�A�A�A�A�~��6 �666=׽�2ܺ�4fkR��]�<���%��߮����`n��,�����S��r!�$I��&��$�����z�w��K�m���ww����,:V�r�v��E�S��t؇�8�`��e�X�kp�WFmv[�(hq���}�K��U���U�Ik�/�U�V&�ZkZ{�S|������R��D����rI��� ���	����4��6��MOx	��Z��k�=U��}��,�X�n,hm� Ik�����{���Rݛ�`b�+}
qH�ӑ5Wx��xo_t��}8�����"}��6�7Q��8������ӡx�S�t�\��j���T�::���Uw���v�� n�DB�����~��{�E :�SRRN+1� �n��n�:ns�d�U�uWrSrD�r��X�,�ݖ]mr����H��|�4�!RF�J2@�,��v��f�.�6�ɉ"F2(SJ�7��y�� N$�j	$�C���,b<"E_��� @�b@���Z�&i!F'�Aa WR*]TW6�m�G�t��Up |���b��B)�! N���Qx `�� b
|��xT
i���~3_c�+�{�`en����)$8����w^�]Ӏnֹ��� ~Zݴ�ȣr6䨜�wf���7���zXۻ,]�mJj8�IJ%5�vI..I�X�wY�Z�Ke9�#��0ܒΎ��KiTqF�F!�|��+ �n��n�#��_���UJU*��Ɔ���� ���Z��H���$b�+ފ�R8��M9,�����}	D/����p�� ݩև�񧛸f��&�Z��H�� ���fa����cZ�<m�[�i��]�	-|����Ӏ�~��nk�ec��L\&I��S�8�g@ŬqYv����g1+�0��vbM������k�=k�"�x	��Ԟ�I&n�o�>��ֺp)w�$���*�Z�I�z��=k�<�� ���Y_��iTqF⎤�,<�&�X��π>��ֺp�o<[��`��t]���w�r����������}w$4'P���Db
wv�{����-�n�LZ!���&�ή͎�b!�D�Ñ�s=v駞ح�S�[���;?7\�����ك����-��lqmlۆt���^.N�`���½�A�p�1�v��Yհ���j��\����e�dswmҤ�lt�<��XJ��t�y8x�@��C��[��Y��	5�b��`3!���3�ݥ��MWkv���prn�K����>����ep�4p�ϴ�u{L<ۅ��y��X�쵳{u�5ck��c�Ts�(Ѝ~m���>ֺp�]�	-|�eC�x�7p�lI��zWNyK��k�����ȫ�����oL�'����� ���Z��[�V�x�S{�u<Z���� ���Z���[�|��{֛��N&�#��>z� ��������� n�j��7+��˂i��g0فى�bdmD�9�B3UR�y:�]�M��=ֺp�]�	-|����/$�8�d���,��V�U*��r��J!%T�!DX7޼ �ϯ �wN��ya�n$�`����%��>��g�ޞ,ǾVWh�c��:m9NK���|��Ou� ;��`w�{YJr$���7$�;�4�'���Z��+�=rk����s�g��7��i�Ӟt[68s�z^5;���$�E�-i+�'��[|�~_ϧ Ik����������o�ؖ���� Ik���������W䍯{֛��9�#��;��ܓ�{=74,"5��l"�F :t ���y����I>�f��J�j��ֶ�o��Z��O)v�37e������7}m*�jQ#��7:�U�ꥻ�O�����ݚXͭ���M�I� IJ�ND�!!���g�Q+m=:�:j���X�۳O'��:FI�fn�幮�������X{_�+u���t���9NK��:"dޮ������� �Ѯ��)Ȓ���r;��U��y��r����K���`uf7����
RRRN+�DB�DB�y�N w}����(��ई�Az潙�'����.a�\�4���V��,Ur�w�����+:�U����`F�L���r��C,��F��0r���;j��yz2D%߽ٙ���R�7#br
F7'���X׺�	�.����%\�bck[I7�n� ��:�S#�}8 �u�����*�#p7�Ҩ��MB!	�`n;�xK_ }e|��xg��sq�ph�+W*������w��`w^��s���7���a��ӊG�թ� ���Un��]�	-|m���v�w�oϼ�9�ly����n
��y'c��8l���ɐ4$m��D�ϮClO(naM��N�덫Z�uv���q��NČM��New���w�k�h�G/N�%�aT�흨p:m��)Q.��fm�E���0be6�OIɽ�rc�bH읎��\kF�t¶<�;r�pn�`�ڃ׸ �m�4E�[Mn�:��r���:�����}�������w/���k��nѳ�K�$d�{@iM�<t[����,Yy�{w�����:*�� ��$rh׿���٥�fn� ����Ki98�III8��g�G�	EPw}�����Λ��r��=�{�))��ӕ��n�Ӏ=e|��x	���L����OT�����a�U%��K<��`gvia��+����ߥ�������F�mIQ6�Un��Ӏ$����������u������~p�눜��!�ʯ�ն)���5��Nb_���}��!�o4ם�\�M\�_� n�x�����BQ�u���+k~�MR�M�t84�,u��JB�I]޻�<�\��_����H�a��ӊG�M9,~����z�p���QGD�Sr9,=UU\Y��+s�� n�x�L�>�Ӭ�Sv�J�.���qXݚX��> �o���{���fV�(G%)(��(ʌN,\�ۊ�\C�5�d]M��'l��M�ο˻�������6!jx�g�����W�z�w�����ojM��7�w[BM��w�
&M���v, �n�&Ni�cN�$i�ԕ���?yX�۫6�@ �+"C�55��nI>�},�f�J�Jd"�V[���`�^ y��B���V�e"�N���pi9V��,�Y�������������lˌo7Lli�޼X���烙-��f�%K�;]u��m ��^��u�~�ͻ����M!	���'������'���	-|�n=ưlI����M�}�Q��`w�^ y��i;I�#�t��N+;�u`���RF{},��������$I�m���}׀ϯ �v�
���"� ����+����rO�u��k.��]�Uw�z� �BI|�$��~�����`���Ÿm�jEI"��0ӎ�\Y�w�<���p:Փm�ɒ�[�\)�X��K[ǭ�ֺp�Ӏ37g��s�{},��[J��DIUf�v��&A����׀y���UW9T�����j�:n�JB�� ��x|�!L�u�=�� ��+v*qT�6�6%$���r��o�����o���B�o��:�WH�$��o�������%��>�}��yt�`$ F#F��,"����j�t�1+	d��7�4&Zl8t�+ �AB��E��X Owi��7 h��@b�bDAf�$�#+
�	0I$�6B$ĉ1	�FI# F$�V)Aĉ�J�)��A��^$�th���	Ԕ RYH`�"�@!XU%!B	#D����% !P��%����6�[tRmN�Q���;:�˯�/XmM�ܑ2�C�ͻ���\f)-�1�]��v����*������+�F�j�8N[N�)z$p��b[M&�d�t\Y
T�rϖ ��5qP�u�#�O:�0��s���*�ӥ]�`�+�Khk�j����t�+��xM�a��м�$;j������OEI���;i�Ea�J
׋��kp�\.�`��]��y
�b���)�eױ0*�-���"`��[C�=]�b�͹��k!�QU�-M�n�L�1��+�Ke^ݲ�k�>K�{K<���^�.��.�,��q�M!yI�n5J��S��g�8
ֹN]��x���T-�vLj`1��mG���2����j�mEb�Z�"��Ki
�W�W��)ڱ�j�t����i�7]0��5�8�[<H8ι�L�¼-�Z4\`X�DIUl�vP&���Z͜�/JD������ �d�� R�

��:�Z��R9����ڃU�ljj�\ 6�nl ��m��I�1���mm*�W��itS�;,u�wm��cSn�q�*�F��^X
�iꀫj��A���Z���4�T��.�V6*��V���פ���k�*�iv�e�У���6�l�f�[%[@,2B�s�q�lk�vZ�8m�9�{ �ъ�մ�$*m�3Ȏ���8��	�vl6�e�m��m����L�+��&M�r<�m˹|�MI��D`�]��K4�mx��+�&��clZ�[&�0��"ځݷl����R���@Y��mmJn�k�����m�EA�ۂݝ��zQ3��Yv,m�U�h�wi^x�M��` �e��X�t��+�U�WM)28��A��أ���m�&⭄�S!�ҭ[�U:��e��[�\�ҩ�M�e:X oY����v�Ġ��X}�����ҵ�`{dt�͎�7=Z2��m�c52HC1�Mk�`l1@#���A �!Ÿ�@�|���9;�j�5.]I�2�K5@��ϝ2��6�m1ś9y^����vQ���5�W����xu�W�Δ�����)��[/hs�9��Cի�t;u�V,[=�#�d�`�X::uq�q#��Rg����(���U�؋��>�t��n�p�ո��≐������&�vI�ί�۝W��yx�D����#�Md�(E�uux��'��};�/n�pޕ��z��3΀z<��x��g2l��ٓ�5���s����:~c�6��o�wwb��� ?=w�(_�7���;���RT�Q')�*�37e�}�� �v�}�rJ��wd�U՗w*q�kRo�=��|�t�'�� Il�7��m�N1�ԕ��ܪ��z�`_b����L��^ �eL�Ckf=4I��xK_ }evwf��s�y���6F*�i��P�1Dk��FN��x���X��̽6Ů�v�{��Ӗ�L�T8%$X����,�͖�t�'���{�2׸����4h�37$��}��S�?�����r��� ���z"mǸ���66��7l�7ծp鑾��s��?)�6�LloLԙ�OGN ���Y_�]8	��cl׺�'V`�w�t��_�7���7�l�?O߿K59:���jsڍ�{[�x6:e3��l�v.z�8�Ɣj���P��c���M��W�z�Nz:����>�˿�%��i&���[|�t�'�� Ik�����	yn�Ckf=4�� �m� 7[����Q)!,��IE��� ��}��{��M�=ӵ�!VT������J}U��׀�ߥ��٥��ɥ�ް�ة��n�4n���+�=k�=8K����z㔥'�b�	�pRPN=)H[v����Ś\��<Zj�W/CgK��y�3Sci�ֺp�Ӏ$��ϴ�},���:N�BpM�����9)�o�����:ns�25:>W6A�)A9N8X�,�͖z�\���S���p}���M�Y7b�j���� ?=w�y�s�o�فq	}@��qj+�^"�������������t�Q�RTRK��U���f n�x���QZ뤵S2�]]]���i�/+t���Al�3��kTWK-�)tw��{[W�:u<�h�|>�� �n���x�78�%�VT����� 7[��D(��P�Po�������7�l�=���W*9J��Xۛ,��Vz�\��6x��zX�bڊ���
NBG%��M���f n�x���>��e?#Vkx�a����=8K_ ~z� �� ���Q�ؘH�����]��kq�:��f�Z�gJ\t��eY���B7-�g���p�ρ1����m������P�>n5�R�%�h	9#iF���p�:�B��mY��V�l�tkmn'����`�t�Ӗ�S�;aM��d������}[�����d�����4[gmp7lJ�"�۬i�E��bs[��H;x6u��[cj�~����v��t'V�%���3�=�;8�«���s�n��ak,t��R&�DI�qà�zXۛ,�ݟ�#�J�>���������n�Uu5Wx����S&�wN ����/�_�\��l�����t�Q�rTRK�_}8�m�lDɭՀ~z� �lʩ*d��*�ÔDD)�n3 9�^ }e|��x!��f�L7��v`�w�t(J"}ϯ���8�o����~?����G)4���W��ۅ���l��B��m4<;��qՀ۪��a�sD�����:np��>�Q
>��UWX�����3��EJP�9	��78�1DDB���`�n���y�s��q#��O1���� ����{�xK_ }e|��x	��V����')�����W����w��`v�w��R��ֵ��l�x�ԛ��]��(��}����������qu[D��랥4��m��a��l��b ٮs7`%��1�[�B�D��%E$�;�uXܚXf��Us���o����M�d����BqXܚg� �u����t��(�P�������/�(���RNB�=�ߥ�}��nE@�`�oB �]^����rO��4�;��
qTN1�lJIa���U%�}x�wN��s��J&[�]}QR�#T��$rXݚX���[�|� ����}�����)[$PQ��Sl���$�1qml��G���ݲ��l���Z`�Ѣ���lԙ�O)w�$����}
_�7�����\��.f�T�� n�y�P�d=ϯ ��� �V�Έ�P�IDU�����ՓV�.�i�,?{��;�۫:�U�w�����-��9nFܕ����9ř�}[�{���$��{7'�ڐ� ���|���Lo��^���p�IN�u� �>��^,�Ӣ���^�O>�sc�h�АۘN��*���vs��plh9�9LU۱��㫂����n���x��\�K��}8���Чi�%Q�I,�͖w6���V��6|�g��/�$���t��T�H�!9	����:�U��\�KV{��;���>��5�Ԓ%%
AI*������V ~z��$�y��`j3}�Q8�
JjE`b��9%	}[�}~'��+ə��n3�陟�����www�y����!���b���=�-�����j�5��\��X����g����v6��<u��ck�a�rF5$�ٙ[N��%��#nzm�=��،j�{<k���6H	��Gra��=�*�쳭jT�۰�3�ҕT�cY�������gs��y��掎��Q���c�8��k�	�Ě{W@��d#u���1�4�tn�N���o�_����g{�R[I��L3��wPN[��1imF�Lݶ���[8ܴ�خ6��h��%����H�۩i$��5~�r�֒^��$���{��9nFܕ��H�۩����Kro��$���Ei$�ۛ>��W9M���=MTd���F"IR�InM���[�b��K�͟|�F��KI%��[�(CN*���/�I%�6+I$�����$nmԴ����7�{���%��p�i�%Q�I��_nl��76�ZI,��_|�KrlV�K4�E�Q&��<��>�&n��H[ul���cJu6&��'�M��j�9ʪJ�)R$9��I�]KI%����InM��I/�6}�Iv��X����MH)%KI%����+y��R�T ��? 7{�~���I.�}>�$�ͺ���ʪm����#e
@ ���_|�K�=��_nl����UT�=����Kro��$�v��Ԏ�'*q��V�I}���H�۩i$���^r�����g��eݶ����.�k1F�m�QI>�$�ͺ��K�r�/|�Ԓ^��$��sg�$�����;qTs���|��YX�n�f�Sc�9۱;n�#�Rpʾ��r7ʮU])wMTqGRT#$�Ԓ^����InM��I/�6}�I�u-$��	oȡ8�JJH��$��د��m������=����K;3W�$�rmQ�"J��+I$�����$nmԴ���!� �!$�EXVR$�F$I�HͺF��4C��*hC�v�h�]�:h"�d@�	�L $BDB���
(UX��h�ȄbA@"D�� B �DpI�U���"H& �'D�D����D ��*�/*��@��y�^r�o}�˻m�w&k"�*A�' ��_��9�ܪ���v�����~_|�KrlV�I}���K��f�h�u�X�_ ����� ?������?{��u$����>�$�ɤ��[���pݭ��Lta�\�ۆ�-���H[�9`�Zg�oa.��C:]ح�����KrlV��6X�l�|�q�S�F�j'8S�n�s]�gwe�<���:p�v�z�oM=mp����R��8�ڸf��*�F�8�G%���f�X�.I��{[��C:�.�{�f��6���-l�ƞ$���:pm�`���7k\�BI.\t��拙�[T���K��9�݉�h�kX.ƮMmiKs/Kt�JU������Ģ���4��@�����־E.�GN���k���I�owe���|�n��m\��X�׫^<y���|�\�vه)�OwV v�^�w]T"n��n�M��|�(�;�8�==�X�ݖ���+����H�G8R�uf�[u�}�){��n�N����s��6���r��� �2(�2�Kәure�Ml:�`�`��ݤ��Ut��t�y蜶����ۮ��QЁ5��p��������]�8�oI=:����e�u�7C��pn3�Ӥ혖��e��3�Uzk��l�)c����CX����lq۶y���У�p[�p�F�7D����lgY9���[����٥��<�Ӻ�]���{��>�ww:�ش�Z��2ӎ�\Y��]�^�:;0s�6;Fo*hKu�l�ٝNZ��~��	��z�N�ٲSwm$��7�H���:pn� ����I����I�R�Cr�q�?W�����'�|�Ӏ�@��S�E#ITbR��� ���H��z�N���4�Է57�mp������dt�=��p#�y_�a�+��z��2�%�<����2m�ng]�Yge�)�C��-�6�� ��� ��f��u�� {�� �3ބtȚ�E%H�`fd��V��*|�D(�%����t����^�Ss`}��cR:JN*T�ۅ����`6���3�]Ӏ6��ڪUeM�hI�i� ���y[��Ӄ��qc�y�K��*�F��$NK�z� �6��l�u`���>٧D�$c��Kh��J�j6z���v�8KO��;e�\����L��;7���h�m��w���u��w�D(�!�]Ӏ{�+�T�QHЈ�RWw]�}����vi`gri~�W3Y�dU�!����� �>�ަ�	����m���]��u�	"�ܩJ��rKW*�d�N ������>�׀l���)���E%E"�3�4�:����͖z�U��o�_�78�"c�;Dv�;U���5^������r��0+6�����q�(�
T�ۇ@տ�; �se��+w������IV�m	=M5���Ι7k�p���=>n��
!BFR�y%Q���D�I`f?yX�t�=��p���\�)��X��&�mMU���l�=>n���x��/�	�"�TO}�wrO��!��k"�F�F���:����͖z�U��ɥ���4�N��Q8��q�U���6=:۵�6��d��n�cW,6pd���N�J$��>��`w�uXܚ{��9_ Ş�7o�#�9	II,�����f��u����D|�PouM�M66��<X]� /;���^�;��cR:JN*T�ۅ����`���=�np9Kל`���MQr^$������������OGN �����9�r��h���R mҨ8ʺ�@��n���R�]v���Z�=��v�����/KFf��=�{G:� ���-�#�:!�UX���bKő�e�9:b�nq�e;`�#v�����< V�08C&�J�R��vP�����`\J�{�W,:�q6�z�[6-&��ŽX�^��Mn|9�h���kcd��ѕm:���1���﻾=�5rL�
��6�hza�j���������l.�i[�Ë�r�]��cm�������OGN �־ ���	��9�9�"R�r+;�K ����>��`w�5_��H��=8��H"4�� =�׀����J&wi��]�w�Ȫ7���E$��UĻ���$W���Ӏ>����Y+m4�x�Lm��{�Ӏ�����W }e�m��������NoP/���n#9����s�5�4v�68s�73����s�|t��c��π�����W }e|�xLR����n&$��}�U�O ��w�=����~��~��w�Ӏ�ˮ�=Z�5�6���Y^��s��
e�0O>��^�"��������n����B������0�� �se���i�L�)I���7�l�>���D-������^���`n��TӸ�:N
p%E@�%ۅ��{��6�%k��;���ۮ:��Χ��mkw[8�ʸ�k�'��$t�=*�6=K�֚����"&G���w��^��7Ե�wwDqJhp��`gri`fd�����W% �+ �j~:*"w�\�����������|t����p�$���e\����Ӏ�b��WH�������?K�XС|�V����=���3&�����Jr"(��5Ť!k�㭜�ًn)C:��3=s���R��h:1�y�[Z�ԛz����������9B_�=<��S�t������=8H��}�U�K]��9��3/Zj��R5)9!`f�� �/]a�'�u�]�~�E�k5�M��4n�p�W�K_>�znH�D�Z�T��_k;��J��X�K566���������t����&{nV޳ZR��3��A1��K�������4<����֢tp��+��zI���~��� ?=w��~�<�� j[�.��=oL�=#� }e|��Xܚ_�UUĎ�=�i�)9¥8�l�~�� }-|�t�=#��E�Cdn&�##�Ia���Iw}�`nm�{vف�(�>�׀j��H������ަ�	���zGN �����ٹ" �OH��$�)��)&	U��J��))R��J��4�!rt�
Y�a�8|y]:)֊����w��
�"$��+ �i! ]�D�0!"�����q4+	�0�N?EyǾ���_��i֑�7f��m��4&���SM�� J�ٔsc�����t{Qָ�ݎ۵����1�pJ�8�:ڪ�	��啴���c��yI�Pa�nG,�Z��x�����%�p���hWdA�S�'R��a��������#�t�ף&��	�3��kdnuӶyN��]��ě�V��Ǔ!��]��E�qrM+yD#2��<vz�vļ��ٜ�g	Ûe���i�u܆��X2�q�-(����8��wS�awH=��aI��a�n�}fM�q^q��1u��=hB���$Hj��p��7O:ɵƸge�˧��V��8�r���ٶe����(x[�7�ƍ�`���`&�iZ��8�Z"����<�˨Ҹ�T��Gc3�N�0���ݾ[�M���mw-�/V�ki-�+�R���Y����`���+��Y#����e�$&����ճ�NÎƱ�vN��"�&�3����i��:��Ws��Kf�:U��U��c u.7
��kpp�Vx:rYf�������׀lm:l�ۀ�]AK,n� cT���9��*�]��f�q�V�|[���逺k�*�@U@R�U@H-��I�m ږ�m�%�q�l$�ɺ!��:�Lҭ@T�gj�C��Mۮq&�[[,� ,1oU�i0kX6�ȑ�T���Tj؀{<��ۍ� ��-�zx����æ�h�l��V�9P���7\���]�&CҴ�xM�)�-�iq���Qt�"��4�8j9[ʫі0,�`�7l�;eE�SV�꠺�nYPds�)-תl��r�훤r���;s�]��U��:�!��L����$�!4�đż+j�qd���K�W+���/y��i��s����ۧ�V�v6�a��kY��W[/<�f���nq�%���(H�*�q�t�3eY��l��ѷnЮ6�lf�m���]{t�fFm�C\mm'	��WP����z�-������ :<(�NEO�S�=(����ʠ>D`����}~��TO�A�͛����+M�Ӯ����i{I<��\O�����ud��c��s�b˚:��M<��&yٮ'�uƹ��f�f����X�ܶ}x/�V�;c��M۵�tvεmK����LÓh�˅�t#��t���K���8\�-��L�����$�ƞ��:�8ۅg�����KvD̂�U��p�����oe�ݓ&7\���w���ȿ0��}���(�JSs[ɹ8U[i錧i���І����Bp�t�[�������l�������Q脔z��_��pO�:QG$�dbR��� �7e��ɥ��ɥ�������o����6=m���π����8�[,��I�G*!�G%��W9\��y������BIL��^ Ի��Z�ǆ6ē8	#� }e|����Ӏ��eǚ��=z���ɹ��w]f5ڐ�.�X۶$'tg����7�us�T�q��J�p���K �[�}�Ϣ#�n��<�>
���d��e���'=�f��. ��Ch����۶� ���}	Dɫ��VZM�ǏS|��8	#� }e|����v��ē�ŋS�M���[0��x��x�Kל`�����z�m�n�g }e|����ـn� �(Q��J*�"�M]+���ϵI��rkn�ۆ�I�p6�t��ٲ�*�O=sۿRP�ȤR5��������3���I8�+�'�J�޽ǏD��|�t�$��������L�*��i�1�$��I8��f痯�5(5tI��y�'����}1J֦�m�f�bI�������OGNH��}�J	-hi�M=m����OGNH��Yo�o��~w��f��J:qeuƤ������.���V("y�4�7��C\5�=m��Ӏ�������W�}�ն���n�cr��w&���ă��K ���������T�(��JmF����6Xۛ,�UU%��Ł��Ł�f-��REi�8����7�l�7�l�q�J��޷�X�X�ש��ѱ��=8	���Y_ }e|�iCF�o5]���*9p�.]l$�k�}�m
�r��t�m�c:�١�3N�6OI??_��������+�$���)Z��=l�R�*�� �ۼ艐�>��|`�_�UUUI�{^��ڌRSQ�$�s��7vه(Je�0��x���Rw����I%���T�v�X;0�n�9BJg������5*j���m9M�*������s��������'{�lܓf
�"��}�xkƳ%�d��n;e�,ĸ����xj���n!� \���jE+R�����##���]�����WlQ�gQ�����rl�苗����;W!-�2�=���n6eN�݀���Ͳ�ṗ64�n���	��eSn���v�C���m�!�j�;u���\cu]i�*yT֒Ӭ+�k0�K++�x yIٓ&��Z�Im��!8���uWW����M���j���Z]u�̖�M�[h�Q�]7ھ�T�Ι��s��U��B���g�π/�|����t�=6��,lf�66���_=/g}8�+�'�J��kOE�Fě|����t����,��6J��=m�`�ƛ���p�W�J�	%��%�+Z���a���&p���J�	%��7�4�h�~��B�5"�Q�#�-8��M�Wq�mṁK��uؑ�e�0��uˡ#�b�������oq�����Kı;���ӑ,K��nzT�Kı/=�fӑ,K��OXk[�kF]f�32��X�%����6���"���Mı3�=*n%�bX����r%�bX��ײ��X��#�ޚ���&�ui�n9W���#��b{�=*n%�bX����iȖ%�b_wّ7ı,O��p�r%��n��~u��2V�:@�{�oq�X�%�}��r%�bX���dMı,K���6��bX�'�sҦ�X���~~[���2L�������ŉb_wّ7ı,O��p�r%�bX���J��bX�%�}��r%��ow�99�~���+���Q����������ɶʂ0�Qn����Wmo:�Y���Mf�"n%�bX�w���Kı=۞�7ı,K��ٴ�Kı/��ț�bX�'ƾ�3F������.��"X�%������~ ��j%�~��ٴ�Kı/�~̉��%�b}���ӑ,K���5u�&a��MkY*n%�bX����iȖ%�b_wّ7����ḛ��{�6��bX�'޹�Sq,K���t�L�������fm9ı,O{��Mı,K���6��bX�'�sҦ�X�%�y�{6��bX�/�z�Z�kZ2�52\̉��%�bw���"X�%��\����%�b^w�ͧ"X�%��{[���!���}��}�R1�8��N�եz�;YM�Z��f���'���9�k�����j�k5��%�b~�s����%�b^w�ͧ"X�%��{[���%�b}���ӑ,K��鞹��fL�ɓ5m̕7ı,K��ٴ� �I��� �	�{�BE$N�{"(���X��O_�[�5�-3Y�.fm9ı,O�����Kı>�}�iȖ%�b{�=*n%�bX����iȖ%�bw�k�30��]Ks5�2&�X�~DF�w����Kı?z��Sq,Kļ｛ND�,��!�B@ 	 ]di���9H�#��Wi�k$e'"TD�ֳ�"X�%�������%�b^w�ͧ"X�%�}�fD�Kı^��B�B����˙�uMX���Z����$Gj6���v�\ez�:�\�Rs��3i���������+c����{��Ľ����ND�,K��̉��%�b}���ӑ,K��nzT�KǍ��w��ＺP��f����oq���b_wّ7ı,O��p�r%�bX���J��bX�%�}��r'�uZg)綼�n�n�q���9Vr��BX���p�r%�bX���J��bX�%�}��r%�bX���dMı,K���ܺ�ֳZ3Zְ���iȖ%�b{�=*n%�bX����iȖ%�b_wّ7İ?MD����i���������O�S�B����X�%�y�{6��bX�%�}�q,K��{�ND�,Kݹ�Sq�r��G+]Wt5)C�AƠ��I��;Y���y��(9�x�]� gHF�۫��K;���,WG=C�m]�<ƞ����v�Γ�h^�v�I�Y�[ĎYj�M��.�66� `G��4냬�����.������U+n)�[�q���8�(v�1ݗv�N�3�wm�gG9`o�w{�ou���ui�X.��
�����Ȧ�7m��I.bJ�42F�{���{��w���|��-Ն%λBN���Nlzv�ݥ�����'`g��nf]\��V��h�k2fk3��Kı/��̉��%�bw���"X�%���������5ı/߿~ͧ"X�%��a��32��d�k�fD�Kı;���ӑ,K��nzT�Kı/=�fӑ,KĿ{ّ7ı,N��}��jkY���.��"X�%�������%�b^{�ͧ"X��� ș���2&�X�%�����ND�,Cw�9��#=�`�+c��{��7��y�{6��bX�%��̉��%�bw���"X�%�������%�bp��<]L��k5��.fm9ı,K���q,K���k����Nı,K��Ҧ�X�%�y�{6���7���{����-�C�؄���Ιx�R�q �5�m)��0je:�]@���ݭj�fk,�f�"n%�bX��}�iȖ%�b{�=*n%�bX����iȖ%�b_wّ7ı,O����uK�f�f����5�ӑ,K��nzT�8�`5"�l��Wb
� n�}Ĺ��siȖ%�b^��dMı,K��m9�DSU57{�ݯ�xdj���w��7��,K��߳iȖ%�b_wّ7��*�D�O{߸m9ı,O޹�T���R9H�fCV��!��$r_+�,K?��k��fD�Kı=�~��Kı;۞�7ı,K��ٴ�Kı;�5왙p��[�fk2&�X�%��{�ND�,K���Sq,Kļ｛ND�,K�����$)!{��*wwST�mX�撫��0��nx�s�kK����i�T�ib&�m���.f�3Mk3EsX]fO�X�%��\�*n%�bX����iȖ%�b_��ț�bX�'�w�6��bX�ߜ�}����[��oq�X��{ٴ�Kı/��dMı,K﻿M�"X�%���������{������~��Mr�E5�����%�b^���q,K�����iȖ1����B�'B ]1�P$,H�
4bE��lPee �BQ�T�c@��a�T��(D(E(�i���
I)$JA�F�KZҬ+��(��ZE�����H�؅R+�Z�)��c
����!��3dt��$Q��� �R,��� �D6�-m%H&�&s��iF��QN�	�`
��E4�AvxS�mD<u]��ȟv�Mı,K���m9ı,_w=uL֮j5�a�Y�7ı,O���6��bX�'{sҦ�X�%�y���ND�,5]��2&�X�%����˪]k.�na��ɴ�Kı;۞�7ı,KϽ��r%�bX��{2&�X�%�����"X�%������r�0s�ooV՞2ݮp��;��i��^�:��ܸ�Wc���#T�f�nd�Ȗ%�b_���m9ı,K���q,K��������^�Ȗ%�����Sq,K������W3Y�CZ̙s3iȖ%�b_��ț�bX�'�w�6��bX�'{sҦ�X�%�y���ND�,K��^ə���5��0��dMı,K���6��bX�'{sҦ�X�V����߿fӑ,KĽ��2&�X�%��]��s5k3EsX]fND�,�F�{��Mı,K�����r%�bX��{2&�X��ځ�Mn'�߷��_�r��G+��Қq��J�p���%�b^{�ͧ"X�%��*�w��Ȝ�bX�'���6��bX�'{sҦ�X�%���n��53Y����.֐�������������s�:�@���we�Bk�R"������oq��fD�Kı;���ӑ,K��nzT�Kı/;�fӑ,K�{���N���c]ow��7���x����!�����\��,O߮J��bX�%�����r%�bX��{2&�X�%�����]R�Yus�k�"X�%�������%�b^}�fӑ,������fD�Kı;���_�r��Esp6�T���68ݹ���X�"(�D����6��bX�%��ّ7ı,O��m9ı,N��Mı,K�����]f���k2e�ͧ"X�%�~��"n%�bX�}��i�Kı=럥Mı,K��{6��bX�&)C��@@�[ٯ��ѻ�$!f�d��Z�i�S�N�^'�Wn��,�uӶٍ�ӷ�Iź4m�
���霓h�I2�R^�m�)! h�g]�:,���B&��I�#D�X��:��[��j|�,�M�h6C�[n�<a[�
5 ä����$�'
�o&�ֳ�ݸ6_3su��#јѕͧ���i���-��wD�S����/�f�D�ڮR�pz���i��j=�o�%6dy�k�K���E�Ų[l�;QqI����1�wjN��@�]-8�O�X�%��}��ӑ,K��nzT�Kı/>��a�(��蚉bI
w�셄)!I
HZ��T�Ъ��Lf�ֳ�"X�%�������%�b^}�fӑ,KĿ{ّ7ı,O��m9ı,N����jj��
fMkY*n%�bX��{ٴ�Kı/��dMı��5Q;�~��Kı=럥Mı,K�������)�ۊG%�9H�#�TU3��ސ�n%�bX���p�r%�bX���J��bX�%�}��r%�bX��zꙭ\�&k,�.�"n%�bX�w���Kİ�QH���ND�,K��߳iȖ%�b_��ț�bX�'{�>���Q��\��!�ś�ɹ8^Pն���i�k�4d ��#�	�ø+��ND�,K���Sq,Kļ｛ND�,K��f@�'"j%�bfﾫ�|r��G)�hz�T���68�nd���%�b^w�ͧ!��(� | 
.���K��"n%�bX�����"X�%�������r��G+2�nH�)������!,K��fD�Kı>�}�iȖ?ʄ5Q=럥Mı,K��߳o7���{������jx��]Mo�bY�T�E�D����6��bX�'��?�Mı,K��m9ı,K���q,K���}�\�CZ��\�Y�ӑ,K��nzT�Kı/;�fӑ,KĿ{ّ7ı,O��p�r%�bX>���\չ���2s��\�f˺�1�ݨ	�'b6��ݮ�(����v�������dg$[qՕ���o%�b_���m9ı,K���q,K�������&�X�'�s�����R9H�v�mz�"h��m�#��_D�,K��fD�?��MD�;�~��Kı=럥Mı,K��m9� WU5����uL֮j5�a�Y�7ı,N�߸m9ı,N��Mı��$��(��Mĺ߽�ND�,K��fD�Kı:���]R�Yus��ND�,K���Sq,Kļ｛ND�,K��fD�Kı>�}�iȖ%�`��{w)r���3.�̕7ı,K��ٴ�Kİ���w��Ȝ�bX�'}��6��bX�'{sҦ�X��$/�����"�ȹ�ԅ��
���7`�-��m��u�#ncI�jnM��t�L�˙���.fq>�bX�%��ّ7ı,O��p�r%�bX���J��bX�%�}��r%�bX��Y��.kh���̉��%�b}���Ӑ���j%��\�*n%�bX��~��ND�,K��fD�Kı>5�{W3Pֳ4W5��a��Kı;۞�7ı,K��ٴ�Kı/��dMı,K���6��bX�'Mw^���M\�!Lɭk%Mı,��DF�D����ͧ"X�%�}���q,K�����"X�PC�S���Tغ7ȗ�=*n%�bY��<��L��S���K�|r��G)	~��"n%�bX�w���r%�bX���J��bX�%�}��r%�bY�~o��GNdc���讞Ҧ��P�x����*\�ԅI�z��
ݿ�{���p��/Jf�3Yfu��%�b{���M�"X�%�������%�b^w�ͧ"X�%�~��"n%�bX�~��.�u����ə��iȖ%�bw�=*n%�bX����iȖ%�b_��ț�bX�'���6��bX��'�r�.f�Y̺�2T�Kı/;�fӑ,KĿ{ّ7��S�i�2'�~���r%�bX��\��7ı,k2mG�I
�B'%�9H�#���{2&�X�%��{�M�"X�%�������%�b^w�ͧ"X�%�~~F~��-��+��������ow���r%�bX/�!_߯?�O�X�%�{���6��bX�%��̉��%�bT��P�D��"v�n��ww�����D��f��E�ٶB��kf݌�a5г\"�aq�T���۞"�Kɸ�"Z�:��+���c�M�\�*渊N�ZX����][mv5m�!��^n�9j��	�Cۄ:�G�͕v�䇋rVk�R])UON&�0=S����8����܆:�V���.���g*AW��$�bض��}��m�~�ls�[\�pM� �//n5���w{综���K\6�͝4��a���[�ܦ����ĎM��\8�nîin�T��Zx��->O�,K��nJ��bX�%�}��r%�bX��k�C�g"j%�bu��!~!I
HRBj�qSV��])R��kY*n%�bX����i��GQ5Ľ���Sq,K�ｿ�iȖ%�bw�=*n%�bX�>Ξ5��Fjk5�k.f�6��bX�%���T�Kı>�w��Kı;۞�7ı,K��ٴ�Kı}�nkFkW5	��0˙�7ı,O���m9ı,N��Mı,K��m9ı,K��쩸�%�bu��ܺ�ֲ����6��bX�'{sҦ�X�%�y�{6��bX�%���T�Kı>�w��Kı;5{�k5-іW$�����iu�S��mlJ�g���b���..��و�)�uB�w��7���%�}��r%�bX��k�Sq,K���ߦӑ,K��nzT�Kĳ��6��q�LrB'%�9H�#���{^ʛ�C+���b}���ND�,K������%�b^w�ͧ"]�7������ޚ�t��Q����K����6��bX�'{sҦ�X�%�y�{6��bX�%���T�Kı>;�r�kT�f�au���K�� j'�w�T�Kı/���6��bX�%���T�Kı>�}ͧ"]�7����>܌g�:��=�7��bX����iȖ%�b_��eMı,K����r%�bX���J��g���{�{��~_���3F�5,� ���(�����vѫv^65ץ�VQ\��m�f�"p���O�]9H�#��R�?Eʸ�%�b}���ND�,K���ChA�I���7�{�5�5����e�e��$�H����n'�X�'{sҦ�X�%�y�{6��bX�%��عVr��G)��tߓT���'#�ND�,K���Sq,Kļ｛ND�߁ �<W�x	�D�Kߵ쩸�%�b}�o�iȖ%�bzt�~�0��V=�7���{��?�{ٴ�Kı/�ײ��X�%���ߦӑ,K� MD���J��g)�r�`o�)t�$"r_+㔄�,K��쩸�%�b}�w��Kı;۞�7ı,KϽ��r%��{�����#��M�n�^nB��u"�X�w6����l��A�Tt�%7(�X���a���7ı,O���6��bX�'{sҦ�X�%�y���ND�,K��{*n%�bX����fkT�fɬ.��iȖ%�bw�=*n%�bX��{ٴ�Kı/�ײ��X�%���ߦӑ,K��k�WY&����dֵ���X�%�y���ND�,K��{*n%�bX�}��m9ı,N��Mı,K��^5��X4��#��_�r����r�y�.U��ı;�o��r%�bX���J��bX�EP��]n&�f�㔎R9H�;�X�F�e�J�H�V%�bX�}��m9ı,N��Mı,K��{6��bX�%���T���oq��_��ＪF8��n[)c�k����D�Nș�x֯&�=i�sd"4{�i��kE�Y.�2m9ı,N���Sq,Kļ��ͧ"X�%�~���?�Ț�bX���m9ı,O��g�l3��hx+��oq�����߷��Kı/�ײ��X�%���ߦӑ,K��۞�7ı,O��w�Y�g�ա������oq��������%�b}�w��K�5Q<z��Sq,KĿw���r%�bX��g�KN+�#uT{�oq�������~�ND�,K�nzT�Kı/>��iȖ%�b_��eMı,K�{�܍�rJU)7�|r��G)�;sҦ�X�%�y���ND�,K��{*n%�bX�}��m9ı,O���J3T�*��F,5$ �#����%��H�`�$D�K+t�I�Ϡ|��H��QMC�:E�')�T�{1Gb�mwa	�5[@P�h%M�W���
@�i:D(n��8V��s�ZTQϪ�FvòInH�����t���ϙ1&ѹi�<NH�lF���Uti�8�TD�0��]�xs��Uбt�����Ҩm�y�0Flܪ�zr��6ڋ�X��bzx3�Ҹ9��t�:��A�����.9	nv5u����q����!�LS�r����$���A�\ttvE4?��>;�>Tnld3�uۧ($O2˛���Kg	�ll�[��'��u�V���
����mV���*�͂�@ݓ<Q����:;&K��;�l���`��9�݃^�T�jv�������WZ�7��>|ɼ�=l���m�Z۰՛��Slŭpul�`Y��6�ڬ�s˓=D��s��X�PNS��bóm�Λ��:����2:gD�v�b�j`mcq�R�j;:�M؞�<�bv�Y�ڕn����&��@W6�!�����s���
Yj��[�^Y�\��W���4+9n9!�rծL�y*}�j\$�b9�趔V�V��ճU�xƇu��l�3��cS�[d m�����l �@j����b�j����#t)�1�HJ.���hڭRpT��)�p n�i�'N��P@V�ۭ[�Am6�Lkh�Ky��9��b�m��F�Nr'�ҭVXL��<��`��Ye� u�-�z���aSl�4�P�
wjG ��I�����W�i�f\�A�:�6�ma�{h�<GVQ7&�\	�n89-�����y�B���/-�$U�!�
L��Ʈ�U0۶mm�i���g\�Ϯ1�ij�V��e�v�PS!��iؗ	R�n1�z˵),l��l:
�Wͻm�kj)�L�v�0��ҭuJk��� ��,�6����Gώ�#��}[,�a������HC�d6e���+VQ�|�zCY6�֐@�@ns�M_&h�����4��YeӷLM�[��՝:kףƥ�P�Sѱs�[<�v���nz�WBj3v1���Na�_��@)�z��C��Q�%W@���'�/¦"�S^��Zֵ�%5�35�<T��KҚG�\��m:�h��[��!wq���ۑ٫�s�Z�;'�'��F�ˎ���i��e�:���jݐ]X��#n�������h7��㘫�xW	f�����M�nY"3���k��lcs�q�k��N3H#�M����oY�Y�	`pA�����F܏A��NOI7"v^��_�v�w������1G$��3��8�	���ϳ��C�W��v�ʼ�d�Mo��|���#l��=d5�d��ı,K���ٴ�Kı/�ײ��X�%���ߦӑ,K��۞�7ı,O�;�xֲ�a�Y�ֲ�k3iȖ%�b_��eMı,K﻿M�"X�%�ӷ=*n%�bX��{ٴ�O��L�dK���sZ3Z��L�Y�\̩��%�b{߷�6��bX�'N�����%�b^}�fӑ,KĿ{^ʛ�bX�'_���8Yl�a�|�7���{��������bX�%���m9ı,K��쩸�%��	����m9ı,{�}5��O4<�w��7���%���m9ı,K��쩸�%�b}�w��Kı:v�Mı,C{�?��6^O�'��׵Zt6��t�k���l��c�8{1���Ept= l�f)�s��.�6��bX�%���T�Kı>����r%�bX�;sҦ�X�%�y���ND�,K��5�5��f���u�f�"n%�bX�}��m9�4���Uo"dK�?�Mı,K�����r%�bX��{2&�X������߫\�Pu����w�{��,N���Sq,Kļ��ͧ"X�%�~��"n%�bX�}��m9Ǎ�7��ܕ�<�nVǻ��ş�A������fӑ,KĽ��2&�X�%���ߦӑ,K�Bj'�U�\�9H�#��Vem�Sq&�NFܹ���r%�bX��{2&�X�%���ߦӑ,K��۞�7ı,i}��|��R9H�#���ӌ"�I8m��[fg4�Ƶ%fۤ-�-v�a���2Ë���U����c]ow��7���'�w~�ND�,K�nzT�Kı/>��a���蚉bX���fD�Kı<����Z�h��f��fM�"X�%�ӷ=*n%�bX��{ٴ�Kı/��dMı,K﻿M�"�oq��v���t5�,��V=�2X�%�y���ND�,K��fD�KD4��$"��(@P(*�ӆ�n'{��6��bX�'�nzT�Kı>�I�5�3Y�SY�2�3iȖ%��2&{��2&�X�%��߷�6��bX�'N�����%�b^w�ͧ"X�%�~~F~���g���=�7���{����~�ND�,K�X����S�,KĿ{���r%�bX��{2&�X������>q�ڑz�4��r�F�86���Ngz��Ơ�V{j��������Ӝ��L��Z�N'�,K��럥Mı,K��m9ı,K���q,K���ߦӑ,K��k�W1��\ѣ2ֲT�Kı/;�fӐ�c���b_���q,K�ｿ�iȖ%�b{��Mı,K�޼kP,f��k������oq������Kı>�w��K�!�������Sq,KĿ{���r%�bX���5�5�f���h��ț�bY��D���iȖ%�b~���T�Kı/=�fӑ,Kh�`>�)���{y�7ı,O>;��Z�h��f��̛ND�,Kݗ=*n%�bX(��߿~ͧ�,KĽ��ț�bX�'{��m9ı,Oz�kZ�������.(1��p۲�L ��U��L�qsp�nֻO�c���(�Bb�����%�b^{�ͧ"X�%�~�"n%�bX��w��Kı;�sҦ�H�#��Vd7Z��G1�ܗ���bX�%��̉� ��MD�=�o��r%�bX����T�Kı/;�fӑ?�U5���_�ֲ�k54[�35�q,K�ｿ�iȖ%�bw��Mı���j%�߿fӑ,KĽ��ț�bX�'ƽ�kY�MM\�L��Z�M�"X�%��˞�7ı,K��ٴ�Kı/��dMı,K��~�ND�,K���M\�Mk.�h̚��J��bX�%�}��r%�bX w߳"r%�bX����m9ı,N�\����%�bA�������jE�W
��q���/WX�F��i�tQ��c��u����t��9���7m2���9b�7���j5˘���������3 7u���Ou�c�]���P����y��#�p:,��GR��[mf4�������}j��ͷO9����̮·;��r�6^g�q[(dу(���[ �OcG+L�Im@���n��������wv��_�Ӧ��9ծ4�-u<u��x�ۧ�M�諭7����ܭ��YH�������d�/}�2&�X�%��{�M�"X�%��˞�7ı,K��ٴ�Kı{�n�E̖幙f���Sq,K���ߦӐ� � �DȖ'�������%�b^���ͧ"X�%�~7ı,N���K�f�r�f��̛ND�,K��=*n%�bX����iȖ%�b_��eMı,K���6��bX�'�鞴ˬ&fj�ffYs%Mı,K���m9ı,K�u쩸�%�bw�ߦӑ,K�P?�R�Oߥ�����%�b~����W%˫�Mk2浙��Kı/�ײ��X�%���~�ND�,K��=*n%�bX����iȖ%�b^����Z)ϚKng�'"�$���Ƣ��Q���뙔v�t�g6S4�np/���bX�'{��m9ı,N�\����%�b^{�ͧ"X�%�~79H�#��V3scQ��#T�)��|%�bX���Sp�"�xC� �aRB����_�RB�L���wm�Ͷ�[�I�X��	3�>�� �J�	#�<GN{#W{�=����X{�\�%��Kwg�:d��>��`v�6�uID��u����8�k�������5~d�sg���H�\�,����<
��m-	�×�&��Z��/��ㅖ�V*���m��[� ����Q���0�=¨��H�$�	��>��`I_�8	�:p�mZ�z��܊'%�}����d������Ur����Ϧ����zћQ��$�]��$�)m�����x���6ʖ��V����$��OӀ>�� �J�	#�ꉗ�z�c�:�u�×[Z��Dg��S�%8�c�ݴ>��o�{�۟��J쌯=Y�o����ߟ }%|�Ӏ�#�=�]ůu'�M-z���I_$t�'���[_����Ǻ��c�����|m�J�=�׀}׀{�����mK[5��B:p��ܒs��nN���D!�d�(��]�=7$��s�֋�&�4\��i������W�zGNx���UUs��o���*H��)���n��I8;i�q�k��<��5�*��m������W��)5!LRG#���~�fM,�N �Z�夸��#su�����f�6ـ���ۮ��S&����i���6�`n<Xٻ,�U\H�論��Ł��6����J��Rg }-|����t�'���{�5�Z�$ГK^�m��W�OF�|m� ?=w�5��ZQ��K?9U��]��Wf���C����gu��/����m:�ƭ���0�C�8s�]R\QEӐN�k�tk6��5�K:�ln-+��^T��b�m�Wnܛlv鶕�^z�h�:�N��sv�U���P�|z�Dl㰠��u+Ԝ�9��m�g<En]�S���r��s���ŧz:�Z3� U�nun����&��d�ə��#�@�T��|O�̌q���2��ɶu��l+<'����f�K+��eЗk����V��=~�o}��f ~z� ?n��=[r�RR2�䅁�2i�r��}����K;�K�W9I����'(r46��S8߯��K_=8	��3�j
&�)���rX~�r���)�7׀=w��6ف�g���ړ}Q�d�%!#�������UU�m����K �7e��^KR��RRsh���K������9�]8̜s۪n�i�����cnVRAY�nn�ͷ�~?u�:z> �D���p�=�-ŭ�4�5����rI�wٺ�� ���)2L�����HGN����I�_�Z�$ЛI=z��_ߟ=8	��Y_����b׈i��o��:pӀ>�� �Z�{ۋ7[dNR�B��2i`z����z|������K:�kqНH.A�G��ė\N�b�v'�V����n��#;�+���;�G/kc��	��u��>�� ���	#�2GN�m�Y�V�b56�M����I8	�:p��߳�7K=�:�@�)	���Vd�����
��5�GDKH�H�+a ���<�#����~W����I4���0"�!�'Q����	�1t� �B��h��@ E�I�[�$ B0��' ���	 	��UC`0J���$����a �5 �!P!RT`P��HP�aD�B(@`Q!@� ��	�FIY@�A J��*��#SA� �*�B� �D��"BP"����	#RRI> w֣��
��bB��@��D�@�eF�%�X1&�:dA��JĆ�.�eaw"y F(�Z�@>Uv(��
���u�@Wb�P$�Q�"�.�� {�� �/]5C�Re9M�X~�R�ݿ�{��>��H��L�n-o��ı?�Uf ~m��>���n��5n�3m�>��34bY�� d:���7=�m	(�M;��Y�Ԩ)Wa��+����׭� ���	#�!?���~��2�}i������D�32i`n�l�ͻ����(��
�p�t��IH�6��$����� �we�}-|�Ӏ�%3�����P�Zk� ?6� ?kw�n�#�C�3JAk,�B�$�A�HD D�"D�"A�Ҕ�!h`.�4E��A�AH�b�@"<��g��nI�j���K������i7�K_�3?�-���K<Xۻ,�ٴ��	Rp��7���U��I͔#����t��<:�vbn�3cƞ���ci�����2GN ����k�&m�-ktM�j1<I3 ջlϒ�S!�� �w^���f�qkx-Mn%��4��[_ }m|�Ӏ�#�=�]ůSm$ާRK �se���K+�4��+�K�������mԔҕ�)%���K|m� ?6� ?n��>�H��	@QX!'��f��5��u�L�[���Y�KWR�س1�j�g�*Xnz��y{�R�v���!�ݲv��rIZd��\\E��I	�g����X�Ψ-�"2tÀ�q�*v0��2�[sXWv.YΎ��8c��-)UI�kq�X��6ì�r��Ey����v��N��۲�[@$��M�O�H�l�{���� n�`����n'�6뭵\U�ﻻ�>|�)!ݡ�7)�5�R=Qn�� �//c���|��~Cӛ$����<,�Q�[l�{?��G }m|���GNp�*�JT� �H:JB�>��Ӕ�w��`n��`ew&�q�5RE$�)#��`nl�32ig��*��-����;�zX֌ڎ�q��JBI%�$t�&z:p���Y_3l��4����ۅ��ܚXٻ,�Z�H��{5�c[��61<{� ���Q㸑�g�amQ�t���j�i�͊��nF�zbX��I����޵��Ӏ�z:p�5�Z�6�M�M6��IϽ����O*�Q6��7�����t�����Y���x��z�=m��Ӏ����K_ }e|���7M&!'���g�� }m|���GN�%3����lX�n�p���Y_$t�'���߽�������rp��z�b�6�Ғs\�m�ӹ\ۊ�v�]:l�N1�TUѭ��o�[��GNx������Iq�mkKww[m�GNx������W�L�*M`$=U1V���|m� ?6�I%BAz�{���7$�����t����&�Ʊ<bL����>��H��OӀ�ɮ�׫{�I6�]���x(�Z�q���0��6ߟ~�}�:���'S�3��Ƴ)s ����sE��)��
i؎ۺn5�r慏[|�t�'���K_ OJ�	�R��I��	<M�p=8�k��_�8L��fk�Ǐq�,�l����/�|�t�.z:p�Itf������z����ܓ��=7$��s�rqx&���_�\��UW;�{���Z3j:���Ф*�� ��fйk�? {�� �ߤ����u���n�6�l�:���ڹq��S�\ه/Sô�6�vYg�Y��OL�.z:p�����������6�響(����F�`n�%|�Ӏ����Od�qkՍ�ֵ&����_$t�.z�p���{,��q�x�m4,o��:p=]8�k�%|�����ēi���6��\�t����,����M�>@�G_}2��p���FAE#c��F�90�R��Rk����Nt�GgG/k� ��s�1���s�f�2Pv�nL��xl�[-uhX�̭I`��������v� ���A.�[K:���8�3Ou�uR��&�^2�����
h��m��Ý���m�o���T��-����8yCg��\[G&��h+�|��n�6�22DAO����!�NkV��Zh�d�3]�62�m�&�0������+�b5�!�����8�"�!��F:JC������,̚~�s� �g��5�|�)"�T5��M�����:p=]8�k�'���X�i!i���|�Ӏ��láD$�Owu����5K�Uu�u'���<I3�����[_ _Z�	#�sm���[�����L����/�|�Ӏ�#��=UF�4ι�t�,�<���́�6��UT�Ϫ���7�憐܍�	�jb��a���7vـ5�l�H���5jJ���:#���ɥ�W)󜯹�(R�B�۶`������=�ۛ�6��f���\�t����,��GN�i{^�=x�B��� ����_$t�.z�p�Itf������z��%|�t�.z�p���\���4��`�ms���I+3�@����3vs�j�h�۸Z'�ci���$��=#�s�Ӏ>�� �W�{6ʓX-Z�bx�gs�Ӏ>�� �W�zGN��qkx�m�ŉ�$��K_ _Of�
N���oz���rN�znB{&��^�m�$�i� ����Ӏ����K_��K��lM���m��Ӏ����K_ _Z�m�����_����ϝ��ZW�"��ܛg��;d��5�4��z�S�K�����PM�p$t����/�|�t�3���(�i�N1�R�n��s��L�ou���5�l�=�&�,��!
�E��7����d��Us���vx��,�FmGQ��&
A�w�ВQ:�q�rn�����L(��2�N���n˖inkj&��)$�䎜���������ߝ�����8�M�7B��Y�����}+bL�\e9n2]{-���+��9��Uf ~�� ����gB�!�]�nV��j:JR�nI���/�ʮr&Mn��9o_�[���n�WV&�B�&�H��\�Ӏ>�� ���O�Gp��z�kbm���+� }-|d����7ok��⌊�c��,�ݖ�W9O۾����N��vnI��
����ª
��������"���
����tP�UEb�+��TW�ʠ���*����QZ ���UE�T�uPTW�UAQ_�UE�T�@TW�?���PVI��EdBk@�WV` �����Y���    @t          Ƞ   �$)B�	(*��E"�I@�!UT   �@(�P� (@�R�@I*��E()T%V   A�
 ( U� �`4@>� � 
DR� �f �ܚ��������Ϡ�^�q7Vܝ| '�#Gg'�{� 
��L���Y�f���ɥw} =)��ϧ�T����NZ�_  8} �!@  d���>�7|�ݷ�w���ӛy:u��Ϥ���R���:r�湝�Z��S�@  �    O��|�ɥw} =)��şZri����k� s�{�9V��z���_O�\ ��)I  	
͔ {ϭ\Ϲ��g,��+������ zS�>���}i�z�\��` 6�i��jq���W�ƞ��.@�%�}ΞN�\w:���e� 6q��Wϖ��t�qn�W���  (U �b ީ3���n}i��շ69\ u.��YO6���˽��ʖ}{��\����,� ξ����{�}��w�T �,}�^sy:��x۷��'��{� w����jru�9w�� x|�
 �E U
�h]�\��S���.MWO����p �k�� � �P �D ))   鈥( 
 :����@��iJ7@H�(A@�@ -`�( ����)T�4h*������*�hL�"x�T�P0C L&"{J�ePd21����j��@ 4 DH�z��R ԡ?��������\�j�ffS�o�nޯ�TW��AQ\@AS�� ���
 ���(��� QO��?�D D���J��HA�O�1�D�O�dJs�!��?w��=�<���2~��,zw�%�.{�g ���x��p����
8Ç|?~�g���?~���+����dX\8#��1�'?xs+/����|��ļ�g�����̹��ƽ`�!L��B7��L:'���b�'�߉�wń0���;S?s'	zQ Ї_wa�g��5�k݆���=u݃8K����S3��ý᝸ˇsxA�����N�s�	XZ�Ֆ�$�)�)��5H0 ��FD��N�q��j=d�\9�0��\�ƾ=%�^����y�^=�1��w��s����"��P�!�o�o}�fsуy����y�*�_ޞ~og�'xw��b�<jz! ��'��<aą!��{;�����D��Kx_��	�YL	L�B�y�p�?C��A�!
Bė��
�cǃ�p��Ì�s�����@��0!p�Ò��(8<� �zJp��H�i��	e��r7����rR�
��-1�T:��8'�x�>q�!!����Q���
�#Id���~Ht�!zt����fB�B�$H�Q����H\�� "4�2H��5�s$X�F���I$ A��@��)�,��#RS8�0������^8�d�ys'a�9��@%�=�_�CЁ}�y�~�ܧ�? x1h�J A�&rW?~�s�yK3�`B D�bbA�g0�^�rS�G�ǽ9�`B��� �����R���<���Xz�4���E*�õ�{�F�	N�珌b��<�08'(B�C�����d��O�=|O�)�F$h�aHZg����P�aRS��^ZR[gB'r�� �r�w=!BW�
aƤF��rw�|�%��{/��՗�b�01�0cX�"G�5���1	�h`�`P�>>.=Ǆ9̾���:����K�
��Ռ#L9�x�I�B��+�D
!�O$��B1�*ab��0*e��E�0X@
_�B����R�^��[��9����¨���;�cC��RK���I �XҠ�hţ�A(�W��cU��"�E�P`�D`!��0�F@H�"5 � ���XA	D���%B0��$��L���ȴ�`��e�>�w��ȴ��m�u�6{]��{;���^�S���7�%�zxy���y��<k盲�^���=	��%G����}���!�'����Zl�"R��(�g��8��m�@�R,#X�dD| ^�(0
� d��@�1"�$b�1)��-^�� F/  P"�%	���H1
@H%P��
�
b �"pR�hV)��#�+�D��	�cL+�1����<�cJ�:�1!<I%!����F	��ΐ�1�@k��P��>8ˇƜ�s�9� ��)�15Ξ0�ΐ��d�B���gl�H�?Q�+���&B�dJ���BHR��F����Ȳ>�ó%�aZ92Y���@�J2�8<�Γ��fs!�S��XaW3�'���ٜ?B~jB� Ӿt��!&A��G�������>��s�ɐ̖ \�S;�O!L�HRH�aX1�N$0�,*؟��9�S�zHq�w�)�¾�q`�0*�FD �(D�a��K�1�I��h���LX2{Br��0��6Lx�$��r' ������x�18��C ��Ñ$��[0�	r$ HQ�$�S���8�� 7���Ȝ���H������r2	 @��`s���L^y	"�������"���8%q�@���B�-��q9��IKA�#%L�a��,!$RD��dS�-L�D�J`�@:�*� 0
��=�pX1����Ct	L8��C�K�B	�<�vNaǳ1�\?��3�<c	8��ԎF��BH0`���D��!*A�� �D!��H�0� �IBDN+�� Z��H\�u��-yh@Ç:�%�2����F�&��H��4�9�<l��d,&8�����ޞ8������,q���N�a�T#P�)��H����0
�O;�~���ጐ�:���y�B�A�<JU��(Ā��K?R���^�p�V-���|0����%�$�Ʉ�\Hw�I�q��������y�2=p�@�(�(	�dEddx�F$����`$!$��"��@ �=�b�$`�B6^��:>!
�zF�@*�!�@	�		�Q���q8���FҬ${�pW�g			p䄄+��s�D�	-ib[ZF�B��	\y
�x�#Ȕ1�0���Q�H�4D��qAE�Q �peBX0XW��,#d0:�0`A���Ъ| ��,.	����HS����9�����r�JV!ÖhY_9�:{3���q$�/�så�睼:?�R)H����1��B�(a��)G�9û�?0��g��B�¸�`Ăx�k�F������
yUï>�(q�ZI,�`0�A$��O����}�/<��y�����a�/��{�B#X%�H)��D�p��q;�$=�!\��a�|�羜�	)����*�)	�vvw���!Nw�(S��T��'��Շ{�|��e�ÿ������+I�a%@�C9��{k*?0B��t�Po��kw�VF����ī�U3��0Ngd�*��s��u?��Hx��6ČX-�<I�O4���H���̦�"$$��'���Y��E�e+�1~B�����s���2Oml�I��ܚ!��|,��phBK���?s��c�C�#D��I.aB2������-9�)�2�;¬��.8�xִ�:#��Y ǏI�yC�r$$!��C������ș���'@�-�Oa�#XS�DHָ~쑒�<�Q�.4"Zq���}�@0xydK�ń��C��P�0卐�ı�a'�y�d��<��:�8x��!�Z�&a�X[�F���%�����:t��s(�I�cI����=	�}<"C��a ���r5Ì.rHQq�01��`<Z�	��c��rYԡ��:�0�`d!d�Α�f P"�	��:w9҇��aX%)�g3����êU��
Yp�Ҿ%0�S<�b�B
D��E�̰��V�F�D��K��� Ō	,�,�! �`��aզp�)�P��d�Y!da\B��*xN�H�$	�ôX��+Le9���q�L!bR�$Z�B��a� �J@�
@�B�%	Z�#�p�1���� " �(@�,�P�@�b-!W� ���Z�R-#µ\H�� �2F��\
F�V8�����"Dd	�a$�@�c$a��#
E+���'�#@��",`�'�%H�;��9�p � 8  vɺv�&�哮�Z��x�R�]�Å�ۦ��O��"�)D���֦ʃUz�� $�ͳIx�$�E���$-�����UU��UJ�*�����Q�ʪ���Be(l��2KJ�P�����S����#;��ժ�q�m���-�igR���q2ZEA���!s��6r��2U���e��ݖ��-9�j�sY��ҬUR9���2iV���U+UJ��v�V�j��Fh,u5M�*�0��UJ� �-6�����6���BA�Z�Skۢ�H5�m� l6۝t�� ��$�4��ݰ[@��}��     ��!�i6m�gF�      H@     kh  $  m�  �po  ꥎ6�{V�ݱ�`�c�zQ[��ڣe3�7�|Ҷ�/g/j�h��Ԡ 5J�agnv�֨gZ�J�(�j��mΠ <*��fa,� 4�-���Ϸ��8 h�V�qi�d�*�,`��]���m�n-�$$�% �UUF�uH�;�jWg;9&� H ��t�v]U[*�x�'`n�,H��z�km�m�j�&�V
%�ڐ�C����  si6v��U�@��&9�I/M�k3gk%`��;n�l��m'`�a��p�l� �     r��k0�kD�Pu�d`. X�,�pUUe�Wj�[@(�BsH�m��H�]��t�ݶ��W�n�j�8��zؘ�%�T$   6�lu�m�� H[�K�	6�#n�$N�sm"�*ܴ�|����i�N3f
�e�49���٪��X:s�.-�mp�kk�0��Y�m�����U�<�jN��[T�Hm�Hj��UW*��U� �s�Y�$kt��n ��9t��zlM�ݳ�im�f�� 8n� -�f��v�z���e�*L�Ҳۀ /�}l�.p[�i4�m�F�g�+���6�X%j�Uj��*�|���]�U�Vڨ�C�S�`��p6�$$ 8 i2�,]�  � �[�o2$6ؐ$/[a�u�VQ�����5@T"�l �{n�����$���Zݪ��tU<�ܭ�{$�� �ր8�[F�Am���E  H��j�`-�nI��\ ���5U*�Pq)-�n�*���llu������)� id���m�v�	 �om��$;E�U��6 =p���Q�{?� � �  �m�^����LpH�ք���q�׬��I��Z�2@  ���:�NH?6�|[dHm�l �6�I��Mn-�!CrBڐ ۗ�ӓ��>|m$�6� Z��}��nq5u�ɑX�媀�H �,���� ��n�4��۶�m��� ����U)8̪�� 5U˹�R��R���U\���J��R�m]*�vF��jyn�W#�� ��Z.�-m�UC��l�f��enH�e����H�� �m2� �  6�mͫI���vF�mm��j��S���   6���� ��Hք�K��E������UU&�:��aͯ^��9z�v֭� � *��lqg�G�M� � ]j$�V�F����+<ֺ���m� �knhڕ怪�۶����UnHHp-��   ��  б%����8� �,�l���Ѯ���m�mme6[xm�@p8��:@j�� 	קY R�n���`  �6ض� [Cm&[Cm� 6�Jm��6�@�@�mvHҖLm��ۤ��p����-��I&�d��@m�� �1����"F���6Zm�[��[i%I�� Xe���K�  �M�iD���m��h�m,�Y���%�� � �� H�           m�H m�          Ā�  �  �M� n��-�p�<��5P
�R�!6�q*�PuF��,Ԯ̒��E�l��6ݛv�А�@��Ͷ.�6�   mUr��U@t����(G7m� H6��ԝl�YA  $-�pH;E�2�*@km�cm��`$ 6�  � $� � ���f���z�ֱl�Hh-�  |}����`CkA5Rdm�*�E/1��N����  ��`9�k�� �m����m8�v�xV���ʪ����V�T m�$��4ۘ Hڶ"�*=�� ݶ6�  6Ͱ	����[pH     $       ���	I��������$om� j��u���@ ��Kkm�}��}�p��&p[�崺m��t-�[x R�P`��UP*�V �|   h  6�-�  �`     $  l� l m��� m&   �� [@ �cm���xpګi9�6��m��y�Fݨ��G-ԫV�Cm�8հI ֲ޲��Q�-���m�M��� m�@ l�-� � ��  �  	8� ��8$����^�p'mU�E$�c,���$%�mc	�E #U` [zImm �Z�@�����H[@B�q��kn�����-� ֲmrj]��-��v����v.�� �֖P��i0�  H�m�  [� �mrCm�m�8 [v�q��&���������X *�N'v^B6��l��66���*6
���е<�R���Jy��sh1r�pϳ�l�qs�J�<�YI�r�˙����<�Ut[tM��$h��7-�^l6� $�[p���h[@  ��WYo��m� �  �vĀ 6� ��m�l8  Ѷk�8H H6�k̀ �  m� Ӏ�m��$8��X�e�[p�lDзUW!s)<�����&��L�K.���`H����[E�@ $L�\	.�v������n�Iͥ\m� ��mZKn 7n��T�˱�HNQy��#e���N�9�� Z��nu�[��!�m� ��[C��!�  *�@A8j{\t5UUz�$���6��/G9�C�8k�:�"��Gr�mU@�UU �U�Cm�7]�8m�]l��-Uq�*t�uUY!Yv�� PUV)��cm��h8q �m���K,�H�N��[�m[�o����[E�*۶����j� �cax�n��   �H�H X�f�J�(li5;I���� ۵��-��4�m��   v�  ��}I�i�����h0�	�  �$    � m���   �8H   k5[Kn��a�ݶ�f�� �5�V���� �I4Y,s�mvΆ��U@UNUUZ��ԟg�>��*�ȡű�����    �f�     ʪ��BEW&K���0J�ր,hy��T��C�ڪU�pb;��M:J�gn��մ�8�lgf��j�j6�9�k�)�a�kpsN�ZT��`��eP;c�[T�e����6B@^mK�e
 �cm���_Y)!���E��WT���;kcm*��)m �-Inm�sm�l�l�Z�E�����&R�J� du�v@�ڪ�]ŵa�l�F�;���Y��c*�[Lb������%jBK@��-�@86�nv�*ځ+Uj��C�N#��]�j�F-"i�J��v��*ؓ�����@   m& �� � �T��s��@<�UJ�Pm ��n� $m�m$ٷZ۶e� <�I[L���HI�ـ Bõ�_Z 8Ĳ�=i��iUV�Cm�$  -sI�  ��6m��8 �l �e8�%�f��Cc�ey��Z>��� �䶍�� �@�I�D�m�	�V� �����}>�Yuڱpd)��ؖ�eR�v����6�[]�6����d^�&3v�k6�a� ����m� �`Zkk��m����m����
�iT�
���[l�]6 m�������  [%   h�hm�l�$  m���  �=;l� [�7k�� �Uu2��P]G��\K(Xe�[G� u��ܑ:�� ��V��@Y�Fej�rҜݳ�m�m�X�l R�PJ��\Tu�W��� ���m��6�j�C6��u� �       �6� ��5�M��$U��Ͱ�-UX冧�dJ�R��,*�y( m��]�`U�[<�u/@p*ʻ-A@    6�UV���Un6����%���9��(���(B � ��?���"�:���1�D>���$T_h���P� � ��@�zN�� E�C�^ {���EN��:cE�4T�#�� 0<����EC�}���~P��A]C�<W�瑱�@��07�~hb�������Ѣ)��A"��E�	 �5����ç�W�D�2EWC�
�"���}`
AC�b�t� ��<��A�X�q0:���S�(�z�@�Â�#�4h
uq�*�]^��x����A�OS�D4U�PȺ����Q%�"g�p#�B$EWPQ|��D�� �EqPb���<OTG��ŀ�WC�=�ׁ'@���O? (��@�*Ԩ	�W���({T=UJ�(h�*�o�?��QE ����"�E����S�ű؅��MLv3�;X��K���
�I]�+�+F1�55\B�N�<�m��Rw[����W7:ZT<-T$��i��@�6�v sCT�^˄M�)�J[���D��ہ�$f�c��:��
]ڂ���u�©���U�Pn��\f�Cg�S<�m���3��gmnѱ�h���Z��(���mt��HO4uET�@J����A�K�z�ny��Ҩ����[�!7K����-i#�.������s�`���h)=�3�R��c�݆��Uj�"
N��N�6��@Ʀ�!���V��݄��aݷn�L�@tlkPlmV����鶼u7Vz�	�m��3�v!C�EYhTT<���W����^�����m��IJ����8�bW3�n���ۑ��Z�;*��C�!�UTM�H /]���M�F�5�I"-��t��2\��;�$�Ϋa�.�Tm��v�1���.R�����;C�l=�ļ��Kt�ݜ5@UWWK�6Gj�냭�h8�$�fع2ʴ��+UJ���+T��+*���HN��^�r0��6�t[�H2�s(q�@�ҡY�;q��r�n�M�.��K�Evn�B'"�����mڅl4ZdD����Ł�s���[WI�K-*�H��s��L��'�b����+ �#���A<��ͺɤ0#�,�֪W-��#=������U�T�����oMڠ7,��uM�P�k���P��` Fnim��#c��Y��ە�0�CJ����UT�9=�1AU�����1���F�+мWT���G[�P�b���6���K��|Ō�9��6�ȕS�ؕz4��IZ�U�:l�����gfRB	^��������dn�l���Zd�[ l�0ɩ/%����Z&��FF�z���av�r��lG;�̼��K��di�0�&�ܞ�u�v@&E�g=��
���k3 W�@8��
T@�U��0�"��G�E�S��@ g�o�9gl���<���6;.�*�᮸ia{N�S���-�Y[�h�ȶup��#4l�rD�;��U���ڄ��S�5��.[(�Iwa��H[[�v+S�;CWOlC��+�m��L��y��wC�M�+lm����-;#m�;�g"�NP�#˓��Ϸd��Kʜ���RG[�n���5�f4�'�*�.�l:;u���:�^�<ɖfL�2\�Y��r<�l�Þ�;pg(g��a�e��ñ������z��I`�6�С��۷ ��y���	�L�bX�o�y��%�bX���.d���[-����;ı,M�ws��>S��'"X�}�y��Kı>߾��Kı7w:D�Kı/��{�̗r�3�/9�O"X�%�f��ؖ%�bo��u<�bX�&��H��bX�&绹��%��ow�7�w���9��W���7���w|�yı,M�Α;ı,M�ws��Kı,��q;ı,M�{gp��y���s���yı,M۽*v%�bX����SȖ%�bY���v%�bX���O"X�{���;����e��sM��ڋ�V��n:�I�����ųڠs��f���¶�7/9��\��,K���w:�D�,K����,K��w|�yı,M�Α;ı,O}�/w�^s�s3s&g9�O"X�%�f���j�dA��
G*TJ"M_C�"~�b~�߼:�D�,K����,K���w:�D�.�����b�9a�w��oq���w|:�D�,Kv�J��bX�&绹��%�bX�n�8��bX�'�7r�幒���/9:�D�,Kv�J���ș���w���%�bX�}���v%�bX����:�D�,K�m˙$��[-���g
��bX�'��vu<�bX�%���'bX�%���{���Kı7n��ؖ%����.�&�R$�88�F��l�M��Y�����I�;�Z�3e�Yk�(.kw!L�[�^��,Kĳwy��Kı?{�vu<�bX�&�ޕ;ı,O=���yı,Or�s!sm�,�s�9�s�ؖ%�b~����yı,M۽*v%�bX�{����%�bX�n�8��bX�&�=��ng�Kl�99���yı,M۽*v%�bX�{����%�T�c ��AA�EQ$@X�A �# ��Ñ9���ؖ%�b~����7���{����ߝ�a[k�5E7;ı,O=���yı,K7w�Nı,K���gSȖ%�bn��^�{��7�����鏿$��^�x�%�bX�n�8��bX�'�}�Χ�,K�ݻҧbX�%��ݽO"X�%�� ?o�[��&L���9�������ێ���V	ƭ�3.½W0�`��\��Z� Sv-q�X������{��7����:�D�,Kv�J��bX�'��vu<�bX�%���'bX�%��Mܹ�nd�!y�K�N��,K�ݻҧa�G"dK���SȖ%�bY��s�ؖ%�b~����yı,Oٷ.d��-	L��fp�ؖ%�by�7oSȖ%�bY���v%�(C"dO��ݝO"X�%��w�Nı,K�n\�3y
g2�r�<�bX�%���'bX�%���{���Kı7n��ؖ%����D?'E
�� �+�|"���L���{��oq����������'�f�UIؖ%�b~����yı,M۽*v%�bX�{����%�bX�n�9��{��7��������b�/'Dz���J]4�Õ׍Я0Ϋj�Mi6|�J�3��ww�ۗ���)m��'9��'�%�bn��S�,K���nާ�,Kĳwy��Y�L�bX������%�w�������#�B���w��ou�by�7oSȖ%�bY���v%�bX����:�D�,Kv�J��b�ow����߄�T/S������7�ı,��q;ı,O��ݝO"X�%��w�Nı,K�y�z�D��7{������FQ��}���爫C�=����yı,O��ҧbX�%��ݽO"X�%�f��ؖ%�by�w.�&f[�%�/9:�D�,Kv�J��bX�1������ı,K>��q;ı,O��ݝO"X�%��'�Bt�2;�o%�e�s���f"n�i����4���1��U�r5۱��q�\.���9��-�0���Dչ��k�<v�aĭ��}A��Bcc���Ɩ6�{�'i%�۵��i2��kk���-K�n;lB9+��V7��w;���u�[t��s�m�*/(�Y�8�dЗ����.ջl���M�bm�����R6�}���}]��`���w�?H�6y�\��m���m�M)=q�ќ�l��s1�#��ϖ��͡l6�%���g
�ı,K~��z�D�,K����,K���������"X�&�s�Nı,K�n\�3yÙ���O"X�%�f���r&D�=��ө�Kı>����,K���nާ�,K��)�B�Z�TIWwE�������$/n�gSȖ%�bn�t�ؖ%�by�7oSȖ%�b]����Kı.�=��y�fB��9s����%�bX���"v%�bX�{����%�bX�����,KP�������K��{�?7�|0�g��7ow��o%��ݽO"X�%��.�1;ı,O߽�Χ�,K�����,K��O��>2d�r�sg8fa'dT�Yӎ����R5���l6�.�`L�j�0�R�+
�=����oq�߮?g��Kı?{�vu<�bX�&��H��bX�'��v�<�bX��m���L8󙗙rg9�Nı,K���gS�e��p�������G��blK���S�,K��߻���Kı7%��'b`"S"X�dݙ��3-��/9:�D�,Kv�J��bX�'��vu<�bX�&仼��Kı?{�vu<�bX�'�sST*�tL�wuV��������ou�ݶ`[ŀ9sJj�ЬUJ��p&�xRQ�����빠y�S@���I��La��z�o-�z�i�Lk�7bNu۪�[���u�SJb���H�$�=��/[��y�S@��f�^9,sf%�H8����:"!B�<���:G�x�m��'SN!�m(�L�<l�w���E�����Wࠈ{�O����-�)cmE#M��ov��&�<����� 9Ԕ�$O�6�LrM�zS@�n��w4
��h~�u6�8�e����z����m��e�졷^X��\��t�o�����3`�!6(Pb����s@�޻�G[4=�M�UM�����V]�U����ϢL�#����x��(IL�.����.�X����Y�}d��@{�����@;c�1W1��$�RM����^{�M��;$���Ӳ �``�'�T���-�x�,�L1,RA����J#����H�� ��`>6��ۦ���s]��ϜcX�ݴ�)�F]�<�T�Jd�:9XV���n*���H	c�P�@G"���ٵ%]]Uu5%U��[��	TD(���gƁ���h{Қ�RQRA��#7s,��@{����� %�I�r-�M�JNf�z���m� rkw�)B�?����B�s��	#s4;�4
��hwJh[ŀTjB(Qs0�f.�U3}ѹ�=F��\�v[����1ن�*k�����WƘ�tȽ+kJ���HlFe:�u�ܓ�n��R9۩�l=ynn?���kc�M$mCw"��x�t���k��lʖ���m�Fq�(G������J2��.�ŝNĻ9�)mm��Հ��ƴs`�ؼVɗ��ף�s���{m��[]x�h�n-���$~���g�{�폾��Z�
t��X�v�n��Oa
n1F�,��:�k��Ƥ���<�2yre�w��<��/[��y�)�r�1:F��
I�y�`��EH7 %�MW_�Uv���9����p�/[��y�w4�Q
�H�� �w� �꺧5UaU5&��������ɨs� #�s@����EDmF�rf�Q���J=�8�>�X�m� �1�NmM��25�Es��`eV�e��z�s砚�������l+�S��@�DX�#���?Ͷ`[ŀ~��9~��u�NꞵSRM�L�Dݘ��e�Т���N��<E�4=�M�Z6bVcX+��ݼ�@{��,rj������T�7�fC#��p�*:٠{�����@;c�+2^�PIwwtM������$�.}ߗ�=�|hl�>�����В���G�F:-��ы�큪րZ��J�i���>gC��a��9���BG �����)�Tu�@�ޔ�.wdn��iG/wv��@K���=�9 -�)cQFL���M�@��f��͝�y��|P�4!0),���0,Z�)s��q��GTtg;��0JV�`�����g�'?u���ԑ� �/�9a	�HFD#���d ����q$"���W�L^�a�̏�� HB u� F �R8�t�8�	 D�H$B$�((qZ��*
*P��� ��D��
���>H�@B
�������,�{��v_�Q|E�c�h}�{�~4��nh{ҚG[4E�X�ئ
j�욼?ϻtBS$�^q������u��|t(���$��Ϩ�-]\������۱ϣ�c���[t�f.ɞ5�\�����/�.1]���������������J!.��_�=�����)B��~�Ł�(�Jg���5%P}b�U+��� �u��	}
%Tk����D%?w�b�=�>>����x��V�o��DrD)&�Q�y��(P��~_����P���u�i�J��UTI%��DN]��}ذ��f ���W�B�Ģ����T/���'d���?�n�Mɚ�����Vuz�����������F��#&8)��k�vFFӹ\C��v�me۫��v��;�Y��F�16F�n#޳@�ޔ�/[��y�Jh�IEq��c#J4�7P�@G"����&���cb�!�18h���<��4
��h{Қ���f5�L�5�Hs� %�M@{����ʪi�ya���i�hl�<��4���?{m����#e�]\�T.&��id�+�;���K��r[%�2m\��%�2F�Ug���:[8�q�`8�[�և.��ONK�ҦM����W��|�$:�:ڀ�ɼE����j��e��17�ҽ�㸬f�CnN��S�c#[�9y��D+�����=I�"��a�m�����wX6����jR ��%������d*B9�-��n���n��\��瓱�t���:4u��WG�p����y��K�ܱ/lm�ݲ�w�}7����@K�@/�B�\�؄BG�������=�`��η2^f�e��Ԓ)3@�ޔ�*:٠y�Jh���-�G`�1FF�nGY�s� #�R��p�ܙ{�1��c�h{Қ�w4=�M���[mIq8�F�I�n���ۆ���2�����@ψ�6ϟ&?w�m�}�Ĕ�E�����}~�s@�ޔ�*:�����zύ���6#�2<��3@��b�J��u�����`ʊǉ�co$M�@��f���$���y�b�=���6tڡU5�DrD)&��)�^�s@�ޔ�*:٠ҡ`���E!�����@K���=������q@�ݬ��h�v�1��g`��;&�Z;��+�u���m�OK\�Y�k�s����95�{r*@H��EB����4
��h{Қ�w4=�MޢQ�D����wx�m� z�,=	(Ȉ�
@
	��U�vs��gd���w��جblS��Ln�w4=�M�������⪦�d�L�7uUk ��`
!GP����|h���>����E�D� ��b�읱�f�][a�5ɴ��\x�\��k��^�����#�O$M��>E��y�Jh���<��4\scq��$�NM���T��=�X��8�,.1���#p�/[��y�Jhl�<��4�أ��1�7rI�Hs� %�M@{��~UˑR�Dv%q
4�M�hl�<��4��h{Қ��2����.�F۷�� �8"q�kL��W���5��j��	�I"���'b�@�ޔ�/[��y�Jhl�;-��&�1,on������@K���=��⪦�Y���#nf��)�Tu�@�ޔ�/[��*+d_�7w/4@K���=�9 ���ߍ�V�O�($�I"�@�S@z�,�� rkw�S�Q�N��۠�-ǃk�ݬ������D��G%�Y���6�����(]uT�9��ɜ4vml��ڳ�[p�J`noe�hp=�Tͳ���`(�-���D�-�-��v�2�=�4���>�N�-c�X�3t�m�b��u���evzWy�*<4Cq��C��{s�,�z�3	���+��wA��rY�K[��[m�T��saK 3�����Af��77h�۟)�.��
�Ʒnj�Q=��>�&�-�юG�!G��}�}��y�)�TwY����>4����SmƤ���x��,nj���T��ٹ��j6&�TwY�y�)�_m��<��;�J;��d�crh}W�/��� <��,nj�MV1���cq&7�n��t��Q����M���a"���I��]v�N����ZBu�[d�9&;n�Y���� ���b�E&	�R6�hwJh�hwJh�w4�EuLq�~o$�>N�6�}�w� ���������?{| 8��{�<®m�]��"�@�ޔ�/��i���>4�o�@/�B��q�B7�n���l����9D%	)��� �jm�ۊbI�)&5&hwJh�hwJh�w4�>��1<�F��It=��y���=@qY��ÓY[��tsd�j���
DLM�$p�>���<�gƁ}�s@�ޔ�=�%�M̍9H���?{m��2v�b�=������{*��4�LX�M��n���	�j*B��\ɺ� ��ـzZ��Y$sLR6�hwJh�hwJh�w4�Eud� ~�����<��:EH7�@N��W�A\Ok��l�u����<�cr��d��ו
M˺��N�SK���lb�׻�7�@N�R������X�*1���#p�/��hwJh�hwJh��m�0I���W7k ��l�����|��v�nh�#��$�rH8�TwY�~ݶ`����G%
!Fo������!G��ML�9HnM��M���}�����Gu����[P�m#���;���gp-';�0k��m��b�7c���[PC��3T[�DBƢm�z�����?{m��u��Q�K���0'���Iě��Nf��)�߿�1��}����0��gB�]'WM�7a���j��o� ��a�B�*���b�:�?��ي�#BX��
I��D�^q�v�b�?{m��z�������c�HF�_m��>���xH�^��l�)Rqp����&�L����}d`8ɀu��:��(p�P"<ޞ��CC�D�e� ���c�#�Y�B@��F1q��{�M	�� �b\	<�Q�SOxe���� 2�B$Q�݁9ӳ�J����!=� �@�$O�DsЄ��đ�d"Iu��q[S�FE����DT��`FBI$$$V`HDBH�dH�I0$!@�!$$#!d$$�	��0�I		YI!#� j��*ES�C�(���p!\J`��bDq��aB+BSS#q�a\�o1@a{�9'9�IK-��Sl��q���I\U���n��g�8ݝ���Kv'�nQM��u�����ݮ k��tOn��붰��ި� $���pmT���ym�G\��}�eJl�n(40&��Ȫٚ�*��R�Ø��i�gZ�m���5`4���b۩m��
�m��&)U8m��v��GT1�i�PGC���ƻ)i������E�؜Gi;v�F���6�*���ui��˂U�%���D�f�;6����W9r�]J���‎ڠ��LvX�\5��na1�MM��"Yn�j�S)��]$Y<�Le���&��m����!%�y�(�ot�^Ŝ6��D�s�+��y2��v;m���_}�|ь皫j��n��T7#�ʦ�lF�.d�yvf� ���Nq��Wq��]��ږ��I7Z�ջ4k%�� ]�@ �5ں!�v�s<���+gWuG �����N�msP7J��S:��0��6,�XD�-�ٍ���q��݁e�l�4��M���k���e�iZ��*�WXظV����e��W��iK���W�Z�;uD��!�{���Ե*�U�)/2�s��3�M4v╃���#9Uu�h)`r��AX���D��x�/<�;�� ��ъجb�۔��N�&E���?%Y5�]�΃n]�F�nQ�{M���9��n�A�,c\��luW�f,�u��v��;s���+��� 6��ۨ�l�Pm�Rq!�X(;n�QIyG��A�UUU�/��f9�fT[��}+���uUJ��i�n-�-	�-W�,凳�V>���;t ��cq����n��)�����9M��c��֊�F1*�s��5)�������ȅnҪ���UԷ	Uیm@WZ1�����j0��j8 mJd��Sg+m�1uAvn�Y��Ai{g vʆq�wX���F5�nʲe��`G%�:�m@�*�DY�5��y�������"�Σ���_TD�'�@����%˚�v6-�lhMk��[�$nV�%������������k��5�,e�9nmmnDZJ�ѝ�ʬ��15M+��C]���^��
2�#�R�V�r�Q�ū����Z�������rkĘ��p��1Q:yeK]�VlP�v��k���v�ދtL���k[gZ�ϡ��y�8�7/nα;J��	�m�U;��{�ӟ=u/w��6���]��ts�g]>�6�z��h��-�D��8�<�S'��|��)�&�RH���>����*;��<��>����ۚ�� �Q$���I3@rn���"��*�}��`��M�1#����Ě��q6!�4zό��XtL�]�t��������"Hj&ۆ�߱}�}�h��s@��C�^�ߍ���i/�����#nb���U�}��߄� =�o���I����7N�压�'#h�v�΅.M4�CH�<92$�����}��Г׃ov��I��=�`��"����ʐR��}0�	brF)&��)�?L��Ծ#�� �$`�$�XE�XH��B!(K�D%�����`�b�������Ӥ�T��R$��.����R�����s� %s�̗�I�&���I�����*;��<��0:(���� {��M����U�YwwH	csP�@N�R�������V�Rc58:��w&��g�;�=����y�y�����6&`K�q#�� ��`���?{^.P�/�#}z\�E�`�$5m�@�۹�y�)�TwY�y�)�f~ĎG����U*��7uUk ��� rn��SID�Q�f���� �Q]#$��)���s� 'H�U��h���N�hK�1I4=|@;�����s@��@=�΢Hcs�8�ʓ��,v�t��m��	i��I#;t7%�5�6�7�<K"���@�۹�y�Jh�h{Қ�{#u6BbȤy{���=�X�����T��r�L�@I6���Q�f��)�_m��<��4z���� ��Uw��"}�8�;{�`������!AR��L<�)���fniԓH�+/o33D� =�`��75��Mޱ\�%YQ9�����c�cYA�շ*RZ�WgC�nz��)�w�ŗ�=&1�ۙ����Q�f��t��}�s@.TVU19���$���*;���2{]�v�b�?n�X�;5L#BXܒ
I�y�)�_m��<Gu�}9�C%����@�"������<��+�nd��LCY��3@��h�hwsgd��w�d�E*�� @RPb���f��9:ų�BYۤ������ѵ�=4^!���΂غ���7^_D-]��~�՛�˘ܸ+��@7�pi.��rⳎ�w��
jU�6���FY��s�f�1k��-'b R��<91kC�T�xݮx�|��$Zݮa����.����Er�����s�V�G�ms67HۓG�\���j�;9�hx�����d�ў���;��+*}��Zꇛ^գ��z���5��hg�e��v� �V�<D�SgK!$�rc�g�|���@�S@�۹��3?�Xw�nh��Q�8� D�cr`�m��(��;{�`o�`M�y�$}~��Оj&ۆ��}���u���E�M�gƁ�-��1�jh������|�~XH�^�vف�"{{�, ��u6�옕Wv]Z���>�ǀ�����H	Ņ����u�>���6�o#nD��F��9�ɩ�H4��u��nDO��#�=�!�$��=�8��ŀ~��\�Ht���i�J��ŉD�p�/��l�ϲC޿nh��� ��g�}T|�W5�Ҫ��.˹���k�`M�xtL�]�v�fh�X�H��5�#��TwY�~��0��`}�kＰ��}E�݆�m�fn�=�`�������s�*@TwY�^eV4(��≵Jd�aûY.qq��호)�=���m�ۓ���!�d��0Ƣm�x��ۚ����*;��<��4Qh�&G�&)s4=׋>S'H�^�w� ��, i��x�9���$q��*;��<��s��^�s@�۹����yr4%��!����{� <���W�}��*$}ŉEI�h�w4;�4
��4;�4�+�'i)���[u���ǵ����T���1#�����y��j 2L��&hwJh��<��:EH�7!F������f�	csPo`��"���߿bG_�G�L��nM�g�t��o`��75.��SH�*����0:!%���`n�����5B��J?+���`'�T�ڴ�1�ۙ�yϪ�*;��<���ŀr�^M[멡M\�U�WsVU��gd1�l�rk��5˗i����ּ���5�5��^���I �^�-�hwJh�w49�Z܎�B4%�� ���	�*@y㖀�s���˰���S']J�3dݕUf���vهD,������=�|hӰ����b$Qn������sPo`���{�:9	��I17�޳@�ـ?kŀ~ݶ`	D,�B(�K:{�c2�p�X �K!��D��_��tlά���Y�oC���ڭ��ַ\M�#4l�3Ӻ����L角b����urC����nt���6��׬{lF�f
��[Z��L�۝��u�ztv�b[���l��e���<�
���1dr]��l�m��d�\�v3�g�w	�2]Y ]9��4�)�⁁�.e��1y�^c��2Fy�˷��m˔�f�3��̻
��L�3��LOe�xB@i��Crhw��@��ŀ~ݶ(�!�k��9�3s\U%�T��UY�?kŝ'��XI�� �S@���Ʉx�b��3@�����xrQ>n��;_b���U"]���˻X
E	GQ��$�۽�tA�666?{�xtA�66"6?�~���llln�f�3�9�K33���s�|�������: ��߼: �ۿxtA�666?d�~�D �`�`�`����v_��[ɜ��X�����i#�D�8-�n�i�yd�܊]W����b�c�Rq�*���������� �`�`���xtA�666?�~���lll~���΢>A�����~�|������'s�d�$��9y9�: �ۿxtA�#�h�S�A�ly�|��|�������tA�666?{�xtA� �66;��s�3��N�/9��rtA�666?d�~�D �`�`�`��w�N�>A�� �A ���xtA�666>���D �`�`�`��~��>�rs�e��̳3���llln���� � � � ������ � � � ���Ӣ�A�A��A�=߳��A�A�A�A�~����0�8C/.fg'D �`�`�`�����D �`�`�`��w�N�>A�����~Έ>A�����~�|���������?�6�g�Qru�����ְ����2����,g�x�������?n�ے�s�D �`�`�`��w�N�>A�����~Έ>A�����~� ?���9���â�A�A�A�A�����a.H�9ə��� � � � ������ � � � ���Ӣ�A�A�A�A�߾���llln����
Dr9��}�_�9�Zfg9��3��A�A�A�A���: �����>A��zH {I^!�Ed	HHN�)
xb@>1�6���E%0�`PL<���&ϼM�@�F�ABb$Y1ba��@#�B�@�#R!����H	�8Z 2
��2 ����1��a����|�H�L@�B z8 �. :�`��B��<@}@�+�@�1C������A�pD��#��Pxx����lwy�ވ>A���s߾Έ>A������)�d��e��9y����llQl~��: �����A�666?f���� � � � ���Ӣ�A�A�A�A�٤�}�fK�NNs���D �`�`�`��w�N�>A���G���: �۽�tA�666?{��|������]3�!p��2�Z����O!��+hu�+�mr�b�U�lj�ծ�����t��Fo�������X � � ���gD �`�`�`��w�N�>A����~�à�C�r66>�wՑ�w�M�ԋ-Z��������o�t���� %�1}v}>.��ѡ�a�D�p�>���<]�����[��=�|h�֛��LR6�h�� %�1���\�=H�,��'C1cr
G�U�^��t��}�s@�wW�}����1G�ǀ��뭼����ɍ6���3�v�9{[�]h�M��Z��!�$r?@ﾟƁ}�s@�wW�U�^�_NB�ZQ�$'"q�:EH[sۘ��{�إB�)�⃓4uz]��wJh�w4���B`��LQ� ����O��o�t���� 9�Qׄ&Li��MǠy�)�}�}�~��V �u��B���!@�G��T��h�)G>.�e �ֈ�h���'�N�-��lܭv����f�^�v�8{3��fem��O����ʟm'g[t\l{���*m�89���Bcnů�Lm*���)s���H	���g;=I�c����ގЎJ��Q�c�����ܩЕÝmq+��1q������$�Хrm�'h:p�u���	Q�m�A�z�y��b������=}����3�uW�ȭ��y����0m=�mו���v��g]j2NH)�������ۚ������;�4QkM��Q�I�F������� <��:EK�]���>MbO�̘܂��+~z�Қ�����^�w#��ZQ�CnH���� 'H��nb���@2���i		Ȝp�/��h.��
���<��;׊�7r
c��ƺ9񳮟l�Ob4B����]�9gD���(�3�	8�S�&h.��
���<��/��h�5h,���b���&�}���J��� ���'�}?�������^��P���ɍ5e�n <��:EH[sۘ��D�q�<S5m�C�^��uz/y@�yݴ�9����	��y�H[sۘ��{� �������R7j�,d�j�ݼ�ɣ��9�=)Z�l�$����.ӫ�]m��c��z7q�W{��>�>��� 'H��nb �G?δ�i�$�@�S@����<]��{����^bBCr7uf ���w]a)EA�BQ�BM{���=���@�����)�"q黴���1/���� '8���V�!0R9&8��*���>��������x���&z�wU1��7
KuW͡�k�q��X{=6�Yu�70��K�O��
8��ɍ�i���zS@����<]��{�����1'�bƶ�34@NqR����@}n}�7�@z�Zlvb���r4�h.��
���;�4�]� �QSyY��.�j��
_W����7��0�x�3��0�[�@/"�δ�A�8�R=��|�ޯ�'؀��bLww��nk-�̵�ln΍r���Io$��%�I9��:R\�����|�l���9����	|�~�zä߄̩)�J,SDㄓ4u{��#����<��?kŜ���T�"l�-W{�W������o`��������GXE2cmD�n=���Ɓ��b�?N��=M�`����	�Suu�����t���� %�1�����#vI(nES7qeœkN�u�ٚ1�gVrQ���ιQK�O(mͺ��n��"��n��	p�nH�8]����;Z��i�*����yo)�h��mJ��9��u���8��3��F�46�z�]�&���{RNd�b�ql^��
��c<w���m�8��v�MnL2�n�ד�oT�*�&n-���!�����L�/w{������DCIum��pkf�WE�HE�N�M�����y�����ܹ�s����Z�ͨ����@Knb���T�r9���MvM]`w]g�K�F�_����X��u�	D�7#�����bN8ԏ@���_z�h.��
�W�=�"�q��C�����w~X����n�>K�����$��J(47��x���*�^��t��o]���`�PNLUp��=�g[E�^���m1ɰ��oS�\s̓؉��w����73s3��~�����?{m��x�!(_�=:���$�uͫU57USWu�~��0^�JI�(���o^,��]`|�g$��τ�[0C�1cQ4�4��s@�{����˾��������f(�nEUk�ID���`/����f(����f�}�&���39"R=���(^ל~�v,��]`�˪��Xud�W�m���;p�d髫&Mx�����[�;i����}��N$��P3���ٿ�T��󘀖���f�pQ�$9#��@�n����#���|��=�zS~��R�O���M�Ԓ+��zu�`u���+��!B�.u�xhw�nh��:�q�Ҏ8�8�>S��� ��� z�,�DB�Vߞ�o�Q��"�1��m9��)�|�7ߗ�=:��>n���T���"
��wk'J[���9^!
z9+�j�ɷ�<��"��������m�m�߾�T��󘀗�b��Y!����x	7"Rf�篪��?��6+����O�@��s@.r+O�,ō�G ����vه(S<�b�=-�`�����A�H�N=�3��Ɓ��t��ﻝ�4��(r���s�F���H'�]����ft�������@��S@�mO`�I�ΨStmm� `nt��v9w^2��hp�5��-<�m@`�1Af�VJ������~? �����g$��o�`�������q�1��W���3�bG[>4��X���>P�)��I7\�ɵj��j�n���Ň�!Dϥ�Vӿ|�xJ��ca1cQ4�4?�}o�f�}Հ9�u��S����UQO�7�I�&h.��{k�=��}�zvI�`�p��)$j2#)]�⌊�b�J8:�
�J��H ��9Y�2����!�7�FN����xx�~$���D!"Ba_'/@O�#���BX@�F��ĐRm�O�X,h%�y���d��T�$�H1^~���JV�J��b�,)Da"�JD�� �H��R�0�B��1���aD�H0X<z"R�-#8�(��{��յS�T�!w:����cڡгl�nh�U�ffGt�d�$,7@�mԮȩ�8���ѭ�u�@f�y[���9[�mUJ�֧��� �Hm��f˞��tem���t�v^�W�5X���]��p�����çktj�ψ<�,�De9e��݃6�\q�N��*0p��X6Z��.<��|ln&sɍͱ���p��bݜ5a�d��k�����(��\d3�X��!�LHŠ�]��<��V�(�le�+j�ݳ�s)���6�+�l-=�����l������j�4�+ldi؎��(�blYVbu<lN�tH�LF�Us�BA�3n�J�]�J:�ݩ		�ܽ/K�t�R�3ʻ�>�Q<sխbZڬ��k��"�,���a#�2Rb��'Hz��[nY풠W9Hb�(�ve�@��l�� !����
%����/`Ir�ۜù.�\��Q%ju[���s��,[W��[��f����np9�8���lr����[l��Ks����rd�v���<�$�M�m{KhݢRY����l�U+r���)+*ʪ��T���(\X��ml[R��ezIbۤ�L�v�ljn�;������5UU)-�P�cҫ�u#B�#��i�K� ��xrix�:��'D�ˁ�#��G'k��Tñ�]���rg��ht\����UN�Nq�cp�*[8�
��Dvg�����/<�n+u��]G$�Y\����8�N-��U;*gFn��*�
�vZ���c�YQ��,j^�8��&��r���u�ƍHs�V{m%�$�<<d�6[�d-��=���C�(璡��m��ڮ7D�x�UA�*��۬N��Ґm8�I��[�S�6u�--^�ErGY�-�Z֔�B�bT4J֥l�죔#�]u���n6`N.u�V^��uٗi2����ɜ�D�E���n�s��f]ĸ�@�qI�����{�w{�G(����@W�:x���:/�%�>*���3p��#̥98K�vM��^a�X�#r�N�Ȑ�^���2���.:�� ��:��.��.G:�RsS^,�t�'7t�;C���\�����4���U�6�!����^ܞ1�T�Ʀ�,�[�N֓���vy$�5�4�n��d�#��\ Z����؞MC�[tq�����/��q����Q�8٘j�Uن���aا��랱����s}���s�=K϶�gd����<k�8]��oc�nε�x�����G��;����{� �� z�.��!�]Ӏ���)�4�$�@��S@�n��;V�WZ��߿$}~#gё�$�7os7D�� <�K@Krb�� =�Ȏ��1��m������|���X�m�������u���U�q�0N-����Jh���<�np���|EUқ*n��]�A�Qͮ\V:Y�Va�in�&���gj�?������L�Q����/�O�@�n��;V�WZ�xJ����ōD�p�/��;�C�@��AC�Ǚ7���{$�w� ��>��L���UEWT����.�`u�8��a�L�w��݋ .r+M����F�ZVנ{�)�[�s@�@��s�ch1"H^n 9��G <�K@K�b��C��m��5m�r�q�_��x �n]*�m�F�̋����J��	T���-.9����	&� >��'�� &�jI#��{�߳�G����;���w4}åMF��G&�쪹��u�{�ل8Q��DD�I)P��(Q�"#39�,����hQ�qFL�(�RG������1w}��O� ;�K@K�b���x������33D�*@wd����t�h�ܺ�y	̒)�"L���F�V,p��>�|Ք�ak{b��ev*�`뮜�[K���ݤvIh	q�@t{�*@�"�<t�1(��ŠUz��Ҙz�`�ns�(��:��&�BBn웺�7z��o
P���wN�����,q61&���C@m�X�M� �X�IQ	z�PA^>��>�9��;$�f�\��B!4�9Rf�ﯪ�*���l��o]�⿹!��Iy	&D��1�"���X��^�k�;<���r�����n�d��B8��N-���{e4z�h�����Q�qFH(�mI��ٝ
S's�X~S;��p�}X���cdı��n�w4}}V�U��=���^m:H�$�p{����-.9�t� $qR �ȯǕ��H�n-���{e4&�ӲO߳ݽ�u�u�:T��!8)�,�D+���RS�[���X��Y�=�ـ�Eå�5�R�ɞ+����:ask�G6��i�î��r'��O]0���$�=Kn��3�o �R����rŝ] �z��u�CV���/��{L�y뢚5������8�^65rs��w������q�td�-�f ���SZ�!�.۟����%q=�}�鶶�F5�1�,4��� �:�h��F�d��}#h) �~�����o]��_U�Uz���#e�&�&���G ;��.9�t� $���i4�7�f�ﯪ�*�^����H�w41wI�x�PO� =�`���H�r����+5Lr8�RG�y��-빠{��
�W�~�����QɒI�?����n��y::�aaۛY9��n�=r�\LcWbn]v��Q93�>����{��
�W�y��<E������L�=��Z�dr���;f ޼Y�NN�4�s3�8�Z����<��h���=��Z/C��1�� RAH�?��}���*@wc�����f�7L��4����-빠}�/��>__���S@��j�r�2AŎL��g^^�ے�W`���mvd�]Qh{��m�5�e6�$��3@���h^�@��)�x��ۚs��q�2�܃qh=u�~�`�ŀ{ծs舅�Q��(���1̒(�RG�u��Ɓo]�?���X"�� !�
���}��˻�{�%S��Ɇ&≸hf.�ߖ�O� s���>��� ���E$��%$��4}}V�����}���=���/u��<I"Cqr�t�.��n�\=)Mӂg�K�<������]�gLH�Ǒ��H�n-�mz�۹�=׋���Hn����:��Ss �^�t���T���-/����%Tr|]Q�]�!JUM�V����v9h	|� =�*@F;��) 6�$q�&h}��~��/�@�u����,_B���ٚ�����h��QusUvU\�}���(��~_��}��{��^�E2F�71�F��Iǳhm������y��hv�n���z� :�ZLM�S�"���z�۹�_z�h����Q�N��_L�M`*��%U�MU���X�Z� s�u�~�g�D(���ٍ����褑��R8ԙ�Z���ϵ�BJ!)�o_k�X �˚
T˔�nꮪ��I)�o� ���_m���]�����^?��@�Id����ـrJ>P�|����7]��wW�vg��3�ȩ��g�ci!����d��\�Kv#M��-���V۪q�m1�v�lh�3����I��ę����7R���`�N��:�u�ˍ�4��t-��8!P�:���%���Px#&��9��N���,���f�xo^Fs�f��p���s�����M�]�cg�{3Z�klWG$�6ٞ^K��T奎۬���nv���R�~�w�_m�N�ݧ�i,��\�vZ�5����х�kk�����k�������l��N��o��� {�� s���_�=�|`ÛO�I�m�)$� �޳�~����{z���şBQ2n�Or$��T]������O��� �&��
X�&9�EjH�=���x���x�Jz���5����S&%���p�/��h���]��{e4/d��5�q8�F�H÷k��K���^sd�Ȩv�j7Bl�Q�y���{��6_�I#m�$r'3�~��]��{e4�s�Lht�1)�I6���x�pD�@/ʡ��|��`�ذ��y��%2�GK�T��)���j� ���?7��(�2n���o�@����d#�Ƥd���ŀ������|����������#�16��G3@=���*�@��)�_m��?�+��jD��"��m{uY	c�n�^Mحc�M�u��w�݌�����{�����:XF�ͷ�~����6	�*���y>�Y{���t]�UsU7wX�;fw�	DU?�ŀZ��Z]���IT�1�`��i�`���=��88�aAs
��BW��H^��P��+�`F��Q��� q������9��B��$�$H@�D�H����$dF$H1d�HD�� �A��@�F����A*�BB E �ߏDC ��N�Q�*z)��~�?' $%q	%�~����v��J�swwUUSe��լ��	*o;��>�� ��)�_m����c��bn5\�w]`(�Dk��ǀ���,ޭ�@���'!�A8�h�&%1�	;n���e�0N�M�͞�HGhsM-���&�n;U�BND�z��MW�|�<I.�w��?x�K�o��J�l�1F��q�ȵ$���3�K��ũ$���I{g�}��{����|?�n�U�i����J���Ԓ\���Ē^�bԒ^[|�<I.�
PQ�	Q���-I}���ߟ�[m��}��m�n[t;�T�B1����g���|�Nũ$��B��L�m�ڒ?<I%�-I%���Ē�wqjI.}���Ig��߿_�-ϱ�n(��&k\v�ݭ��Έ�ݬ�E���K��ݷ�}�?}�Z���HݘbdMD�r.I%����<�$���Z�K�u~x�K�,Z�K�^�9�j9$�<I.�w���J�~~x�K��E�$����x�B�U1<uŘ��F�-I%Ϻ�<I%�-I%m�y�Iw;��$���s�1���$�I��/��~�RI}����%���ԗ�cO����I\t��FFĒq�ȵ$��i�%���ԒU�_�$��������2{�{��o�{���8�[�lp۩��gFX�:ٓ^ٝ�MŲi&��(�����9mВlusZ�� ���{7[��ױ�&��z��ũYY#jRw�qpl�ʙ�����i;������ɓF��m�;�U>ݶ�y���}�Y���\mq3&˴�=f8'��Vۂ<�[�����<��mn8�j��snxA�A��b�d�;%Is?�_w��wv���'��Mѷ^iA�6���N�n.4�8b�X��64�c_�w�d�~�݁M5w�����qjI.}���I/l�~�I{��y�x�V�S�%����cs����_�$��������y�Iw;������D���Q)��9#�ĒW�E�$����x�]��-I%Ϻ�<I.�$n�12!1F�r-I}������$���ũ$���I{e�RIx��;s#i��G$�<I.�w���>�~~��K��E�$��|�<I/x��b�1��$l�b���=�cqN��:��&0���#�nJĽ���xպ��f&�Q��RIW�_�$�����~o��%�T̷]�r@ղ:]h�RMs�˜��'��y�a�Sȝ �>�H��H	m�@:�a7ܴ$���I�_m��;޻�}�|���߯�@�r��bI�)"�����u��t����]�|����=auҒ�A��n1��^�z�/~�O ��ۚ{�s@��b��5���"�b8w&�ʜ��+0�a;m5)/H��7LJ�G�$i��yz���s@�z�~�˯�@��>�b�1&�m759�H�*@K�1 z9�ꪻ9|��8�F�Y$�9����W�^�o�^�@�n���U4�7a��������կ� =ϯ ~׋�	^�y�#�^}0�!9#N= ���������`}��J!s�)���%�%�[uܽt�={4�ndH���8�q�vK��?�վ]��N8�V����H�*@K�1 z9��q��9�&���G3@�z�o߱#����~�����$^��
HӉ�;�j�ӯ� ?=w��)��ذ��4}�R��&D�nG�^�@~׋ �kŀ�/���g�(�KR�_�w�}h�,�8�ۍ���/�w0�����:����x�5o.�WU֬�.CW^�<Hx��%��1��l�rnY�g;m����	)#�A��)"�g�^�nh}����}�^���ذ+�马M�#16����*���/Y�_z�`�x��rU@ӓ�R��EMU�{���=�k@�sT����@:�a6�D�$܌�M��s@�z�hwW��b^�~�����G��I�f���H	m�@�jt��?Ǆ�k�V�cu�N�ǰDK,Ja��6�ٺr�ZI��ų�mk��ή��wnq�9x��&^1Y���Q�q;;LGA�[�N�� ��<&gH!W&n��[g\��ܣyrC�44w5�������b�m�+�v�����3�c <�0l֮���Nw!<<����vݍuS<�[�Q���#.�I6�kZKض���w����[G�}��P�j�ێc��F�q�뭇ki��:ۂ�V�GO�~��z���H�#�Ng�|�����@N�R���ٻ���x^���� �sP�T�|���gBJd{��}hR�䚪�����;{�`�x��(Q3��V {�^�G�Tʪ�Wwuuk�>Q	W>�� �{�� ������՜�i�n�16���H	m�@�jt���T���ϴ�H\��Em�r��iv���t�l#!6s���6��������羻Wfn���;���'H� ��H	mǠv/Nl�"&�d�h�w5��������ذ�����x�(�r8m�H�s4���Wuz��4�{�Y�)dw$լI(���������`#}�s@�څpY2dLQ�$z��4�B�D/��yx}�,����JZ�N�[uW�_o�XZĜ�=*ٳҞ����+Z"#Y���sVQk��� 8�-����@z�����m�jB9�{�s��bG�ߞ�������9T�Bt3j(��d�}�s�O.����(qD<�b����s���w��yӲO���ds�s�0�!'"N=������� 8�-��W��2f�E�Wjn���`��%Ͼ��OwՀx�W�z�.��29�d�8��A�3:�ۍ��� �����d�l@Orf�¸�u�mʹ(�L�;޻�]��+���� ���s@�r7���iH��'3@����9�	�*@>qR�Y{�4Y D�rG�x�W�_m���߿%z���|����%�b�6�#q����7��`w]`[��Q$���?���G�6����m�)�h�T�����9�	�*@zI��Ψ2�8�/N�r��ƺ�<1�f�,8������tv��-����`����9�	�*�����ϕ ���鄘�	�q�+���w4��X��Y�$�����⤵",�ʼ���� 8�/���:��(�r9��B�)���������:u�`���B�����=y��n��'0Nf�W�^��^����׋ �0�?E$)ݛD	,$;�~Nu@�u\?��`��!8�����9�
q���A�$�a-�*/U�1�� pC�
�H0cDb���kj�G��(@��]�;� ���������մ٣����T�K+�)Z8
Z��"�6q�$`�ke� �� ����i�l��E�o^�����J�&3�,��^لq�����3��s�8m���,�˓I=���gR�[��=�Tps^�Q�=�ָ6���1έq�l�����b�<�B�۞+T��=4`R�$sk6�R*vzx*^3<�C�A�t��s�
��rl��3��y`#`��lU�I�<e�!����.�
�US6�f���:�f�n����	L�8��+mŲ�(8��<�+��]/8}���M/`����y�]b'v�a)����m�qP�wKU� �nS�k�U��v���z#4�1^VJBq��tʱ�޶�m��p��,�Xjx#͑��t�ԤȘ�` 6E�	 ��*��w��-gR�:�v�pnԨ5R��ii��-\�T ����B�֑���f�
iy3���In�=�;Y8�z͛8��$k�AUհ/��m�ƺ:�(��gY4�	-��` ��e�䘉�(T-���9��nYuc���Z�,�5mV�U��%�ŻAh��p����'gv�d�U�U����q��dӹM�Q���Џ3�J\��̡�Ay�M
���m3O!+�S�y�7;�	��ZE�Wf�w8�H��U�w�
3YLj��ZF�Tt=��p����:x�PN������Q1s8
�6*����;p���k�hh	 ���i���V������Mi��U������*��gE���S�n���>����l�2\���x�^C����X�3t��ݫ&�3���2Ж�J�]!mH��mY�0��ס,���4^�Pۭղ����b@4[�^�8u��+��r[R��m��˸ѧ�	n�[��cG�:��� l�m���	e�t�.���l m}s�^�wHK0�=Bς��-��'2�g����㿅1Dt^�w@�"r"H��|A�_PE=N�t�����t5��os�P5��H��v�q�X�\[�jm�- l��W9�M��LF僙
��=�F\�k��,��-�����ȣ��k<�L8zϤvC3m<�K��	Y[�GL��'B;r����9x*Sm� Bsf�%S�bv��']m��W���ҹ��3��ZՔ�k��v�s�q���]v���qfԏ;�6�r�Z3~��{��]�7H]E���-��۳hz9�8ɬ���C��t���*�*�]�I��[]#S��~]`���7��|��_DD(^��{����$O�,pHj!��}�s@�u����?K�Y�B�='9�빚�m�nB9����Wuz�����`�e�R*�)J�.j�Д(����O>���X%������郂'$mǠy_U�_m��;޻�]���eC�� ��I`�v��6yj��]��х�i��Wl�V����~�(�e�TV%�%])���ov,}� �u�Т�O>��suG+���������o��ű�BS�!�D(�^H���Հl��`��Ϣ���#<m�r8��	��>V��.9�	�*@>qR�Y{�4���WSWwX�z� ~o�׋��<����'�X���M7&�}�s �kŀ9�u����>�Q��Fcue�MI']�G4��OD;q�#�mzs��:0������'���~���҉�Z���￱`w]`���?Hv�b�gMc����7�������h�w4����$���郂H�	��$�����7��N�P׀R���&���s@�ޯ@�^���B��I�ڛ���"{{�,��X��X����(������%#R9�{�s@��Z��4��h�+�I�f"�ӭ{Z�&���M�`�+��k0�e�v:�ɉ�M��Ǎ�G��9�W�h���q�H�*@wK/rf�[�w��W���=��*@>qR�����1c�I���z^���^,>�Q
e�>��ϫ r75N�8�m,nB9�{�s@����z��	/�(�J2�_���*U4�(0�6�i �9h\s8� ��Z�Z�9�	��ԙ� �H�{xlXBur�ƹ�����ʝ4뇙�&^�H60n���=q�@8�� �-ؽ9��1���H��w7�������@�^�@�J�e��co����빠u}V�fb^���@��b�7ڮ��VswEU�j�BP�S�o� ����׋�(���,z�G���@Q�O��<W��-빀o����s�Z�$�B�DB_��|��`$��N��Ů�-������t����
\ZyCnmv�:���� ����5���sk��l���Qv���=�H2������jh
�[ݺ(7g�*���c��X�6� �������>�[h���������HtY�X��(/k�짱mij�ۜ�r�H�WN&�@������i�ؕќ�U�u�����k`vk�O{�޻��w�)�\i�3�f��ێ�X-H;d�-(����|��ӣu�A"I�,pHj!��{�|h�]�����z����QȆ�U���� 8��Z����x�����p�L�<���<Q�@H�� ��eM��.®�oov���$qR�c���^��`�#lr-޻���ߗ�;����k��j�'�򪲪זeStmזQ�f���'.ݺC4�s$	Q���p���	6ɑ�Ǌ9�<��q&9hLr�8� ���L�3C���˜'3�d�����:C�!��ʤ��r��T�|�s��&iu (�'�qhW�h���;޻����<�.�X�Ēj!7�oUH�*@I�Z���K�������52G3@�z�h��@�@����v>�6b�1�ӄh�b��y<g9�;��ʯs���Ϋx�Kq����ް��6�i&9hLr�8� ��� �=Eyf8�HĤQH�+���L�ϱ`_b��s�j�4�0S�69�o]��빤�37�(�(P�(�����5ֹ�7Û��M�QH䙠w�w4_U�y_U�[�s@�NȪ���4���$�-�ZG 8�-ԫ����`���\�4J�M�Ѹ�ǳv�Q���5��J���(F*�j�^'�������@H�� $�-�.�j�c�$�Bn-޻��$wY�_U�yω�~�߱"��dqȆ�X����|�&9hLr��T��w.�	�$LUYsv�9B�I)޷Ӏ{��{$���N�� �1��k30����)74��s�1���JE��hLr��T�|�Lr�{߿����e�#m��tTC�۫@�&�E��f7f�o��6���Mj�8��f߀�|� ۊ������>����G�$��Oq7&h�w4+�+�h�]���'b����ͤ�9hL���T�m����K$a %<MŠy]�@|�n*@zc���w-me]fݗ��y�h�*@6��9hL�h��ʂO�����F�#j*�X��Fd�=	��]�y�C�P������5N&�g[�S���DZN��Dƃ����g�)=��#�pt�B^JVH4C�Xۘ�u��d�vݶŦ]ʲ+�m���kpj�u@���j:�����K����q��[vv�G!��ښ��޴�I��e����6�l���N�PK�]{rq�r32N� ��󓹅�9�V�ٛ�c�%^`ض�ޗ��y)L�S!�8�c�cf�F���NJ��ߒ|��Z�$�� =n�� �G��"s4+�+�h�w]� ����jbA�H��hZnp�x��(Je�ذ�}8ύ����!G�@�m��;��h��hWj�;ҥn"k(�rE�n�ŀr�Kz�O�=��p�x�
����R
22$Șb� cnQ+�Į��v�������;a�F-��3h��@t�-�Z��T��j�FaQ<iŠy_U��~���\
"PR"�DF�DS�S�y�{���d�{������~�߿~H����lǋ@��QŠ]�ŀo��ÔD%3�O� �S�����d��Xԑ9�+��3@��hW�h���M��K���2'���Z��� 8�ϒM].x��v��8��; ���F�鸸����!���ɧ��0c%����- �EH�*@t�- �l��#�E�@�m��;޻���Z��ZzT��BdMc�N���׋ �s��S��K�e7(EČ�*��Y��D �o�`	�B�i�	���1 �a����:� b�"Fb�8���+�B�4��8CČN��9�8���+E-Q�
s�7�!�U�����S�A�i�@@�u<��y�7<��I��N�=�=�ĔQ8�ӘG3@���@�@�m���3�~�4o���F51F�G������ 8������?�~��G# �!$ş����L�4u_^Hr��/Qӫ��kRV��+�9��F�����`�x�:�?G�D/Po���@�G��o��21���i��;޻�Lr���H���^`� ��W5k �s�~t���
"e�v,�������j!#�E"�������v,w^,
J#(���W����*�l�̉�bXH�qh��"m����}8�M��m�w3i�:����w^��,�-�LPඝ�j�6H��%{�Vʣ� $WNx�f������R�9hLr��T�|=/&���\��K�%��~��o�@?�W2{�]�����׋>�2y�M�ݪ���T�ҩ���]Ӏo�ŇL���W�y�%V�x�łj!I��f~���z�O� :c����-,��&E1LbLR4�h�w4k�+��I��ޝ�hq���N�&d{~��Ķ�f@�rq����BKeqQi�HJrT[NL2i�K&j�1,�&�48R�Jj�x*�S�ɴ��ɞ$��R�:dH�V^YLsN��=��\�X�OE���;f`���3��8ݝ��m7`ӷ �(#��3v�����v �n��4'���V�XD^3��v�4ۯu��Ɠ�x�^�N��Ѭ��@�.V�Z�@B�v��w������~t�tDL�=�˺�4�5y�c��v^�d��׺���ȓM��C1�2'3�>��h�78��_�D%�A�ذ������X��QH�+�h�w]������6af�ĲG�8��x��x��
"gz�N���7�Q��11�x���3C�V���;�~Z�ڴ����蓱$�N&�!3v`u�p��u�O��b�7v��m�������nh��Uǳh�K<dIy�k�i��ŗԆ ��V��r��Qr\KW�W�����- �EH����Ω*�cŎ,Q
H���͞��� =@}QO��韷�N�>�ߖ��v���ݑLs�����wm��k�>P�g�]Ӏ=�ŀ~��5B%;�sV\ݘ�%
)�����~����� u�<��n�ue�i��hL���T�m�1�@ZX�9���㍨%�q(�$Ͷ�n1mvy�O4ZE�:2f��w{��t�����bXH�qx���;�S@����3����h��O>rcx�<�F㙠n�ŝ
"dާӀ{��p�x��Q��ċKD��q69���w�O77oe��  UE�{����;��h�B�HƦ(ډ�N-�����*@6�Lr�r��ɴR��IVws�o�ŀ|�DBP������pΛ���Z��n�l&nuջxv�X�ˠ��F�%�p��m=dɞ�����`��<��a����~����w�t�- zI��*@z����iB(����`�k���	(Jd=�׀=�nh�w4���	0X��QH��M@>qR� =1�@;��C.�\�YNg	��vO� �@3�����'�}�ӲO7=��1ЋԠ��AP���y����f�\79���an�jn����(�u������7�w4�
�)hn8���h�%dHlm+;�[<��vĜ��V�6�}����կ��$�c��H�s<ߝ�h�٠w�w4uB�HƦ(�(�7- zI��*@6��9h9v��0x�$)1�$�;�w4}�
"��>� �w^ �l�wT��I3�y����m�H��I5 �EZ��M�����H��h��h�В�J�﾿��`��`���aE�"0!S�;�-����h4����rf�݈�M[�t�j�7tdYg$�&^Ѽc�[.��4L\)c�{W'�F�^4�Ã���P�>�wXT&�9��雔Ã�y�;Ir�۷j����:\��vM�aįӌ훅��[�Goq�5��M��.y��Uv�3�ո`�F���:(d�e�V�p�Um�-�<q�W;�����=��z���h~��6��n���-q��y��]�̯JFs�]=���.[k���Ǔ$�b�E"����w�*@6�Lr��y�e�7*�mWx��Y���P�U��,�]���ٵ"�O+�bǎH��4�T���- zI��*@6=�ɩH�"l�$����� ��4��,�
����5�Oe�ګ�n�MҜʹ�&�8� ۊ���#��w�9t��ynn�ݸ��Fu[q�� ͘��
���'��0k�]E�
u����s5w�{݋ �׋ �s�$�������?�ls��Ĝ�����y�UU�t��@�j��r��]�2���j��Z� ?6��2����-�nh�x�H�"�hD(P�}�׀=�ŀn�ŀyֹ��sf:�S�a&&��;�w4��Z�hu�߆��o��/�n���Wi�ڻt/����Ӟ�x(�8�����߳$��[�lX�I�g�}��ۚ��Z�y� �f@;��;#��3ow.�i��	���*@6���1#��/�(�HD�7���߾�h��a��%������o�Z� �JVLȄ�NI�w��h��`u�p>�Q�߾�����k뚤�1'�9�w]���� ��4����a�[L�����ȣ�b���y89�v����/r��pq\�8��qXwc�?D̑���<���-�@�z�h�w4G#�<n���D��-�~ċ�������}V�$�l��Q�bnM��s@�빠y_U�[f�ޕD�pi�y#��3C�m��{�����.}��	B�%�)B��Ｐ�;����n¦�o7ͤ�9h��@>qR�����9�N�����bW	�17]Fp5����6̽%VÊ�1QVe��MU� ~z� �kŀo���G�u_����%��1'���6��@�z�h���Z��4
�D�M�1�5sW3V��x�ε��B�7�^z���z�TمyA��bs4.9h���|�� �ǕyYR���3M��@�� H�I<��od�<s��#��Vaa��$d�+�?"@b�`Eꐱ�A���#�m��*%`����(%�X~p��TA�N0h��abQBP%������ p,��a1�HH�n0`�Y5�S�� :)�Ș�	���+b/r�9'9�f�=�l��c�����-���/;2��F���qyc�����5,N1gM����X�ɀy6��3SҮ6�ޠ� ��i��j����:�l�'(�zF�%�Ģ��Q2p�[�#�u$l�7C%�&�K���`l���]\��zݸ�Yڕk;��s6Ct3qK*���(c\��ul�}	���7u�v^@u�&�݃�3Q��P��.e�A�gq���lۚ$]u4�ۙ�i��Y%ݻZt�=k��Z�7 !�d���b"�k���&D��n�v�����v�(�K�a7j������qEf{�j.@�H;sV��{5�NL]
�x�Z�G3��i{k9k=�m�kuSB�v�����Wu[=�ւ�xv�F��``����&��׋�:����kN�"f�Fi#Ȅ�����e�	 	�"�t�!�j�A���n�Tcl�h�/]Q�9�WUP� [z5K�e9ɢ1�]��'s�����>y;���� h��� 㭺u�2�<�gaZ��f����W\����[<�֩U8 *�,Lْ�� ��m֣��q�	Ѷ�A4����;�=9<�3�jsn��<v�۬�CT�)�]��'�@x�y���t�k�ک0T@70�ҡ�(�TxL�r��˓��6��b� ���s�s��S�U*��L�Ir��Rkb���lj�Y�b���'I��+�)�΃�:��٭hn�j1�2�5��U�@p�R�*�m#b���L�������u�e�6-��j���0벑�2ûv�:[g�6�;8��N�œ#�]�q��x�ns;��NԚ:,�%-��NQ��F��d(����(n^����˨�j(�� )Ux3���R eE�!lV,v�*��m�C��]J��r�.![m�ؐ�-z��<�F�C�@M� 7+�A����
�$�UU�x�4�M� �yS�r���۶rs2	�. DN��zC��\A ������C�_���Ts���n�g99x��lFɦ�ʯ��.�gY;Lvq\�l����z;^zGcs*��ؚ�M7,iֹ�{�C�����^zI�zc=YTl�ی�R��F�1�z�nl��+p��z��]�m�� ���'	����F�j���C�˻bV��sYӳ��8�#��v�'�(q�,� ܺ�{N���ڛ�SX2����sWM���Ar��>5�G��N(�/���_B�8�*�[,�뭼�tp��h��^c^n�#��`��k �����'˹���uwF�^n����T�|��9h�l�;Ҩ�W�4�ǑHӓ4ε� ~m��׋?��K�(UG�D��#RM�#I��;�����l���~��-�nh�
�QLsL��5W8��x�^,w^,�����������Q1FӒh�]�������}8��x���UV^��kj.=�zD�A�$v􏒲�5�MY�k2%�$��2"18FۘĜN$�h�v���I5 ��H[�y����]�5k ��\��,^Q�$�Q�]����ذ�x��d�UE2�I[���m�I5 ��H�T����w��1:Fб,$�ܚ~���_�H	'ʐ��I5 ����37x��6������}V�ym�{�s@��mVC����I2&l�-��ۜ�thr۲��\��\��YGh��d��q8��hW�h���;޻�~���}��[��S��nG�z�>�2s�ŀ=�ŀ9�� mȕC�n1F�rh���;�w4�ߟ���B�QNc��� �Q@#@H 21�	�b�`�����m�7; �޳@��̉�1��R$�h}��B�{��`/���]�[ŀzv\��\�&�ueU�ηX(P�{�x��4�w4�u�F�6�5��t��Xڞ�琫c�1�j������]v}�k�����jx��k�9�x�}��/[��w[��Uֽ �\ٕ̈x�Av��� z�,�D��v,��V y�4�(�V�I�ǒ8ۓ4�w4:�a�S&�u���`��4�i��cs4
�נ�f�z��� �@�����N�7�l��^)�d��7#�m�@��}~���~�s@��z���Hڄ#�$NH�:��si��.�*�8���a�:w7m:nF�'j�H��b��$�/[��w[��Uֽ ��4i\�jA�8�I��7[şDB�:_u`�u�[şD%2z��6`�"�(dpnf��|��m��P��>�X}ذ�gf�Je�*+37L���M@G"�r*@Kr� �\�I�ł	19&�z���=������ <��*T"(U����Dј��RE��,�Bdie�$��:;]m8��r]t]�8�;�}[V�B|C=��C�����̎��Z�(kզ0�i��Z�;n��v��;t�iR�����m<��6�hz�8uq.N���8�gl�\on�y�vXp�����v_GOn'�5��`���m��d�n��r�Z�kj��6fz��yqNm����Ô�.�����o^��~��p�i��{�uƈ,CVC	����km�8�qҾ��7*�#��<����~m���R[�G5�����ܼ5Z������� �[��DDL����9�b�7���舙�'��WT��j�q ?�ڀ�EH�*@Krb9i*��n(��i�4��h��hu���P�%T�� �>���ʩ�(I������s@��z�h����??��$�Q�A2��v^�q��*��-��� `)9���v��Y�hwG�[�fm %�1 t�Pȩ ܻ�#�&�N��N1H��l�A������vg���;'������*v%�bX����SȖ%�b{�{��p�Bd��39�'bX�%����u<�bX�&�ޕ;ı,M�ws��Kı,��q;ı,M�{{p��e�a�9���p�yĳ���;ı,O�~�:�D�,K���'bX�%����u<�c������>�Iծ���{���%�bn{��O"X�%�����1<�bX�'���O"X�%��w�NǍ�7���������%�n��Q�q�Z;<×i���dz4���s�+x��'Q��ɜ9��9�3�Χ�,KĻwy�ؖ%�bo��O"X�%��w��	�L�bX�f��u<���2%��?����-�yL����s�,K��~�é�Kı7n��ؖ%�bn{��O"X�%�v���,K��&���nd�K.Ng2���,K�ݻҧbX�%����u<�c҈g�P� �tO�<�gw�q;ı,O�����,K��6�̅�yK,�9�fp�ؖ%��2'�߾Χ�,Kĳ���Nı,K}���yı,M��J��bX�'�=���˷��&K��y��yı,K7���,K��w|:�D�,K}���,K���w:�D�,KM��Y�r��yՒ�ݺn0��umd�kc��B�s����qYk�uo�����_Z]��gEٹ�'�,K��~�é�Kı7�Α;ı,M�ws��Kı,�l��O؏؏؏�x��n4��8����,K��w:D�Kı7=�Χ�,Kĳ}�q;ı,M�o�����#�#�#�^.���$܍�\��,K���w:�D�,K��y��K�@!�2'���O"X�%����"v%�bX���]�ɜ9�̜���3��K�� dL�o��v%�bX�o�xu<�bX�&���'bX��>�iA�}���>���gSȖ%�b}6�~�	zr�3�.g9��Kı7����,K��w:D�Kı7=�Χ�,Kĳ}�q;ı,O�~���N��0�s���÷Ek7�x�ض��t���g��������������. z˜=M�bX�'���gH��bX�&绹��%�bX�o��'bX�%����u<�bX�'��.d��9Y.C���;ı,M�ws��Kı.�w���bX�&�����%�bX��ޕ;ı,Or{g��e��d-�r^s:�D�,K���'bX�%����u<�c��"dO��t�ؖ%�b}�����%�bX���Ci��2^g\�1;ı,M�wé�Kı7n��ؖ%�bn{��O"X�%�v���,K��g����[�&��\���,K�ݻҧbX�%����u<�bX�%ۻ�Nı,K}���yı,J�p1_{���;�������M��,�=.�c(�h�vh��:<��a'g2%�)1չ�P�t�v&�v\Φ�Fn���q9��`�mi�ܥݖ��re�l9Ḿ��O+*���p����=n�V�=T��8	ۜs�˵m��wpm���Ӷ�䇅�ǭ���C��� [��9��ɱ�ޙ�|G�7XLXQȝii]nЄ�$��s"��!a�y��8r�3=���P?�{�[?���e��sU��ڈ�[�;�&��y)8���nQ9��\�Û#����L�6%�bX������yı,M����Kı7����,K�ݻҧbX�%��e�9�����fg.e�s:�D�,Kf�q;�T9"X�o�xu<�bX�'�_�T�Kı7=�Χ�?�G*dK���ό%��L�Yy��v%�bX�o�xu<�bX�&�ޕ;ı,M�ws��Kı6n��,K��&�.d���sr�SȖ%�� @ȟ}~�ؖ%�b}�����%�bX�7{�ؖ%��L������Kĳ��D\���Pݽ�oq����绹��%�bX
~�}�'�,K��~�é�Kı7w:D�K��{���?����'q@�<�s<m�.66㍛T�sk6��6�S�uo[�0�E�K���2Ys�/9�	 �&�v� �	��}��$BA���<��,Ks���yı,Or�s!��	2[̹���Kı7������B��| �"v%���:D�Kı7?{���%�bX�o��'b|�TȖ'�6���g2��0��2�8u<�bX�'�~�S�,K���w:�D�,K��y��Kı7����,K��f����\Mq��{��7�������O"X�%�f���v%�bX���SȖ%�bo�zT�Kı?{���d�J?{���oq�������,K��EH��}��~�bX�'�~�S�,K���w:�D�.��������s��B���]�t��j�ϩE�f�&e�W���O�o�}�w�kH�g�����s9�'�,K��~�é�Kı7۽*v%�bX����SȖ%�bY��8��bX�'�7m��r�r��S�����%�bX��ޕ;ı,M�ws��Kı.�w���bX�&�����'�TȖ&��.d���V[��9�§bX�%��o�gSȖ%�bY��8��c@�&� 9=�c	�J4�WIq>{@��_�E8��(|;(Ő @���"�����i8/�3���0���X�=IH�G𡊘`E�A!���!`a	c�FMG�=��J����a0R1���$m B��
%"Z#	*D�F�"�=��DJH�$,���$bD�b��)!!�$$I0�� �1 8�Ĥ���HU� �@�� A�Ǌ�
�@���1ȰR	$#ȱ� ����<G�bp�$�e� �BTeT�H��R�0��DH1� ��,HF��$,@�GPV�� �����
��@?,�@�zA�QC�j*����6&o�xu<�bX�'�n��ؖ%�b{��=�3��K.s%�3��K��A`dL�o��v%�bX�o�xu<�bX�&�w�Nı,Ks���yĒ���ڡ�E �f������) �,M�wé�Kİ�#�߼*yı,O�~�:�D�,K�ݯw��oq���?�e���/,'Dz���B\�mӲ�n��>&5�ѹ��3u]�&Ù��s$×�˜���%�bX��zT�Kı7=�Χ�,Kĳwy���DȖ%�����SȖ%�b}���4���h�[�w��oq���~?���yı,K7w�Nı,K}���yı,M۽*v'���$���7��������Z��~�7�ı,K?�����Kı7��SȖ%�bn��S�,K����Χ��7������>�e�a�w��bX�&����yı,M۽*v%�bX����O"X�4�V�q��L�y��v%�bX�d�r�̹e���8u<�bX�&�ޕ;ı,>D?s�Χ�%�bY��s�ؖ%�bn��u<�bX�{���~?H�6y՛�=�73�㫭��f0�7�7v򕬯l�c6�\G�'T�
��bX�&���SȖ%�bY���v%�bX�����&D�,O��t�ؖ%�b]6��3>��d��2s9�O"X�%�f���*�r&D�>��:�D�,K��*v%�bX����O"X�%��Y�d&��p�%���s�ؖ%�bn��u<�bX�&�ޕ;ı,M��Χ�,Kĳwy��Kı7g�w��.Y,��-�8u<�bX�&�ޕ;ı,M��Χ�,Kĳwy��K����'�����SȖ%�bO���ul�e��}����ow�����O"X�%�f��ؖ%�bn��u<�bX�&��H��bX���D ��@C�~��ܼ���^^�kvvuҴ��ܭ��9��)p˰m��������M���h�nDZ�i�[p�춗�n�˞����<�c��vs4�v���HX-�-�w<�(�Pu�6��U�;1ɜ���$�oE�WN��ŵ�,S��N���a۾��^6{tu���Tm��j6�����:є2�nk�b�P^���S9C�)|��8�n�BZ���w{���;��8�s����WoU��(d�M�Q�������]��BFL��l�����2�Χ�,Kĳ��s�ؖ%�bn��u<�bX�&��H��bX�&���SȖ%�bl�m���f�fr��s�Nı,Kwwé�?ŎDȖ'�}�"v%�bX�g�}�O"X�%�f��ؖ%�by�}˛&d�巐̹é�Kı7w:D�Kı77w:�D��TdL�g�}�'bX�%���}���%�bX��n\�%�Z�r��.p�ؖ%�bnn�u<�bX�%���'bX�%������%�bX���"v%�bX���=��n��:g�w�{��7���~~~W�ı,Kwwé�Kı7n��ؖ%�bnn�u<�bX�&��3/�5Y]s�ɞ�����N��7vv�b����5��նy�X\Jiwi�=���jNı,Kwwé�Kı7n��ؖ%�bn�v�<�bX�%���'bX�%��=��m�r�I�r�s�SȖ%�bn��S����QOQ} ����؞ı9���^��,Kĳ���Nı,Kw���yĻ�ow����r��45������bX���gSȖ%�bY���v%�bX���SȖ%�bn��S�,C{������>��%jV�}��oq��%�f��ؖ%�bn��O"X�%��w�Nı,Kovu<�b�ow�� ��l=c,#U��{��,M����yı,>��_�*yı,O���N��,Kĳwy��Kı?����\���0�^^C�9xW�*4�l��x�T�M��#�����V�t�d�)�o!�����ı,O��t�ؖ%�bo��Χ�,Kĳwy��Kı7�wé�Kı?fܹ�[���fNs��*v%�bX��{���Kı,��q;ı,M����yı,M۽*v'�TȖ%��7���p���2�9:�D�,KϾ��Nı,K}�|:�D����W�� �A;�;�zT�Kı7��Χ�,K��,�2�9p�˙�y���,K��}���,K�ݻҧbX�%����:�D�,K�n���$)!=6L��쩩	���p�yı,M۽*v%�bX'�_����:�ı,K����q;ı,M����yı,{��d�C���]n���{:�ݱ�Y��IC���u)�d	��h;%����Mi��}����D��ݝO"X�%�f��ؖ%�bo��SȖ%�bn��S�,K�w���1��+R��[�w�{��7��f��ؖ%�bo��SȖ%�bn��S�,K���ݝO"}�2!�߻��u�z�XF�����ou����O"X�%��w�Nı,Kovu<�bX�%���'bX�%��Mܹ�.YN[NL��O"X�%��w�Nı,Kovu<�bX�%���'bX��!� JTT�� �.���SȖ%�b~͹s$�yk-�9�fp�ؖ%�bo��Χ�,K��c���Ȗ%�b}���SȖ%�bn��S�,K��>ݿ?�I�B�&P��v��E��7e�-�J����K��mu�2�ɧ��{Gٜ�'�%�bY��s�ؖ%�bn��O"X�%��w�Nı,Kw���yı,Or�s!sg3	,��Y��8��bX�&����%�bX��zT�Kı7}�Χ�,Kı�w_T¢���&R�*jBB���p�yı,O��t�ؖ%�bn�ݝO"X�%�f��ؖ%�b7���_�RB���2�j���Uw̼�;ı,M�{���Kı,��q;ı,M�wé�KıM��0��$)!I|�v]����U\�s���yı,K7w�Nı,K������%�bX�}~�S�,K���ݝO"X�%��hA����>�� �g�[vR*��;du]��;oV��4xK�6.�k{-���p�i���]F�wa�:ًBC������n��Իݍ��LYUd�����1�`����x�&��m,�n��v�1ngb��'wn-u��-n�Ec�x�cr�m���5�B6�vX��֩KoT��>R�$�{���1N��Ў�go�}��?Yn�9�'���
:~O«��=�3��-5Es߇�o���t9ѴS��&�H��׫���]H7>�a�w���d�?�߼:�D�,K}�ҧbX�%����:�O�2%�bY���'bX�%��'�eϦ\-9�����:�D�,K}�ҧbX�%���vu<�bX�%���'bX�%����u<�bX�'�ۗ2Iw��ٓ��g
��bX�&����%�bX�n�8��c�+��>�~��yı,O��t�ؖ%�b_O�{�f]̤�.s9s���Kı,��q;ı,M�wé�Kı7n��ؖ%�bn�ݿ{���oq���SWr��4i�'bX�%����u<�bX��~���SȖ%�b}�7���%�bX�n�W���7���{������krܷOR�G]�:�'�p4�����] &Բ41��٢�X3�/92�%�9�s�:�D�,Kv�J��bX�&�����%�bX�n�8�<��,K����,K�������V����}����ow�o��O!��_"b�� ߆4�?D�,����v%�bX����O"X�%��w�Nı,K�v���S+̍O�����oq������wbX�%������%�bX��zT�Kı77w:�D�,Kݶ�s���,��˜�8��bX�&��SȖ%�bn��S�,K�����yı,K7w�Nı,K̛�\ܷ�2ӓ2���,K�ݻҧbX�%����u<�bX�%���ؖ%�bo��O"X�%�����y��LtD,=>ݗm�9^�К��#5����u'O�9���2����c�=�����ŉbX�����u<�bX�%���ؖ%�bo��O"X�%����S�,Kľ����w2���K�gSȖ%�bY��8��bX�&�����%�bX��ޕ;ı,M�ws��x��{��������������bX�&�����%�bX��ޕ;ǹ������x����=�����u<�bX�%�����,K��g�w��˔���%�8u<�bX�&�w�Nı,Ks���yı,K7���,K�dO��O"X�%�~�o��0�]r��&�����oq�s���yı,K7w�Nı,K}���yı,M۽*v%�bY��?�����Z�B�-\�][���V����tv�m&z�ôa9]9ݹ��}}񏾵Z�2g2�s��~�bX�%�}�8��bX�&�����%�bX��zT�Kı7=�Χ�,K��m��圹�%˜̹�s�ؖ%�bo��O!����,O��t�ؖ%�b}�����%�bX�n�8��bX�'�7r��e��yL˜:�D�,Kv�J��bX�&绹��%�ʩ��,����Kı>߾��yı,Oٷ.d��-e.^s��*v%�g�
��C�?����u<�bX�%�����v%�bX���SȖ%�D	��g"}���Nı,K�{�f_�)�I��y��yı,K7w�Nı,K}���Kı7n��ؖ%�bn{��O"X�%���N��r�˚�T�݈�݇���d�d�rDWG$�2K�Й���Lew�2Ӧ�w��oq��&���SȖ%�bn�t�ؖ%�bn{���~��,KϾ��Nı,K�gp�8^e-����:�D�,Kws�N���DȖ'ٿ}�O"X�%�g�}�'bX�%������<oq���~~o��0�]p�P����Kı7=�Χ�,Kĳwy��Kı7��:�D�,Kws�NǍ�7�������ߓ�H�̋O����bX�%���'bX�%������%�bX���"v%�`}2'�߾Χ��oq���~~�~�o"��W���,K}���Kİ�|#_����H$�����I��}��I�QE�QE�AQ_��AQZ�
��҈*+�* ���J ���"*��"�b("� �"�1� ���H��0��� Ă�B�X� � ��("�0"�� �AQ_��AQ_�QE~QEj�*+�
��*+�J ���(����
��҈*+��AQ_� ����(+$�k(�3�`{�0
 ?��d��-�D�  	���� $�{��PEP�� J �" ��@�!**��R��� (���H��AJ�J �BQ �  � D�`  @5* B� 
d m���Ž�S�h���9�� @$��N&�R��R�Y�)A�}mԤ��ΊR�YJ J7YҔU�R�& e*��)JR�)JR�R���R�� YJR���14�)n�Ҕ��R�� �8�  
 
��.
R���)N&��,̔�LM)JX iJSEJ��g�qսǢ���zf�/�X= �
 �}��}��gA�ǡ����:�� }�zO-�U������Z� ��)E
  (
� }_T���˻z���oO'U;� �/\��UͩU�J��{��} ��q>��=������+���ּ ws��l���]73S�p@s»��^9�|��w����qK��>�   
(
� ��7�>ܾ�y�q9U� �$�d4bt��0z��w)\���{�   ��ͤ��wm�� ��K������f�{�G�� |���ӑ�bi,l��x �   (�*� >��K��N6Qci�95K � �z#��7ͻ�����$˻!� �sɥ�n op>@w��݃��u�7�;� �� ��|0x����L� 4�M�%R�  0$�JR�  D��RQ�T���LD�*�F�j�  ES�Е=�J�� ��	��	� ��t�����W��?���r��Oxs�����TW�u좊��O�QEE袊���**+PT��O�Ц��L��)#HB @ �b1#C Q��B��H�H��b��$H�"EH��`X��	4ԂA� �H"�x�����}ωu��HA��~y>���F��̄��_�d���჌d�s>hk��f��L))�!P��A�D۵�� pO�gE�
�Ve�Z��c5L��)��5��h��3L.�d�XHI~�0�b���p5�4#X�1%1���s3]����e2�R�"j��C�`L��z�O�e�'�:S��|�b|�<�B�e	v˄(@HB���Bs�j2Rq˰�Ħ����MRLt2�8�\tj���h@�
A���A����NQ�9Jr�Y�7?҆��Bs$�D(J�e��k5��Ç~��߈��Ff�s|�l����K���$X�����$C��/��8�hc�gS�S.�1�E����4s�M0˷�/5Úto��!a�X2$ B$��4�6|�5�B|�S���r����o�����I��B�Ϲ.y]P>g>�o٠��X��#�a2`@ ��K���:!�WS�9x�沐: q5��V�	u�� ��K�g��u��l`1+�ʑ���m�X$�>�)�c��M���7.kM�@�$K������<GJi�\4h�_�L�E��,c��5�q)����a���4�4t���$>9��M���aK�)���đ�ۨ�"T�*`e�޷#�톳 �H����aXۯ���!s�i�$��棃�4�A�@�VK�4�϶I$5����'�� �bP��F�0�ċ\'�c)�	���}�+�$¤)�
�#p��35�ճ(Mj�).�1�A��2�[��޷��ϓ�K�p?���P�)s'��F\�f��1§��(��YHF��i��2��C��v�淾%~O���Y��w\>�>�J�����ͩXp�JV[�� b�#�d�w��(!]�{z>Yq�3d��kfB�f�3�eIXT�0!BX�P�!:�)��8�d�80#�9���!�8av�/WL7���F�}��9�N|���`	���	��xS\)�(00�.4��C�xR ��)�߸�W�;�-��}�g���N����"A ���"$A1�0@�P"�LR+� j@��#q1 1�8i�
b�)�q�a��H��_��4�����,FXB �1$�D6�n���0)�F�}�2����> �
��2�r�8S�5��
���A��>aO0�:�3dY�*�^8X�aMP�p!���0�aA��PaV3F�!�i
��B��K�4)hee�l�i5sG�!���+��!':���̇�̡\��xB`3[���f�Vn5aJ�f�M0�h@�	�$Z��|��@�a���hC�q�#cBT���b�b�E�!�Ũkf��s:��	���	/t���HCi
�E�8@#
}�����S!qʒ�)�).�)�*64�bă�4蒛ae��֯4|��kA)���kd(@����sF�h�n[4xVi�zaL��S#����LH�ٿ���8B�C{	����"$B!F� �c��8f�n��a����dp#RB�3&��	!��k[!��8Q�H����"V��FE>����S���BH6�=N��,B��cB�幹�k|7.��s��t���!p��\ZdKv���.$�,��\��@�4�N���
��'&��eQ\�r�}���ɸ9-)�8�)�\�`�
9Fp+�s��g���1!V �F�n�-0ѳf�|��7�\޴sF�>�˜4/�l	�(� �%��O����h���v�4sd.`͛�h���F�����`������ħ7��0�
gW��$M8����4�a�	+�3H`�E�"�#Zb��7n���	 �j`C�k6˽n+������łE�3j-�#��mS7���Bp���B��[ؑbJf�`a�0��f� �@E��\ֹ�W;S4�K���������+�Z� �(:P\�\5f
iN5 �'�8�c�	��nx�nswe�ڞ�{��q���0�r������9_�ト���1�)�\).}Ņ٧a�8�F�f1�j���(J\L)��s$e��� \�Lr��1!
`��橉:Q1��$\bZ�}�����s�3�`��c���(�%IB\%�S5*�@�2��ݤ&XII��J�*J��E�S��gĹ�}����4MbK�#�6D�(K��f�r��,.�Y���R�S\	q���S%aJ2���Jb��K��\5��,0!B$��-26K�\�aL�S	B,%(F�j�!�l�0�#�X�#����XST�$ �c�:P�"]�H��$(I#�3f�a
�����0�	l�hJ�S!L	H�8�"F��JB$�%2���i���.5)��ο�����a,!�8�`$*M����{�/�fJ�c��\.�m�9���s���>�*�!�8��/��i �)&2B��oħ�� �X��!M���."`PC�BXH\q!FRH�$�0H5�s8��M�$�	.E��� D��k��I+fѼ���t�T��΄��$@%���}�8��BL`$�&�>�R�E�w�Bb
jZ�P�	Ǐ��`Mk	T�'N�Ϸ:B�q�Z� C����b!֌�CH�>��χQ�.gÀ�0��`Ipp>"Ɋ\���`}Bo����ߍɻ�����p�
�|��\����P���B��(i
�7�����Ve2�.B�	hB���%�*��)��u�M���Ǒ��a��O0p)�	�y�{�o4�3�R[�%���#�pt1j$H+]`G���R�)R�&�����9ߦ4F��&ɚ�VMRh�$��t�V�X�'	5;u����~61!1b�b��
�F�� @��k����0XE�K ��C�)t��	.�Wha�ǐ)�A�9�.�BM]2�1ٱ�Ѵ�7�	L�2!�R]D����j�����ܣ���>��LD &*��01��>��j��%�¼LhJ1��qYs[��T,�2�uH�
1`&,)
�*O�$�N�J9Ȧ/�����߲�rt.i����v�������}�+�8;�[?y�� i�B$`B�))�;�c�m"�����"P�0���58z�͒�D� `D�Y�(ʒ�lX! ����@�~�|k���e����X	�[<�u��)�(��3MpP�(>��'S������~����sr���0`NR�>�:�s�n��v�9�%����LKNg-n1�D�~̜q.V0>Î�P��̄Pu5�_��9ˇ��P��8<�8S@'s�NL=�М���99�.�*L	�Є�����T%�ƸR4n��(�����
�Ж��!� @#$`bX, B��D�c*�� J@��R��`�\�3�	���@`���+�6���p��6�XD�51CIV�:P��IX���!�X\�*�v��lB0X�`�����B%1��
W W5�Ґ��ϳ%��&iϴD*j�a����O��٥���=H�$�`�#H$A�b�0h(�h� ��R�5�AX�D�1`i8�*8�514j�,	0��D���tZ���[�4P�a��:z��Ou������ m� � 6�H ��  �m�� NM-�f�Jn�,���=.渙P��媩Nt��C�/I�?������N�"]V�8I��v$H��k&�Q�-�����N8^�V� s� Ie$�n�m�� ��� ���Ŷ���jmUW 6��
UѥZ�(
�*��������-�m9Ҏ��T� �ۀ��M�@ 
���@As�;5T�0$p ���� ^�Ԁm��` [N   �.� �ٶ����E:@i��n۝�6� I��ր�[\	}(�e˦��[B�  lt��դ���ж�m p�zr�J��Um˲��x�R��4ٺE�$Ǡ�L�	�k^ʶ��#�FDj�k(�7`� j�qP��J�gZ[c�����-6H 9��īv�m»�ϒ���4̷m���i��ɝ�2�U�����SY:�驶j��� �hٺll �c�n�Z��,�U�MnY��Im�m��s��uR��V�q@NSh
�ܜ��Uu��K�3.�K� K�R�q�,m6�u� jۍ��^�o��OJ� � H -� -�l       -�      $  �v $ �O��䀶���ۀm��@��{N�f�n�5�  [B۶�6� m�f
�ɽYڕWe�8��(H�\*����mm�$�鷴j�(H�U��$a�-�gF�QڙV��VÈ���3�<ꐐ ��۰ 8m�[% m     $	     8    �     �l6�� 6�  ���	$i �m��  ѵ����m�%��n�qmg�6�'H���rf����ر�ضIn6����@ c:ݺ���CR��u��{rI�Է 8$�-���z�ۧx�e ����?C�| qm[@ڐ������l�� ��\L��Ko [@��N\K�����0G]�.�uR�t�ml c�س�p@��U��x��i��  �^ɫ�qiÜ6�  6Ͱ� p-+kh I2�)yJ\�UT ҭ<�4u�Lq�4�l� ��W-Uu�l$+����E-Uu�Γ�m�kj� ���v�{]Q\�4�@zҗN^���:%6�cf� �usK�%�PP ��n�y$պkj�lLUQ��6�Vۀ�g&�t{H����!�\�ĵu�o��|˫=�u�-�R�-��KFy5%Uo,��3�ҘRR�;U{�VJѳ���MҼ�� ��	�G���7!�n�lY涫j�%�� z�\�M	m1��e�w^�mp���1�ݒ����e9�m�[�2E�� 8�����ڻZ�)�����%�Lfݤ���N��l�@��W�6�`�j�
��2)��	I;��66` :AmvI l��*�K��(l���^Z�ܰ��ZV��k O��"���8kCH��`�Z����+v�p6�t  �8[sm�qǻ���蚪�;��0�JiuѲ�d�[��lH��m��JçN�M��&�YƑ�7����Z��V^Z�۫�]��� -� 9���yc�r�WT0*��m��mi$�$့Zۖ���ضg��|c���MR��UYx�Z�m�d���XH�f�:.�u)  ����ڣ�KoI�$ 	mz�m�N [�k�Uv�0m�$�� r�(o����6�H � G�Ӳ�.մ��v���9ʁ��Y`�z��u�����M�m�8p$H	� �r�8ɣ[�GN��lƷ�׮$뮌�ZmRi-�&�R��Ai�� �eN��lIu�M�9.��)V�Β�`@Yo[e�W]!m��6�@��*ڐ� �%��`�]��۴�ͮ$����m&�6���� ۭ�ֻyJ �� ����rIe��lNlK��U@�.�b�"P��$��l�ƌ6Z[�:�ζ�i�*�Tu�:+��Y{!����]&�B��$r�Umm�6��  �l�sn�-�!�UT�u*�UU+���_]��R��m���*���5�ٶ��P3�����ͭ����IɆ�N�*]Jʾ�j��h���q��H�<���nE�H[[M��ݐ��m��M����J����(
�UT8�k���]:.�7t';-�-�Ԩ
��HvM��m�-���N���[-��lf����X`6��Z����]�i�ڭ��15���&��{����]���8V{d�]�d�e^���v�Xvo:6��^���sj��Diҝ�g����v��;u�դƒ�Iߧ�����᛭���ʙ7dѠ�R�a�r�ذ�^��@@uK��U�*���8�Z��$m۱���1R��Jnl�Q� m�/.1��UR���{l ����8��^k;P�&@Ƹ �m�Mn��m�4mc r� r�s`4���e�_n�@	&�p �mR�@v�mpI7j۰$�m��U����,n@j�'76�<�t�k�]�lHP�� �Nvյ�pd�BBA��t��U� :d�J6^�e�$ ��m���1k!"�Ö��]���-f���pN�Հl6�Hݶ |m�8�6Z+���6�]����7���$m{Yu�  L�P�Uke���|]UPhRа���&n����g�4o�h h� z�+��[p�m�m�[Uu@U)���� 6�j���y��},*��I�h-� ��!"޸;�6��+� �O�l��j�ArW	V6 p۶-�l�[����m8�5����� p �    �%��؋�6�  9�Ͷm�n�[$�5������knmml�i;�nG��`��RKyoN�k��h   "@	 m�	ew˺'�b�um���A!5N�A�X4�h9Ͷi&�tۖ����Jm�Y�:v���۷m�8� ��n��[,2�Ö��ע��H���n�X�BGl h�A�$�Mv�� 9�Q�e�=d��&���.��R�9�9vl���MPʻR�um*�
�ju4=���8��iV�8y����v�ke�1m@�&Z�S�k,�/[��� h.�Z�H$%��� 'YGI��d��Z��3 �8   ՕZN��;`x6�f2��J�*�	/[�e��Hp�=N�$�m�gm���UT�V��N��g�mJ�*�Utu��!�+��*���e�<�p�i�۶��m"�[��%��#�� 7m�	6�g^��Սu�ɷ'�0�t��@ ks[��}�& ;l�$ M����rLc�z� �5J�;t�Z���F�Yp  ڶږ��]�U��V��g�!  m����iiۭ�;QrS�[\m� "@�����86�l�	�$�L9�n������   ��   $  ++UR����U*�U@T�6�f�:��PP��� � ���H�m�	��8ɶ� 8-�8          %��h�[A-0M+[@�   �i,�Q��[C� @�m 88p� �]��-)�m@++W*���m��qÀ 8ڶ  H�-����c\�  �[V�M�i��`���l��-� /I-�̑���d�ր�  p    6�X>>�� [[l��l76뜒D�"Ӥ�m��	���:�   m� I��V�[�[@[x�jc4�CD�-��6� �;�nհ ֻ;[�Z    $�@m�K��m�6+*Ӣ��t+J�ʵP  $;v�m�m���V�	$u�&����Hm㄀ �˓i-�V� 6͛`�νp�n���` 8l �8m� �m�	$mڦĤˇ � $� m� �b@�Y:㍶���� ^�l6͂�ɤ��mIm9�   $�XI�	u���� ����[gH  z�������ƚ�f���	d�
LEv�q�ޥv捍��c��W;+qJ l��͞����C[.��� �e��  6�cm��"����@��m�e�    [�� �  "@8ֶ���#m��(Am$I' Zl���ڵ�m�U�\��Է9涗��An�	  [[l�$-�  �� �	���m�$    ��  m�H    Ŵ�-��[M�Ӂ�֙� �m�� h m��    6�`    �   $	 Hm��  ���m�ٶ �m���+T�S� @mU@U��J\z�&R2uƚ�?�PAAS@���@?n mG��.�P1������� �(A0C�A��Pt�P�TT���B.
 QG���Z ���]*���`�i@����EȀ��z"p�QN*s��O�[�����<���1�` EF A�H 0(�m~@J|��:E(�����A�T��::Av��P�*"�8s��PL@T��mx�H��W�v��D��τ��ƔS��Ȧ�R�@U<&�Z�.�E�W��&i�*� �$X1P�H!@'��ms�O��@
���(���A"�AE�~M���ZiA��EU�% h�<uE4 D���*+��D��Z���fw�^Z���A�ӆ��K�٭<� �!�-���+�lĻ�ƻMZM�w<�ʦ����1T���V��|-	ĥ����xǆ^O���m��!ծ����i+	��rnw�YM<�vj�\A���u'	��`����!<�i�ÌR\O����lh6^n,�Ua-I�����@��vܶC�$�[W.�C.�8X�RΌ뜒��rJ�������u�ގ�$x��G7Q�E�=s��a�늡�v��BwF�d�YJ]L�vb7��0,�v�Y��Z��j�[����Srn!v�q���6�������r�c#=���6��<2e��{bWv8���ґ��,ugV�\�;N��Ւ�vs�m9�bQ٨�YS,�(�/Q�r&GZ��e�s����6R5*�h�R�-�Γ$�^7i6�U��ZVͧ��@��V^����ӫ:$6tY�tV���ɞ�k����.x��#�F�dk��ܮcq�`%wn�a��[GlqO.�q�^��;s׳䒳�B��;u��-s\��v%������և��N�9���5�q	ۑ'SD�GɄqgZvܹgk��	�g�U�l{eƱ�E�	ۇ�)�7S�9�	�f�"<��66���R�t<i稴�u�jyEEgV5)�E�v^d���5� OS�/\��0&�8'=f���(�Z%Ӱ�Yq��� �]R�@�n1��fU�2���2;�' q2[�,��G������pݙW+8N8�k�
mn.��{;WR��/,��%;rJ��KךrVp �����G$�[}iҭ@�cbY��B��θ�ƻ,`�
�UE^5��.�]��QU��gjWn�r��V��r�6HӝI��e�ح�rh�*;V۬֩��X�{e Шgcl���az���d���dų֬������@c,Lp�ۍ@���F�;f�kf�H�$��(� -�i],Ꝑ(8�i�0�@%g�^x�:��{��� N��4'��'ȃ���Q��N!��?Qa�e?_Ǖ=� ,�
.80�u�r�u�� �(0�1ړ`j��dƹ�9��K�闝�`��8�r��s�O0M�n����ۤ�ۘ��]��8qr��3
�@���k׶��k�Mۖ��H�d�V�`��\��4ڡw*P��;P����q�-�]��H��J����ǲK��Q(�׳4��E�+Y���{�P��&�u��l�I��7e7/8��p�;�QNO9@����'M0�I5��j��`��`o����%����X>��ɺ����a��X�_ov�$ �����/}>4zS@�����RE�#�M��h�)�[Қ��h���c#(��8����-�M ��4;O��=j/�[�G���[Қ��h��@�YM�{�?7�n��`x�Jp�P��t�R��z���ۜ���xS5y���zt��z�����;�S@��4c��4:�R���-Ė��4�;�S �b�@R
Q���%	F-ID~��_� om���4�=pN��d�cm���;�S@��4�٠Z��֥+c�&L�
�`�:d7�� �Ӏn���^�ErG�8�X�N��h��@�[��[Қ��;QbEF9��(�ԓm�F�[�w�J�:��.�1lhitWb[i��:9j��~~?�Šw���-�M ��4zPsn1�	��@�[��[Қ��h��@����n5HnF���oJ`�]�D$�F���V���@��ܩ<x!�I��4׬�-}V�޲��)�r����2aB94_U�w���oJh�Y���������m7b�^i�열]���`N��]�=�ݐG][e�
�%�<�v{]�[QŠw���oJh�Y�Z����]i&I�`��$��oJo�}~��;��;�S@�Tj��Q�c�	�@=m����;���oJh�Ût�ȱH��-}V���{l�脗$� IBPE�  �� �h�������?~��A�6�(��8��)�[Қ��h��@�p�nclx&O�>�G۳<�s����7=��١me�k�p��1��Cr4�4zS@�v���h�S@��ܩ��C����hVנZ����h���A�<�`�2dO�G����@�)�y^�@���&��a����@�YMޔ�^�@��Z�R�$�.�)*����f�
'y�������D~��J P�$Q5B	pH0ȡa#"aZ��b)T(H�P�F�H�UG�v���6H�m�M��BCML2�rQۑ��Ia�NY�Z�H)֡�����{[6�v!�{P]��z���N3�8�X�X ��,nv��oF')��ek���ڬܶ���v4 ��u�5�t�=AYv��r�w�}�g�|۱n�j��ˬ $��K� mj�Uf����R�Lu%�b�<keu� ���xd v�����{|-v�Q	�	�ki�2u���A�Cqԝ<��E���H[�)�bR%�k'�U��[Қz�h����\9�0n&�o"��@��4���-�M ��4z\ě�x��D��;�S@��4+����@�.Vb�7HnF���oJhW��-}V�޲��em�I�I��4+����@�YMޔ�=�.�cP�Ns����-qmӋ����l��ƌ���/l�a}vh��hI��L��I#�-}V�޲��)�y^�@��𓸞$I#��Iw���ψ$�YĶ[M �l�-}V��ԉpo"�I��I!�[Қ��h��@�YM��,ڬM�؊0�r�X_�@DF~��kiȖ%�`�=��7ı,O}��m9ı,w^�Mı,K��vM�I\r�+�n�CD4C@�w�I��%�a�E������%�bX?���I��%�b_w��ӑ,K��Ƿo�ļX^��0�У��=�ݖ�z�m�A��۹�K�[�p,g��:����Kı=����Kİ}�zi7ı,K����r%�bX>��H�CD4CD}ա�|�K+jKc����Kİ}�zi7¨șĽ����r%�bX?�߮�q,K���#���h���S������[��f��q,KĽ�}��"X�%��ﮓq,|P�x _��7���6��bX���M&�X�%D>�5�4D����Yn�CD4C��ﮓq,K���ߦӑ,K��u��Kı/��kiȖ%�b>�'48�$��]#��{~�ND�,K�צ�q,K��w�ͧ"X�%��ﮓq,K������n��b��Ƥ���F��޻�p����\ñ�v-�A�ȋQX��zk���r%�bX?{^�Mı,K���6��bX�s��Mı,K�{~�N"!��śU���6�NUH�Kı=��i�~c�2%�����Kı?w��M�"X�%����b#�dDCD}:��J�ݕ�X��k6��bX����I��%�b{�o�iȖ%�`��zi7ı,Og{��!�!�{ۡJӎ��*l�M&�X�%��w~�ND�,K�k�I��%�b{=�fӑ,K
�D�E�E3p}�ni7�!�;���k�9emIl�U�q�X��צ�q,K��{�ͧ"X�%����I��%�bw�ߦӑ,F�h�5�kB��r$�D$'��*klu�oMG+s͌v���qs-[��	M�ꚷ5��M&�X�%�{��[ND�,K��]&�X�%��w~�ND�,F��۪���h��|5�4D���.���Z�r%�bX>���7��,O߽��iȖ%�b~��鉸�%�b_{��ӑ,K����[�3BbЄ�;+�b!�!�7{���"K���17ı,K�w��r%�bX>���7ı,N{Ի�nje��q[V�CD4CDj���CIbX��wٴ�Kİ}���n%�bX�����r%�bX=�5�֮[Mj-�j�&�X�%���}�ND�,K�����9ı,O����iȖ%�bzw^���bX�/2z���ۨ��^-�;2�V;r�}H�˷�\�<������}|���D;[���Mې�&��@<V�3w]b���9�lC`���p'c*�9�<s�i'n�y0vScTc��ۉ�It s��f����rt�m؃qԡ��=N|+H�I�Dݱi4��J㕷b�x�3���������<�t6L�:�F�:m�Wo`��:n7���Ϟ]R��ʔx�[���I1ڲ�z�\7!�#�<ꍫ5����� �D��bFUepV�Α���h�����H�CD�,O}��m9ı,ON��q,CD4F��f�CD4C@�n�+N:��.�\��n%�bX�����r%�bX��צ&�X�%���}�ND�!�vw]#���[\��-2�D���ND�,KӺ���Kı;��iȖ?� ��~�Mı!�>����!�!�>��odi7��%��F"!�#��لq�%��ﮓq,K�罿M�"X���uB1��~�"Q[5%�5���r%�bX>���7ı,?���߾6�D�,K���LMı,K���6��bX�'���\)+e�Fr���D�q�l���<��a���l����8Y�'f��u�eRb�}�X�%�ｿM�"X�%���zbn%�bX���ٴ�Kİ}���n#D4CDsu��#�K[t&�v�#��ı=;�LMÇXEQ$A	��P1�Mı=��iȖ%�`�=��Kı=����K�h��D�D�J�T#�'���m9ı,g}t��bX�'���6��bX�'�u鉸�%�Q�&�mJ�ݕ�Xr�0�"!�,g}t��bX�'=��m9ı,ON��q,K��w�ͧ"X�%@�n�+MJ�@�WH�CD4CI�{�6��bX�'�u鉸�%�bw;�fӑ,K��w�I��%�b<A �{�IJ"���V�M�ܡ�n�M��hʀ����wZ7o0��=��Bp�CЬ�p��������ı;��iȖ%�`�;��Kı9�o�iȖ%�b}�u��2�l���ʩ�h��h���f�<�DȖ����Kı>���ӑ,K��u��Kı/�=r��V�ԬK0�"!�gu�1�X�'=��m9ơ���?0��)�X��c\�&�"@`.It8�E"E!��iU�hҤ"@4ŉ�D��@� �� hŀFBB@�K�\LB\)�+�! BMhY�,c�m�Ɋh`D#HP"@�
�K�`�DBAB1�?Bt�:G�����@��RR� �
���!�a� N�֡#�:T!�P2$c��-�V�"rkHQ� ��ӂ��~T<�� ��V���G�/�!�.*1g�G"~��k�I��%�bl�zaD4CD4F�X�� ��(RL��]&�X�~`dO�~���Kİ{���&�X�%���}�ND�,�
 v�#����y�D�n�u���Kİ~��i7ı,?}�{�m>�bX��߮�q,K�罿M�"X�%��(=�n��q�.-"N⻱���֧=�Gt��-5qz��lu�v�;�Կ�t������ı,K�~���ND�,K��]&�X�%��{~��>��,K��l�1��N����-n��9m���bX�s��M�����j%�����M�"X�%����Mı,K���aD4CD4{t(�jT��AM��&�X�%��{~�ND�,K�{f�q,K��w�ͧ"X�%��ﮑ���h���wcq�D�1-	�F�,K���٤�Kı>��ٴ�Kİ{���n%�`T("n)ϕG{����ND�,K��ŮQS�[i�h��h��wsiȖ%�aP���pI��צ�$;�E@��uG��$R[;�\\��`ӷa.��v��wZ-����;e��^�*�9(u�UQ`�لj!�!�{���n%�bX�w���r%�bX?{��n%�bX�����r%�bX��Ǣ
��$����h��h����iȖ%�`��ޓq,KĿw��ӑ,K��w�I��%�b}�Yw�$�H��7U�aD4CD4۹HȖ%�bw���ӑ,K��w�I��%�b}�o�iȖ%�`�ھӫ�����U;i�h��h���#��İ{���n%�bX����Kh���w)�h��h�M]�mJZ���XrK0�"!�����h����ߦӑ,K���ޓq,K��>�iȖ%�by��й��V	h�=�U�r�h����hyz���!0l,���r�������������1I�{c<��U��N�jµ4��dW�$;&�E�pv����8+����]��g�l�{�m��w��:�V��;�`�����Px�>n�tZy��2[��w/V�wiɞ����5�Ś79��&n%�(���ɱl�J$��w�__q��ԉׯf�]��Vx�Wig�#�>nb㛶��P�h���ƪ�27!r�J
T�+�|�h��h���paD�,K�{f�q,K��>�iȖ%�`�;��Kı;��-�o�PĴ7eXG���
F"K��>�iȖ%�`�;��Kı9����Kı>&x�̘L�J*r�h�b!�!�>�wf�CD�,�}t��bX�'>��6��b4C@�������h���ײM���VɆ��ֳiȖ%�`�;��Kı9���iȖ%�`��l�n%�bX�ϻ��r%�bX��r��E0�33.�WI��%�bs�ߦӑ,K���٤�Kı=�w�iȖ%�P=��H�CD4CDs�w�!d�Z���c���g80lk�.�/0����6���g�CV
�[NJ$�H��6,��D4CD4���&�X�%���]�"X�%��ﮃ� �DȖ%������KĨ�~�;$X�J�h�b!�!�{�w�i�p@�DȖs��Mı,K�k��ND�,K�{f�q,Kh������-n��YmxG�X=���7ı,O}���9��j&����Mı,K��~ͧ"!��܉�$u�(qSl����ı9����Kİ~��i7ı,Ng��m9ı,�}t��a���N6�$��%��+�8�i,K�{f�q,Kļ���ӑ,K��w�I��%�bs�w�iȖ#D4G���c�6�"RQSq6��/�Gnm��a^�6�+�;�S.�&���3W����%9e�R8�h��h�N��CIbX=���7ı,O}���9ı,��Mı,K��޼����WUaA[�Y�>D4CD4��b!��,O}���9ı,��Mı,K��}�ND�,K�n�/�h�
�;+�b!�!�7��xGİ~��i7Ɗ?p���Q7�߽�ND�,K����q,Kh�w[y�Y�7BlY+�8�h�����٤�Kı=�wٴ�Kİ{���n%�bX��]��r%�b4v��;"�+iT��D4CD8��]��r%�bX~A׿]'"X�%������Kİ~��i7�!�9կ6U!n�婸ЮJ�Vtq1a���Q,v�v���M�7���9.�K �YmxG���t�D4K����ӑ,K���٤�K�#~�ׄq��=��MQ#�CEɧZ�]&�X�%���]�"X�%����I��%�b{�w�iȖ%�4gu�1��w^�|YZ�����r%�bX?{�4��bX�'��}v��bX�s��Mı,J�߯u�D4CD4G�=:�b1����kF�q,K����ӑ,K��w�I��%�b{�w�iȖ%��Df�b!�!�;��lrUiCYf�WiȖ%�`�;��Kı=����Kİ~��i7ı,Fϻ��!�!�_���a)-NUq���$��ۃ��s�g^v͠w-v����L�Hr� b
�;+�b!�!�7�w�iȖ%�`��l�n%�bX�ϻ��r%�bX=���7ı,Nw��ح�H��6,��D4CD4ۻ4��bX�'��}v��bX�s��Mı,K�k��ND�,K��́�#��J���D4CD4F�{�iȖ%�`�;��Kı=����Kİ~��i7ı,O�Ӵ�Bv�%�V,��#���h����bX�'��}v��bX����&�X�%���]�"X�%�{�a��݊
T�+�b!�!�7��xG"X�%����I��%�b{�w�iȖ%�`�;��Kı>�����\>��\'O:��1���9����ff�ϟ�;��l�t�x槓��g;#�_1��Ɍ۶�	`����<�X�m�;�!&�{7"Y6*�*'-��ch������A.s���u���=�������ݽ9�W�M��vu2�gWNJ�猖V��ą�$]-��<�m{j�hv��u��lv�֭# ;Rqu^�%ve[e���I"�p$���J�q@�i���t��ފ����r^��^vG+4�,]�5tGD�KCn��D4CD4��Mı,K�k��ND�,K��]&�X�%���]�"X�%����mlF ����H�CD4CDo׺�9ı,N��&�X�%���]�"X�%����I��%�bw��0��J�҂�\��!�!�:�u�n%�bX��]��r%�bX?{�4��bX�'���6��bX�'�%�0�)"�W�CD4CDo׺��D�,K�{f�q,K��}�fӑ,K�����n%�bX��7�K(�F�M�%xG���
F$�,K��}�ND�,K�;뉸�%�b{�w�iȖ%�bw:K����8�IY���ջNݛ^�>Xޫs٬�tGkn`8XHV"����ġ������X�%����ͧ"X�%�ٝ���Kı9�w�iȖ%�`��l�n%D4CD}:�����kB�m�aDX�%�ٝ���>)b�[a�_�ѐD�U<�4��&���v��bX����&�X�%����ͧ"X�%�}�a�D�Y��EVW�CD4CD}����"K��}�I��?�ș��߳iȖ%�b~���q,K��g|e+���Z��ݯ�!�!�w����,K��}�fӑ,K��w�I��%�b}�w�iȖ%�b}2���e�-�9m�R1���n�#��%�bzg}q7ı,O����9ı,w�4��bX�'>Ծ���Z���˼����;�����rb���2�sIˋ�h6|N�g��~�[�D�,��5���,K���{��r%�bX>�i7ı,N���m9��Pt'4@����Y\#,K����Ӑ���r&D�{��&�X�%����ٴ�Kı=3���h��h�����vQЛ�M]�"X�%���f�q,K��}�fӑ,t� 
j&�zg�q7İ������8�h��h��n4�ve�j�h�n%�bX�Ͻ��r%�bX���\Mı,K�k��ND�,C@�w#����hN������m9ı,OL�&�X�%����]�"X�%���f�q,K�;>ݘG�� �c��V�t���.=lY)��DY��/4r˫H���3ʰ��K�Jk�\����{��7�����]�"X�%���f�q,K��}�fӑ,K�����n%�bX�uwba>	(��hNʰ�"!���Mı,K����ND�,K��]&�X�%����M�"X�%��DSb
(-�9m�R1��Ͻ��r%�bX>���7����;�^�v��bX��~٤�Kı7����F�u���f�CD4C@�;��Kı>����Kİ}�l�n%�`CDC�ի�Rn'��ܘG��oRs�!$��]&�X�%����]�"X�%����߸i9ı,Og~ͧ"X�%���F"!�#���lBCT�pY{]1����Ԟ�����l��s��v-�k�݇f��66�+�����RW�>D4CD4���&�X�%����ͧ"X�%�����?��MD�,Ok���r%�bX�;��i�썥[�R1��;�{ٴ�?1ș����t��bX�'k߮ӑ,K��}�I�����!�S[��IkB4���#���h�'��q7ı,O����9��C"d���I��%�b{;��m9�h����JP۲5C��[��1�~H����iȖ%�`���Mı,K����ND�,�2'�~��D4CD4Gڷ�0�tJԴ&�xG"X�%���f�q,K��}����O�X�%��g�\Mı,K�k��ND�,K!�Y�� ā)�X�  D+�(J°��W��� :�e������H�H�:�8C �� ���,��a��h�6�F0bD%eGP�)�1M@��}��} @�a�0@�A�D" T�*J�"F���x$��(�T��(�$`A�a��f�eSD� � @��0 H���
sa+��1�p��jTGE�BW�@��H� �)$B m٧KWh�Z]0X�F�dMl�Br�s`p!e.�KR�HB1R�Љe1wr�-�Im�Ԓ�T�pB�r��n9su6�I9��RxX�b��$���Ӯ�p�]�*��J��U��mX�r��c��=��G��S/[��zq��ٌ�]0�g�c�u���wbL=������5��2*���<�UUR�J�RI�1�v�&xp)qBų�Z�J���z[�NBݔ��m�$,0 �6��K-��<��7M�O��m�&��u��9�F�-�"b�mW�3=a:��+���1\t-8�����G[�dL`8;��"��+������ٍ�5�x�^�����c�F�@l��R�v���;tb
'4�u����՗v`�..%\�E�Vު��A���7,�f.��P��:j���{u����qs�:-*8�Y��cV8-��D� ��="l��`�F|�v�����A2;��乄�� ���mHS�.e�9�Bݵ�5�8j�;rX���NU:nxL��;ðg���\�( U�m+s�q�FLu��q�B�ă�GF���,��؛	�*�{[c.U浜&�u�j�L�u��UW �e��GDc�V(���Q��Z@���[Q���T�	x����"��3��+�Tt'���۲H�%S�o��g��/Ţe�e��J����&��l⒀�+0�lq�EY.6�A;;�y
r����^^w�m�ӵ=y�n/4��1����h�ݶ۶q;T��sZ���R��a���e�hVz����wd8���qwD�)r�����������T�Bz�e�]9��щvC��O� %�v��@s�O[z�1��m�e�TT�.��|W"�+m�UTQ/�p5UU�F���m˶���%V��F����5���#=6Dí���b��i�R�ۍ�"P��k�(��r��6�98X��I5�q\�(4��\�l�\u�88��M9-5�F����: �[u���@��J�k8��`�5m�r��V�Mj(��n$�!!�;~>o%QʪQ+Ui���x�[��X+�6��$�$��jv����OV�6�d���g۫�&M��j� �@-Aj,��a��Zۜ!�s-�sٞ���{���p+����3�%ɣZ�E�V�ze;6��u䛪��$N���� �=n9om:�[,f�\����T6�e5�M�vӥMr;��;+�Eʿ�H����*��e��}�w�߁,s9�Z�b��R%Z�e����[Doq��hq5��x����-�sE���UN[m�Ȇ�h����ߦ�CD4�'�w�q,K��u�]���L�bX?��f�q,K��������5uL�V��Y��Kı=3�����溉��'��~��ND�,K����&�X�%����ͧ"~L��,Oe����CZ�)ep�D4CD4G��Ȗ%�`��٤�K��i�������ͧ"X�%��3����Kı>ﯣ��ځЛJ��"!�{�4��bX�'��{6��bX�'�w�q,K��u�]�"X�%��]e�\�֬a��v�F"!�#g۳iȖ%�bzg}q7ı,Ow]��r%�bX>�i7ı,N�Rz�֦ۋk��6ûs��6Ѵy��6���HD/K͍��gZ9�c�;cN�A��w"X�%�����Kı=�w�iȖ%�`��٤�Kı=�{ٴ�!�!�7�B�F�QeLJܮ��%�b{��Ӑ��!�;�����Mı,K���6��bX�'�w�q?� 2�D�>���a�˗Fj�֋n�v��bX��~٤�Kı=�{ٴ�Kı=3����bX�'����9ı,O�����R���-��F"!�#g۳�!�,K�;뉸�%�b{��ӑ,K�2�~��Kı=�k�~�6�u��n�f�CD4C@��F"X�%��뾻ND�,K���&�X�%����ͧ"X�%��2�ْ�z�7\�\��fē��e{nŅۋ ma��pX0.��y^rn��pm]�T���o%�b}�w�iȖ%�`��٤�Kı;�{ٰ���İg�]&����ܮZ�P:uI^Ȗ%�`��٤�Kı;�{ٴ�Kı=3����bX�'����9� FDD4�����El6�nѤ�Kı?g~ͧ"X�%�����K�JX����v��bX����
F"!�!��whN�%��k.kiȖ%�bzg}q7ı,Ow]��r%�bX>�i7İ"h��v����#{4)Dn��T�չ��H$�߾�pI��Ѥ�Kı=��ͧ"X�%�����K��ov&-BKC�Wjb�[���q�N,q��u���������ς��Ob��5�sZ-����Kİ}�l�n%�bX����ӑ,K�����n%�Q��ׄq��kNͲ@�u�S��E#��n���1"X��{���Kı;�^�v��bX���M���TȖ'��'�I���N���G��7����ı>����K���{��&�X�%����ͧ"X�%�ܳ�/�LiZ�)ep�D4C^ DwپxND�,K��l�n%�bX����ӑ,K��H�,�@�H�"��!�, �C�n'��ܸ��bX�'�z���̵6�t&꒼#���h����
F"X�%��#�w���}ı,O�=��n%�bX�{]��r%�bX�����9(8�5DGv0\[Z�l�F4��Xn.����7n�����o�:ٱ���'"X�%����ٴ�Kı=3����bX�'��}v��2%�`���R1��GV���[�+nk6��bX�'�w�p����j%���~��ND�,K�����q,K�;>ݘG���h�o�)Dn��jS5nj�n%�bX���~�ND�,K�צ�q,K��}�fӑ,K�5N�b!�!�9޷�H㢊�XKsWiȖ%�`����n%�bX�Ͻ��r%�bX>���7ı,#�ׄq��kNͲAV�Vf�sWI��%�b_}�kiȖ%�`�=��Kı=����Kİ;7]#��պ�RF�uc��i���S��l�����9L��w�7}-��n��5Yќ@�ݞ竞۸�q�m�ǭ�c�쐴�\��h��;Gmƺ�.��듎�n�Aj-�Y�g�����,�ul�l
��c���Hd���4��ۛp��gnƹ����ٸp���n��k��WRQ��c�܋=pض�����'#��`�}�{�r|m���/=k�����v����n;���Pt�'��8�fPv��N�C�mj��v%�bX�L���n%�bX��]��r%�bX>�z�?�aȚ�bX��}�[ND�,K��g��F�I��F"!�#~�ׄq��,����n%�bX��}�[ND�,K�=뉸�%�b{ݷזYZnBn�+�8�h��h۪���%�bw=�fӑ,K���z�n%�bX�����Kİ{�a�iZ�R�J�j�b!�!�;7�0�D�,K�=뉸�%�bw��ӑ,K�����Kı;���ԎQe�Ҷ�0�"!�#T�p��bX�'��}v��bX���M&�X�%���}�ND�,K�{^�jc�we��!͍�0]m��:z�������۲V\�E�7d����00���bX�'}���9ı,{^�Mı,K���6��bX�'�{�p��h����m�\��E�nW�q%�bX>��4��")��,N���m9ı,OL��&�X�%����]�"~C*dK�����-2�WV�%�UH�CD4CD?���G�,OL��&�X�%�ߵ�]�"X�!�wn�F"!�#{��M���$��p�"!� ""y�����i,O�k߮ӑ,K�����K�4C��ۄq��?v�$�J��]f����%�bs��ӑ,K�����Kı/~ﵴ�KĦ*���Ҧ��A,x, !<��8���ƭ��Mg[2�vM�Y�t8���N[@f6Ҙ%����S@��zWj�-}V��R!a0�$I����L���p�}8�l��M
L�FcA$q�]�@���7�31���l���zנwtpj'�`�1ĜZ���S@��^�ٟ���>�h�%���#�a�@�e4
�k�:�V�y�Z�"Ru�8+
�x�Z�vi�n{,�g���^xҦE�E��j�,�8g�W--��o�������h���l��{���Ƃ(�(B94�ՠr�W�u�������E���M�8�^���S@?^�@�mz�k�#llja#M8��S@?^�@�mz��L��H�ϻ�[�ګj�P�ǉRC@?^�@�mz/uzn�X�� ����z� �K\jD�U9����:wO	��]$��'L�6z]�FtN��hNO�_��-�������@;���"'�`�2D��*�W�u��}�h��~�Ď�b\�fn&��Y5u�>�� �:"��z˾�������p�LnF��f����^��l��{��H6D�B(��9[^��ֽ[�`�]��(��ܙZ�nj�r_w<��>�.����i��wd��!��L�8Ds����q)��z�u��҆��q�w1�m��l�r�{=cÂA[Z�^�G[9����Eٺ�Y�ݪ��[g�LsoCu�n5�#(M,�np��Y�=��zN-�/+��C&��ν�t�z{<���nD�*��ntS#��Uz{����2A�]�������-��M�j_�I�ǁ�K fEjV:��',�9��3�����f�����J�7���,��q�8��ߞ���h�Y�r���:�n6����F�q�l��|�ߡ/�{��;�X�,v]L�&<h"�{��9[^�W�z[)�r<s�'"rC'&����
�k�-��{����tI�H�H�z^���M ��`[u�r�P��<M��f����l���d��v�P���Z퇧O� ]B�,\�O"Q�q��N?�}���@/u�VנU�^���r'"pm��u�I	A�"a%#��`~n��S@��c�aO�6��9[^�W�z[)����F*(?�����z^��l��_u�+n=��]$m�$i����h�Y�r���*�W�y{�6���k�n�鎐��X|���v�j�]��5�O�y���b(#�M��<�E[��t���6[j�?k�$�!%�A�_G�	Ɯ�ƃq��n-�uz��h{�����('��(��U�9�]`k�a�TC�IdZD$�) i մ��ĘԈ֦;E��dS�$�����-$��[P�1T*�C
�)P���T�	�1�Č!�1�R�KZ5�L��� ��FDd$����!"HH"E��X�$�"�2�*�.$�	`S��V�lP��G�.���m �(�)� ��h )����|�	��ky�n䞿{�nI���5F�`Fd�@W�hV�z+���G����7r7��.����z|�_�Ɓ���~�q�tw':�팴f���[�7�/p��pⳇ��]�)9!��a�SDg�\qh]n=���u��:��� �`�`�`����J~��u�jk\ћyg�~͈<����}���A���ߵ��b �`�`�`��k���A�llZ�k~�@����n9f��������b �`�`�`������A���9��k���y����6 �666=�������F�љ-���yg�~͈<����}�ߋ��A�A�A�A�~��؃� � �(Q 2=���6 �666>�;}���uu��-�Z��lA�lll{�~�]�<�������f�A��������A���ߵ��b �`�`�`���ϸ�~�8���e�ŷ.Q��(E�ܚ���݂uї���������VN�u��v �666>����y���y~��M�<����}�ߋ��A�A�A� �-�O���W��0 ����y~��M�<����s߿��A�A�A�A�~��؃� � � � �������f���ֳZ6 �666?��~�y�~3b �`�`�`��;�ٱ�A�A�A�A�~��A�A�A��]PzI���Gj�@<@�\l_�d}����lA�lllg���؃� � � � �߿p؃� � � � ����lA�lllw�ɇ�aL�Z�WXj�؃� � � � �?{�lA�lllP�b��|lA�666?��o�lA�lll{���͈<����6 ��`������?i87Wawv����n5s��d͜%�±Ș *΢u�RUqmlp,�8B6��c6a\\��r��S����i��cI��qύG�,i����9���8��7a�\��Zn�k�+�rv�9�DL���w������t]=�Z;E�x'��'��/�i��H�VX�͹�sQ�������,��c�D��:ے@��H ����8�!������u��C-۵��d����,�[�{j��M�<�ځ��w{�w��߿�p؃� � � � ����lA�lllo�~�kb �`�`�`����ٱ�A�A�A�A��[�~5��0�r[5u�6 �666>����y�߿؃� � � � �?{�lA�lll~����A�� �b]{<���eA��v�� � � � �߿~5��A�A�A�A�~��؃� � � � �����<�������f�A�����x����je5L5u�[y��~͈<�����߿p�	G�"!L�y�`wr����e*����A8�m��9^�@-�&���zX[���"�M1�cj��$Ƅ��q
����l-ާ��b�J�=���6�rf���zm�4W��-�s@�<�6�������mW���
G�Vy�`������|���� �s&����m��9[^�[nMו͒H'�E��5#��V��+k��� ���^��$jcɉ��f��ڴ�rh��@��h}�*_50���q�|n�6�۳�v͸Ə0)����q�jܻ���-�M��k7["�I'����>�r���)�uv���Ǖ<��E&M����M�Z��rh�*���h�"M��@��i'o}���;T�!D(₅6�ɠ~]����,1���HӍ�@��^�[nM��z�S@�>*�DS�7#�@-�&���z�S@�z�g��]SŌ@�<FV�;����Ep��b��,�Y�X\�:漯4�j'�� �s'�?+���f�m�� ww+�7��.��M"��D�q��M���r}��U������#b���I!�u}V�[nM���l���=����G�$�@-�&���z�SC�2
�A �wٽ��=~'p�9!��Y�4W��-��W�h���/4�+�JD�5!�(̷�`qs���6��N͎����x)�6)�	���25�R=�)�u}V�[nO��
��=ݟ}��q9�I�Šu}V�[nM���]�@�>hU��S�6�@-�&���z���:��@�T�b�E��x�.��`��8��`t)���x|}�G1�0�&�z�S@�� m�x��XB����%	!BB@� ث؃���6,���'��ة��]�ƕ��
�Nd�F�u-���'F�g։���x�����ž��N��ɶh�`娍9]i��pĩ`�)�qǟ ��cJ����,�n�8.�'q/Vv2�.��\cC�����lN}R\���l���[��u\�Pd�S5 ,R�r[�R���'�R�&M��e�S��y��\�A���=�}�_7&��AӶ�calM u�u�ad�OYm���
�,��q��>.���;4�[ N�� 6ڼe��l�6C��	���J�jĒ��?��e>�V�{ذ{l�J&C�G4�]���X���4
��=�w4����W�~nZ����\Z��wX=�ߖ ��N 6ڼI)uϫ �W�lx�N1�G�L�9^�@-�&���z�S@�5R��$h���$��w`��Cdg��tz��֋.S�9�W����b�-ikiD�7�nG����+��ݳ�I/�����ºiLLڄuWe]n�� �@ 	ݸ`:�8 �j�DDɼr�����UQ�6��>���z��@-�&��ֽ��!rFLq���g��-�`wr�g���!Owg�:�0S#JH� ���mɠ�������|`=�`��t:�U7jj���.�,p���v<V�n�u�,t�Ǟ�E�z��j+��Ff�x-r)k@��^$��ޘ��)�z���[nM���7@Ȭ&�˫��l�S&�wN ww+�<�kߒ=����$c��7#�����w$���ksh ��U�ݻ���?}���-b9�4�S�$ZS=������l��
wo�pGp7���$qG2h^���M�v��n=�Um�xf��jG�f�ǅ�TS�:��j����Є�r���j����&�6���}>4yڴ�rh�l�;����P��6Ƃ���>�����*���yV 7�^ ۔�<�s�S"JH� r'�U� }�w�(���� ݮ���'fZ�����uJ�n�`r�3��xw_�Ss�q
>j�y������j��m+���v���v���z��8��u�~�[7N�*�SJ�U%{7,���ñ]�yƛ�=�=n-Ҽd]���2f��c���ԍH�yzנZ�Š}?7]	G��0�$tt�M��R���� n�S��&M���������[��s��v�U��Cč���l��"!)�������շl���v���If%�� !���x�wN �6��DN��V �L]vE	�bA�@���@�ۏ@������ q�K�P� ��=��&2#%v`V��HH������R�(�`Ji
IP�&�C���E�Wb��1a�
K�n
ؐLSJ�٬�`#�"r�a��m(d`AM���1D0���L�%!9�D�	�2,'�&i	��cb��9�M���*�yk!!��T���@ $`��D/n꺀��ʧ%`�U���f"-.�JΔ�'f�0����Qs���[�Uy�ɓi
VBlb}�R��k�)�:ɶ��D���Oa{/7E O`[O�t)�.�;ฐ��Zp[m���v��Y���86=mٴ�5��ր��a��4gl�×���jg���+WQ�( mi6�������	ٶʷ��]��Bul;E)��;3�Ê�P
�Ӗ�h��8N��g=�N�f3��MVy'�À�֍����+��J�Lѩȹ�����n4Yfv�n1�N���n����iq��K:{^!�c5������-vư�bI^���r1M���8�sb�+�VB�dq����l\�]��]���1Nfµu.�OF���A��&3(�A�k��n�kI�QYo]N;D�4�,���H�i���8��<�Ը<m�S�{�k��"����[[f©CJ�O;]��s��t��oI.V�i3���	�<v8��PS����g(eT��ٵ�:�n�@�s�{x�'f�8]�t�E��
aΡ@"Q�r3�v�i͎��0=�ʨ
s/lcVW�s�6�mٶ����x.n�������
Okɵ��:3����s
��:�5vM�ŵ�4�[!Vհ��k��5�+;�gg�-)�*v)3v.�q�=�Ov��Uԛ�\ۙ.!rE��V3��f�=7��X�+��խ�\���W1�&V�!s<�wWLv'�r��H!�'A�]a���YPNk�컵&�!:I맦8 [RM|$�U��m����Pؕ��,�m'S�5�D�8�l �UN��sN.m�Ί�d9���'�R�k�ԁF�.Xn��TZd�X��l�^U������HZDb`�.r���C�9��k:��b!&����KbU��4��kY�m�]���]@t�V�-�r�,�6��-�
$�6��`)`�*�Z�Z��k{v*tT��8�"(hP:��Wg�<�XN�f����c��ʌ�d6��S��W(��Y�[�·9���� ��oY��й�ٻ��7����ƈMRK�ѡQ��s�ۃAʁK�p��//\Џb����<ӵ��\s�&�s=�����A�.�\��mt�y�$��5t����%��cG=Yç[����*@[��g�693m�lP���4��̓�-�V9E�F�H8c��Y�����d�7l�km���	+��jNJľ �sd���$x�9���o��/Z�]�� �4���<I/u'�xZ�V�,��hz��z�S@���@�ۏ~���'�甆!Z��L�Ywu�wu�}�:�
���/Z��˗cRc���SwV`r�������`O��$��}��3gȉE10�E�UmǠ��@��h�h���6l�m�.�<�Ź���չ�k����88�(�����=��ӥ��m��[4l���;V�U��Ա�uȭ	Y$��In�Մb ��AF!Ge��t�=ܫ >���L����X�FE	$4���@�ۏO�Gw�M��s@�/rʉ�%$x�9�@�ۏ@=�f�m��=�j��\;�&�!��"�&���^�m��=�j�mɠ����(cM�2�y�'�a�@Y:�S�������P�;D!%?�$z�S@���@-�_��薽��bK�?~�S�KUWd���>����)���W�l�u`�fk1.�Q(�&��zm�4/{ٸ���h�
D`E� ��[f�.���S�����B8�Z�N��V������`m��:�:�H���F�n=�)�yzנۓ@���@���m�&<2e�$+HϫJ�&�y#r÷Vr�[qݡ?���
Ĥ_��,��G��$��;��- �ܚ��z�S@��Y�D)$āȜZm�4/uz�S@��Im/�6xX�V�,�Wh��׾��v�:?��Ͻ��{�W�}�"5�E�O�G�m��<��@-�����"P�xl߿~��=���'!28�n8hVנۓ@�ֽ�)�}��������MG�{\�nm�D@��,����g@=<s������)�LP���n? ����M�Z�l���mzw)���_�L!��W�l�u���������.}�V }��d�/��q$4�<�nG�[e0��Xz"d��W�9}Հn���d䌊<l	$4+k�mɠr�k�)��� >�a�R�&��L���� 6ڼg[��l�>��`У��z���[uf7D�-�5���t.vs�X���<l�6*��M*�OVʵuYs7���U�yv�m���ܼG!!�U�;�n5�C���餮Ka.2[r"{8L��f�Kf��\<�M9Ȝ�cҾ5f��d�����i9v�;�����l�◧��s�er�d+��姂�ۜh����q9�r��(Ol@���g���+��K�w����w�����#Y�⛔H���=��Ein�{pJ]��Kr��FL�U�c#p���/h�W�K��l�>��{��������^FHZ��L�Yuu�6�䒙6{����^���y(����U/���⍸�r�[nM;��#�pl��pqɦ,x��i�D(��m�xK��l�>��`�t9�@�v�-��Eė_wf$�@"!.��?��Հ�� �G&�9.�Z[]����hUb��.w��v�Nn��3��ѹnGȔ�7�`F�r=�)�}-����z�%����z��M�����6��Չ/����A&E�m��?N�Xnٝ	D(���I��VDG$āD��>_}�=�Z�l���mz@��q4�$27�)1�t$�!K��Xw_�۬�mV�@ԔD"ħ�#�@��hg�B����t�r�g[��5ˉ����a7���.�Kڱ��&�J�Ji,m�h���'Ƥ�()"�m����-�Xη\����w_OԺTxB!�#q�[q��נ[c0��Y�I%�G>�UG�"I�B���V���`�f�RP����������n�L� ��nJ��IB���0���mV�)t�����d��A��$��<��@�(���ʿ ��V ۶`W�s7Ԝ�>�ѕ�2�t�������r��;I$���Eͷ-�WN��M\�����ʰ�n�ݳ�B��=�X�Z��M6I���JLz.�����::���6{��-�YВ��%T6w��&�˕3qe���z�`Kn�
���]k�?{�Q�&% �qف��v�����U�l�u��(���P�{��ܓ�����XMe�U7*ꮰ-�XBJ��_����@�Ѯ��f)DiL�6I�J�2 �n�`�[�Y�kpN�ɗ5�W��ϙ7�$�$qG2h�נ[e4+k���GK���ė�~x�	HY�� ۶`Kn����:�g��P�	H��~yJ�(��J�V$�}�V 6ڼ<�\���;�����Z �Ym��b_� ����q%��V ۶`y%;]�X�n�ȩ�.՗T���x���
!yD(���x�>�� m^�Q	~!%�53<R����vwǌ�˦��\�	vn$�pJ��V�v5����KӤ]u�2rY'76�%6�>mn�[�cu�-�1�۰uڰ�Սԍ)�-ݻ,roiN�NuWNp��.k9�䗉�Q֮�!��d��,2Vb6NwX8C�6˻�]A)kr�m�ωԮ�ڲ����Y��pu�(�J�m�^���X|j�MZR�p���{�k���d���{b#.���;�[��y���iq�;��9��!��F:�S7]]h�l�>��`m��@Ɩ���$��<�;hn�$�U�6�<�Jd;���_u`�fy(�P�N��#��S4�nl�����z.���M �[4��Kqᄘd�(�M˭z�ՠ�f��H�����E����
�,�I^�k��[4޹4.�������k�j���l�=g͕s.׍�Y������z��n� \���5��{����y�g�7�<��= ��M˺���h�.0��"I&4
7�[�&�?0Q�T@�
��u���������pӭ�y(Q2&�.������sv� 5���l��")���V ww+�7�SFI*՗*fһ���l�?N�X�ڬ$�(�*����:���<�I1)ێ�ֽ����W�6[��v��o'O+ک��	=�kn���j�{q�K�N��O��"��@3*��� �W�V7��,�#��yV���v���u�o�-�Rv�uj��u�tD$����� |�� m^��-�ͩ.�hW#�Y�-ݺ�%��ً�
H�G��D$!F@X4��4���e-] �J�P�Z��P�H�!H˗u��$I$�L��b�c	��`7Rt��f Rl�*�F1F��(MКh��*��������!DP,E"���^���Q�"��|$h��+�8 ��_zw��M˭z��\dx�G	$4<������ެ ���xӺ� m�0�\y��@-�&����N��_�z�`�[������Ŭ��q�v;	�VC��]Z�7�C�NɌs�k�nr�S)fN7WMv��E9�N��l����(�� ww+�/>�BY2bS�G�[e4�[0���N��Q
d�Wv\�\�w`�J54�呂[nM �u��ـ9�9���EҲj��S=������ݳ"%1	8J!DUz�4��x�����ɠywZ��� ?kw��� �%��s�M�Ĝ��mzS��V�|i���C"a2u��ms�)5����V�����:sk�o���ޜ ��� 6ڼ��u�~�r2X��,
$���Is��<-��{�+~z�ՠ{��*DIUUw��� �w]a�
g��� ��1$��У�[P�]��_�1
'i����� �:�`y$����W�^/Ƥ%�!%?�$z���?�ؾ��_�;�+�>��X$��߉�&�un���磞�"��.���c*��j�X�[���lF�n������ɧnƎGk�-pd4�����Q�"gvq�n���d���=�\�ptM��\{lq����ջ������ծ×�N�=���+g[�6�=���Xyp��2u�=q�u¤7V��U�kn:5�`讔�cZ��L���嵎u=�ڰy��<�[�k�[u��3�����'lι�:n���l����Kgn�����O�����
D�I��9}��= ��M˺���u>������E�\�� 7�^����s�~�n��B�^Q
�;�┞T�U�����W�9��`ֹ�<���_�;�+�?=Eӫ��U�ꦪ��=
B��}8��� ֯ ��@��VkS#�28�`G"�?-n�/%	BU�{���w� n������C���ϐm�� �u���Q�^�ns��m��]�L�+�q{1F�gPMda���rh]���V��u�u&���`�r+j@��^q���pLc����R~P޹o����[m__�ԒJ��?~I"�t�Bɐk�U�Lm�����m���n7�H �#���󍷯��1��~[��XⲤꮶ�|�m���q�����6�^�	�� I��y���>j�\p7]NYq�����6����m�m��8�i�k��I{��NģI,�6Lm�jL]f���Z��w2�c�1��䋭ؠ��0.��{gBV�ݢ󍶻���m���|�m���  rF�����ٵ��I�(�ۙ5$��j��$��dԒJ��y��]��s��7�w�r:,���
$�������m���/8�k��.$��Z�~I/&���Ȕ����nI��2O{��m������n��� �7޷m�w`�x*�V�,�Wh��m����ov�q�����m���6߈?P�ߔ���.K$��t�l�����R�}v����ؔ�w������ʶ�UXn���|�o�����m��ۍ�����m�����o���H쪸,��_8�m�v��I��xNq����&6�����~ H�?4�*�7lpGXv[1���{�s���w��[w������|椒�媥�Ld�Q9��׻�cm���|�m���㷀b?�$,�"��	����'8�{:��������IE��}ۺ����H{ޗ���{��i"۹5$���Z�mxC���#�}[B�,c��Xe6:�Ѹ�П˦�+����Ю��r��m���K���7tNq����������~��>q����Ή(��j�&�5$�;n?ߒH��MI%�Z�q��M�3�M���m/�� �Q�Ԓ>��ɩ$�ӍԒ���Ԓ�������D�Jd"ħ��f��ڴ��`-�X�B��ߖ�{�&�j�8D�)����V�z[w4vn�I` �{5���r��u�T�����#\9��{/H�tALB2pb����ۮ4*�J����k�I<
 �,s[��:��h+��$�F�gr'5)�݅�Yڃ���}N�֞�tu����t�{0E�c�ZmJ5��A$��9�zh�g9j1;7m'T幞��t\j�b�3Z�!϶�a���l��s�mYX�jBE�ب,�S).��>'����3��s�y��uA%fZ��0�y�.:v�۞e�b��������g�~
G�8�˾��m��Wj�*����:�G�O�D�s�m��Wl�[u�l��gD(�����]a!*���UUU��>��n��Q
e�>��v,��1�j�]���������
W_{Հt��XͼX�np�}fF�5#�h1)����[u`��6u��<���(�*KSR�8�����$�']�dc��Gǘ�-�ܾ�أ7+j������*�>Io�߰`]�@�ֽ�����*ĂdU��щ.��yG@�A"���y}��@�n����VH�"yIH�Vנr�����Wj�;���dr;c�XҲ�K��	3����;��,]78�N�yX���Uw%�AwUuWXm��<�DyB��g�?���X�n���r�
�w5St"��H��s�q�vwb�6/gtِ��8�6N5tnGe�G&D,<��i�3@��Z+k�9[^�����꿵̋$���9s�k��9D(S#���������Ȝ��r�@�mz{�ٹ���T!�(�U�	'DO���?s�g�.�g���
rGc�Ƈ"��q�m��:�V�k�h��@��p*!����X�npB���!$���O�t�ެ[x��5ˉ���S(TM\�Ym�H�OV�x�>��W��:��z�s�u��Юɹp#��)��ڴ��@�n��q���Ė��VzG��%�W,��� ��,�78�n�ДB�����9�$G�h���.�s��D)�=�XϺ���j��,y��nf���h��@:�4�  8AU�
�����������]dx�j �Ԑ�9[^�u�hm��:�M�u5$����5�"�6%jKOV�mmָ�l����&�I]�j��*�e�#����h1G���M���[l�J"_��u`����RU��T����?���/�>�� �m� kn���2n��:IE�.T�E���t��9[^�w[4m��=���=��.��������{�� ���`yBP�N�g>&n��h��&�O���f�m�����m�$ê��|�<������V�ٱ�P�t!@t � qdA-� �21�13%�Amp�@`�KkB�I�O��<&x hIHS�����
=zq@��^ֵ�kU��I+��굁�M�-ee�ʷۧVv�k]�jJ�<�^��J�:丹���V�p�
�n\��Z� �M���gt�]`מ{�8��q�.z{n�A�Wi�aÉRJg#�$굲Alҷf�M���y��h5� m����ֺN��y�lq�щ��E��gfۥ�����U\��a ��Bte��bbw0�g�%�Z�z6E�id��;5K���y`���.M]tv'։:[g/g*1��cS$�:�y�4�O�l.�Cj�M��륅TN{��Or�%�u��t��>��y��7mƑFQz�Yl��͜��F��=��0m�"l��x�T�e��/�&��S�&�>N���YvRs����ӦG�ӕ�r<�w<��2��C+��k8�{`�6�w )���ۇ:h�i�F�V'�C>,��ul!Ņͻ<1<hd��eknN�]�eYp�"c\���#ۃ\K�A���A���R<�W�8��X��vS���;;�j��(��bq�SiI';Zű�>�=y�C��;N���j����=��:G<2@�j�JzՈ�8��#�Y�N4��a����㦊6+��{8��vlE!��_:�����I��ٺy�U�pV�am���(:�؞2�ewQ�rWU��6dǮu�N	3͔�gigbI+I����dK��+��!v�7=uz|�hl����T�腧�ټ���V�pX��`��;+� ).w ��4i�u�L��gm�EQ��v$��� 6�^�%@]p;�WH��Ƽ�N���&j�h\F��{nRZ�WU��b� �ó�7���W����M�v���+�\��m���� z�X��j�`ñ# &ˬ�î���×f�6V+Z٠e�����@)�JVE�uZ��v@�"�i�8+�-�'U�2 M�D��a�;a�/3k�7E���΀$j�����F�Ԓ5���*�clE��V0�mYp�h��
���6�m �D�&�8'UJ�����S�"簿������$;v���^�ukZ��v+�U�'m�t[U���<&u���v����&ƇqP�ͳ�cr��j{yb�kl�ln���@��)w��awIu��CZx�G���<�<�jCq3�l���N��մ�^�E�aczc\tb(N��t7H�����n^@C���燗�L�Ba���K�:y[�=4K�DL�{�{��#�)��kKm�ԗI����V��γ�������:{��{EJ<M2a#�I4�j����"#�"!%���� ������&�nf�yڴ
��@/[4��� _w|�:��[IF�����Հ[���`i��7�v��SWuV�AM����>��;��`i���P���� 8-qR���Poܚ��h��@�������G�?G��l���@���]�:w;:�b磓ۧl����Gn[Ic���t���!j˙�V]��:� m���ߠ�G^���Z;�hLK*��,n׀�y���2[��o ����D%2s9J���*�SJ�uw��� ����hu�@��J<M!��%$�/[��^v����}�ى}~�h�ֱ�,��cLM���\�u���� ��X���q��[X�m����u�>�;�:�v��P\s�O���z�R`.�)�������~�Ʃ&�1i'������ ��^���p�O��jI&4��@/[4m��/;V�U��������X�i⎮���=���I4��H">IK�!@�F2ֵe�@-�4x�0��S���78�m� =n�=
!Ko8���c{�8�7�4�Z�mzz٠wt��yڴ�
���E�g��56,�Fs��ƭ���4�V��tr��6XvY�qS��c���&Ǡ��wJh��@���@�]�[o�Q�&��Қ�j�?.���f��^m� _�!�1�!�^v���^�DD)��u���~�^MX��Wut��.�� �:�`�� �vـ��
"�H�+��Ė�)�krJ-���	ȴ��@�t��yڴ��Z�7�~9ܽp�.���\p&�@n�4qβOVC���n6�ظl;�snƺ�4�7&���M�h�ڴ��@�&4�3"J6�^v��=_�, ��x۶��IDD)����VYJ��J�n� ��t���J�3�ύ���h��<U���FĤZ ���>ݶ`i���~w�8R��4�a�5$�=�)�^v���s�[�R�V�J#�F��&�(N8�q�p9n�[�����enc��e���u7nC:-<��,]�A��۶ݟ�����M�W,�����O.�Xl��ݽS���+V9�vޞ����v�k3�W�Hr=n.'�;q���4��=b�=�t��ve�<���RiN�j-�s�7[jeX á��x� 䣑.�����\L�l�p��T�@�2�P
�N�On&�ו;u��m�Q�;j����:ѵZ,E]dq̻�LIHp|��@��ՠ����4�������k#�h�ڴ��@�t��yڴQ�ɍ�	#Ƃ����@�t��yڴ˭z@��pi��,��M�Қ��h�ڴ�٠w�p*i�fD)�ӆ�y�Z�v� ��h��?v�X���C%3D�I��0�
�75���Xsi;����q��[Uv�C�<����qh�j��f��Қ��h���WQ#i)�_[5dB��JL(Qvkw��ֹ�7�np�|V��jI�z���y�Z/Z��٠~�r�f<P�LIHh�U���@/��wJh��א$��,�Š��}l�-�M����li���I16��콫�R�um9���t����J]٧Qu��4���rǍa��}l�-�M��޳@(w%A�!$G�G&�oJh��@-�4��@�5؊�a1�
4�^v� ���h�P�I,��n��ـ~ծ�.�<Q�X�ģ����z]k�:���z�h����1E1<���Z]k�:���z�h_U�~^]b�w=��1iɍF�E�k�棎5�gs���	٫���p�&˩�d֎KO�o��Jh�����ZVנ~�9��G�B	�)�)��uP
��R]�u_� Hms���V����I�m������]�@�Қ�S@���(��ư��Z�ՠu�M���7  uXE��#b�	���m׉%�}��)e�Z�BH��)�[e4���-v�Ix�^o�SRMYSt�bT*�©��V�i�d�[]t��=�䐴n�@<hNz�HS���}���@����k�:�����ե��9���p�:��@����)�[e4�]������&���*���Jh�M�����,b��cPR8��)�Z���X�����>���J���rƔ��m��9^�@��z^��o���;��VfҰ���<s�;l2v	�ЮQW3u̵�cO4�LOa���{F���F��vWf8�KF��=����m�<�ŭ��`Wv��Y�6�7Z4��{<ŧ�XGR�Q��ɷ��cr㓶�,��fMq(�s���dmy�3��YW=�unIu$f�&����{K>I:��N������'d�Ø���[���w��w����;�3���t�Hi8�9z=��h�h5�8�Bw���}Ү�b;5E�Kx'�$������u�k�g��!ϯ�x����#��8�
�נu�M���9^�@.�9��!��8�{l��fԔB��Wz�Ӏz{��_5���Ǔ!��N�)�u}V�WZ��)�~���̓�Ī�L�Y�k�s�z(�/_{����)�z�"�d��?��ƿ����5
]��vN{%�:v�6�{n��r�8�}�d"byQ8�
��@�Қ�S@����t�1�0�X�#�M�Jg֠J!�D(i$�D}���`���wv������]>a�u
�ڰ��X��8t(�;�� |���X�FF�B`�H�h�1_��h�}��:���m���R��N28� 7�[l�:���m��W�h^�P	�0�%#yO���6��R;	�V[iz'98�K3������շ�gWG!�c�I�����h_U��4�[X�B!O�4m��9^�@-�hzS~�ďv_��a��ű;hĖ�o�$���ł�@$h0C����!!!@�&(m#{�l�$��(D�[a��8F���b�����$6�B�����*��F���bB1P#_�-�F/����@��XAӤ"kF�e�	(F�!a%�!k)H[M	!�����l`+"	�!��%(L��)H��gĥ�cKB[HR��P��-%HŒRY�B$X�c .)�6���b�X�10�����5�/'�(J!����C������E��U�X� R1XF(D%Ȓ(�|�CA(�����8}i)Z�aHT�%>AF8ω�� `��*D�#
ĬBr�������h�Y���M
X\�1!���7�"2`�c�)��5��H�d)J����m��D޴M2� $�[IIKacc)V�]aib9hʍ�LF,U��R+B4b�R#XP�R Q�DT�T�$�!|�������>J�^QN����U��(�.��7!��Y�2|��:JU3e��sR]]`=�X��`���%�>��]pdx�i�G�ץ4m��9^� n�BP�����B�Sd\���ܕ�t=��˚2���Bm��L����^�j��,�/1���6���>��4W��m��D}A���ow�I�E�Z.m*�4W��m�^��-�s@��q�srcXA��[l�:���%3�݋ sϫ ݪ�jnʻʫ����Q	K�`�ذ���;�� #��s2{�^޺�J�U�b���oޅ~�W���x��hn1H�O#N	��L��I1E���]�v�=M�Ə�͖�P]99��m�h��4W��m�^��-�sAplҴA��q�,Ē�ݹ�H���wv,]k��L�\�����(I��ύ�w4���*�ى.}�L��F(V�ݫ�H���`���[u�k�f�uʓ-�L�S�G3@����k�:��rO{�ٹ'�<�QB�	A�V�PH,dJ�~w��C'>�����cu��;�6�eg�
���j�;Gn;\Qۀ��m\�u]�ܻ�Nx���\2N��q۞ÛXN����������s�����j�n��g�3Z�n�ݩ��-�^�6$�y����`�m=WU��y�LV|��S�)Y��[W%�K��݄���K��44Os��Wr��68��i�Q�/�^��nw�EJ]����?}���v�v�R\vM�;u�4��V�����.�J��N�,��6H(�ư��_��}��@�Қm��B��HwS��M�Oڛ���k$R=ޔ�-�s@��ZVנw�LYSX�2!O�4m��-|�Q�z{���|`�ZʕX�UՂ�"RL�-}V�U�����m���;�\���j4��*���#�����ŀ7Z� n�sR�&&��<��M
�D�k{;��y�M�s(h|	��8dys �i�G�oJh۹�Z���k�?z���X��2a$�ڱ%����	��G�b��y��}��-�M�uY�4�� �d�k n�� �X��Q3����s@=·OQɍa0n-�/��|����@�����h��:�1H�"��@��4m��-}V�U����]M)�B�!2C@����3���g:�chq�{ uۛ����T���O����Iw$���Y�}ذ�\�u��If~A��|h�cܘ〱ȣ�4�\�(Q
d�}Հw;� z�,�ʨ�T��jfU�75u5s�{�ޜ����A8?��#���M�~�6nI��{�{��`�'�(�7Z/���s�ŀk�s�=�� �;�J\ʘ���f���� �O����wN�m��%�]�꠵rX+�4In��:7�,��Y�1�n�%c�z��	�S��S$��q���ߖ�m��:���m���Q������@��3�/U���b�5ֹ�DL�p����qőcqŠ_���-�sO��;��>����/�1`�2!Ē��U��(S���`y�`���%�B�A$�TR +J �FM߱bK��R@�Q,��-v[�+��]�@�Қ[w4�
o�����(5q�;���[m�C5)tԞ�.����k��O��9�hM3��ՠu�M���+����&<��&G��M�Jhm��9^�@:�4˹cU�_�L$m)[x�����DG�Q�{׀w��`��kPs��q��:��@-��{l��B���� 5�����]�j�W8 �w�y>y��;��`��%I?�w4&��,q��ƚc+�݌U�Z	�rbpbٕ�F�E�� ZkQ�q�؇���a�N�ir�֫ct)����k:7�R4mta��MJ�4�n�%N��;��-u��2|ܜ�`���d���b{�k�Ԕm)��i�]��i'mQ�j{N�ύs[�G�l噉�&��:�Zz��p!�S�R����`��%�K�`��ś\���rVi�)b�o�l��L�Ӆ�]c��2�X�q���kK+����2e�9&Jf^^N��|h۹�u}V�[l�/�#�2!Ē��8h۹�u}V�[l�:��������pX���3@��� �٠u�M�w4իX�	cɏ"j'�[l�:���m���~��r�}I��(�H��^��-�s@�z� �٠ya�O-lۋ:���n:�M.�q��mZ�g��C\[AY�*�kr�ǋ�jRb�-��+���Ͽ �;��=��#�;b�:b[V$���3E$l�h]�@��o�ă��É�$$b��z��}4�)�[e4W����BD��G�d�ɠu���l�6^���3��xkV�OT�&H�O�8h�M����f�ץ4݀uK63�������.�/P���3�ms�6#ȨŨkj���d�9 �9n�����m�^���WH�YA@<�"h�= �s�{�8�/YM����H�?��tYsh�Wswx�|`]���D$�	�E(���;����~Սֱ#'��6Ґ�/YM ��h���!%��w���MZ&�¬�CY$��u�4��@�Қ�)�m�v��?n:�=��= �
;:ks���s�:D�ݞ�!\]s����u��6a�ab�'&�^�hzS@�e4�Y�˛*$I8�2,�94�)�)��_�}X ���ڮ��y"�?�h�M����f�ץ4�UC[���6�����`wu��ف�IRS(B��D(�]��?wM�U�IJm4G�[l�:���m��9^�v߯���u,8�ׂ�Ω�6�ݺd�����Dh�0��Bԩ�چ�)S\�Xx���{l�v�e�BK�O>�˪���� ����oJo��"���@>��4�)�{�u9��Z&U]ـl�u�9z�BP�_;� ��>4�.��������zW��:���oJh�W�­�B!�I�c�G�u�Mޔ��f�=���;�:D�@��4m�,�4iL���V���%͘�bEuXCJ��j�l]q�eH	X��0��5h�A���BB�9���jX�`Ea��֔5��+x	��U^��VH��@�g!$����T"�haF0!>� K6[���E5�a	dA��A�
{����$��Vڧg$l��:�[e�kM,m��kr��O��S+c#�˾�g�6ZP8jU���=�#f�kbWlջ%Quf��<x�
m�t`�E���+7��7lb
s�������˗6غ�qm�Ӱ��HMUU*R�mQ쉍�9���(��Jyg��nɱj�� U�j��Cm��6u�r[OlGl���bBy��h���%�^���o�	�2eW��X7I�Ż�#Q�3�Bz�OY��OiCt:�r`殉mՙ+�"�]���mR�hユ�ΰv�v덵�+�s#3��E�n���J:Z�n�%���vx��qBgK��FX.��]�]������s�e�m\:�@�z��q#�j� ���-�zu�G�2����]�\�t��{s�6��2�G&��n�np�mq�/�,8kmv�d�t��oV�3�;�gb�YJ͈���Hy��Zy��$�ڲ 9Pt[d��D��vOH*����%�����V�'*������t,U���d�su����k1Ի���u���/�CF��<�����pf��5Uڀ�]l��[(���z�ص۷�Ҍp�p �S�"2v�����<�u������6ۤ7L�-��֣@qL��v��:U[�f�,l�aӚ�ε;`st�lEumn�m�}� ��Km#݁�c��髪S�Sɬ���V�K�N�Q��Yg��Uuu�=�\�.�=��� /E,��h����g���q�T�T�\!W ;El�,��� ����۲d��?}o�Ҵj@�r�u��+ض� �U*���f�),4�<���v+��ձf�B� )�cJ��vv�+`�ض���t@�M�$���J�l9����E�Z�1��c�y�l��-�#��6� bb�¹�Q]\�8��X�m���`�,��j�A*���+̫�%&���j�+���:���<&�C|�LE(�&��� "�\TH�Ɇ��c�Ź׮������g�,��"l�y�)r��v��K�)�<d�v�q7\[�v8�cm���z��F���֩K<*gcr�0O7.�����4~����'ծS&�����:�Մ����۱�h�|�ݩCWf�M��t�E�m��v�sk����0.x�X�l��P����:����P.����K�v
�H���p�Y�V�JhMYSw/۝b�D��I�%Qћ����W\�ۉ3^�I,�V�' -U�MA5c��� u�4_U�u�M�q\{���țp��f�k��)�[�V � �d]��jAG�W��ޮ���ه���)��|`�׀{���I1�'�$�@�Қ�l�6^���I(���Հ}�9���eZ������ om��D'\�����u�M���ƙ�a��	�'SűśWs�2qjƎ.�<���N���������DP�H~ �_��U��zS@��h�V㉱����NM׻�8(�A � O8��^,I{�~4�Y��U�qDHԙ9$z^��-�M ��h^�@��@�R�
����$��� ���^�@�Қ���	��6�z����zS@��4;ߟ���Q<玼����XV�7�fn�&� ۗD6��[����==��7x���{l��g%�@|���|H��&��@�Қ����f�Wuz�c�	����ݘ{l�z��$�@�Q�#�?��[��l���uZ�4�"���C@:��]��zS@������x�G&�rhu�@��ءD'	�9����� 5��]��~b�뭖�sh��Y싀z�"n�͹�ŋg��̶��ܖ����rԕ�̎=�Jh�����z]k�/�a@�j��TT՘�lΈIL�}~z����:�����+�`����I�h�W�Uֽ�Jh��$���E�Ur�K�K��u`��=v�	�P�?%
k�s�w���<qDc"��zS@�e4���*�^�h;S���f�ۖ�,�u@���v���Ѹ��p�.n�xYő�Y0��H��!�^��W�hu�@�Қ�uZ�py&@B��0�\�DB�:_u`������{�n6�G'�qhu�@om�tB������O� ��C��"�#�@��4�S@��Z]k�;�1���&<��N�l��s�9�u�7��҈P��������i�׵b�t��k��E���U�ݘ^���21������bw���zX{j������(�tk���-�a�1�፶�yr�چ���W�6��;XMu�4;�n�˺x�l��u�U��g�]����v�@���F�I����[ӓt�>��1q�^�N�Ó=ca�6Qp���7�8�7��t�S+RVųQ9����w����?v̕t���]u,t��qv�m�I�Q�8�n��N�6�憞�<S���D�#p�yߖ�WZ�zS@�e4�v��!�iŠUֽޔ�/YM��h�֣ǎ)�2)�oJh���k�
���?{Ʋ�1b�	JC@������*�@��4�Tu���$�$4_U�Uֽޔ�/YM�R%d��dѦK`�xT��v����8t��!/Jg1ә��F'1��dqAbx7�>WoJh���k�����I8F�Ȅ�ى-��y	 ��$[ݸ�%�-Z]����J��&<��n-��h��@�����h��{��(�J27��hwW�Z����h��Q)�C��ƜZ]����@������-�ִ]��LO\�S�.
]�q[����ngmNw..�}x����b����_U�^�����*�^���#���k�&,R#j8����@��Z]k�-}V��:ęL��$� �k�ηXR��򄖤�!-����w�@��|h�V��m�B���
�נZ�����-}V�_��i'"n<��=��h���k�
�נ~Wu5���X����m.�]q�����v���<c�vύ��n����4��LY?�qh���oJhu�@��Z��c�s���@��4
�נZ�����?Qܩ)�C����4
�נZ�����-�M���H��b�L�]`r��Ӏs�� om�V#�P�DRE��	�"HŃ���2 D�"Կ���́�/��œHm���/YMݶ`u���s�r��Dk]ߦ�I|k'\r��ZM���K�Ѯ���8�7�"rh���f�@�3vy��U������~������@�e4�+pq��!�a0N]k�-}V�z�h���_��RD�y9z���/YMޔ�*�^��|5F��cɋ�n-���-�M�����@�Ÿ�n'�bsmF�[ј�n��\�]� �8�
`J=߯È�%�wOne:8�̎zۇQ����������Bƨ�d:=�^�7m56��N	vy�(wv$�.�v��ƣ��ܛ�֐]Ԏ�@�r봫v� �8�[h����3r�����l��kֶt����*�i1������<��)��3��v�l�V.&ˠkr�R�&X���)�^�c��y,�Aó��_M�K#��	;���I$� ��Σ��\��,%��{v�P�p�-�#B�t�w���\�aKp9mgW@\==�������`ֹ��g���|`��u���1F����@�e4zS@��z嗄�ǋHcm���/[��[Қ]k�-}V��5P����A"��X�%=�8�:_u`ֹ��<��, �ut�sSSrYr��p�*�^�k���h���w]c2!@���Q�Q@�#l�+]g��4%OK�����d�Ըؖ�5�n��Y�X�q��H{�s@��^�z��gB�$�* ��$�[��$��P�����>��Xu�p�F�J�ONcQ�ɚ�w4
�נZ�������P�%�#ȱ��������@�n�o]��sk�x�x�����@�n�o]����ϒx��HE ��MI���rWN�m&��E���[vA.x��R�Iq˅�ŋ$�mG�}n�o]����_U�~�:�L&0fH�h���*�@��Z����&���&
L�*�@��Z��~��v@���:�4u��3�#~�X����#����d/�� 
e;ֹ��a�[jh�������5ߟ� �P0�!V�b >a��g�p$� q�C����äSyLH��7���Jcρ;�R	5,)�a�"=1t�T�C��C��� �a�	XƉF���l�ҩB$�� BAH��X�BF({��?h���@DM$��6L�|�wLH0 ��)(C���pbW����j�Sp�*h:,hJ!	�_�:��z5 �с�;c
�}ևP�.�L��n���0�[�>D� ��C���9�QE(: Q/�T}�s�ٹ'~�1$���&��),�m��I �Ӏv�b�׋ s�� ߫QN��	�&,�͸��w4z�hwW�[Қ� �nL�	���'�Rn�q4�մ\��<nl\yM�`R&�k�N�q��5��[�s@�����h��h���q��<y!�7&hw:��s�?�ŀ7�r�IDL�u�l���(�Ǡ}�-��h���*�@���&�<X�L1��q`�l�׋ s�����S� J�,$$H�$�� �$`� 2P��H��2��,
E��ZF�Z0���# P�Ł� �(�,�={g ��*��T]�-PP���w4Ϫ�-}V�}e4/f??���X����V��^q=�q�I�j}���]r�"��Ii���I�[�خ�/>�@��Z����w4�s�rqǑcrE�Z�����޻���h��:�l�y1d�mŠ_[��[�s@�����h�-b�����5��[�s@�����h��h���4	c�0��ɘ��Xu�p�x����/Є
 ޅ�7���T
X��(�6��$�Mظg�l��ʆΫ��8Lji��GG]�����5�rm�\��V��H�v��v9��p�������',V����xB�
�G6��:��vz�:5�޻NT�ә�nQ�
��*��5��[�Bԓ�Ży�Zا\��ِ(Wh�7G��<�쫂^f�u��k�F����Pn#�c�}�{���]�E�V^۞��N��m��ڋk>{��V��/�u�6�n+P�"�^xխ��g�m�9����׋ {Z� �+榩�ŋ$�mG�}n�o]���_U�~�;�ds	��Hh���/>�@��Z���um\Q6�k�&
L�*�@��Z���-빠˞;�N<��-��h�)�[�s@�}V�k�R�aϫX�s�ޮq��ںة-!��c��)t��L�f5��=yX�m���%4z�h�Y�Z���KX�q�+�Gb�U�-��� ���:���񤾰���^�S��7�l�?h�`%�$�7&h�Y�Z���e4zS@��w ���q���@�YMޔ�<�W�~Y�a1b�0��QŠw���oJhW��-}V�y���0�"'��AͳO6s];ϥy\�s.�9�c��!�ˏ��(�QG-�y	��H~���<�W�Z���e4ܕ�
&�1Db�'��z�)�w���oJo䂵��	��"��@��Zz�i�?� @13��|������o4
�����:�x�4Ly3qh�)�[�s@�^�k�e���*�WusSt]U�z�`�[\�����@�YM νZ�Dd�������{�����o �rp]\4!�h�zw7Rո�]�!�xA�����z���;�S@�����ͫ��0�!����;�S@���z���⃹&�L1�Ґ�;�S@���z���)�~�dw��L`��C@o^, ����`L%�BB^U��f,I.�~M��:�t'nh�Y�[Қz�h���:���u���e-����ų�擞��9�b�%�v��7e�*��݇\���Rh���޲��w4׬�;ϰemb��F2'�e4zS@=z�ޔ�=���7�$����4zS@=z�ޔ�;�S@�Ō�x�<��'p�^�@��4���-�M���W�<2aB9x{l�7�l��f |�� DD�"z7[vI%��d�F��E`S���������r�Q�Fy�m���j;p�;')�+��紼����Y�GQ��\r��n	�8펛nĶ.�k=����Þ;bg�8�,��������,�I��ZW*k
N��^<����㇎�
f��3�8�N��ۭ��;��Nm��t����m�vΧ��7N���P�w�����WmHj�r]jeua�Im�3G��'�P4� '>K��i�`�;[Q�(m��=�3[F�b��ϣ� d��˲9�W���9��=�d�cm���w��ޔ�^�@��Z�R��o#�L`̒C@��4׬�-}V�޲���5�B��0N��h��O������^�|h}gƁ�T��`GyG$����;�S@���z��y�U��<Q�3"qh�)�[Қ��h��@��� 9I�3&���;Nͻ9���3�G\�*rn�	:�/2ct��##�&�#p�-�M ��4�\�(��z��>O��MQD��R��ff���w�ߕ4		# ��B�	*���",��,2
� !R0`��D���i�����v�O�ޔ�9{9���s&�H��-}V�޷s@��4+������x�d�cm���;��h����z���h�JV4�!��#��[Қ��h��@�[��\�������l�=iVF����b;[��${n�2�T�7a���K7V$8�� w��Z���n�oJh�K�W�FH8�,�I4_U�w���-�M ��4zPjciLx�	��rN��znI�w^��tEj!�I�!$�߾�����cN��h������4zS@=z���h�)�~�eX�����h�Y�Z���e4zS@�k�q?��6��z匼v-�����=�ٝ��t[kS�О�ܬ�,2<l��b�d�<�rh��@�YMޔ�^�@��qdŒa�USus�o�ٟ�	)������_U�~�)X6���2G3@��4׬�-}V�޷s@�����-S*mV`t(�S;ϯ �Ӏo����Q�LB^P�B����6xuK��$PȲ9$�-}V�޷s@��4׬�?+���M%0�d�F�c�̕B�l؞��m���7�܁�$n�=��d���b��G���Šw���-�M ��~I~��Ӏj$����������7���Jd7�^�O� ߛŀ~��1<m!���n��h��@�[��[Қ,��A��L#�G&�k�������^�@�����b�0��QŠw���آ!B���|Ϫ�߫���
!DB��QEE�QQ_�TQQZ�����**+� ����j(����"�
���W�*(����QQ_�EE(���E�
����**+� ���������
����**+��QQ_�QQ_����)�Ȗ�|�/���8( ���0���  (H  ����H"�   �*�ET(�"�\@     "�P�T�R
*J�B�B�UE(�T�
(R�B��	 ��@D��  D�(   @K]}��緾ϥ����w;�:w�˽��x}�)���l�u������ojp !�v�z����{�Û�����)c�t�׭��iS&��}�<��}i\��k�)�:�  ��E    P ���W6�͹iɧ6���^���
d�_R�LYU)�*�0��Ԫ�,�R�Ԡ*��UJ��R���uU � �    
 @�  ���  �*�D�X: �J�Ԫ����U��*bʥ@ X      �Pr 4�����a%j�*�T�� 5UV3R�bk�uo;u��绫c� ��qo{R��o 7]�z�����| �=[^m��O-��v��zy��U��êggEW&�#qiO�;t��|��  @((g�Ѿ��sq:��sm���nmr������7t���-sk��oW��>��+�r�7<��� i姭95�ow� �R�=9<%}������� t4,�w��ͺM��+� > P(   *��� Ͼiyۭ��}�=�}z��γp z��fޚ����כ#������=�^���O��ͼ� t�o[��M� �<����{yo�[���o]��q��=�NO���י�����U�i
f��"b B*��*R�  �'�UJ�LFFFL'�T�6�H  )������  �!�)" ��>D����O��i�{w����^�w˥��g����(��C7&_� ���AS��QQ_� ������� (*w��H��4�+���	��1��&����j�q	�N�04�:c3��(e1�N!�6o)�V����m�A���)t�F!��i	�$����z<6�%�-�h�fFZ̭ �Ը�a�b0pe���I�J�F�SB��ً!PfL��Ec�t���e���aS�#qRE8���K�l�"?����z0��eI ���-��o����ߗ��g4"��Z�1H�
 �,��L��4��NФ`�C�KI�kZ:)�8�-(Bz0�.�Bh�zz0���ӌ`�$����,��<�y��F,�,-,dig�3ñ�;H���#���di�'CHLbl���M�8ho>lԾ�H�o���A�җ%�4���;|�MH��F�L�V����A��f ��lf�m�&�݋�l�{8�ᤌSK��7�s[8&כ��qӱ�ÊH�̴A��ɍ�|4zym��z`N8h�q��8��.ki��9^xN�����9L�sXY�4���ǉ��Kk���l6��A������>�h��5��BK���J�T�I��_ܟ"U�_?w�ll���L��q�,��L4�Մ����&Z�.E-����1AU��"_>dO��.� ������'AQ������{M���fC�/�!�ɏX٠�5&�ӦѶH�}�6g>&�G�n0ݜno���Sb��鴷�A��涱���s����ٯ}ovp|���0:vo��4y�Z�z�a��=�<��XLW0��A�n��f�4.�y�O3~���W�u�0���f��^��=C��� �	o"�7�����Y�f��4�Á�N.&�G� �t;�����v� 0A)+��q4�B�xA��������k����\�[��3|��~�3�6�G���FÂ@I�bx1���f}�������h6��z�c��7��3[	 �7f����Gc8����D��UD������
���pJU�M̤��J����f�㍽q�h�����=�����`��	��9������6����%pи�%�F"��sx�q�N������8�[�����lÐZ$���{��TeG�U_>�bJ�hQ^��x��ĜL&`pt��7��O�y�k���q &<J p "d�!Hd�lc�!&�I]����6�<9�Y�a�<N�SGF�o��.6J�D"�\�d���u
"��4p#lߥ�m�j
����N�5�|8�=<4l�4o�aVoIa�8�i,tFe�I�XC{�&��20�K3��Kk.D\՚�:�z;B�~�[�z�5���^,`b����lMT�����k�of0���k$��c���8N�6a�c;��߄h#H4a�k���{��	O�!�ӎ��g��g��)	ň|%�t��D�Ei,o�*�BB����T�3k�r��|�ه78�q�%0('D�/�A��ol<��a�I$���#5��#4��6p�!8��<�3[��1�8�a��46s�Yoō�bPG<煚����8���[�bFa>�:D�X!۴%���?"i6;!�M�.&����ޑZc����"�hM�M�\�݅"d��}φ+VD��zR�9(�بR�"E^�����֜~����4���!J�R!X 4���)iY�JHB@�b���bʐ�2`��� ��`l<fJ pt������ԃӳ>��v<|}<p4x��y�V� ��Hqц�$�k��FB	�K�	\t�u:�����8j�K������K�&)V��j�U%m�.2*N��3,���H�K%�E�|�ٿz����ͱ��Ą�p`��Bq�Lp70��4��vg<7��c�a���R*�f}�)Jر}�C�M�б���(�s�_�F�<	"
1toy�#�����)X��&b?�e�HXy�c�d�F�	��F�s�歁OK-	�f�C4�x�a��l3Ë�O���}#A#-'��=�b}��l-h�|[�SLa�n��^�����Ձ�1 )����L�����x�df$�:6�-��P[�N�Æ1���g��Wtvs�Y���fj���4�4��o��j�Z[�!8q��4h=�RHXi�jsn�[��|Q<�=�����o|�kd����	�<X�&o�����M
qx��Jh��<`14o�h<ŌKћ4�1�8`����F$.f7kx����G"�xj$��,8�'�� ��l�t;|'4m[�>���ݐHjL	�A'��H�qW�>�X�*rq��4$�ԓ��ow�+��(֣\޳�> ���u��ͣ�O@�9F�4Na$�`iқ1b|7���$�H`�e�#e��ѧcÔ��<*�.]_Pt� Br�4�kQ���5lў�">*1fB�W)�1���*�%gs�I3�j1l1&z��G��5l�a����c����fFc{�9�K�Q�A�N}�Y�ϼϛ5�}��}i�K���x�X%H��,�P
TV*�k�v�t�c���]��"D+��.r�1�ʼ�#���ȋ��P�<a��8�02BD�g7����<c��\R�QRD�8����X�ԓ!��l>#5x�1A8���]�R�Z9�_	q*T��J��1�M$ N�1��Z�_$s�+>X,K����T$R3��Z�&g�=���\f$1��i�N&��g^��q��sͺ�s��R�&���\M�R�Ϲą)�bFs�$!|���5er�_5��RϧN�|/���K�+�g.^|�\�f�l#5�1�5�ChѶ#3pDTģa�7U�$�
v��	�(�P# �XX=K�.Y����1ћוf��
+U8��q �X��Jd�)�dm�` ��#�|5��l�����#�F���xs_o�#�<1�k�`!�o�`h����縐I�x{�;�������V�7Ͼ��"D�h>�}*���h�l5�|���h~Q�h	�}�y��a��k;��F�s�xi"  RVA��B��I�2�	�iL��Б�D�C���f�3���I�BH=�]�@`��Sa�eh�"5�	X�Wy$tH(+ň�x1|q��#c�ŉ��!0�%<M�(dԱ%RSF3�D�1��dF��ܑ�j4�����:0�3Ai�8Z���s�ka�����&�6��%��5��i �R�xG��11���q|:1��.o�;���<"�n\%fq�	�e�J�w:��8��]�����#�n�I@NN�24��rM�8��9����G�|����-rQ�"�Tj���Ŝ#N�xN�F:m���.��b�+m��>*�-��Ǚ�*�\_	I�DQ�II�2!41��1�F,a�c6N���IkZѤ�]�5� �6�23Ѿ$oZ#Da:ƈ�IEB� ��	S�J�<�I"U�h4�a�h��J�:Y�Ӥg

��D�$f���ֶ\֘�p�4٭di'+[5�nF�ČHcA8C��ѣzծ�fQːD�!U��ȳ�1Jb�
*Sh�A��2ִ�Ii�4Nhb��BUI
$*� ���+r�����H m� 	 m�h  6���� �  m�  pj��$v���>V��a ��mC�r��8�J���,R�Ѩ�:��µJq�]��� 6�h�v��@q��m��n[x!�nh�� � z���m�2�3j�  �Ԁsn��[@��8 �۵�3Pl��t��ݶ  �D��c����ɫ����b�1m $	k�Hj� -08�[G)zԲ�l�� �   -��$�"�-���  �!�m�m -��m�����  �� [@  "Al��l [v��m�` -���    8	i� qmI'm�p�� ㍶�i;  6� �   8 �         �@ �b�-�Hsm� ��8 �    $  �l���� �i�b�lp�� � m�      ���tm� |m�8$�m!mq ���@ -mT��]m�M[T��D���   H mp8   	  �kh �� � @ � ��7�|m�!��@	$ -�mm�"Cm�-�m�        m� ���@� m�� [Sv� �t$ m��$8��@k&�5�5*�Լ�~����3ӉV����`          ���-� �6ٶ� �#m�[Am����@mm    ��[� mm m�%h@	$p�s����Y2ÕX�ͻ�h�����#m� -�� ���-�Am-�Kc�,`��3UHMl�̺� � sm�[Xh��I �]ζA��9�Ā p v�&�Z�/i�z��s�7'a
��+)ekk#�@U�W#��gWR���7C�孪�̩V[v[@K!v )�v�3CV�F�䪨 �	�n�h��-���g��d�nܝI�ճ�l  p� �Lm�@8-� �eֶ�l�Iv��  j�<h-i-�k&�8�֜@ m� H6��R�J��OZ��ݖ��  H �8�2{ѭ(�Ʈe���%�� p!4dZ��,����UUR	�kmc]��:B���Ycb|�M�
Wm�j�8��ݶL.Ŗ��V�`1��m9�[tՓ[pm�v�wl  �  @��m����(�m�[�  �� I kVܚ&� UP�
 r�����
6�r�&kh�#]3y���� m�id�gN�x��TUR�p0lTuU�p�s���j4WWd��j��
U�T'vڶ��l � [\�j�;U�^� ��ym+m�N���d�-��suI�Md�n%SSV�R��plUN>8�_l�N�����K��	0 �t�6�m�ԮW]�6f���E��]���=r��:#g�Y:�6殒-�GF���NM�7����t���m��I �^M�8�eRp\��+�xj�v&v�c���[�~~T�F� f��A��2q6�L�!�[�v�H�]20[Vq�in�vȻkh 6Ȳ� �$�uIm6��n�d��lI  m"�rI'e�vL��j㵓@-�6݂�6�-�ּ�"Igm�c5�Kd� $[@������`�UU[]������뤶�� �� I����}�ʲ��T�qg69��Cb�e���`�.]d��v �4�����Z'A"���t�(��j��)<��HH�@�n��%Vŷ)��V����7N� �gI"H���ڶ�-��/Z .��m�tˣ��q�d^���r�6$v�at�{kg[�`�� H[M7gMN�n�`-���H @ l���-��/OLvշHh-����*�����TJ\�nS�����@uV�UP�T鱱&��m�-6 $ �m�� � �'���&���@Hm�  n�F�]���jv^nV��yz
Ci�H����N �Zl�vcn�i6j�:�v�b������s�s�U� ��:p���p88�.�coIRm����s�� 	�Y�Q�V��' �Z�]�n�Jj�:��{N�eVUU���-]:v���ۀ1m��I�۲�8�[$%�g��ݰ����F� C[�l�]�6 �K5Zq;K�x�Pʦ�l�K��m�(�����+L�vݸni� ��Y4�2��&ٶ�l�H7m�[V����d��հ�UU�e��qն6m��Á���+d��k�6�U��ط<�uZp$m�e��zT��q[)9��V����U���ڪM�P,������
V�F����-�= ې��V�ڶ���,� m��k��ŷ�����u��m��j٢�  -��N��
V�H�v�lH/]r��`�8É��N�m�g��E�[5J�mU�s�,�W(�bHM/"�h-�[A��n�m���K��U��9��l��P� Nݮ 	��VN�I��	�WV];`m���Yd�3u�ڵo9]X쇕�u.�t��L��.88%�J�ͭ��WJ��R� 9�e�-p�)���U^n��lx�]��%ZU����;*�P�
�U�6�ٹ\php�*�O/5l1Ͷv�<7ceo#��@T�t��wm�I��� ���US�vZ�U��1�V��U��Y�٪^$���!NҪ�h���-���e�����P P�]���r̤�ی�Pm���c�[u�n�` $�X�Y�� �d�]m��@ R��ԣ��ckķ�p m���$��UP��8q�v8*�K�+mm�u� %� [d���M���8��ҮҠ5T[(��!=mƵ�$$m�U�@ �K�s�N$c��f��I%����M��]��wD�o`6�K5�K$�y��$��t�h�m�h -����c^�NͲޣm�@ I�n�v��?�>  �a��t�$J�� ���m�@[VҼ� ��i��[)��H9������KR0��M'�Y����  �[�[zt-�$l T�+/2�#jUZ�T�۶���ŵ�   m�[�� � 趖ޛ^�Z-����-���UTͳT��4ԅ;--�D��� m�  q�jA��$��-�h�� �ڶ�ɶ�����5�.�gf����į9GR���3f�6�Yym��� $  �����o��l�Ԫ�r��-\�ڪ��v9-$���t�n� Xc��XlĀ6�k� ؔ��.�e�j�z�$�xn�qn�Iv�P/,���[:*�(sc%bHɺ��:T�9�m�P�m$p[R�$�d�`Hm�[M�X����"�am� p��9���>��~8�j��!6����w7i-�	*�=l��������Ʀ�ռ� .���U@h8�����j6�� �� ��m��{6�]�켍d��V���-�ܼ)���ך��jRZ�TN��gY�pȼ�v;/̴��WR~�~���x���j6�k���k�  ��&���<�h       .�+�˭���V��]�n�$RC�����^�P��d���� ���I��l۶���[vKƷ�k���V����l(�|$}�Ze�  ��Kւ
�4�ҫՌU�UpR�UU�*�+cH���m� �h   �6��� 	
�V�oY�l�  ��f�&	� [��I�[v^�  ��6�� N2kX6�HI����H�& qa�$�Q�b�*T�<�e��YЄԫp�P+*� Ǥҵ�ph�J�^�i��ֱh�6���6�tu�\�P�)�:�-ɲ ��`��o��  � ��I��z�� [@�8@ p l   $� ��P m�ШU[mm!4�T*���	 u.�@�kh  	    m�H�z�[@%�sl��m�-�Ĝ� -�    m� ��    �-�-� ��E��mq     H  �I�	� m�m�  6�   �m8�g�ƺ`qm� �J�B��ms-�UT&5*�Yi(�UZ���K��`��յbYV�s��� $: �m�|�    �@S�U�#����y����<��(~�� L���` �l��6��l[�ӥ� $��Hll$H�d:β�l�H U\�mk���*��U�/*��Yv��+UW:)V��AR �B,	��J�9� �����
lP|�@�."�p@��J��~Qz��N �1"�/U���6(z0"�)����t�"���_�
��)�)�j���4z�T�7�th���� ��
p�'�D � 
� ~CJ���𲰁(%(�J�`��|P_UYD41BĐ�UCP �
|���H@6m^��0A>PTqE�� D_Q�D<W�$�l�I�"�$��`�P �*�����U
�����=D^��DW�D}�1N��P
�*EGS��p8|	z �DC�>�h ��@�| ����ASa� C`|�{���ʨ`��8cE 1=U�� ��A�oj�������YD }��U<@t uU!RD<���ڏ���HF!�{����q�ۼ~?��������m�e���ai��WX�N�&���2�1.�؋�j;t�;Sb�îwT�Rڥh��̬��I�U[���&���U�&�&m1m�3�l 2鉍\ԫ�ju0��»<5WP�aB����vc���Pl*�@����UmP��"���7����2�sUU� �jmuk����hlr�v!�x�8��:�5� d�Kta�grK:�s�`��Ι2�9��{v�qwHB�Z�a�SIxH.�g1��6C�sEWs^�K����sa�۪YT��ѹƽ����L��;[x�r�Z{Cp�����.2��Y!�%�mR������/�^1���92JX}���۠�T��v�)C���-;60.�o��c8� U��;t:����s-�8�g"��s����Jl��³Oiɲ��P�ne8m֤�,�::z�&�5�X��V����3�x�mƮ���Ši^؍�C���#qێ���QL�kg' f`�삩�.�Q �v��X�tU��n���nx�n�M�ɍ��pl�[�]%.-�r�8�nn|gOE8����dV6�M��/=q�/>z܇b�x�ݻs0�ۢ�,�����\ݭ���#N�3ȓI8�����k��c���#���6x�NA���;<)z؛����6W��YE�i�/<rm�T�e�ڭ�LV-��r���e�UƤ� ���;2ۻ8�9v�-�-m�I�����#�=�o=��\�K��phnz�h��b�H���i�{���`�a��{Vά�i�Eʜ6E]]��3���cm�+ ��&�/j+{0k8:�x�������[B��n���q�+-ljB�vHu�8ħ]�m���<��y�9��V��'.�!��TlU�+�2�6X�����Ul���d��N�$���u�N�:s�*�u����m�9�E���ĳ�;pD��Vs��7j�j�h�|��P
���aBF� W�l0U�G�qT�}�b�!۶��[.��l	��� d8+q�����=���%\7F3��l��f����ok�=�c���[�f�ۙ�W�)�n+����u�՝i�c�\d��G��o,�g����g<�����mݟ:�q�js[!���WC;�q��έܰ]�'7R2mZsc;M�V{I(�n�]���MR���6�B�J�,V#������&�'m�8+�)
 ���E��2��Gq�(a�ɹB)P���*MP��>���,��X����ɴ�O���, ���a"U`������g�m�v�� ;��`��`n�ՒE(�ؔCs��@nj ��=m�@>���w��Dqp����͖f�z�U�΃2��J�I7�9�@zۘ���Z �sP���o�"+� �ְ����]in<T�G8���v�^T�u�I�M7Z��1������r����'9�G�p˵$�	R�� �Wve�I$��l�_U@x*�  �ך�'� 	�j��b�-������7v��sv�� �j��b�VPjݢJ_������;�,_9�Lr�� 
py3/h����
3wP�s��=�*@��aEn��_7A�Q�6�	��8����j�z#�vKӧ^�΄�����Ӯ�ݳ��@zc���8� >sP�s,�n�^��G �o�����1�Z���9�����j����Z�����{��&���b`H�*@���o~�\�r���xX̃�H1�QEQI�f�������5�Ojf^՗���,�����9�7 �j����'�I�^)T�˔Z�j�IVz��(���u�]��.�9�휌n�-�y���a�U$T��>��]Xw6X36X[���	n�"�8�II*�3�5 y��\sn*@��f^Њ)S�C�X36X[���]��Հno����VI��i(��rX[ݬ��q`yݼI�6�CHJڒ�|��� :~�_��o�y��+�%�&�N��8�w}u`��`��`qwu��7��W�(�S�����Z�a��@7������;����䎎$�Ʋ���Q�J'+���,��,�7k�m7�n����.�T�sn��w7P��������qR �rX��Z�i�!�%����`y�� w9���@;�9X^vI(�����Ի��U�fo��s3e����`n�Kv�$�%$� �{��y6�����'}��>�w��FߩT��qh%!3�6���B�/����]It�P*�oi��@ݓey�[Pru�ӭ����@w�����ġ{5�v^9���rg���<#D��;�f�rB[�;B�Ki'0rn�ٱ�zh0�:������3��nqh�����+��0Գ�[O��/��
q�s�����*B&Ɩ*<�:����ʅ@$��srLP��Ej�pM�x���,���Ĥ��V��nݾ��[��IŸ�'b�$����[1J�Ł���g�������A�ڔ"�T�P���K�����qR �sPIKow6��2ͳ2�7P��n*@�j �sP��W�.	6�v���;�� �se�s3e����`s�̭bTTl�����@�j �sP��n*@s���T�F����K �f������f�X{�,�O�h�7"����uݹFz��t�<��*�������z.���G#H_
��$��=�`s3n��͖�͖*7tbb$T�k{�*��Ý��*����M�j �&�=}& $���ܦ*N*RJ��6X36X]�v�����;[U-
��Ww��ܾ��@u������s��m����i6D6������=�Uwv�p3},��,}������4�"|�y�n_92�V��*O'c�@k�d�voG2�m\KK�M���#q������ �f������F�+X�#��R�wo?6�I������� ���0w �����7E$rX36X]��-/�����Gz�}�ʯ=���\��Z� _
��$�w]��ͺ��6X36X�wH&�$R�*�������s��<���sPmߝ���~7jy[��$a�Wh�����+�Ƀp���u��հ�)���]s.�;�� s����b �9��� V���jQH)S�C�X����͘��� }���m�n��B.�R�������}��� {���������\�&�ӱ����/���.�߻�|���{�V(u��RQz�7�[^�][	 �J�I.]��sP�L@�5� <ܢ�Y�� �F��rk-�[�>�ڗZ�'i��D0]����HsXssG/bc����~Ԙ�=�j7�@�5�Oja�dWd"*��wo<�i�!������5wu�en��Ҥ�REHo7P�� �9�	}& s��o�Vӎ��8�IG�������`�5� 
�O.a�U�]f�f� %���=�j<r��s�����띋�g��p��%ٚͶ��xT�j Z��g*����ď;cQ\��	��yݦ�� y�p]��gf�v�;�ϯ#��s˥Żk{<g3����5ɠ�ㆇt�룩�яN{I�^D�s�AQ��������q��,�l;]Kc:� �o!Tl�g��kv:��P�Q^W�p��v.��x�=����{��Q��f��[TE��wq�����͏���!�&{n��64�2�v��k��v�7@�۷k�o#�Υ����FӧR������X㖀�󘀗�bߣ���,/3���y����@u󘀗�b �I��)�%ED�:IH�:�����,�U�RGsޖuμ���T�
8�'#��9���9��`sj�:���md�d�/�$�$������i�o}>�����ݼ�{$�����"5����)7(u�l���7��9��+�ۭu�D�gi�"���2��y%�:��@�߿~������I=G��
R�"I*����f����&a )$�J	I^".�_I�@ɨ<��G����*�t7q ssP�M@y䖀��1��S\o�6�:��NK �we��{-��b ��=�9��䬻̼�FFܜ���`~����y�| ��K �wo �I5���B��]ը���0�\t�e��]���&{]�V��[7�C�x�n[ `��t��E�1f��s6X;�,c�V;�{NEM���r8���W�v��P3���b �O*a��!�!�%�s����<�gk�ϕW�
-QD4�5����bS���A�g8'6��2�0�:XE�� ��%�K4hM:p҈�:��Y�OxJ�8#�34��޶9"�I��E֊a߂����P\cH�
���@1_G�*��hA�� �t��Uռ��^����SM�%JH��,fM,�s���=�j�.�7s?e�f�w�������t���{�M7�#=*�(��%]S,�+�Rx�u����e�{r�١-vۣ:�+��=���6���� t�j �I�7�@u��`gpS\o���6���9��~����,�; �f����j�r�
64�q�' �z~,�͖�͖����
yZ����t��B���m`��� }���R�x�R��Z�m���i�i>K��0��Z��*��]+�w7���u|� <����z����~I���-Ѣ�$����Q��5�Kκܝ������dƺɋ��s��� �I�7�@z��@nj ���4�BT���ܒ��f�X]�v�͖���j�$o�T%{�H_9���@�5��[��B ��H)�s3e�s����f�X��Vw5�����if� �9�7 =��75*�kwD,Rժ%�\Ub(�.�TkUd֞g�Gm�]�"��4��=���۵��ѹHv;k`�
gs��&���x��ʗ���u�:r�-�쯳�m7g1�<u�=N��.�`��A��CcQ9n͎
�nRe�A �q�y�+;X���c�H��h�Ov�R�ؔ��h�z.�z6�g"a��h�e����m6��|�}r�.)f.������ԨOm<���ӵ|z����ƨ�e�2�y�u�\q����[و��Tc$T�whQ:�Q7'@�{�����s���c�eҨ��)%��μ�`��`�l�9�4�9܃6�)*#q�I��s��sPo`��c��#.7n��HqrI`�l�9�4�9ך���,CwJi�$�I!�%��{����s��p��m�BPs��yPg�����@�]m�jLn �#vН�ts÷��=��}��Uݘ�{��s�Ͷ��9�~0w఑
+��.� }����Zm����6X̚X��W�H��O8�Ѷ1�m'%�w7���d��UW�w�Xw},a��59`�`�m��;��v9h��@�5�
���$:��R8�u� �f� �se��y���_UV�f�g�PR0q�$�+ְ6plbC,t����a�ͷn��e��Ru��
8�&㋀���wvXǚ��� ��t�EH_$8�9$�t����-ݎZ �sP�HTLi%JH��,c�V:�U�����D4
�@w������{��Z�Sl�AN:JE`s�5X36 s����- WB��6���t2K��w�x�I�9���6�� ����մSw#�Jd"���E'����s�����v:�c�n;^�6��%�e����y��=�j������9������m88ۓ�w^�X�r����=�j��wa�y[�w{����c��9����<����r5Zȩ*qA8���,��<�����8��+�VM۫�!I,�ݖ3f�z�U�w3e�V�7����A�DS��q:zN��y`�)������Ψ͎۬y[]sG%n�)%JH��,f�,�� �f� �we���[��|0�	&�`w��@���Ps`�+Ыr��!R��"��l�wvX͚X��Vf
k�ҍЇ����ɨ9�@wc��9��1��7<�j6�G�p溜�y��;���>���4����*�$UW"�,�{��^�lr`p����)���qlH�n=!���D⚃���9�c�ܫ��8����ӯ7%�8��I��5�W;���\�Fv�,�I{N���k6ݝ�k9M��!Z8݇��v7:�[Ÿ78���o�>ɷ�!7d� �:e��=*gu���;�A#Eg�:v��2���ggH�X3Y�p];��+��j���e��{���<H�ė�ͷv�Rj6��7lװ�����ѡ{�Xkm�#��71�����p�`����;���9���_}U��Ofƫ̊��G#�H��l�t���_9�WL���WvUٛe����=�j�EH�s7��3Q�P�i��R�X�۫��b ��s��ud�s2��f�w�����9����<��X�F��Oi�@�j�MP��A�[��g�M���\V�s���=7X�M7h�+t0��@���sPr*@z��`f`���#T!�m'%�s����	��� �}Tp<U�\��p�]Y����,a��8�`8�N������*@z��G�~��j �>��j�F�Q!Ԕ��ʰ8�����,�͖��w}�U����y�RUrafnm�nj��>��� s�`Y��i�N��J:��2*r6�V�R�jq����=����붷%�����S�G��e����=�j�EH��@ܖVj��tP�J�ے��n�_���UW`��P��@�5 ��r�dC�*�D��� }���;ݼ���iq������9��X�Ȏ��]n������=�j�EH��X��64%
hpI�`�l�<�T�=�j ��=�ͅe��ͽ́�{ny��_96R�u=�s8y�
��[=�noG2�b@Q~q݃���HӒp����9�5 {���sP�.����2�K�76���@�5 {����H�J-DT�F�R���`�l�u�@{�T�=�j �&VM۫�(�Ͳ���@�5�qR �9�7�~��R��@>��Ce�W��}�;�(z1�B�*CnK�ͺ�s��=�j��b �ReKͫ��î�!ɵ�n���-ی��$.C�6�:�޳�Z0�ҡL�(��)�BQ�V��� ����>������;�ŀ���JT��(rK �se��$uf����Հs���I��=�48��:���#��g9��s�@z_�����m�R������ܫ ��K �;���Ԝ�x:T[�,��J�
�X�wo �i�M%]�~� w~��w�9V��IpS���@��I����pD蘻�0љ�3�2��ҔUQ2@0EX����a&,A�<"	���8!�$+ ��L�����$���~�"�ᯑ�xD��9�DAIb8Ɋ�;o�[�Aa���,!,��2�F�E�AD�! $e�@!>B~LҚ ��2a$3F���A�Q��a��6L�Ĝ9�$�����Ap���"�q�z��&#�8X<�#o �,��x <��X��Y �MELl������9���Y�he��������eh2�p�
H1a"$`�$��1%el �#3đ ����uU�U��ת嬠���Z�)Q�����z��ˡS�ݐ� ����wWU���UM�����V�̧N�U��خ�i6;t���l6݂@�m��*Lͫv ��d�����8·�X���2Z$���T��^�nr��M��ڠ*�x&���aGZ�C[6�-��[��2"����uv�ڎW'7[��#�����ěRn6����Ĺս;�ӕC=`݈!]�ݸUI��WYN�%�*��&�T6�
nG��g4S���sۜ��M��� �)^#Ab�(
_Q��]م�n��Ϋ�nm��8�7cN��^ۙU�����k�o}��,��67l��G]��7pVHɎ--���\�4���+�J��6��=�ʷ�1WKk)��vv0����U�/0�V�|��MҞk�9�A@�3�#�P�]篩�w��!�v�kJMr�!v05��Ue��pn�tA&��+�u��6L���>�q�t
��W7�ԙ=�'�nn�ܣ��q���{F�g�(Y��.U���l�K��سNR�:�__}��j޹q�wV��ml�O$�9���٠9�s� t]B����<1mۭ��M�9,C��=�1�Lu�-�b�n�m�YS�C9Ѵ��q�]�5����k9����7ۥmu�]���3r�Ԧ됥z�ٶ݌�.��l[�Jrbk�v���@ 0� �7C-��"� غ���ѬL�T�Xu`ǉ���9���;k+��b{t2ꚡ���c�N|j���C-��ā��	ΎKdK�jmz�c�`�ٴ�)��ڷ�Z��r�譔�Qfn�q�]��:x�ѡP;�)K\j5���-�x͌k����t��%��xx�����XT�t,*�<lͲ�]s�#eyZ�<��k���W���[;�6v[�KH@<]Ur��t��8�T@�;�,�%d֍�e��޳ZӡA����#� ����6��|y��F�-kfQ[�Ց���rnJ�`�&�b�b���i��]��{:�V{,�Vy�n�kG�6�d��n����kvè�}k��#j^�.����-�2�mu�Z rR�N���c��[q�p�<v������OcؼC�f�;��q�V�x�n:9tv�RM�����ZMr��D���fU�EsqN�j�5\�n�1���h��i��d���~��n��K�P'�&N3����v�¥��'bB�6��.�����S����Y��P�6�t�nO��ߥ�s����sn�\@fo��o���B��$��7o?�i��U�~ŀ��x�;�~������ �J����zx��6Y�����,�]j��
j����w4@�j �sP�M@{�i`Ԩݢ�NQC�X{�,�&�=�`�;��2K�Y�y�����u�.�O9�WN�͉�$8�2sm۵�7�=)P4�$hJ��6���9��`{�� w9���@z^��@�ʩJ�U��s��'�>���5Jýͼ ��� }����ڐ�J�|�r���/t@ϵ w9�\s鰰;�Pz�T*M��)��;��`z㘀�M� |�yW3n���6�3wu�b�6�;��+q%�q�%4Ӑ�5D���C^1�K�9�V�&���{u�NE�t��ݛ���.�owq�qR |�s����1�ѻh�S�ģ��;�,�wo �sv���ŞI7 w�y
� U+Qwx�� �sv���M�ľ�G��V��,��Ƅ�Pu)��u��1�qR��u]�z���e���H6��͕ �;0�{6X]�vv��)*6�#Bp��o@&�Wn�ܻ��&Mխk\y�e۠��o2��FJp"&4�!ʰ;ܚX;�,.��ͺ�3���ĨT�q:M)�sP��� ;�� 9-:5��B��$�w]����X�M,�͖w`=��N���R��X��w�,���s�x�K��6&�&�	6�_w+ ��;��PQU����� ;�� {�������Vt�&��D�18�:"c��7K�nsh�s��#�bci�-vۣs{aX�@�]�0m�[Vf���=}& =�*@{��`w��64%
hpI�`qw5߫�~�����R�߄�sPc���m�V�mԍ7' �o��w&���� �we�΍Vh:Q&$�!ʰ;�`�=�j �9�t� ;��m�&�N�ԅ�w���9��`s�4�9�ޘO�m$�߆b��%+U���;ko%)�l��vڕ�8c��C�-�i֓$S��ۮ@W�W�ѥIÈ�M��I =y�,뮹{u�ƹQ�]q����]vݍ�98�b��N��9��B[�uk��k(�ўe�:������Nt�9�s��+���B�Kmt]z�+(t<z�#��^�U��۬��=[.��Ē�gKq˚uk�b�6�ԝ����9�p}񮋧-:h�p�݆�[��s��!�ku����s�^����[0=�;m��1�w`���=�`��{ꪯ�������z��!)�q���/�}�}I�<X�|�.���F�0T9LJI*��ri`uw5�]�v;�u`5Rݢ��Rj8X\� =|� =���?_8�˺߶�M���Sq�]�v��Y��ˠf�~,.�0+5���N�Jm�_�#������yt��\u�vݺ�f56��������M6�A������ri`�l���@w7���j�תRi�'R�R�`s��ci�%T�����^�6���o�j���)��J��U%K� $��P��G�Uw���@s���v�a@P��!�%����o�����}�ޘ���V�^�����U�F��,wf����ߎ fo��%�;���mwP�و�Et]H���r�.�@��C�%Ɯ�cx�O<4vܙ��G<|�T���PP@�P�����k���%)K�~���)C�wi�����;��m]����$%�K���){��� ��1ԥ'���<��>����)JR{���<�����vE~�.J����*�@��}���������8�;D^�?��5���O�6����h@��;����0W*UR�*U��ms����'�}���JR�߻�)B�!d�۾��mk�����UAT�I%ٍ��'�}���JR�߻�)JRy}�t<��<����)JOCߝ]�v���`���:g6�@����Đ���=�n��G[P�V��³�%n��������w�)JO/�����}��6��nׄ�mh�l�����I*��@���v��y�4���}~8�)I�{���R��=��⟳�i�o�V�IwqB������w��R��}��%)Os߻�)JP���h]�&�uT��
�	.��R��H2O{�~������k�R�>}�v<���@����ݘ��5�H��+$!T�J�V'��������)<���JR�{��8�)I��k��R��
�{؋���=��hǦA���O'�z���%�֭�ݸ��ض�s������H�Nz�#?Ҕ�'����JR�{��8�)I�{Z'�h\���6��}ӻ/�*�"�R���R���mk��zbK�@����%)K��|R������y+��'�{Q{�]��T�I.�ch�����y)J^��w�)� �d��Rx6���׽1��k��R�.)���RT������w׍�m{w��<��<�]�qJR�Ͼ�a����씉�Z����@�$����y)Jy��┥'�}���JS����R���<�@�?��ߟ��;�:��<0 :(A�p6s�
�[OZu`�	�e�p�pюm���r��x9+��*���=#�R�霳��^���t��Y1����KѸŴ�ן��@��ݙ٪.^�.���|�}���Z�r/5�;`��n��q���8u����wZ�;�n������=�272�n$%�;y���å����6�IֻE;fUT䲵n��o	|7<*���pe�ʁ�z��:7OX�o,X���I=�V�IwqK�wI�6��ͭ���)I��k��R��=���K�����Rx6��o��\���(��$�w1������y)J{���qJR�Ͼ�ǒ�����)JP����Hݙ�Z�.�O�6�9ݬmh���O%)O=�{�R�����y)Jy�dW�%�TR�EJ���6�?�ݴ�R���w��)JO>�]�����m�h@�yݗ�*�"�R����*�?�)O~����)J?�}�u�%)K��|R������y)J�������.�M�჻W��m��g=��[y����v�I��ݻ7��7:�6��)�z1�?�{�R��ߵ�%)K�~���)I����_ɴ|6���׽1��k�إx����RT�������$�'֖<CY��	����[��%)M�{�@���kD�kͱ86���H��RU������k��<T����)O�	�8����C�JZ7}���O��芹RK��\�އ������)JRy���<��G9ݼmk͐k��<@�=�=몡Z��.�6��}�։�ڠ? O�����)JOn��������ٍ�mKWa�j�Z��.�]\���%�v��-�W^�+4�=n6�݅�C����;�L�+$!T�J�V'���gwՍ�R��ﻡ�)��s�����@�}��'�h]�Ig�u+Z��޸�)I�����R���w��)JO>�]���������3����/�*�"�D�V��WI�6��ݯߦ6�JO>�]��
�}J��B^+�%
�W@o��0q�AM�xl �Z@��� Nk���'LR�{(g=3ۂ� �X%f���rHH��Q34g��<BY$b	!&������hK)�5�PG����ȏb�R������ �*��*s�	�D�+�PGJ�H����|
:���U:����S�O�e>��+@����h_r��e�%UR�B��6��}�։����w�┥'�}ݏ%)O=�{�R��s���E���WJIR�O�6�s�|R���ﻱ�)��s�R��w�m�����MT�]�U�*��tι�!�FM�"J�Z����5��:�C�N���RU������k��m<@����s�R��}�v���/}��┤'݆�r���w����mk�V�qJR��~�ג���w|R���{���m�mmTRDU�Ir�b��'��ݯ%)K�~���)I�{���m}�ݘ��'��n�Y$��Z�]�x6��s����6����i�)��s�P��I�~�ג���;,کuXQR����k����R���w��)JO���^JR��;���m_#�T�dT\��˧-�=:��M���n�s	�kru�lvݹ��l[]e��Q*��	V��m}�ݘ��5�~�ג�������)<����R���m�d��J�����5�{�^JR��w\R���ﻱ�)�+vch@�9إj,�EJ�RJ�m�R��=��┥'�}ݏ%)O=�{�R���ﻵ�)}���k](�*�J���m����<@��k��┥'�}ݯ%)Os߻�)JSZi7DK�QI.�)wui���ܭ�┥'�}ݯ%)Os߻�)JRy����R��t� �
	:h1GH�.�#���Z�FΘ<�,��i���� �&�Ķ�C��Gg�J^�tɷe݆`�s�f�����q���W���t���wn\���Y�n�+[��әь�ʥ��ugK��u���c��ش�nsٞγnz��IRV�8�^3�%Lm�͈]�ΎR��η.=�]Y�<��^2�b����JR5�XVv�g*F��r��S��;����S�-�<���vz7Ch����K�4��n��\[�y�`\	�Խ�Sr�Z��.涁�}��o�6�9ݬiJRy����R���w��)J�I�rB*�jT���mk�����)I��wc�JS�u���)<���pmk��mT��*��(�WX��'�}ݏ%)O=�{�R���ﻵ��Nwk@��ΛR��W*J�j�5��)��s�R��}�v���b��(J3�(J��J��(L���ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP����pJ��(O3�(J��J��(L���(J!(J��=�w�YV�*��+�W>�4	�MhD%	BP�&f	BP�%	�%	BP��%	BP�'���<��(J��(J��"��(J3�(J��J��(L���ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP����pJ��(O3�(J��J��(L���(J!(J��=��g�	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP��G�/,�8�n�&�h���ʤ�W���cs�Rm��d��z����vFxo|%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP�����<��(J!(J��30J��(H��(J���(J��=�p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B{��~�<��(J!(J��30J��(H��(J���(J��=�q��%	BP�f	BP�%	�%	BP��%	BP�$BP���&��6���)*�]���e	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B{����(J��<��T? �<@�D�/!(J��(J��0J��(J��(J����y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP������(J��(J��(J��(L���(J��(J�Ͼ�����%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP���=��D�u%���h@��&y�%	BP�%	BP�%	��P�%	BP�%	BP���߳��(J��(J��30J��(J��(J3�(J����ÂP�%	By�%	BP�%	BP�%	��P�%	BP�%	BP�����<��(J��(J���(J��(J��(L���(J���8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�_���oY̰��,����x%	BP�%	BP�%	��P�%	BRʡ(�>��� ���||���A�4~��(J��=��g�	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�(F���ArB*�jT����Me	By�%	BP�%	BP�%	��P�%	BP�%	BP�����<��(J��(J���(J��(J��(L���(J���8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	����<�J��(J��(J3�(J��(J��30J��(O{��8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	����~�a�\�{m��t���=[.��l/c/h���k��j�a���ܜ�(5��rP�%	BP�%	BP��%	BP�%	BP�%	��P�%	B{����(J��0J��(J��(J3�(J��(J��=��g�	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	�{���(J��0J��(J��(J3�(J��(J��3��~x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP��ޭ�VUȮ"S�A*�4	�Mj��0J��(J��(J3�(J��(J��=��g�	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	�{���(J��0J��(J��(J3�(J��(J��3��~x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'���pJ��(O3�(J��(J��30J��(J��(J߷�~5���f�[��o[�<��(J��(J���(J��(J��(L���(J���	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bg�w���J��(J��(J3�)4hG�+"��*�M�!(H��(J��`�%	BP�~��	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�����P�%	BD%	BP�&f	BP�%	�%	BP��$&�4	�Mw��"�DW��[��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg�w���J��(H��(J���(J��"��(J3�(J����ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	����<�J��(H��(J���(J��"��(J3�(J����ǂP�%	By�%	BP�$BP�%	Bf`�%	BP�	B�4	�MM�M%W�%]����IBP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP����pJ��(O3�(J��J��(L���(J!(J��=��g�	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP�����J��(O3�(J��J��(L���(J!(J��3��~x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P���&���K�)W*)u*U�
Un�H.�e)69�q�6��M�n��A  �۱kFY���3{޶pJ��(O3�(J��J��(L���(J!(J��=��g�	BP�%	�%	BR��	BP�$BP�%	Bf`�%	BP�����J��(O3�(J��J��(L���(J!(J��3��~x%	BQ���	BP�%	��(J��"��(J3�(J�������(J��(J��"��(J3�(J��J��(O������Z��3[2��oy�P�%	BD%	BP�&f	BP�%	�%!'���%)K��|R���ﻱ�)��s�R������UJԩwm����wo@�y����R���w��)JO>��^JCk��mT��*��*���m���{��JR���߳�R��}�v���菊J� T��{�7�)@k�7j��Ep%;V�<@����8�)I��wk�JR�߻�)JRy��h]��+����eX]��/o%v��˹��)��ڌ�w<��m���q1���*]������m_w�m����w|R���ﻱ�)��s�R�k��R�B ����*�������$�86��n�����v�鍠m_w�m����	�UjBU�
��|R���ﻱ�)��s�R��}�v���/}��┥'n��ś�BEwQK��O�6��n�mh�ﻵ�){����)<���y)M����ꪈ���BJ��@������R�����R��}�v<��<����)JN <E�N����t�cM�V�>��-Җ�j��\rkA�`�6۲�'YM��0cZ��ˌ{c������"��2E+)��ϭ��k*v�:��;gtvM�䌬u�*��<�й+�L��v_n�s�!�T��e�Tݶg��vcnf�s�a��̣`�� -ĚIxw�����4u�ƃ]�9-͘y� %dV�چ�mg��96�=��͟f�wGH�f����ԃ�ڷ���g��m���5n1���cj+���M�����gn�o9x����+v�8�넫���%)~�����)I��wc�JS�{��mh���o�6���f�Ir�"�ֵ���R��}�v<��@��O~����)=�my)J^��w�)@k�ګ��\
�Z��i���ܭ�┥'�}ݯ%)K�~���)I�{���m}�ثh�)B�v��U�iJRy����R�����R��}�v<���/�o��┥'�w��U�$�V��m�v��g�}ݏ%)O=�{�R���ﻵ�6��~]=�U�V��J����Y�m����N!;a��gZ��1��� �ƺ��Y[�����]��͠m[����h_r�s�R������R�R������)P5����K�)wQJ�v��m}�w��9�'!G���JL����)y�{�)JR}�{��)��n��"�TIR�ch@�7v��JR�߻�)O�$�~��R�����6����7DXEU��wm�Ҕ�=��┥'�w�JR�{��8��5�ݶ�mk��mT��"�6j�kz┥'�w�JP��~����)>���ג�������)����6E�#�H�e'NT������ny�{��,��t��f"l��SL�.�c�JS�{��R�����ג�������6���v�����F��\�T�U!.�mh���x6�����\R�����c�JS�{��R��w���@*�)%J��mh�;��R��}��y!�?J�4R�w��@������h]�WJ۸�K.Q����6���v��������)JO{��y)A� �>����@��x���r� ��)U.���
y�wۊR������R�����Ch�wm<@���{R���[[d�fM^Mj���\s�y͘A�����tsg��nLE�%�H�*�U՟6��w����){����)>����R���zch@ޮtE�QUXJ�v�JR�������JRw��ly)J��_�mh���x6����{R]JE+URU�6��w����m}ͽ1�ɱ%��z������^6��}ӻWuuʒ�Z�*�<A昚�}�1��k����@�9���e	��YD<:(�%m^Zx6����Ҧ��*B�Ԑ�f)JR{��k�J���w���)I�����)��n)JR|wW`з�����6S=�6{3��ݸ{#jN���vۢ��@��'� �c�F����iK�~���)I���ǒ����}��m!�6���޶�mk|�l�]�Yr�r��@����O��i7Z�������)I����%)Os߻�*��m^<OxD�B�Wu��i�ڥ=���\R�����גʢ��gwՍ�m[����h[5��@D�Q%]Y��o�I�%��z��JS�����)JO��v<���Zho��x��6�?I���*�	������=�~)I���ǒ�����)JR{��k�JR�#, IA�y�Td�@�Shpm|X>��&�	��Y�I"Xz= 	�� �8/6R6<��" �|E�M�`�	�H��oA�J�0B�ؠ�頒H&`��ij!	�*A����'|� t�� ~����6� �ϒ�ԒCD�R�D�L�!�4xI2h5��L|HC���R�4���	�@D`�8�,�ddM�mu�_.ꪄ+��@U]�-u@�T�Zj��u������:56�-����g�6%ܲ�Mۆ�5�UT�J�I�9�%�s�����b�v)UWj��j���d$�cC�R�ee�T�c�2���UV���+�=�r8f��]��9j�^^�:@4��UmPKn��H���^��0UWj�YYn^fƪڢ,dz�:A\C����Lr�	n;r9uX�0�U�ƞ9vm�M�������R
X�X,8t�/�b��Y�ݪy]��[D�3�l�j��֣��69�iȘ�����0��̗s�C˗xp�ۡݐ�\�ld6܈�n�m�3�)����ٹ2�Z�^wD'���	+���V��Yrf��U�1u����z,З7<`a�����R ҙ	1�Gl�;�F�6� �kI������	��>�Z-B��Cc<�P��	�true՛k'k��I�kr�b��՗̕�S6m��cqٝ�cgE���oV북��(�\Xȯ�)�`�49���+Z�1��mѰ=+��s���WF��`�Ξe��ܻm�Y��tЖy��KbŶ�9��w;�-���:�c��)3����\i�[o�1ꔤ�>�,����2��v�m)�·W�RPgts;�5��9�Y��tjC��`�j[�|c;&��'*��j���;oY�k��<�:whAC�v�U�D ��(^�㍃�ݥe�+�k0d�C�80R�9��u�/vQ�t�Kv�ۃ�eo��N��K�{����� CuEY�;�q�i�$�JZ���7�V�� %���i6�v-�B���A�f4/i ���vv����dʠc�04@H;�+�=�1l9un_����R-�d��[��.JP�H,���MB6�u�mFH�^V���*�Y�+t�����h	nN�]ju*8/K]@U]J�v��\Ke��duF�)�i�oww�׀2���P8���^�����E�:��{ث�ެٳz��MAХ� ���"����l�v�
-��$U�2���k�rs�̶��n8׺pn��D㌳��cf�6M�n�{Z��/=mŹM�Tn�v��<����Fn�w1f��@x�5��n�v���oF;H� s��W@q[:]��=���N���ݰ�@Dg�u3b�t= =7B�k�<���z��m�ä�77VJ*�n�N;�����ӹ��,���d���R[6�h� ()�%�ڲ�_�i��ё^T���+TT��mh�֞�m}��s�R������  /%)O����6��sM�]�^\Y(�KYWv��h\�{�@������mrs�XҔ����c�?� !�O��~����*B�Ԑ����m]��m���3߻�)JP��{��)��n)J]��+nBI��T�o�y4�!3��|R���~��R����kɦ���z����򩲽wIe�!wwx��'���x6���6�┥'��v���/}��┥/�~c���1�]�rc�8�J�.��[�>�pY�l�޲1�γk����X��؇pn�(UU��ms����5�ݶ�iJ^��w�)J��v<��/�gz�)DJ�D�uf6��w�����"��;D��K�w���)C��<@���zck�H��'�"�(��%�]��hG{��mh���x4�1A����ch@��m����;�I.P�R�U%]�h@���v<��<����)JO��v������{��mh�Oz���.,�J�����O��w��@��1����Ҕ�����)JP���c�JS߻�?��ė����<�Wa���`۞l�$un�ܺ�vkm�7����i!Ԑ%r���R��}��y)J^��w�)J{��_�/�N�mw_�@����J�r�U\D%U��hG9ݼI~hpm}��i���;��m]��o�186���U��"�(����hP����JR�{������D �`�LT�G@R}��m����wo@��t��%�!"���UWi����������5����%)K�~���)C�{ݏ%)h�t%�R�J�	*]�mh���x6�%���}x��'���<@����1��I|�hˢՑJ,-�pVN��p$�DGny24�n�^��p���֗b,����\���mh�;���l����ǒ�����)JR}��kɴ�qv+ڑK��)Z��������y)Jy��┥'��v����wo_�I�@�4�������D�X�ʻ��@�����@�����$?�2R�����({���%��T�n��UJ�j�.�ch@�w���R�����R�?w���R���� ء�"������8�6��oT+n@����U[x6��{����(~�{��)��s�R��wv����$�q��Ǖ\���!Ug{u9�ם�N��Nӌ1�J�D�"k�i�x������WW#�(������'���>JR�{��8�)I�{ݯ%)K�~���6��&�� ��(UU�y)Jy���������߶���gwՍ�m}��O�6��7B](��P�����6����h�=��┥��v<��<�]�qHmz�M�HEUa.]�x6�������(~�{��)��s�P�� ׷޶�mk�[��r�T�aEMo\R�����ǒ�����)JRw��k�JS����R������������W	"��Yp��!ǢŶ�p8
�;�xڍ�㳼�9�� %��	�R�]'i�d.^�^۴d�:�����]�v��fF0��ѓ�#qvێ�n�g�IV��.uq�m�CLIsm�w<ͲzGW�;V;���t�]�k��qΖE�Wrp�zy{l�����A��ptS������ɩ
c%��w$��c���Y�;! ����������族��k����Ӯ�|��f��ځ��c�3�[�n��̶�[V���}a��������R�����┥'~�v���=�~�Ȓ������)�����IR�]���x��5�ݶ�_�FC%>ϻ�\R����߶<��<��ck�I����(W�@����U��%)O�����({�{��,�����|��M�u��#�UUZiy������%)O~���R�����h\���6��	���A.�R��2ֵ��%)O=�y�)J? ���z��mk�����6�>�v���o{�~w���]u�mC�׉�v�8�n �����Xs۲��gͺ��qt���へ����)=�{��)�{�u�)J��v��	�"��)����)J_���E�UXB��@���v��Df�����ǒ�����R�����~o�M4�t6���_�B�IUp��]ch@��~�i�������)JN���y)Jy���qJR���ڗ�yS	EU,Ue]����I1'�����)JO���k�JR�߻�)M�O{�i���9SM���UV\����R������R�� �����┥�����)�w��);����UO5�,Eӓ��8�&�a�;elO�wi�m��d��z��8�����+��%)K�~���)C߻ݏ%)O=��8�V\����߶���;���W�e���mh���x6�O=��8�w���*�����*����PF���"T�ܖo�]X�#�?UW�����5 NsP���)Z��WkͶ���`;�� �M@{�T� qriv]fhY�v��wo �m���޿��wذ��Ձ����#DMD�`�O�'t��<�q9�u���9�u�AF�k�턮v�̇x�2�7Prj��r*���~�X���;�^�Kj	���prN��Z���r�{ s������I�����l�k��51�p�ʰ?{�� �9�95�qR��6m�]�n\D�����NNw}x��� ���X\S�� ���N���]���M�(�v*������k �M���ޯ�R �9�Q��+6����+rZ�����m(F����5/Jm({z�
fJO����$j�RG`s��Vw6� �s�^I������`���K�2�mYw��H�*@z��@z㘀�8�~m����mU��?~d�V������ =q�G�~��s�H�ʐ�MiR�Г�Ɯv�ꪥ���9��,������INWwՀs�<V^T�T�����u������_ɦ�����;7߫ �ov���Mu�6І�����|v���+u��܎����V�������kHZ�u�\�:��v;YܻQ�ݗ�zv۲�L�D�d�}����v'��5��C;m�$v����e��\cu�9WU륜bbNV�r�QhE�ޮf�=�6�ţV�W.ń�:���F���݋i�y�\���XQ��ٜB��n�hx�;���ѳ7����ZRZny�3{������������r�{��s�����M�t��h9��a7�i-F��N��H�W@�ﮬ.��{�������`�P�Y ����UV��;���I$�o�x;�ŀowqg�Ӑ�"�T���d%˻� ��ڀ�8����s�n~73?eY��Vff���r*@z��A�4���׀�{�J� ��
K���k�R �9�95�qRҥ�	:�����Ϋ�깞l�k]6ܧ3cSIۣ:�r�u����i��}�X1�lf��9������H	�`��^Ԋ\�IVRU� o{���V�LBFT~XEpU��oW���U��<X;�/�U}�$wڼ;���M��tU��w߱`ݽ0�i�!�� =���;�'��t�"Dr�͚X��� owo�����N���ŀo���ȉ]\D����s�x�N{}��;��sf���zz�J����Bf_dv�j݃iy7���jX������uzN���z����e��B�&(�������9܊�͂��b r����e`Y���UWx����Ϳ�$�Q�߯�vo�V nf� ���"n��!�RM�V���ʼ�~�|�(�|b��A�W�T�[D~�6�a������q̽8 o��޴h�v!�H��#��"d0b@br\D\ؐ#�=�M�T�Lh���z$Bn�a��t����<�1]hDڧ��8 �N T] �( z���<Ө�(�����>������ 7��HEUa
��ɶ�ϱ }'ڀ�8�:l�͙"�TU�*� 7���?6���k��ݮ��OŁ���`ni��le�:���L=����Lb�^�'��5���'n�:fVM�8�#�.8&�ut�ܝ7߮���0�;���M} ��׀w�t���IS+3M�76�͂��b �M@{����4܇}��������f��؀#�P� #��]�%�).�Y����M7'�޼��b���wە����$B!��h�:md�wo 4�UR���Ww�{�T��6�������~�[�>��*Dc%R��4��¢�E��]&��=�2I�x,�E�
���]~M�Ŗ^�!҆m�w��\���� {�����9u`�҈�J���,.���4�n��w}� �n��8��^Ԋ]*R��EJ�����s��&�R{}��7����������i��c����jw}��{}�Xӝ���M4�������ty�	6�%D��X��X��K���|��� ���X�k��$����Y%+�EiKU.����9x=��.�j �]��@[�-�$\����Q�^�� ]2��=� =H���\h��u�ip���<b�m�����+���s��/I���϶�dT�v��Fbُ��S�N��Xl�+�����V L���h�V��s�qtX��i�92��J��ݥ��lܺ���\\�\���sfĎ�t^��5���_��}��5����8q�z�=����n�=��zr6ݼGI����H�;��I�"�
��#���9X���`�5�qR9 ��a4��ͽ/owq G&�=�*@G"��sW����n����R�D.�(UU����R9#���[�b �}��
p�6��*प�X�M�o���9;�� �ݖ;�u`��DI%JD���@z��@}UU������9ϕ #�R�QX�P�V�A�K��Ri���2����4�.MM�m��]�y�:̇�-fy��#�P� #�R �9�̭��ۃi�WM�I�;����ThX"p� &��y��Uw�����`un:5�	6�%D��Xȩ {��}U_�U����@s�*@v�"l �8�(ӕa�T�s},��^�;��?$�S���o�'��
Q�I$���`~�����po�� �se��Zh���EQ%RT_FP�cU�h�@��tb��AQ�em��k����
�	H�!�%����X�4�w6~�&��o�x �{��C�
�)*��9�@�5 G&�=�*_W��Uv��QISp�`���͚��U�=��͂���2�s��IWxi9=���������UU|�s},n׭G�v��i��c�ps�H�� {��������������s�-WU�v�n(ݰ��&0T0d��B�;��' �z:�_绺���1�+��76�������=�j �M@{�T���"l �8�(ԅ�s���UI�}x;�ŀo6���I�o�'���(�$�X�},w6���I{=<Xs},�L��H��CrK�wq`ͽ0�wo��M/�&��ĩ|��	��߹������C�*�RU]�y�� ���w���}x����?6������jȪ�k�K��H�Q�����![m&��R�n�^��p��KHQ��Bp�s},s6X�n/4���\�����n���R+�H��l���@��s���� {�����uG��u_�U!�����b�;�|�K,��9ĒǊ�Z%	7M�(�+I%��ӜI%כ��[��蘭�IWv��$����Q�WJK�!�$��͎�I-���$�q�Ҵ�[�ߗ�I%���4.�����U�.���.�ӷZ4��T�,�C�� ']B2�� K�c�X���vVl�/>����tAt�JNَ�;���i��Xۦۚ����� ܆�nJ�>FN����.z^�+�*�g��Cgsl�[���]��gj{9��p��kgi�6��Wn5l-�h�c�%U��y������:W.Tu����h�H<�x�Ӭ�+e�337w�����_k���»n�\]q�J��G&���b����$om1ێa�z��������Ƥ�QAI$�^���K���ZI-��+�I%כ��U�[�&�BJH��9Ē�=�V�K{���Iu��i$��l�=UU�6ҥ��	����L�I���/��I���d�ɦ�UOn�_�D�k�Ҵ�Kp�[�@H����)<�_�I%{���Y$�~��+��$�kqLI%���s�$t0�5Q'B���n�I-�ڜ�Iw�+I%���s�%��[� �Z��^,�Z�k���']���\j�g����%�:s�{1%���w{�WӾg�a�WM�ʙ�%��������Ē�y��I%��S�I,x�U�P�tܔ9.�L�I���}��&���iܹ�Y�I$����Iw�+I%��E�����9\�Iu���$��I.�ۥi$����q$���k�J8���Ud��&���i��������M�~�2I&�7��$�[�n�I*�7@M����R*����$�kqL�I���K�i$���?Ē����I$����IV���r5@� ���ZcoH[� r֕��lv��zϫ�y:H�BB(���E%��$��/Nq$��kv�IowI�$�q�Ҵ�Kt�[�XH)WU՟}$����g�m4��%����$�k�Ҵ�[ܽ9Ē:��&�Tq	'#��K{�Nq$��n�����FRA&
B  �*�������y�������I%��W#��£b���!;Ԓ�~�V�K{��8�]o5�I$����K--�RM�)(�G)ZI-�^��ﾦ��I4��{�����/ ���0�tb�(�[sh�c�`������#���<��:n�^���X�5������o�����6ovV�+vy��@�v�`]Fy�_%��5njv:�U����s�ݙ���r��IU$�K��\�r�v��o;za���R��X^�'`m-7H��@"��E`o;z`����{��5&�LmZj&�x��I4���r`�@�a ��,��s��$r���-9�,��*kDj�R�L(��&���Ջ���,�����M��^oli���a!:��܈�w���xܭـo;zy$�_ �{�`{w�\s�8TlUt�S�u��Zs� ;��@9z���ꪪ��[��lRTH�+پ��;ך�w5K�{����"l�����k����o}0��K�>�n�ʹ�S��|�.���PH�]�Yus $r���-9�H�r�YU���긁!���5�h$��:F�Y��B$U��)��$82� S=�(iN@b�+���Q}T��#<�=cbI%�`>g�т�4%��}d_$��Z��{����p[��lpm�z�NݙE�h�[i�%ޝOS@v;teq��öcC�ˡ�t+�6]��q���m�jl������A͈\v��*�vؕ�]��U�ڪ�`d�U�(�Pq��˳�UJ�=�h+��.�\"ګ�����WWV�n��iXd	�sh���d�L��,�j]�Am��jR�20MTkn��v���xm�G;]-�7��vv�y�d�A��G>t��\��%XŁ��c`z�:���k2�s���v)Wn0�ٲ��F�q��κ
c�=�2��	���)u����A.��{E�eNd;.kGO	��3>��&vѦ���ǐTdX �Ż�q�lxjeT�z��k��H�Tc+�ہp[2�ջ���M�õ{jIi���;{y�)���m���n��ڱ��U�Ã��,v&pV8����vzSl�\b�$6�N�s��'GI8mػ��ڽ�֍Ͳ���nK�nwM;(�k�sm�C]t�=y�ٛ�כ �sہ �"�	�2W;%A퇗�n��-v� <7/+��l�F]�7E�^�evX;'�<A���l9m^��%>���v�ֻOVk9���\��a�ƶ�3��s<rNz���9�u��)�o8ڪ��E���%���dySv�\�2Z^2�\S�ӑe#��mҮ�;��kv�^��C�y�,��^�^�[v�j�u�؁V�nK8�zB9Q�m���By9����xtE���L�sΟ81�ɴZ����ӒX0ͣr�6�[��}X��kWA�qm�f��p�rݚt��Q��Tݜ�aN�;me��w1m����v�G�C6�"��t���m�K��
���ve��Wd�e��m���Y�na䫫8����UY�5��Ɲ���
[4I]Zaôו%�u�gf ؕ��&FU,�Z�V�#�\uۭ���A�ǥt���^P�َq:s�-�BI�f3�v�ky�V����;]*���U\�`�Q�Q$ _� 5$�i��P����U��rYT� k��*��ܡ���I��'0tP��v�7��l*��v�[cԽ��qּ�B��-���e'rvyk$E�f�v�Ӻ�q7�M���Ncm��r�7=���.�힂���,��+��G�;Z�{J��ڬJgm���3�5,��x��.{Y�<u�1vTN�&3�V��l8���6&���)u����a"�Y�ǽ����>o��t�0[��P��1�tҶ�G�:�OoW�aL�ksf�`ب�E�o�� �wq`�wg�I���{��x���"��S����X�۫�y��7{���]ٞI���=��rB�3B���@s���	���c��������ͅ*�+��IW0?&�R{��xf�Հo;��?6�nwoޘ�|U�?��F�WM�Bp[�;{���$�:CP�.�f�V�m�tg�����gj�99�җNkR�۬�!͎����v�S��}U_'j�m@m�)��G�=��X;[� 7���&�O���V�j�ה$B�WJK�v`�n���\i�6ۻ��������韛M9.��<�*H"�qX��%�՛�������=�`�n�QЀREH���& '=��Ih>��߮�|m��^=�(�EH�(��������kv`�t�����~i%�^G���n�j�j��Ϋ�j��S�,s�&���v�НͷJ_����*.����C�}��ր'Hj�ɟ߫�9��}��2$�TQ	'�owI`uf�7��0v�f~m�{w���wb��,UD�/�6{���7��0�4�I ��UU�<��r���2��mIMTR;ꯗ�oŁ���`��Xy���n����`����!\��%��y%�	�V�:ܘ���w�����[-�t̾쾴V��;Kɭf�ׅj^�®���n���'mu����?;�`�ⱺ���V�:ܘ��{<����A(�@)"�I%K�7]��ɥ������<�����.����uu�s��X;[��6���|� ž�Ԩ�����&��`w���t��wk�km�����, ���!�&
��I8�;�K�I�G �- �T%�a��6����\s���c�i���7>�u�k���٭75��.J�lUtؤ'@����`r8� �Ih�:;��6��3-����`ssn������+ ���`un�g�M�{T.��@W*�I.U�v����xy��rv{ެ��b�>�Y��JHH"�qXy-�x�/{�@z8� �Ih����,��ۺD�T�:�u������+�n�yX{�M�.�T $RQ5�����eע�y�ų��:�d��뭻+b��C۶s�P�{�{b�Nܛm�'oi�Ī׮r�g���v�4%���КmjxB׭���[�鍧n,s�[]n74�uvVx����۝[�w0�-��ն|q�U�46�����n�5�X��]&Ig�[�^�+�\-ۛ��9���C����U��ڪΒ�:^����RE�{�m؉2�5�[8�g�^����j�A��poCM�h;ke.��'��\���*(�*Q)�{�Vc�V�ͩ`un�Ԩ������JIVy%�ܭ@u�1�"�]R\C��B��N+ �ͩ`uf�9��Vq�34�S�%A�[��9S�;�}�G 9䖀r� ܸ�qm��T�;��u`~��͞��w|� ���`m�[��E���F�{kg�ᰋ�sٓ���q�W`4Xխ������h���R
_4㤔NW �~��mj�ɈG <�.ՙ��{�
��`y�W���I6�i$���ͬ��Hy%�@�̠,7n�����[��*@s�- >r���wH��TQ"T��;��u`s��V�:ۘ�*B�@�.��2��wi�Z m��[s�*@QEn����#�%Pu)�S�����X`�=6�+��۵����3Ř8Lh�˼�@Iz��nb�EH<����Z��J�c�Bd�N�w���R���^�;�̡a�^e�WWXۻ� �;za�n�HI�+i�û�/ ���`�e֨
:�uWw��H�@Iz�������U����D��B$)��,7uK��b�EH�@u�*]J�+on���ݞ7c�ge����ˍ^�.X*7[��=���G�U��`�tP�"T��S�ug��I ;�� 9%���p73�Q"T��;��u}�6f�}�)`}9��6�rފn�$�
�ʕ%�����@�j�����t3Rn	��#p��W�U����~%��~��*��W��|�|�2

���F(&�7��K3w�S��&;t&9	�:��v����� 6�j����W~��Va�hz.���]�v�۱���ـu��1����}�k�۳z:�;_罯��󭰢6ܔ��O��� =� m���9�	�񹴂��8�%�`gri`��,-�v7v��U�$n��($P�
i=� I>�@z㘀��R�� 	Z�����$J�ܕ,-�v7v��v���M)7w��Qn�.���n����� =$T�|��+P��� &�4f���TV���T�(�Z:v������Tv��.^(i2D�c��:����磑~��Ų��'Lv�ƺy���λ&�-����Y;;6�<�mJ�^�bB�W����M����T��۷G-���^no�=���ɇ�w,P�+N��]�n��7I�Ѐ���ĵ)�ΗH�7i�Q�gk�+�����o6���ZI����w�������Cvm`9/+�)�>�1	��učm�q׫l(�D��B���E7�RJ��M0���>�ݯͤ��9�{ /j�$�)4 �$n��R����`swn��M,�j��ܕ[���W���� �wqa��m&�U^�����T�;���t��i���v7v�ݒZ nCP}& 'J��V�FU\RK�k �+v`�I%����{��t[��9��V7>R��D�%�G��8����=Vr��dX�x��tv�{� 8҂E��8���X]������%�	R�J�ܢ��v�y���*�=�u��%�x����d����� ��P~���~�ʾ�~�ӽ�Y��ڐ���]S)��K�wX7}� ���0�i997|� ����wE7DZ"U�*K�X�I9���Z�O�m�@y�� T���d�T�������vVf���u`s�9��֕!��$O�R��TE�<n��l��v�=��K֔6ݝzy3�����{O��rB�n�4�>�����fmՁ�{�����vf�t]8�n�p)Ǹ��qR�$���X��nb���_�76����/�⤔NU��~�8�����#�����a���4'b|p.D1��,k�A��S��<y��!1ą2��Č,lH"p�ۈ�j;3[BG��9�1�X<��8��P��I�*b	�%p!ׇ�����	�$���af&Xc�A$��#���C���8r#��c8g��M��If�V�\�"_�1�%�2�!��Xb�12�2��`F`��
�`����&g�sn��Ae�>!���tFc�h�mC���A��4h	��S ��zΉ�f;�2����0�{�2��`2HLE))H��!1,,���A0IH���E��!��6���
�>T}D_G��t@=�&�~
#���w���۫�`MiARHSqXY�� ��v���Ł�Ӝ��� {����TP�"T��S�:�5��۫��U�ř��諭�z�K�r5J4�0�^�z5��m�5�8��t���u��z0�'N�*H������������=�`};�U���k�=�Հ߅?/ȵ%�iI*��=�`qfm;�3]��ͺ�8�v���i��@�8�,�X��nb>�UUw�|��>������� ��n�4�>�W�}K^��;��Xܭف�6����U�n�m,�\�m���v36���W�}U�m���/{�;������>j��EI�QATg';!����>^�O/`���@��K�<Þn�ʁK�8�%�`s�uXY�N���k�9��Va��J��)�8��{���k�M�Tl�~����Xܭ�� ���(��"D�E$�`b��@y����-�nV %]Is+ ��*�?6���X;^���ݩ`uw5�f����E*n4&����&�?�~���� �ϱ���ɂ�s:Q�� uFL��I'I:m&�Ѐ�V"EUp�Yr�@6��h��8+q����s���6H�t��lK�lQ(�؞��탳��-s�5��u�Wk�-	��v��v}�t�g��i��0+֏��㱷}�6
�9�`E�=M��nݻ,g�P}%�w/:����7�XY��.2q�L[o	�ƁbϷ;��K�CBl��νQ�n�f9����j%��.� ���4CP�2�ߝ�}���.��0�C�ݤ82v�R�X�l�A�yH8�]q�k���70����۫��#����b��_�~�U���K��:O��b�m'*pY�v����M@nV��2���e6�SR;��u`���U|���T�1f��܂�
_�I(�� �d���X���1��c����	HS�9,,ͧ`z���ɾ\����wvX���q�Lu%'%$�Y,M�L`;���mu�7lUn5GB{z�
g�Y��J*(T�j�RJvz�U��ͺ�wvXY�N��U��MҡR$i���^}�xs���Q�*��k�zX��S�;ך��J[[D��7JIV����3i��UU�RX�|�������z�q�E*�*'%���������>��� t����󓍈i���9O�b��9��V����3i�2��Z$�4�������[N9���)t�/K�;\Z^\m�f�K���~��_G��8���
jG�;�� �we�ř�������1f���?T.�$�V��n�y��IHrn�V���`w��?$�JCtпܥH��Ur�� ������é�m$��iEG/�� s����j�%�DRF�E$�a��<�;��ŀs������vҭ݉5J����A��fM0�4�;~��M�*�9����m*����"M���%D��i�8��8v\o	oE�f�s:���Y:7(��<b�ێY5����}��=m��v9h7�@qV�=M8ۢ�H'�ř���UURFc�+��Łν�`s7]98؆��Ӕ�,�;��K�{�����vf�uhq&&�|Ԏ������m���� ���� �w��[I�i ��\ԛ� �UM �(��������5ʽ���k��!HTJ)�{���U׻�|o���ɥ��fm��F���3�/Z�F��^Mi�;Yt���T',I�rV��H�������H�:!Hq��:�}N���k�9�4�9׺��Ԟ�EE$)�����_9�7�@{�K@zە�ҭ݉5J����Q9��ɥ��+va����۪���*�6o�V�#M���КQ���^�8�6�����`s2i`qV�=M8ۢ�H'�ܬ@}_��g��7���-��P�\ ~�}���5��o7\v�u��v�b���Ud�4�;vw\`u���Fw��p�룜�_���۶��=�v�6�f竝�vnv��C]]�t&��+y�=�ً�e����@�Y\�sY^��R�A��ez��9�i���%�tn�p�[&[�I�����`vm�)��u����֧3���D��ڮ��o�ēqD���̇9�KJKM�{��s�m�}s���_����}%�ri��&�Ϯ��vw����MY��=���\dq��i�x���?���ɥ�ν�`qfm;3V��8�I��O���̚_�URG<��@u��b���祙+B���*�E!`s�uXY�N���k�9�4�3	�"t��"G�ř������KR�OyX�䟐��	)�������`s2i`s�uXY�N�0
3V��UU>n��c��lfj��N�S��5���v�%�z�r���F�D�v3&�:�U�ř��\A�7���Q�z�n�:n4&�p�9�%��Wꪬ�jV��1��*�P���H'�s3jX]�vz�.��q����n����e*E�Iʜ����}��ݞ,u� �f԰35k�C���&�}���d���d��<�5��b��^�/�]u���pX����G�t��9��vݫ������;���Q(�8q���<�5��gW�9�4���yY�)8���p.f;�٥����~��H=��z���"H�8K���U��o�/ x�(Jʓ���K�4�2wr��j�wlL�@���Q���ɥ����`���?$�_�U���0D/߿!K"�Uue���vIh�CP|� <�U`QEf�k*48�J�S�gh5���Nf��j��gv�ϛ�ں�7<Y�`v�n�����CP|� <�T�����n��rq���[���' ś���!��b�9;�V }����)�OR18�M�n��H��������f�,��;�*{P"8�%�a����wެ �������i���4&�}i��Wݿq`�B���E2]����@r���1�����XQ��S��Hڒ�2�K�$N��#)r�NL�ڕ*ڣu�[ny�mt�R]���f�i��sn*@z�L��_��`v�İ=J��A1 /�j�NG`s3n�������s�$�U�t�КRJ�9׺���R�W���b�y���Ձ�]ѽn0E
����<ܭ@u����qR�$���_�N6St�t6��8,����ͺ�9�ݘ�{��-�u!&4 mF�m �1p�\p�0,����$�fd�H�#�9�� ANb�2c`F`�i�c9$fc��i�b�X9X-���z"��ip�	YHR�t���4-�M����zA$�@�2�If&F*l 4)�L4AdJRJc0D�p�D�	�p�a1A��BA�`1�K��$�2I��`�HICDc`��Yca�����K���_�� I N���/Zn�����:&�5��=�+��ڷ]��:3�v���,���\��]��n�j�fΆ����,��\: �ܶ�J:��˳.�*���Z���YKF��W�
���ٙvx j���Y�2�� ����v���K�W�i���eX�V���9"��T��8ҍ�R̠?ʯ��Tᖴ4�V�')/M��t<�/=�v��ʴ���8{i3�m?_�3(�tdW��T���W��.^'b��.muU��������k[����W7Vp���5[G䲹q"oKl�}�H�ZFqH$v�h��l���a�]��m�#	e��l�D4�u�ۘm����F�1�<<�.��8���um.(�kUq�s�5��)��su��v�&��lvQ�qݶ�S���v�ggk�\i+g�k��:�l+&�>Ę��z���qm p*�i���/]���!�  ��n�v%�P�pͷ+��ƶ�a��{C\��lNCC���:s�M����\j9g;�m�r�,�#��]�iۮ��Y�k���v㪀��f���^�K��\٤��Qgs[n���Д��s�M�w�|�i�ǂ*�8���.�C���֔�MBm�:�h ��0T�X�pOc�����QsFG�.Ϙ�'G�9�ZoY�z@8�`kN�{�`s[@�YN(6�h�Ռ�J��&pL�ۧҠ���E��ns��2S���pMW���M�#�-�l���=[{��6�O���&K<)μgp��n+��y;csp=`���T�$n�Ԟ�Ŧ-׵��\�0�Ѱ�D�r�mlV$�nA�M�UUWBw^��Z�9���XP!�mt����s�n9g-��l�qeڥV�Q��;ca zu�Jx��w�幵Z��XX]�rȴێ��h�[��q;sd������F�fԪ��?}��uUi٫(�v�W�s�D��ѻ[K�+UA�  fƛc��@Iy��m�f���������ߙ�C��)�*
x|�y�D1�� b�:E�|��� ���vzͭ�N�.Ō�f�e`�*aM�T����H����������#^ �Z����rHrEn�Ix�ض��.s�^k�B2�=v��n5�ı�M�ö'ea77c؋]Y���=o=���БݪH����ث��[jS(sWZT�F����������.��Lg��c����Usў+����w�����6��]-ɚ!����{޽��ܮ��q7\����^ݍ�x;/�+\]�׿�}+I'L��lH�;���N"�t��Q8����Ձ޽�`�ږWw]��ȕ=�BB#��[y����- y�j������߿$Ӑ�إ�r�d�.�� sw��Nn��$Ԝ��,��z`�ڭD��$�j�#��:���fmՁ������i99��x�^��J�B�*����ŀ~m���_ s}��N� ���Z���t���1O���u�|9��%s����H�y�u���5�v�v��<ہyw�����1 y�j����۫���zڔ�§��`��_��IO4���M���� ����ڿ��Gw�u���7L�CiHN�~v���}& 7+P˙B��*ꔪ�W*��6�S���`��� >�mK�s]��ȕ=��NU�����j�9�7 =*~�>߅s+��2q�����Sp�ym�1)`K�@���tv�=���}��fg���U��ݬ��qy���6wެ ����F�bJF�IR���k���#����:��v��%���wbM"�.��*���ŀ}9�X|�V�I+=%E�� Ls�g��Q՛���V��)�S��BiI*��}W��������1��ķ��)/�T�18�]������o� ��Vw]�Ώ���B�r�^���0�q�d���ӬZƛ�c��9�v��rG��q�󓎘�2���}V��9��Vw]�����37Sӈ��&�+�u�}��Y��M�rwެg}�,�v�"T��	��J'*���րw����1���u{(ݼ	HS$q�z��Z�|�[�v76�6�m��tWwk ;�6�T�$��ԑ�Y����}��[�;s]���n��DD�:�Ls�	��xv[$�<��rj�v�z0�%�8�Cv6�N+��@z8��rb�9��� ��ݢ�:n:RJ�8�u��������u~� ��_�R���N����V���a������b�93�v3��N:cl�`� ś�`z8���1 ��Gp�Y�U�U�ha���G =}& ���v�
M%i&�G�D�DT�vYU��Y9�� t=9,?����L�y�6��!�m�d�j��5<k�/(�8�����9�v]�f=�N:T�'\,E�K(L��r�ݟRv�M�i-��ǝ��c�n�W�W��:��j��iM�h�Ƨ[<�N�[lq�ezX�O���9��j��,���ф��}Q��:p�ݜPK-�����
�{53?�{���w���������X�vw(z�,�zM�n2��u�9�ұA��ټK�s�Ї7[5�NV�}�����`uw5��۫;���$Lt%!L��`b�k�:��@z8���1 t����̣�j�RG`uw5��۫�������`m*�ؓH�������۫�������a������!{�Tb�M�CJIVw]�������k�9��V�m��"q86���؎g���j�sa��<�n�O]q�k��2O<s�e./�WY�����9��s�*@qwu��Z~Rq�e+M8�,�Vcm��M?��o�`�������;�Z;�I�M�dn;��u`qwu������{�T�� �7�o6�}W�����m�@z8���Sh�1Д�H�1w5�X� =T���1 孼�ڲ�۫k��d��]��peC�/�n�:��OoW�"�k�6(�J6:JH�5$vVf���u`qf���@ww���*��i�D����wn*@y䖀<��_9��R[�Sb�M�CJIV:�U�y���.����9���~�[�����Հo��X ��kj�����ʹ��:��@y����-�ŧ򓎘�)U�i98,�;��RݒZ �sPtS&`�����,.뱻,zb4�:�N���D�'�����ٹu/��W���!�m�dn>��]X�������1 ��u��,7/3M��ͤvIh��@u��qU���)�H��JB��qX36X]�vy.�����?yX[��JQ��REH�Ia��RǛ�`ww�V:�U�tI,�td�E�4D �DB1(J�)��SCM2%�4b�a2��q9�}�vҬ݉4�_*�*Q9��ͺ�9�ݘӽ��99ݬɴ�[�x<Q�ض�N�n�Tg�ێ�N��2^�:/+-���&�1��猛��r��g�w�m�>���� :��@y�� q-��R���NI�`qfk�:���fmՁν�`s1i����E:�cN>��؀�qRݒZ���BKf�	����`s3n�u��3]����`gp����6�"M9V;$�����sn*@J��UY��HUN��;�5���݆�٧�E�	���h-Ãe	���pqlH�nY���i�D(z�5M��;e�����5�B�i7I��]Xykd��fB���*v�铭��H��H ȣ�TR�����	]�p� ��[�-�N��[��gZ��b`�< �a�d�U��X���ѻb���!��P,0��'�z�r�b]��q��q%(f��[N����3����{�������Ͼ7}�VaFZwa�������Z]�%�ܣ�:N�%kۯ$J�t/m��tכ�~ }5��b��HvIhn5�$�T�$�Ws]���;�����`��`m*�z�B]���� <�T��d����1��f�B�u
��WH�.�`y��;~��:��|� ������Ԁ����_*T�4�Vf������f�X��V���5�:q��U(���:���)�#5��m�����q���"+�nb��%�M4S��4���� ��a`s�����M�hqn�u����o�=M"D��
mPع{��u�:�5�]�vw��)*#mԂi� =}& =m�@u��qR��=�"��%!CR8���,����u`qwu�� k"$'"M�@u��qR��b �sP 7G�iUDT�T��BuQ�"�����t]��Kgnh;k-n�-�y�\�@�=���������:��@I�Zݢ��%$�����9�����v���ş� .���T�GUaD�� �� ��v��cIX&�Hi���|���!� 笸J0Fa��16)��3�|g#j;��<̈�[C�:�^�Uu�hݫ�i�x.��[��G�x8�V4l����ٳ.h,ؚ^��E�;�F�>@A��+�6�L�^DGϻ	�Y"qf%����H� l0��J�!�Ya'1 һR0<S�$�(�lX�N��F"'��C+j �p�W0����>L�4'�`X�[$&��~���� �mqd��	�KN �)��)
����A��������HU����E��x�qP} C{Ͻ� fn���O�N:M4S���rp?Ϫ���}����H���<��2��(�6��!���ͺ�?���[���w},������52�IR'({b�NX0�p&GW�R����ss�v�GK���tT�����NU�w���9�������_qw}u`w6��)7BR�����:�L@y�� �����m7Tw��k�R��ww�v~���7 �1 y���c��{v*B�*M9��ͺ�1fk�fl���đ!��24X1��I�H�۶ٲ���{�)<��T��U�*K�Xg{��~m��7}��y��۫ Ҋ+4�YQ�Gň�p6lέ�Z���Iͻck���]g�����B�R�
G`��`qn�9��_���V��+�I�HN�ut�Uw����?�I�swذ��� ������[����6�;��f� �f��w]�΍VV�ID��iʰ1fk�fl�8�u�~���wwܫ���H�����I�s3f����>�w���`��miL� ! 5����Do2ֶn�ބ���˭��˺)�ۄ�7X,\@񱞨g�j=�p���\�4g�gG��qS`q<Ç[h�:��e:M�v�x�n��,�nFT��\�֍(	̫���n��8� X[�{m�z��M�C�ӞFY����u�+��:?Čc}�qlv�9���Y]k�Kb��F&']4Q���Ѷ]էM�̲D� t���!�Y�{����6��~��CЄ�W��Uv�Y���=��A)JN�nV۞g�]=�Z4c`T��I$�<��]��ͺ�1fk�fl�;KډD�I)"�����Y��r7}X��^����:��V�m��t4��`b��`��g��U�]^�������+�c��B�R�w�����1��?���\�>�����'!:)��i98W��`s� ���@{�8��0�t��nu�p������x2�y;\�O/�~>�g��ގf�kh�I�Qm�Cn>����;��`��`uwu���ek�i�)�k7��^���"��2,�"U��k�O�mrÜ�/ ��X���`s���T�%!QI$��͖o���� �5�X�y{��]n�^�������� �5�n;)i�Q(��%$T�r;��K͵��_ɻ��99�X�J//z��pO�`�yڮ��.݌�vJ�Cӌg�ط[�}[ar�]ch��ۓ$�Bm��~��؀<��_I�7�@Ky3/P�T���fl�:���fM,���_URF����'!:)�6���w;���U��o�/�ŕP^|�T�v����V킈Chnf���}& 75��b�um��J�\�.�����~M�;���1g��fM,�gқ�H�l�N��rk-�[�>��ۉ�����b��5ێt�s �R�j��*'$��9������9�4�:���kĵ���R�7wP}& <����b �sW�4�5O�.B)%��.U�`ݿ�������1 �%��e45(�`uwu�36X]�v� �� � ��P,��ܠ�����J� n; �f�����������������p�͒QT^%�s����.���6Nm��q�n���[v�׫r=Ju���KbT�Ӱm'' Ş�<�� wI���@s*D�^^f������{�&�75�������3k�DN���R��K �f�?��Ş�;�<X�F�������K �f������d���U_%��K�z��Q�(U �9����߿WH�< ��j �sPZ�M	��$�e�Uը
��]��Vp %3i�N.Z�a,�)��.u�yc*�V����Ŭ��$*�Ҭ�'d��4�um��leu�{Aʺ��S��h���<��x���&=�6:wn�Ai�\�c<�E�˓�r����V��/hHj�^��ml�\�{L�P�u?���8�F"�v)ի7gH��t�P�+:UuwUv\���wr�i�4�m4����]����������\��p����n<!׌q�l�����X�%�y9�k��<H���A�H�D�|{�ŀw���9������ Ş�5K�	�CQ�Ҏ�����:�L@y�� �[əz!EV����ݼ�����M''7g� ��K3w��N1*l�i98[��@y�� �sP���}��b�M0nq�̚X{�,��,.�34���DԐ��p�������s�mÐ��٤��\���vo2��F�zA$D�:�5!`uw5�36X]���� ���`w64�Q��
(�'#��W�}��0Y!��WS!10�� ��Si��{& ;����b��2����t����@z�L@y�������1�j%J���NG`s2i`v��@nj��b�.��?e��U����s��������{p6���(8�I�@F*Q�bd�X�\hn[�KHuq�k�����YK`��f�f� 75��1���s,�߿)(��+�rp�����{_9���@>�������ЅU]`w�����am�T�m�����M�i$���xf��������Ӓ�MHX]�v�͖w]����]ݿsc^�c%U��`nj��bt��|� >���0g��U��z[e 8Q��7�yչ$��OoW�"�k�$.Cv:����`�}�	�*@u󘀖���[�d�E ��)WWs �n��&�jCӻ�`yn��ך�F��D�����M�*����`j��g�����=�=��, �gkj���QU�U�`y&�sջ��=��Ly��-�6�J&��k���~���7���ws�)TIp��nx�O�:EH	|� %�1ۿ����r��n��BqˍQ��Hm=���}����۶nX����a�lv��n*@K�1�ng�~����<�Z��^�F㤔NU��������`o^j�9��V7 �t�QT�������	��<�T�'9�nJZҔ�(U �ԑ�ך�fEHs����1 ��izU��[��8�V36��^����7Ӡ�p��9W�
*+��
*+���������
*+�@(�������� ����(���
*+
���EE�EE�����
*+�����
*+�@(��� ��������
*+��(���(����(+$�k;� K��0
 ?��d��-��d  P                ���  }�B� (@  � � Q U ���P(�U IJ�(�I�  P �*�H  (P�   aBI   *�(Š��}.}�ﴻ��-{�nד���y�� �����Zz��������;���p����һ���}y5��'��[>�}�+� j�qn��,�׼Α�)` �{״��G��zy=Og5\  >�((�  @� �U.��x�u;���<�^[���\ۥ95��}��Z񻖾� �zzr{������ɯms5v�� �.��=�u����  q
  _@P0 ����^,��Yד�g����*I   @
X�@}Jd��qj�NL]n{u+����׽�髋|�R�M� a�:nh D �  @ " �C@4�t҈� "P D���
 �4  ��)@�J(�(U �  � 1 XҁD@ " ���R��  � "Pd����R�� w��W.�Χ�c�  ڼ�T�eWp ��n�>�&t�S�w�y�}���z�ۍ�϶�_v���oJw�}TRT   �P���ն��}��>�{�j�4�9y+� =}x��nmи��9�Oz��i^����}S��g��  ��:}����� )�T����Ow�^=����s� n��'��O&���z^���'��Ol�R�  E?��S5R�   <z�R���  D�*������F#CS�BQ�R��   ���IIFA��O����b�����?�=��xs�����+��aATWPT�qATW������

��EO����o�`�ˌ�	�!.2���?�����6���nT���&�77��� �HKp$�C3&K�h��7��w��7u��c�^�����ŧ��ySMщP{�_c�v}�<UN�aw�J�:�#���.O���[;�p�-�A9�d+
�"A��r��
Bݦ�j���sYr�La\bІ!0�eͲ�,
�0�������j����80H(`D�ދ��� �#��s�J1-�����q�(a��kG�zp����n��y����Yn$��{�^Sdi�D�8�`P�K]���1M;+� W�>��}�����"J��s�#��am�.:v��#��.j��S¼I$)�Z;`�����q4;
���H�:��	R-�X��}O����-087�p7;��aA�j��}�n$�L>e��; o��z�x��1���1n�rr��
����q�7�L�˼���	Jm��e>�>�C�_��fS+U:�>ͪ/'޿Uc���J>�p���X��X�r��{�R0!���4c�F�Ͻ�Ĝ�a0�)\p�!rR�$7��;�ϨF�0�/�#75�F��!Ԣ��X���Z5i����p��$+��Ja�Q�ih.�����@"A��F��(bJ0t�S�	��@��(āC�t���4�h�
�R b&���m�OΟ�q�����l��K��$���qц�$"c�ؐ���W`$���zbI
a�B���%��m,�0�
R��xD��"�z�Hu��A#��Li�0+���s�&ΐ��ٽ��].�^�^s[5	 �Y��XI*D��a �����e-(Ɣ1�8Ztq!�s��٩	����5̶!!-p$�"�P�Y �Y
��xH|� ����˔ɒ�t�}�����L�kf��'���op;&�5�`]�`YB6]�@��I @�d��MoA�bB�F)��
��^�0��/� �p5�B\�̙\!�.��a��XM8@�x�,�FH
a����M�p����oC ������������maS[���}]\��c
����S;�9l!p���\�k�>�7
�7��ig� �/�%�o��4�+�9���}tF(aM3g��1ѷ�hb����k�Y�|�����0���4f��۶�J�������H߈�
l��7�����gsLM�	\HP�&���4���>	Hdk.ύ�)�}��q7�c�a�D&��'��j���,"?,V�+�`B
�����
F!��F���f�Д�6���a��#H;ֶR\Ѹa�B�m�L� �cHm�d$X��c�S��#e`F� �$ �+�3N�m�"��f�p3q ��#�Ɔ�6����WA�l�ς\�1��H5�	�p���&��1�]��D5�.yB�!�~�ܬ�����O,@j�R	#�J8ġ��H}"HD��ԆIm�%� Y�8���F�4j����ӏ�H�!(5�ƍ�1�B��"G�"P�����hF��+
I��Gf���`S�3x1�
j�(B�j���d�ݺ��:X%*4�B�		�Le`HЉ��K�7�Ks�B0#$����!�N\����,�9)�g9	55�s���|��R[������!�!fo]�5�2��J M�ÌbDH�,h�	6��RB�	e%�M,ގsi��j�dѓ��7���G=��><�^<R(T�E%G��e+���<jB�瓦h�åW�0N��4�Б�������6gu~��������y����qt�揀۱�P"� GA!�F�B�62 i�3ZhF�/��/6�&L��o{H�1ѽ�B�c7�ل.�iO�4K�ֵ���7	��]����w�vY4�&]�I���m�g6q�F�k{�Jf�p.�����,��2�6hcL7���F����7��٣�Lt�+�tƤ$��lcL4ơ
l%�m�F���L3CB�7$�+�aka7�i�5�qas9�Î����̚�r:6���f�1��D�湷rP #�k{��9x��^�,z�H`�4��D�����'8o�,-��f�5�LN\��6I�:��B� �v����5�a��"a��ą4:-6BH�H�|Nh�q�6 Wawu���i��4T�Ƅ�C��$b��!�$!XP�Q���H� L5�kF�i�8����U� ��M�n��B�P6B�B�oE#H������8|;HW�k[.�ԗ��L!BT��G�Q3Fؕpt0�ϡdt�	�)�h�
���od	.�f.�L4�>pÌ�hr�'9�qX3�1�S%�s4@Ѯ	Lѱ�8}����4R���cfVk|�
l�k���[~wC��	�V+@�G�37ɲX�:��kF�1� C� �C��D�Vy��e��;��\e�뾭f��V�d1�"�@ X0�$S�X�)��P�B�z�\Ӹ��01�a\!p�����B��fk|�
c��T��7E�+��M�jlښ�D$��E�<@�[8C��hBs�h��\4;���V�7�]=�|�U��sda�ս��>��ѽ�gXFC �aX�H,HH ��F �a[,V�T�0W0 ���
�b1
$���jY%
� ��6t�F��q8!S�bT0��� �q�qA��kS�1j�"W�b�@�jF� @�bH+ b�"ŋD�@(�b�@�U"R�H�+VV! 1 �L ��L%��P� �q�0 �bC`��@�b�%R4�cP��#q��V�#��p՗3)Kp�f��y��L�H%5�K�{�V��5�y�Ui��W��[���J������t�b��?(��?.��6S��N�Sڬ<�Լ�F��Z+AW��f���,�-tnen�YN��ｔZ
/��:��?PQ�I��ԼQT[���v��;���y��˙y�]ޣ�ux޳r�N؛��+����������p�����T��o��Bߊ�Գ�~��V�y���w�aTZ�3���|6��i2E�D�@�g�O�}>��X24�;'�(+�FH�@�E�(�`�F
@x�*,�Hdd,Y��V�-��7��v�Lf��$��n��{�����0!T��-���6���,H�sAH��T0��tm�!H��i�8��bH�dF5��5�vB�# "m`E�&+	
qb �)��
��e.hM�!Ͼ��8�q�Iv�A� ��$B�V.C!a��,i�"M��4��Cf25����E�ύ��d�
�	7bZ�8�8F,���!\
hӛ8|�������"ILi�Nl��D+���p���	%0+�Fl��0H�����>��$#�M�p����HBD�
�Z��}�� �浽�ښ*�m�B�0�t�á�`B\������������ݷ�wov���UW�UUP     ���    8 8 ?�>       Y^W��B�q�큫f�qFh� 	�m�[[,���F��on��'^U�ɵ�'Nkj�TR����0qn+�ڌ�UE󋇝���qR���!�m�jmH  $����   � }�π�9n�\ְ6��   ����r�(� ^+[�Y)yL���86�,��潵��S�|��0e�SJ�L�+���R Nƅ�m%k�sLu�v��ą�"�hl8��I��'.׷��j)���M�n^M/k�;'.M�q�e^b��8̆g�nm�Y�v���vɹn���p����:k&�պF�N���� m�[V9�mv��C��PU���.n��mڪ�up���;$��Ͷ  �K/j�������H�tֵ�Ͷ� 8H p �m�   �h� p���p-��5�6�H  �am �`$۵J�WU �ƨݙ"����8�]���[x��� �@ ��m	6�6�m����`�q�� 86�m�nܛ�m� p  p    ��g6�$H$   ��   @ ��88[@ H V�)����A�l�U�j��kn�Xl?��v�	� -���  �b@�'6�K-�m"�$ H �[@   ' p ���m"F�H-��D� p�@  ��    � ��m�  H   �� h  ۶�    @��`  6�    �� [@ � m �   @�f�  Am%�H  ��m�r�6��$�l��+Lu���u�I��8u�ݢ�-��A����@-뭝�Y0�R�U[:A��BU��	��\     � H�    m�  m��[V�  嵶�6Ͱm��    À     ���   ����-��       ��    �  � ��h�m� ��[M����8m� ' 6�ڪU�]�y ���ɶ��m��2Km�P�j  �U�����! �m��l�Kn6�nݷ��mm ��l� �	   �m��ۀm�h ��   �����mm�I�R��88-�m�L�n� H ���$����m�-�z��� �:l,5���l�hq�T���[V�� ����@@�����u\Г�mw2 Y�L���f�����9m� r� ;m��[k�\8�Zq��]�Xv'm2��m)/+K���B]J*N[A�m�Fm���g�l���$i����æE��H  8 ���"AK�i �� 8��$l�m�g5C8		�[- :�֠F����X
���v�4� � ��NP������J��v�� %�n��.�n�z��S&�[��	 ��L��_�� �]���"Eɭ�n��#��amp�e��n�6��k�  Mk:�l�Ki��%�� m�cE����: $-�[�V[@�m��F��(�V��Z������un���m��e��k�v�m^-�zl�ÄE	IW���KT6�E��u���V�Ҝ�"��y]���-�J��D�mZE��6��*��l5t��Ҫ����� *�T�lQjۂF�  ���[d�;,�\ ]$�6��kX�!��"B�$�B�9z�� �T�cv��W��l���}�Ͷ�� ���V��WL3�W	;kf��6�Pa�����Uj9݉j�@N�<	U�U<�/ T=�n��=t �Z��u��Z�ثj�6����*�l�b��%[%����V,3&M0���*���m�9ŷ�M�)M1�TJ�T1THH*���jy]�����,����g5��,��2Z�i"�t��&�}���mt��k�흒� U�nkn��k�����$��ր9Cvm���k�����` +Y�@;�����H ���k�V�[8  �t�kXm�W�c�9%(H մ m�6�Ѯ�H�j�ٕ�nt��e��v�ڝ8!��[M�`6ط[�� �� f�Z�W9'mm BF  EH�E�]�[Rj����UV1O.����[s�dv���d�6 �R�!�]6N�l��x$H�#e�H�P��^em�P�nV�S��dデd8�̀x yy�b�n�UR	\�mp�M�v�� �q$�6�^Ѧ�Qδ�g���}�UR���:�l��I-9��lpګ`�f]�ݮ�iT
�P�iv �M����浜m���YKi!�� �l:��m&4VKj��M��`� Sl��I!�� �K�@-�ֱ�[��m&�<e�9��l� �0���H-�l	m �	�sk�$%�rҭ�6ۨ+g�tD��ۨ́�v��
�W��
Z-��m8�AΐmU����m�t�`$�m��pMU@U@U]�R�m����˵i0
&��\P��RD�ҭK��R� �Ͷ	�)M��:UURXȫ]J�UQ2v5�2�5�����װR��y�wM��/�~d��e�ම�����tSG9��������G'^��J�r��V�u*�5Pp�ΰ�[ t�I�n���ۤ�5[*Į�8^^v�r�U�e�v�,�<�EmA�*�s(qU]67*��Ӏ[D��x6�o_l8�ej�묎@V�U�[j���U�LU�<�*�y�i� �-ͳ�.�<qK]ԅ�.��h.��N�f�[E$� �Cm�&�An��vB���tx'ekT�6�Pzt�p��zW���\�T6��x-:%��� 8�[G��'-69<�j�\����@������$����۴�l v�[@	 oSk�����l��/E@�P�.P*�-���H[@���P6�� A�s�ZH�Z^Z�9���+�㗭6�w.ܵ:u� �����6ٶ�ݶh[d�}��  m�m�IoN    6�[�,Օ�`9����k��  H6�e�p8�E�J�V�  6�ڶ���[dٶ�6�٪:]��  m��/-����p �9����}�Æ۰�� ;mfm�ڲ˥� m��v���`   m�[@p       �^��   p m 4���0-�׭qͤ� ��	 Z�=J�v䅶�P]-�P6Z�{(qz�TH
�8��[���@j�J o� ���'X�MQ�� [@�"۶�8Hh l6�9mڶm��@�5ץe���H � q�	  8��        m6�$ H		  �l�Knݴ�H�m�v[D�l  �����[�R�5UT�ʶ�˵R�֛kkm�H[��^�m�!�9!�l��M@uu��$������-�M,��ڤٯMfޠҒ����6j8��i�2PVQ��u�&@�t�$�o�A�%5�u.���%ZR�np5Um����-���p-� ���M���y^v��^�r�T��*�S�ۅ6H�n��#j�>���q�� 	 ���^�5�� �`  $��mn�u�m��     �h$ ����m�,�k��	�AF��#m;9�NR��$���$N�\tU4�;$9g 5T��۲n�ۜ�˰�pٷ�j���n#�u[UUR�lR�hzN��1���m���� �l������ �Y8� 84ӛ۴�@ �A  	6� Hְr� $ 6�   � ��[@ַ�l       $  �  8 ���I�m  p  � 6�    [@���z�6��  -�  e��$ [@   6� �� H -�ijjm�� 5���    �� 8��     -�.f�C��� ��  ���X\��m,e.K�vd�[.Uk3�\� $l6�G m�&���H�m�}�}�Ͷ	-���u���� 9��
�ʨI�C�b�j�N,Hd���\�����bN�Xf�gM��k�ގ(np�z�M��X�hi��ӛ@ ���`M�j��۞�+j%\`d� 	t�]�ն�  �I٢��ݶֿ� QASj�/��D���A �5@H�*�UC��8~��GE��E�َ��!����C�� + �8Ѐ�`���4�T ���A�� ���#�x���/ \E��D�<@�"�x' P�$b"| 7��(�=������:�.�*)� ��G�%'�(D{�G�	�
���!��}�j�H��"��O�Q8��	�����A�"8"WȤQJ �N*��S1��6�5@j�`� �E�|A�*�T4��� A�DqM) @��qT8��.�B(�< �+�S����D�����H���8 
�(�� �,�8t
��`�6q��!� �P�� �$BDHH#,T`D
�G���p�(��  ��8��|�A(�
���D>���ohH|Zȍ��#"uD�E��<
=b���)��C�@�" ��qN�y��AqD��U�|/��8�'�EQ]���E +�
�A���6� �M�G]��U��/]gǒ�K$g`�Ӆ�wE*�8�)��0B׵�wm��=�>��l��mʷs��۹4d��h�ඬ�7\S��:$ƺdf�I�RBݕv�W�ڭ��ck�leI���`ѩ��-IJ�J�:����[a�ѻ=mT�Rٵ�l��-=4�pu�8�M�pk�6UC������@X
���Y��펵�1[q�3Ú�]V�5!�6u������bM���ր��iEӰ�*d��Zư��<;�nH�uUq+l��eՐ�"9��Z�ΐ�N� 6����V�o9�nN3 d�n�N���(���Eـ] fN7.{+�n�B�˺{0j㱎������s��,m�82� ���h�q�St���/j�9�LN�^0����N�l�/*d�p�vڰN0�=�Ny9��2N4���3\sg:���H�g�gئ$� ]��⛇����bf�Wt���j�B�M�':*X�K�c��Ɩ��/3N
�
�sn �j�kT�ܚ�zI뮳ǡ����Ϛ�.��LI��o=\�����1)���g�9vye�̸V�$���`X�huQ� �w#�F�^�8@Eň7k�85����u��a��d��뭋e1�;v"8F��k�rs�yƩ�l��� t�W��X�������
�-hu%�#�u4l��UK.`G�r�{��=.���6�r\M�6�v,8i�����Y���6u���6�&���J�p�efe���h�lH  X���vnf�y�f'<v�b,�F6�Is�B/&\�v��R�[����cb��)zj�! �%�& uh�
�N9�/Q�U��^�.[�7A�ڠ�0�9n�e�j^�U�J���PF$��`�n�%AY�m���G��t���UV�e6��n�7�45N�N�e�#+;���r\V75@�&'qR��ukZ�uh(+�Ċ.T�` ����"��~E &hx#Q���R�����w��ߟ1�[= V[3U�BK�7k:^FD��:t.X�������icU�;i�)ҹ٣\q�5��
r5�-.���޺��N�NwC��ǃcr�B�&۝�|��F.{���k��7���x�����Ϸ.����Qֺ����ϓ��ڧTU�:䎌7^�.�伬麕��l��̐�:�9s�\5B�2 ��P��R+���[9�\m�T3���Gl=��v{r��]�ۃl<�O
�X�����{l���������fLDL���� �ӷ��Wfee�U�z�ʵ�LD�1��+�@\��Қ����A,qE�lqh�%�;fA����:[��1�C�X�q��Z{e4{�4U:�?g�؎v��ָ�����7#V�`ovA�ܡ�Il� ��?���\�
���d����m�Gh.6U������t�^u�Q�%��L*i�\30`må�=�K`ṽw�)���dN~�
,m��<�ڶ�����"�"
��"���\��S157�����;�#@�#@����&5�A��r-�e4}�MU%lf���@�t�,ʸ�̫ʲ�0�=��k���3@�[u�y,F�\�;�#aH��8h�e4}�ժK`l��deƌ��3:Yр�56'�qv�ť����T�a.H���L+�ɚ�mX9��[����~��ɐ`n�A��2���.�fP�pKN<�@��M�zS@�)�y�n�~H��qcY#YnD��N���ܓ���M���h4"!�BD`@���L1~����@��S@�gWb���ĳ/0`N�P`{T���2��h�Z�%�s�m�4���V��b4{�名�EG�:w�u��V�]D��3�%�f�2���[���:��u�-Z��c�ʶ��:�eV�ͷ����07{ ��2����-���_)����̫ʻ��4{��&�i�3@�_�-�����q�l#	x'tʃڤ�:���L��d�Mr	���hz�Z��l���^�� ~QB b�� �>�� �����rN}���4F�������m��=��;��hs�h~�\r�dS$cdDHh���ل&�GUqVۥ8�0�n�T��`ͬ���׿�ތ��5�5�&�LN�~�S@��~�J�����������y�X17���;��hs�h�)�{�)�����%�s�m�4����ɐ`ovA��2���]�AVL�$x�m���f/m�hl���fS@�@�w����ŒD�mI�؍���COa����@�X�$�D �
��� HE	� �$F'�e=���R�.%�f#��l���m���t6�T�q�Qms���]|���0r�I�)�X�V5M��ivqRF�q6�ٓm;��9���I�[<�[Wz5֮�:�b�^�p] ��v��s�5nn9���[+OY�&��a��h�ʷ��������r�GV�U�p	������r:6]��eEΗŹ�8�c����`K��j�r#r��4�}���d�Qqm��ݹcu<'GP�Ɨ��V�sD�����[��HBj��L�6��<���gƁ�ՠ{l���<A�f���l�H%�(��0�?zҭ�"2����X��d#@�Թ0hpKN?�qh�)�{�)�wY��<�j�=G��1���!,�E�ݐ`wL�0=�K`�{n�@�e�b���Q�8h�*r��&A���﮶�.:G���2����`��"��lP��Zƈ�0�l]�]Ma�
1���0l_�[d�07� ��P`t��&<�"�8�nE�{l����}�~��e@�� PҦ��s_�����hs�n�G��.v	�c�I�`wL�0=�K`l��L�#a1�66��ff+~���=���Қ����$��YWh�ҭ�LO���3�&�u�M���q��cɓ��LQLis%����HN%j�۶�5��N.h�y���Mc�X�q��Z��h�Jh�e49ڴQ���%�57"bp�=�b5����P��f���@�X��q]jF� �ڎD�wY��<��w!�@�hDOȧ�AOʩ��<����-�S@��bX)?D�qc�X0=�K`l��d�*��ُ$ȲG�6ۑh�)�{�)�wY��<�j�;ҫ�$J9�DF+�q��B�����ˣX,�m�7��Y�NlMg��1��k�<h$#��$<���/Y��<�j�/YM�,��6H�!%�tʃܤ��`ovC~�ٟ�${~#�"�,qE�l����[t�07� ����t2��E�U�yp]�h9��6���7��=���ܟ�@]�@,�Mi��v�$u��ܻ�{�{Z��k.���M8h�Jh�)�y�ՠ^��6߿���Αh��v +�M�7m�C���w�O�����f=���4��qn��%5pڎD��W��y�h����)�w�kz���m8��C@��j�숙��v4�O��*�<���,�y(�nE�^������^V��]�@�w��cA!m�!�n�A�N�-��R[�}Us��̥�F�c�lM�@/+V��{��~���=��h1��O^��nF�E�l��;<��S���ZV�nu.D�%����p�Z��RK �v�������>3�8��+X��RH�t�mHOY�u��ˏ�M�.�QnY���D9�n]��ƞ�������#�nK��<v������uKm���l��9|��Y�xg`�n�X31���3C��u��7DhT�R=�Rݖ�Q��	�jh�8�U��B�O��( MK�֋tJj��s8��Ys!uT��<�j�����ݣL�9��:�W.U��1X�o�����	� ���r���]��X��8�x7�z�h�Қ�j��]�w33�G��z�dnmō8���ZU}1^�n��3@�j�G$PbmG"p�/;Vhz�Z�)�ػ������0R~����.�+@��J�13-=g�;�3@��V�Wr�q��1�fLm�ș@	���r��c]�Cj�l��\�\ܽ$Ҫ^9Ǒb���Z�)�{�Jh�j�<�ڴW~K�4�ڒb���M�$D "��PE,��~���V�z�h�S��6BG�X0	�%�=�K`NR[w�:�:��,�G����<�ڴ�ՠ{�Jh�j�<�ԙ0hpKW��V��ҭ�L�-g���4޻V��~���gw�y���9"C#M4d�f�:�onW$�,�+�҅yz�In��b��*p���ۉ��{_�-�f��>�@��Z���H��ڎD�.��5��n����uܵ�����)?D�qcn,�<�ڴ�է��� ��`"���T��flx˰��`�!3�]p����t��$R$#"������&b��5�e/zS6$������H�������i��\E 0��b�)ǰ���1����H���JA�J�c͈5U���UQ4����WN/�Gj�*����j#P�AQx
4 �@�!��N{���_�9d����7����7���_�/BZ8�Z>m�����;�1��~�jۨ��D�1^�n��5I�Qt�^]�����r�k�����n���&j���h[t�"?P#��}������+�cNݛn�E9�
�DJ9nAmO2�S6�	7^�S���~��V���F�/.*�~���Su�~��v7_���O�.�>4<�����Q��(����n���b��}Z~��I�ƀp�����2������Kf��\�3Wr|sϾ����w-g�w�����u�Z��~���F���M8�}�M};�f��=�6yND:,A�)�������ܓ���=�֮�ZW�2�{�0=Z���Il}��Wc|@pR3#"�jLNJ\�!F�u5��`�b�gd�r�x��'V-���nI�_]�@�@�ޔ�{��=�)^7�8�,Q�܋@���� ��j���\�]+	��6ӑh��w����y�hs�h+��D�16`���u��Ilr���L`{z�,�V�1��@�@�@=�C�*�'�E}D�8����E�F^e��fT۟��|�|E�r�O�:� �
������ɓ�c-A�m<gK��ccb���;X03��ݹGY�^��܎ս�}D�w+�E�[6�<�l�K��4��݌�ā�J�^��[#��d��՝����n�x�.��&G[�۞�&{\ˋض�ۑ���QE�E��A���Ƣ�������C�
����7eꋫ����{��w��w����橻5�W p�h���ѺNF]e�M�i���^�[;&h�24��㞍וyp]�0�DW��N��x�'��<��1{g�-�̿HbX��Cn&�[���PrO4�x�&Py[u��f"k�}��=�G��#�(16�"�o��1#�{��N"Py[u��j�'��c��̜˺����5�Q�m֟ʮw���~�~��hl��:�x�D�ȱF�Y���)-�ot��d�%�?q���>Ű5���hǄ�++D:D���n�Z���nQv��nqHrh֙J�e�����ܤ��}U_z�c��}�?�ؑ$�3��=��3;3g��Zzۭ ��f���MR!(��qE�p�<�ڴ9ڴ�s$1vw'�o�~�啔E�e���*�`{�����{�=v��fu�ę���M��}��GLj���%�?}U_E�~��g#'md����nϣD�20��չu�u�ڳzSLuqjv<�<SQg
M�0'�`{T���)-���ꪩ����2)?H�q&��?�Z��Z����{�f���J�Ǒb�����{�rO��78�E�����g��s�h����<P!m��l��0����-��R[Uu�H�y&�{�)�}����{��y[u�{݈�?$��̓3"�0N#tV��q�+ƌ����!3���k2Q��3#y�J"#Qa4=v��v��zS@��S@�X�B��-b�,��Il��07�:`{T��y�β�#�܉���)��Y�y�hs�hs��R9"��ZŘ�[ ��j���%���ڪ���uT����\D²�>�J�]���j���%�7WK`�1�W�}���p���.i[��7)]��d�]	����@$t��u�*$뵑�<=�q*�e�=�K`n���7�cڤ�r�u5�L�q�܏@���h��hz�Z��{q YUtH��y]�����%�=}"`n�����sS�J"#Qa$��]�@�u�@���h}�[���{](�Т1�X�K-��&��l��0=�K�������߮����*����<�	�#�{Q�r�5;+&�z�H�m�/5�cp8[

i�jL�ܛR8���gs�6���[�Ս��55E21H�r=�;tMm'e���خ��cnڸ�n����l����ڵe�z�s7F����y�-��ubyl��a���t7/���|z뫠]�<O*�s���v-����H�v)��ݹ]�%�Cڠ���{���x��Įm�$���%��Wi�͖f6���^}�P�u�"ɚ�my7UnfM�@^^��iց��c@��J����A�mށ�?�)�@i�QǠwu�ߒ=��=M��=^�z�
�m���9�t����`{fA��&��L�To"q�X�m��mz�z&wGLl�0	S�e�J���ŉ%���������d�"{o���b6�tflvX���t�
<iY�D�:��`��m�p�Ԅ&�ݷ����бQk����d�"`m�E�w���DF8�B�h{e5�~�Ȓ$h��W"��dҩ�@�wW��f��>uF&��'	�@�[^������߱"���=�Ɓ�3:�bX�܉'���+��Y�~��h9�����@�<R9"��N8��@;������/ �}��@�{��yKX��ҙ"Fba�d��b�u[g��]�ķPଃ1���דu��9WuyUw���v7_��6ށ�����@��F�D�ȱF�r-�m{�ffbG.�= ��4=v� �yX�ǋ'���#�=^�zw���0z�U
 L�����>�נT~�����<�@;��ڤ��H�{�0;d���,�XI3@��j�?�_�|��_����s@��άb�s�%$��5 ���ic�K�iS/6㚳ug<��Z����|�?%F8��n/ �_�z�ޯ@���}� ���-�̿HbX�PCn!��W�^��9'��{���?W%z�+v��H�4ӎ(��:߷4=v�?���w����I�zzU-�̜�������3^�n�Rn�W�^��#�I"�E�]�A"����.���rh�g�?�'&E�6ۑh.��ffs�����hz�Z�ǱDK�z4�Y����G��n�7$��q��x쵔CZ����p�|l��ש�Z6ߧ'z���ZU�L����נ}D���Awq���W���Y�L�}1uu������נz���鉊�����*���/+*����mց��+���Ë�W�z[���>v6�B��PMŠ�bb�i��:�;�=ܶ4>��ff�o���;�}�X�H��6��@�{��b"y'�?��@�\��1���@�����Bx�XA���� 1`,`1a"A�@�-McV�E����1qV(�4P>M���3�~Ў�H�eI�/ɫ��!�bD.�W"�WB<�j֟��D�#b�R�Җ����V%$>6l�'	b1�A)9Y Da��dM�&�@�R��uu�R�H�� ��3a�"�IUf ��i-��'�x���) L4B h֑2!	MUV҉�Q��HЂ���)�%�P��X$Ā0���1�BH�UM�L*e�Q�"�D��(D"�H��*�B	��<���!X���\as8�C���B@aaA�c��%eIFeb��)�w���Ŵ$ ��zv�������.�2���5ͻ;�m�8aj����Z0un��[]v�,�u�c�%i��E0���lX�7=rF�$�[a�eB��7md��5��Qn�AĮ��@;V{����v뢉m����������?>j�aL��3���a;@�UQ���=M�B�n���6� ��OUP皕m�A�"�*�.mF��k9m� �vƘ	X��!J����26��h��`hi�!�v�3�� �ŵ�;&͙��.{Hյt�R�ʪ��ݎ8N��κpF�\2"��\͔͹�%v϶�m�qr�v����A��@�!ڻ0mmM�;��`Ѷ�̈́qT�W[V�7lS��)���u�k�q���@AE�v�3�@�F]q��c;i8�2b *ƀ����w+l��t�\���ػu��`�6�C���4�.��eŕWF�k��v2
�s�j��c��ۂx�v��E9$�Ʒo*lZ�(��rlPL�fHIe�Ӷ�vK��L�n�.�MEJ�8ܷ��mصū��\��:��e����[f�ԛ;u��2sśr��K{tŻm�a�����j��70r�(�I���Np�qcs+��7��˺X�T,�gk����v�@�2��3��a����r�cz�!��'�@v�[�،r �Y���<f�릸=��7mV�n�
^ySE����@�ʃU���OY�w®���-c3+[7��h,,�;*H��UV���;�=�f����ڊ�m�����a˰9��Z��a�|X��۴�`��3KT"�yz��+��!�p�9��M�L�a��^� �c����t��[���6�5�S�j�tmYwa�<�n�-���1Lj�;X���d�6������s��y����iMO*�[UR�����*����ٹ䖠*���$ �j��v*T 6٥�K���;t��@u���[Oh3p(��U�^���[�<��98؃M�;_{��s��wv��@�M�)�Uj�H r!�y9�zt^k�zԦYsWY��4�P��tb����ݹ��pX��&���] Yd�dM��n'h4EU'T^�1��]�s�u����!�a�n1:���E��c�:^��;�t6�c.~�6>b�Z��l�e�]mT;�۱��=[<�s�ė��񸇁K�}x�c�9.t�j�n��v]ӎ.g`�[Q�OeM��u΅8�,ؤ"km��������!������|����Paoհ �&����1��7��?;��]��K�t�4�+�s���w���u$��i�Q�@�����y�h.���O��N����fd�Ww�����~��[������LDfO�@t�w��Y�f~Ď�*_jj	�E�6ۑh�n�W�^�""��h�n�BT�����G#m��>�˟_������~��Zb�i��ݺ��*2�˂�/@�r��z"I;��z�w�z�����J`�&(�p��! ��.��Jv[��Bb�����dqu�/4r�xΟbZ�f8�B�x���h.���z��빠yϝ��Т1�qh.��~ȸ���蘉����*^w�$���ZK�3��k/�ōdQdi��zsN���4��u��h����ի�$�84�jE��Y�y�h.�������U�a$�DۉG$�=�K`z�D��]-�ot���,z���-e���������Ⱥۖ2nm�j[����z;m�Kh�Uh���􉁺�[ �������K`�J�WY�b�I,���]-�ot��iV���+ߦ&j�D!��.�.0���Yl���j��*ꪾ��W�Bێ=�_U�{�]Q&��qD�$�<�%�=}"`n���j�,ܹLJ�B��PMŠx���g���:- ��hz�ZW�\P��i��g3��؟<��D�� ��K��N�gN�[Z%,"EB8�����6��@���h��hz�Z��zz:�ŒH��9x0����-���ut�o�]FL"mģ�hz�Z��z_߳?%�� ���ۜ+��&�(�K2���07WK`�1�U}_}T�(b�]�@uϳ޻�O��3+�'���#�=��4�.������x�נ{���&6���z	���V��NZ�s�U��IX�K�u��anî�w90oG�q�n�u���V���]�ٞ �M�z��B�(�qD�����*�11G�7zr�h���9vu�M%�(�	��Z���0����-��GLYt������ı07{ �7�cڤ�����u׋$���cNG4���?LO�*�?RJ�{�c��qS��c~?�(]IV���g�fl�������*��`�3	��j�˧��[-)r���N7[��1�-`��s��pV:���%�`k�P�]��|�wǝ���r��l&۩4Dk���l��C��{l�[5��d�н�6��:�-��s������>�^�#�Ѥu%�x�=�tnEh�[�&�8��t��pZ�:`X����ro{������\�5Г1;&�N�"ars�i���K4<Gm�X����SՋ]>�z[n�x�`�����ց��W�{݈�f'� �y�s�S��p�JE�x��~��3�bGu�m�hz�Zr��x�~�������� ����w�K`z䉁Q�Wf���<M�@;���]�@�[^��)�w�Mn�(�qe�y����-��&�dwL`wt����m�$�H��������͊i���w/e.ɓ4c���0������`z䉁����=��/T��y�β�#2%�'��)��TDL�v,�?zҭ�$�\�DMP�����4�CnG4���<�ڴ���Қ���*X)?(�q(���zҭ�$�@����$�@�����	�E���"�<Vנ\��v��hz�Z�����%'$V��[=x�8Xs�I���j��5���N�F�F��������G#nH�}�M ��4=v��mzG�]X7�#�8�]�ܳ\�EQ��@�6�@���w�u��J#Q!I4=v���{76�A$ 4p{�;�M�'��M�Y�(��qE�MŠx��@���ܳA�LL׻���O0��FdJ9N=�zS@;���]�@�[^�q�:��M���JI�ƶ�l�]8��ogV�н�4�:�$rK�YiĆ܎8hwY�y�h+k�7{ ���r���>�j�]����IZ�I^��v#@;�f�����{�X&�"6��@�}��@��S@;���v� �jeǏO�9rG��~��k4$�@�֕hzb"f���و������rO&��X%J�V$�`ܳ@�֕h�%z���������������p�qYڶ�N-��u�.�ևI���0fJ4º��ʄnb�/3<����=rD��� ���}f$�"1�A7�ⶽ�z#@;�f��֕k������O0��2�ʬ�ʪ���c4��h�"b��mց���:�A$�2$ێD��1��R[�$L��07~D�)?H�q(���V�ⶽ�zSd��ﵹ"���i|z��.��VkX��:ɣ�Z���P���_ ۰#N���hY��Hƕ���� <�Gf� ��3p:\NIܻn�GO��D�s[���	ȑ`[��˳�h��vM�v�'5q���ܖq�&�<�n�&���i�&�9�kx�yg!���ɰ\ &�6T	�Nd����y�<���Vn��v��Fkf��C�N�,�e�%m�~P|���.��j\4[�F��Y����h�nb6,����g������$뵓�S�I2,Dm)��W�{�JhwY�y�h�S.<x�d��ے=�{�ܳ��A��@�6�@Q
��yA�	�hwY�y�h+k�=��;޺ӈm��(����Il\�07� �;�cz��BQ� ��@�[^��t��wu���Z��?g�W�W��$h�6��=�N�$��n�ɭ���+WYᵴӇk2IJ��D���:���f��;V�ⶽ�uְ�LMF�z�Mf�䓽ﵾ(l ����H\����ݐ`n�.�`��8��(���Z���}�M��Z��%u�RL�JE�z䉁��r�lj��r��Lx�d��(��=��4��hz�Z������Q���DH���L
&�[�Fe:���z6�%�HBj��
�7�#�8�'�����]�@�[[����A�iր�:"�#/*��̬�+2��%�=rD����t�u+f	DDc�,�n-�mz���M:9�d���[�@6Z��ma5��iĠ�����"��}��$���vk����9�vFH�1�N�p0�c�I�F1X��@�i�0�	�D"S J�5�I��/�I��$H�~����S����W0��^ m�8�Q҂P ��� �H*b'DW��@p@!�xuGȨUQ:*�U4|	�{��]��v��fu�ĤMdJ9N=�{ ��]-��R[�$Lr�+�1LCQ��8hϪ�<�ڴ���%�gƁ�ϻ���"2D,m
8�AZ2�͂��l�j���7T��`�7]]���$�)2(�Q9�����-���=�zS@�}V���սD�"�FҒ��"`n�A�ܺ[ڤ�ܨ۸�<y1��J8�}�M��Z}�f��mց�mހ���\e�������%�=rD�>��p`y�_ƹ��DB�Z��V�ⶶ�d˥�7W)���W��R3���H��mic���rQ���rW76s�9Ӫ..��H�M� ��@�[^��)�w>�@��j�<�u�,i��D��wkut�r�lj���"`yκ�)�q��R7�����\����ut��u�Qk+��2��2�D׻��۽޾U�w_U�{uoQ�8�,Dm)�ⶽ޾U�w_*�?zҭ&v	�&}L�U�%U�j��{������G<��U'^0Vl�tԼ^
�`�ӝ�;Gk��VP��-؁܊��,�d�8[�c�OMr묶��/1ñϡ���!�l�\[*.����c��s\	����C	f�76Ү��kS	�u����]O��k����s�RNJҝ����֝�iv�M�l=�7c�I��u�\�x���X��)C����J�V��ɺ4����{ݹ�{���F�Ә��:���]]le�1�c�n
����hm����)s��]C ��m�򟭁ܺ[ڤ��H��)
ő�`��@�}V��ՠx��@���h�_ƹ��4�H�%"�<��l\�07WK`w.���W&+V���Y�Z���}}V�����]�@��8��Y�D��@����˥�=�K`z䉁�ѥv���5��vgI���ٔ��oe�o��ݥz���V�rl�X�+'E�3(�K�o�_����R[�$L����׊%E����֮�kWrN}����*�Q�0�b?~6���9_:�;��hQʯC"q�X��R-�mz���O�r��]�@�Z6�<OL�8�n=��������� ﻓ���$ő�`��@�}V��ՠx��@���hî�)�~1H&�6,����y)uv�d�n��#��4M�x��8u�wF��,�7�H�=v��mz���@�}V��ձ��S󉬂n-�$L��0;�K`{T���#�,�I��D��$��=��4��h��`j���b��.�TϹ���*���9�Zȡ15M�"p`w.����-��&�d{\Ռ�r(��@��j�<Vנ{�JhϪ�;&~ϹEcx�)�WE�
]>��m����������{7ޛzZںX�Ӂ�8�,DlR? �[^�ｈ�;��9�A��@�l��qq��sV��f��,{�{�؃� � � � �����A�A�A�A�����A�lll~�~��y��~�Ԛ�Ma���2��A����׿]�<�����W����v �����؃� � � � �=�ٱ�A�A�A�A�}���j[��i�k0�Z�y�(�����؃� � � � �?f�A����׿]�<�����UKM��u~���A����j�����n�3WTԹ��y�߿f�A�����~͈<����}�~�y��߮�A���}{���Z��r�*�u�q��Ct���X���Kn�ݹ2i��׵�S�f6���lA�lll{�{�؃� � � � ��o�؃� � � � ��~�v )>�A�����ٱ�A�A�{�n�w����S��) �b����~a�������A����k���A�A�A�A�;�ٱ�A�A�A�A���b �`�`�`�}:{/�sF�j�3W5�jlA�lll~��~�y����y�}�6 �666?w��6 �666=�~��rC.kR�f[�]�<������~͈<����s���y����y��߮�A����~�3/��3W5m��lA�lll{���؃� � � � ��o�؃� � � � ��~�v �666?g��6 �6661��"�������6��4��7:9�m��Ib4�/N��6�njd���p�6�c�ba�b�bθ��ͫ�!8l���݆�4as%�v�P�+[w45�۝�&�HM�R��N�*��7`m�'�Wc����N��7�d�kv9���CIr�F�v��wIz�Z�:�%-���I�Yl$=�mq��Oj2��/&����Q�nú2H<��Ե�\۽�{�X��qr���ݛoQf�*�LJ�l�=K�U��Dl��[�맺�;W=fv�?������� � � ����M�<��������b �`�`�`��{߳b �`�`�`���߮�A������s5�l֥����L�M�<��������b"?�(�C ��A�A�~���y{_���A����{��A����{w���3-Նj��\�]�<������~͈<����{�~�y����y��߮�A��������e33Vf���j͈ۚ<����s���y����y��߮�A������f�yd���?5�Bcj$��(��=�|hz�Z��W�z����i)��+2�(�3H�;Y���:Fz9�q2� ��9%��^9}5G�r"����y���<]հ6��`{� ��P�aJ�*˫1+u��'/{��UB(	�����nI�����V�U�j������(�`m�D��vA��R[��}Ua&,� �8�;�4=v���^�����;޸k�H�K$���h�%�?W�U�O��w)����0=������Tݳ]��&5��ɮ��nM;4�6�{4Wr�Y�3#ԍz(���E�����D��މ���ڤ�����cl��Dr$�z�ޯ@�S@��j�<]����k���E�D�f���Y�'���M�9�{�s@ ��L�N_}�@���@==�j�'2"8�30��+ݍց�Iށ��+��fb����;��Ϟ�$�ȱ��Z����Ur��x	�lj���JO1/����ۋ�r+��b��3�ٲ'���nNBvJ7(=���wk���=s������t��Il\�0'�E/	1dy	Ǡw>���?fcgW���_���@�{���Wd��#YU�Z�ZU�~����fj��;���@�; �iDc�(&���3�b���ٹ'o}�7$�s�����AR*���t
=]��w$����k)��X�Dr$�z�ޯ@�3�~�_��{�ⶽ �W;��Q��$��vH��nq����K�t�6H�<��D9%ٯE�D�rG�w>�@��j�<V��~��� ���vV�PR��.�+@��J��L�DU���\��Ϫ�=�L�Cq�X��R-�mz�ܯG31IZu�{���=Ij�M���(������~���_��k��޴�C蘙���[n�.ݺ�2*�V�0;�K`{T������}��qh���%)-	i�,�Q�(D׸�X�R!C�@8�G��!�N P��H�4��H;��`�C�C�1H�F�mi
.#�H�(1�#7��	�@��\"�D�|E�EMR0\��i�)KSs !#>4"����D]�����f��kZ�ff�m։ E�ke픺Ժ�N:t�p ۢ�b�%�uJ����i8���;4��.�"q����Җ�q�0�;���u�uO<����6��]�z��3���UT���caM=l���J�U9t�6���6����IK�Nۥ1��֩ZA��UJ��/R��Kcsi�Ām��H	�ņ�n��@[YF�� ���KnڗkH�� ��Ұ� ��-[Į�`6��h�L �v@-�Xl��v�li�{:�dJ�]�V(�U�Z�ȶ�jK����u���HE���;zv�V8�jS�&���Ť.v�:�m(���9�i��n�^�ӈ�˹���8�.=����<���=��8�\��ʜ�������Ӎ�An�z�-���M{H�Z�<��$5n�۬������g���K�u�GgjN,l[֣����<���� �&�����i�t�m�-�;�Vr뛈҆ݕ8"̂<��8D�g�)T3̨�,��e�l]]�y�s>;g�qġ��i���p<�@"���.�����r�-��Y�FQڒ͹c�<1��m�[8�)�p��D�tp�s��i�lr.G�-�mcq�׊p�<��Z�Ⱦ|u���ttqqd��f���:H[�Gi��lFo9��pm�Ѭ�@�v���c�ѻn��I�k���u�������6y�1��rcY�׹�v��"�Q����U�6�֢�n���:�H/V)f�c�퐼h�`���2�ʁ+UUQ�.��X�2�l����C�uÎ�:.5��q���tvc��y .�b�0�w�"��\�P!�+U8)�;v�aζ nx��fNz���!/n�Tji]�b�%꧕��V�9ݹm�ɵJ��uF�cc��+^ڇ:e:�7kemn		f�J��ɛ��nL���u��K!�tlչI�G/XӖ.r�t�#�U�35f���������8b�� !�G��k�ES�=�iB8"q֋y��HMZ��jkVl���J�D�Wqћ�vx��V�"큦��5<&Z�u���m*�gb�QͻqTxmҹ��� �7'FRu�t�;r#����M%�\�Y�lWb��ue��ԯ7�l\�ku@�۳��^��#�x�L\�ݸs�t�l���Z�媷b��nN��dӸp�6�]-�κ�n�vn���'�qj��Z֦L�]H�^��E� 5ך�V�.�&˷#g�c�v�W� �V%���D�Q�����w����\_*�i8��`y�u�~����r��������o��w�F��4�Q�D�4���@�U�.X�q31TyX�f,M��$G"IǠ_��s��S@�[^��X̉���6�&��s3Ibu�4��I^�����w呂qլ�D��8��ȴ�S@�[^�^�hϪ�?�}�~iO����v	��.r�vu�5�x�����w��H�ڍ���C�3���Lס�8�,Di�@�������@�}V�z�h�F�x�S.�j۬�nI=�{[ᾯ�;�<�~S�;>��r�I��k�nI��^�~��"����b��3�h��h�#O�&��۽ i��;�([�j
	c��JE�^����zz١��غ���;�_Li4Dc�)��?W%z��i��+N����~�]Riِ �uA�
��I�a�c��[ɼ]\��qQ\��;)s��� \�h��Z��f'���S��_����șȓr	�4y�[��CO�z�w�����8�WN���q����|h.��fg�V 2
�&!���߿MϟU�w�L�Cq�X��nD��}��@>}���V��b4"�^$��Pq��@/[4��~^��|h+k����(���F�!���u۵H���.mI��ۏc^��;]1̄&���GI�#�8�nI�w>�@������M�؏�F���9ʬ��;�#\U���M��;��o�3T'cyU�Q���y���mހy%�9���.۷�h��\X6�8��N=�mz�S@���7'� ��@��������;��������7#Crh�M�b4I+�$�@�f"b��U��Ӓ�0څ�h˻6-'mY�ݭčcp78d�X�J����w��V�5H�͓����@T�� �K4>�޳@}���$�ȱD��4
��~�߿fbA�7�~����3@I�4��qUpau�j8��l�-��u��*���s�PI�#�8�nI�[e4��$�C�m怹�s.��*������e4
��@=���=7$�����P`QJ�?6��qP�Kͪ�s{(:v^vXF;n��dۋq��m8v6��m�K����i�T��d����:<:��*���v�s;���\vl��1��qn��s��<�g�Psۢx�.؃ؔ��ucj��YuP��E�!�n6�U99#/R��miqq�\���걶�'�΋���-�2�
N^����l5M���]�P㑌U1�K*H=��}���ϗ���'��D2��J��V֖9�ԯ-
�.�cU���yw0�D���&�$NB���������X��鈏X7�|h;�yP]�E�V]eyz �,ߦ"b*��:�x��m{���~H�U~�"dc"M��O1�"���:d�}w�%��D�<z�i<i0M6������]����Uֽ��Z{�k�Ĥy(�wxh�%z����i��V�h�]����آ�2d�`�����T�ڝ�%���j:%�֋אoC�i�b�I<k'wyyz��u������D}33�������������Ly1�brM�t�ﲪ��H[�ܑ0oL��?g��b>���X�k�h������z���Z�혅�"2� ��A���׭�z�O4��Z�����3�qcL��Dn!8���f�U}3�?���|h�%z��߃�L�
��t��jڇ��1�f�iѫ�/R7�����J��N�R5y��Jӭ���~���33���'4��?�'2E�Q��篪��-�_߿g�D�,K���ț�bX�'{���9��©�MD�?@����[�a�]\֮�t��bX�'s���6��bX�'��k"n%��Gb{$MD�5�]�"X�%��ﮓq,K=��~���{t�2���w���oʁ"w^�����%�b{����Kİ~���7ı,Ng���r%�bX��랒fk5�[��D�Kı;�w�iȖ%�a�D��{��r%�bX�g�߳iȖ%�b}���&�X�%���{=�����4Km�p��mE<T���$%ikӡ�u�+6���oE��R�5�����r%�bX?g}t��bX�'3��m9ı,O���@��9"X�'��~�ND�,K����1�F�#��k��{��7����｛NC��DȖ%�kQ7ı,O{^�v��bX��צ�q? �����[�ow�������`�����bX�%���j&�X�%��뾻ND�,K���I��%�bs=�f����{��7����~�C�sثY7ĳ�02'��~�ND�,K����Kı9���iȖ%���#� 5�3���D�Kı���s��7Qm3-=ߛ�oq������I��%�a���߳i�Kı/}�Z���%�bw�w�iȖ%��{��������cj��C>N�v���Gӹ��tt�\�v�ć/I;�$�M�ՙ��թ��%�bs=�fӑ,KĿw��Mı,K�k���3�ı;�g�Sq,KĿ�O�anS.�k33Z�m9ı,K�}�D�Kı;����Kı>�֦�X�%���}�ND�E�P�&�X��?�I35��k%�kQ7ı,O�����Kı>�֦�X���>����ND�,K�ߵ���bX�'zy�3F]K��e-֮ӑ,K?���~�7ı,O���fӑ,KĿw��Mı,�DQ&D�w��iȖ%�bw��y�٣V���s5jn%�bX��wٴ�Kİ�"
5׿kQ>�bX�'�k���r%�bX�wY�Sq,K������};�뇎�l)��S�.9�P7<�s����UK�G�G)��(������3K��nۡ<��Z��T�$,��:�7:M.m��v�ȼ�k��k���z9���nSc#��E������OP=:�R��3�V�u�T���v+�G���^su�\s˱X@����n��vgS���\kb��ۃ�Μc�ݱ"[-j�w R4�0�"6�33w7^�(�1er4�����i}�,k76����R�&��j�莈z4v[,��{�'��u�b_{��q,K����ӑ,K����Z��9"X�'��߳i��7���{�����t�{ak{�ı,N����9�Pc�2%��k?Z��bX�'��߳iȖ%�b_��j&�*��2%�~����\ѭ]I��k3Z�ND�,K��~�7ı,Ng���r%�bX���Z���%�bw�w�iȖ%�bv��au��T����թ��%�bs=�fӑ,KĿw��Mı,K�k��ND�,�2'}��jn%�bX����/�-�ɩ���ֵ�ND�,K��kQ7ı,N����9ı,O������%�bs=�fӑ,K����f�\���խ�Z�iE��IŦ��4��N3�l�������'�j秦S3Z�ND�,K�׿]�"X�%��u��7ı,Ng���3�ı/}�Z���%�b{����hְ��fR�j�9ı,Ow�ԉ�b�>&��b�C��q9��o�ٴ�Kı/�~֢n%�bX��]��r'�TȖ'~7��m�5a�����jD�Kı>����ND�,K��֢n%����=�{��r%�bX���z�7ı,NwD����\������{��7��������ı,K�k��ND�,K���"n%�`*���]D���fӑ,K=��}�z���\�V�����D�;����Kİ�EH���jD�Kı>����ND�,K��֢n%�bX��3���?M\ՓP���Qێz�Mu��3��3�H�N�n��,�c���5:}�����)�'��u�2��{�w���{�O���ԉ��%�bs=�fӑ,Kľﵨ��bX�'~�}v��bX�'c�}���5K��fjD�Kı9��i�!�(��MD�/���j&�X�%�����v��&D�,O���I������oq�����p=�u�V��r%�bX����q,K����ӑ,h�oLB�f���0*�����n�۠m�����B�ӑ���a��*h@U�	�C���i��X}�I�TY��^�Rd��R���V�H�B@j	���b�P�m��h�� Z�Ւ-���,�fa�RBƄ�%�����1�!�*@h�m�A��(
�^*.*t�i���<D�CDQ�q'"k_oR&�X�%�����ND�,K���{$�k53W.f����bY� �2'��~�ND�,K��oR&�X�%���}�ND�,K��֢n%�bX��Nf�ka�e���]�"X�%���z�7ı,?�?��w���6��bX�%����D�Kı;����Kı<{������=Hò;kn7���T6�[����$��Hl�\�v�]�����X�%���}�ND�,K��֢n%�bX��]��~B}"X�'}��jn%�bX�{D��Кɣ5l�kV�k6��bX�%��֢n�ș��u��iȖ%�bw��֦�X�%���}�ND�E*dK�5s?j��ѓ	u�K��D�Kı=�{��r%�bX�wY�Sq,K��{�ͧ"X�%��w�ț�bX�%��w/����Ԛ�f�5���K��
@ȟ����7ı,O���fӑ,K��w�ț�bX�~*��P�)���?dM����ND�,K�;n�W5R�a���7ı,Ng���r%�bX�q,K����ӑ,K����Z��bX�'����?�/����V��+����l��
���F���g����w_9'������ffkZϓ�,K���j��Kı;����Kı>�֦�X�%���}�ND�,K����p�kf�2�bn%�bX��]��r�9"X�������%�b}���6��bX�'�׵bn%�bX��f�SZ�Y�S35v��bX�'���D�Kı9��iȖ?�R"~��j��Kı=�{��r%�bX�x��5ѹ�����7�����{����k��fӑ,K���~Չ��%�bw�w�iȖ%���"~��jD�Kı>��{?BkSY[�֭��m9ı,Ow^Չ��%�a��1�w��i�Kı?{��"n%�bX��wٴ�Kı? ���K�Г5s4h��-��6�^�!�s�{ #lRi:���ͩ�-9�qg�!u)r�B��\&z�����!˩��W���h��f]tj�u�^n2�m�س�]�Rh��#[���X�t]t.%�!�η`�i���KA	����<�;p��6w<�NN�7<�iM�lj�6���	.�r(p���tc[up�挱T���w�o���Mba6ȅλU��E�ֆ�4ӭ�7���jdm^v�"��ww��^����f�K�j�f�ND�,K�����9ı,Ow�ԉ��%�bs=�f��}"X�'�k��Mı,K��=��a��i�h�����{��7���ߖ���%�bs=�fӑ,K��u�X��bX�'~�}v���Q�X��b~���a��:���35"n%�bX����ٴ�Kı=�{V&�X�C"dOw^�v��bX�'�~ޤMı�7���O�ӅۧY�j~{�7���?�D���Չ��%�b{����Kı=�oR&�X�%���}�ND�,K���<SZ0�.��bn%�bX��]��r%�bX	_���jD�%�bX����ٴ�Kı=�{V&�X�%�ú=�,�dֵ\��a�U����g�O\�]7�)u�$�a5���h-�tu=�����������ow��g�Mı,K���6��bX�'�׵bn%�bX��]��r%�bX�}�3@f��E����{��7�����}�NC��T`R8qTb��PǑ2%��k��Mı,Kߵ��iȖ%�b}�g�Mı,K��3�0���#�%#�������=�ubn%�bX��]��r%��E!�2'}��jn%�bX�g�~ͧ"X�<ow������w=��,ow��7��,N����9ı,O������%�bs=�fӑ,K�*�"w���s�oq����龿�e��i)(����bX�'��z��Kİ� ����ٴ�%�bX���j��Kı;����Kı)��e�5�&Me�k[h�\�������Y�ն�����ѵ���ڙ�J7Ez����oq���~?~�ND�,K��ڱ7ı,N����?��DȖ%��k?Z��bX�{����_�ۧY�j~{�7���{��w^Չ��%�bw�w�iȖ%�b}�g�Mı,K���6���r�D�o���?֌5�ˬ��X��bX�'��~�ND�,K��=jn%��dL��k�ͧ"X�%��u�X��bX�'{�NLѪf���e���]�"X�~��~�7ı,O���fӑ,K�����Mı,�fD�w��iȖ%�bw��y��e�j�5uu33YSq,K��{�ͧ"X�%��u�X��bX�'~�}v��bX�'���T�Kı?*�}��5tkYf��P7�i�	Z`mZ��{[
�F���˺�����{������8�:ƚ������K���j��Kı;����Kı>�粦�X�%���}�ND��oq�����c��m	K�7���,K�k��NC��r&D�?{_�bn%�bX�g�~ͧ"X�%���ڱ7�Tr�D�/ݳ��.�f�kXMeֲ�WiȖ%�b~���D�Kı9��iȖ?�ș���V&�X�%���߮ӑ,K��{7!��:�\�\ԉ��%�@ȟk��m9ı,Ow^Չ��%�bw�w�iȖ%��@t� 1@����yD~z��}��H��bX�%��f{,֦̐�k33Z�m9ı,Owٸ��bX��G�߿]��,K����ԉ��%�bs=�fӑ,K���b�5�����6�9t-�\��70W�n�^ܫ:凱Rj��lu=<$�ow��7�����ӑ,K��}�H��bX�'3��l?�?�����%����7q,K���������.�.�fj�9ı,Ow�ԉ��%�bs=�fӑ,K��}����%�bw�w�iȐ_�f	"w�����0�2f\��A>���6$�H���:�H��w�w�iȖ%�b{�ޤMı,K�ѿ_���4���~oq�������n&�X�%�ߵ�]�"X�%���z�7İ?(L���{�m9ı,�?W�:�Д��������o�]��r%�bX�﷩q,K��{�ͧ"X�%���7�<��,K��;���~���/�9�������@9㗊A���G,�N�}tT>��ͳ���aW.`�v�r;5�W4-����9�hgv��ԗ���Wh��G�-���Vv�]��g �!��ݩ�gj+����\nD��ݲu�,�#�����u��Z=�دKd�.�9PT�.�[�2��=s&�(�]A�:y���խ�7D��p�[+`��Λя��n~_��R�0Ѡ�n�a���� �3��m\�),�����������e�g�)(�=߻�D�,O���ԉ��%�bs=�fӑ,K��}�H��bX�'~�}v��bX�'c��܆]iղ̙sR&�X�%���}�ND�,K���"n%�bX��]��r%�bX�﷩q?/y=���w���<n�fU�����bX�'�~ޤMı,K�k��ND��HdL��߷�q,K��?{�m9ı,Ӷ符�a�.]eֵ"n%�g�G��������iȖ%�b~�ޤMı,K���6��bX�'���D�Kı;�z�����2�ff�ӑ,K��}�H��bX�'3��m9ı,Ow�ԉ��%�bw�w�iȖ%�b w��z&�pI:�VL:)��涱2�E9�n&}���<����WW?�{�۷ϳk7,��ĉ�Kı;�߿�iȖ%�b{�ޤMı,K�k��ND�,K���7����oq�ߟ�o߳�Rc�4fӑ,K��}�H���G�)��n%��k��ӑ,K����ԉ��%�bs=�fӑ,K��w3=Mfk%�W.��.jD�Kı;����Kı=�oR&�X�ș���ٴ�Kı?{��"n%�bX����]L��an����]�"X�~A�V��~��R&�X�%������ND�,K���"n%�`qfD��fӑ,K��}5�˚���d˚�7ı,Ng���r%�bX*��W���ڑ>�bX�'�k���r%�bX�﷩q,K��d�w���I�5�f\�is�=��\����J�X�KW�u�`��:�^q̲�V�*���~oq��������"n%�bX��]��r%�bX�﷩q,K��{�ͧ"X�%�zv�5-5�ar�.��q,K����Ӑ��ș����ԉ��%�b}���6��bX�'���D�Kı;�z�����2�ff�ӑ,K��}�H��bX�'3��m9ǀ��D�����AL_ɇ� ���x�2'���H��bX�'�����r%�bX�����̳Xf���\֤Mı,K���6��bX�'���D�Kı;����Kı/]��4��������tìfF�dշZͧ"X�%���z�7ĿT�
��+_߾��ݧbfTș�?�sR'9S"fTȟk��]�"fTș�>�~�12c$�]�mZn��ɹr]��bt���N�2ZIc���BR˚�9ʙ2�D�w�[��Lʙ2���jD�*dLʙ�{~˰��ϢkU2&eO���H��L��S"gt_g�Yk1�=ߛܧ���=�~�R'9S"fTȟk��]�"fTș�=��V'9S"fTȝ���v����4���S��{���s��A��m�ߟ�dLʙ����v���S"fT�w�X��L�� CZ������ݧ"fTș�?{�5"s�2&eL��=��d�5�����ֵ�iș�2&eOw~Չ�Tș�2'{��ݧ"fTș�=�sR'9S"fP�
�*�W� �;��e�r&eL��G?z~˩�kF���\֬Nr�D̩�;����92�D̩����9ʙ2�D�^߲�92�D̩��ڱ9ʙ2�D�f���5�q�\� �q��7X�b�+\ �u�^ݫ[2\���&S����x���|�~oveL��S��5"s�2&eL����e�r&eL��S�ߵ`~I��52�D�����92�D̩�߹�ֲ�j�5uu��ԉ�Tș�2���s�]��3*dLʟ��ڱ9ʙ2�D�w�K��Lʙ2���jD�*(����G{�~�|��ғ�	�+?=ߛܧ��r��o��Nr�D̩�;����92�D̩����9ʙ2�D�^߲�?7�Os��{�ߪ�:Y�Д�c'9S"f_�P�'��~�iș�2&eO���H��L��S"}�o�v���S *�5����ڱ9ʙ2�G�ۏ��Yk1�=ߛܧ���ʞ﹩���3*dO���.ӑ3*dLʞ﹩���3*dN�{��ND̩�3*ShVw�\Hŉ0�|� Ch�8R��#��M6D����@b�"�I@x���C����kHEj�&+��␈/LШ�B�b�#(���Q��!�M��Y�
��2I$�B�-���>c�ؿ w�߮��~`z�� $t�@1�c����LF��&�I�Ӄm��A(�*��ᒭm�m�a�Gc��Ŷ؄��j�����<H��לt�=����igm�	��u�,���Q����#s��ml�UJ��cl�)GF�V�36
�ء헝�g�Z��[cF�$�mk i���cm5mUH
���W�7`6��-�)H�)�j4��FN�A��髕�fU�)�������>��keZ� �U+�U@R�� �2����)W������yݥi�*��KX�[PI`,�V�e�kv����[h���Ճ��[�<"�JOnK��]���٣VKӆAz�2c6�ƻf�nn��R�����rYfmL�\�鵭���{pH6�'N�	��C���e=`�M�"olRm�dps��9yyAW4�|!���hN�\��Wk\�9����eG�*�T��n1s��gg��km�Xn¶�U%=��öG"HݯW ۦ�^vWm�啲��B2��zv�m`���yC��G�G��2馧`�ikrl�c���-���Ɏ�(�s:�8�*`wn�`�MZR��ã��j-#�Ш�99�N�G�ɤ�Y�mۃ��&�N�wj��P�\�ct�s���J1�٫\@s�q�j"����\��
vu̠m+۬/�Q�y�yy 1m��J�P��r�N�l�n���Up���y�-�Ɓ�Om�5]�v�=�X�t��ea�Yl@f=�]C��<֝c��!�1.�.��6F���0&��� �5U��0�,cF�\=���	yAx�c' �r\:w�tF��3J<�g��9'J�������t�UYXuqdނz�;;#�ݫ����g�(�y��%Z�,��ڹ���*�Q�cb�B��y����A���;P9A��rҬ��ʆ�
��Ͷ��+ �ѭyٶ�Kb������Wz�99Џ\���0B��~w��}�;����D� �ĂA"�"��
��*EOE�0�@_���d�}s5�����MW�!^����p1�+��1lg7m�4n�qYCs�45��+������6������J�C/���d�l�-n�=��v녇v�qqM��/< ��X�<U*�m��ۖa�yڸz�3�u���q�'�ʫd�	v�Lv^ڲm[(����k:��Ɣ�l�����IJ\��fPR��j�p����w������Q�(� �n��Zݤ}9ӱ�qֹι���t�ć/I=`��e5l�&\ԉߪdLʙ�w~˴�Lʙ2���jD�*dLʙ���n��(���L��S��sR'9S"fTw������`y��eZ���{��93*{��Nr�D̩�;����92�D̩����9ʙ2�D�^߲�9������SN���%����nkV'9S"fTȞ���ݧ"fTș�=�sR'9S"fTȟk��]�"fTș�=��V'9S"fTȝ�z�]ST�u�u33V�92�O�R�S��}����3*dN���e�r&eL��S�ߵbs�2&e��"]������NOr��{��}��P;=��Y����L��S"}�o�v���S"fS���s��O���3*dO{{�nӑ.Tș�=�sR'9S"fTȝ��=un�5��S-�����܌�4�Җr��y�5�3��uEk���www����:RwA,b����3*dLʟ��ڱ9ʙ2�D�w�K��Lʙ2���j@�E'�T�Lʙ���m92�D�S�������5�$�˭\�����3*dN�{��NC��|�P��m��"fT��sR'9S"fTȝ������Lʙ2���jD�* &�j%����ں����R�]kWZ�ND�,K��oR&�X�%�Ͻ�M�"X�%���z�7ı,O���6��bX�'c���f�Me�d˚�7ı,N}��m9ı,Ow�ԉ��%�b}�w��K���2'�~�Mı,K���y��p�Z�3Y��֦ӑ,K��}�H��bX�'�w~�ND�,K���"n%�bX�����r%�bX��o�g6n�
v����Ռ���I+e��H��Z����cQ��e�?�w����j秄��jD�%�bX����M�"X�%���z�7ı,N}��l?�	�L�bX���z�7ı,N��C3����5��ff�ӑ,K��}�H��bX�'>��6��bX�'���D�Kı>����r'�S"X��k?kV�j�5uMj�"n%�bX�w��M�"X�%���z�7��V��&�0�M���ߦӑ,K����H柱������b��(�B���Kı=�oR&�X�%���ߦӑ,K��}�H��bXȢ7Q;�￦ӑ,K����3?��d�je֮\ԉ��%�b}�w��Kı=�oR&�X�%�Ͻ�M�"X�%���z�7ı,N�o�g��l֊�v����ǰ�N�ٺs��V�t��T�,���a�&�-�Xb���w���oq���"n%�bX�����r%�bX�﷩�r&D�,N���6��bX�'��~��fkT�YfL��q,K���ߦӑ,K��}�H��bX�'�w~�ND�,K���"n%�bX�x���,�kT�ffkZ�ND�,K���"n%�bX�}��m9��2&D���ԉ��%�b}���6��g���w�߻���\��U����ŉb}�w��Kı=�oR&�X�%�Ͻ�M�"X��Q���ĺ��"n%�bX�g��]kE4d�[����ND�,K���"n%�bX�����r%�bX�﷩q,K�����iȖ%�`��ަe��s	5![M�Pvn����pP@���/NDFՙWRZ�����um������ow>��6��bX�'���D�Kı>����r%�bX�﷩q,K��{�s�K�5����՗Z�ND�,K���"n�#�2%��}��iȖ%�b~���D�Kı9�w��Oʽܞ�{������G�;BP���q,K��}��iȖ%�b{�ޤMı���"dO���ӑ,K�������oq���~���زܳ��Z�ND�,K�׵bn%�bX�����r%�bX�﷩q,K�����iȖ%�bv>���fkT�YfL�Չ��%�bs�o�iȖ%�a� ��~�ND�,K���M�"X�%���ڱ7ı,H�� T`@B�ݞ��2f[u���ֵh86�X6���L����;Qʠ�L�[jl�If�Й�ڵ�6hV�P'Wk7Vzˉ���[���--�snӠ�\4s��i�<�;���oQqu̴�v@8��f�ut�͙3�qY]�۷[	��1<���n S�|�l����u�nkYx�3���;qٶ	�v�1��Vk�5kq<��S�f�f���{�g����.V�#V�/U��C�9�<k�s<���:��<��b��=1٬��kS��Kı;��ԉ��%�b}�w��Kı=�{V&�X�%�Ͻ�M�"X�%�{�{5���a�.]eֵ"n%�bX�}��m9ı,Ow^Չ��%�bs�o�iȖ%�b{�ޤMı,K��fL�k5)�&��L���r%�bX�q,K���ߦӑ,K��}�H��bX�'�w~�ND�,K�׵�e�0Նj��jkZ�7ı,N}��m9ı,Ow�ԉ��%�b}�w��K��&D���ԉ��%�b}�nf~���Y�Y��Yu���Kı=�oR&�X�%���{�s��}ı,O���H��bX�'>��6��bX�%�[�55�����C�F+��������]��MiK�=ZܵM������hJ��|��%�b}�w��Kı=�oR&�X�%�Ͻ�M�"X�%���z�7�q���~���زܳ���{�7�ı,Ow�ԉ�U?LT��2%�b}���6��bX�'�~ޤMı,K﻿M�"X�%���{7!��SYe�2�Mı,K�{~�ND�,K���"n%��2&D�}��iȖ%�b~���D�Kı>����ᚙ�3Y��֦ӑ,K��}�H��bX�'�w~�ND�,K���"n%�bX�����r%�bX7��{WkE.�ˬ�֤Mı,K﻿M�"X�%��?����9ı,O���ӑ,K��}�H��bX�'�{�.6�0������u�%�q/k-���֍X]^�Y��G\i+o��D�,K���"n%�bX�����r%�bX�﷩q,K�����i�����ow߷ړ�z71�[{�ı,N}��m9���&�X�߿��q,K���o�m9ı,Ow�ԉ��%�bs���h�̚�R�fj˭M�"X�%���z�7ı,O���6��c��O`7Q?~��"n%�bX����M�"X�%����2ᬆ�u��sR&�X�@����_�4=���)�w�;$��H�jC@�e4=���)�{�Jh_z��0Q�)��$�Jn�X��;���ǜ�7#��]��λ1�����mő!i��=�Ɓz�h�Қ�)�{U(ハm�!�^X��qv%l�x��_�LDD�.�e��(&�RC@����)�y��/YM�x��"Ȉ҅���b>������@��|h�#C�R�$Q
��J >C1J��7�s|��s��kV�a�(�!�y��/YM�zS@�e4�߳�Z��F(�Li���=���$h���ny.�Ľ����ywR�����~+c�X�$iHz�����=��4�S�����@�Z��"y�"jF�X07{ ��2l�0'L��}UX�y����s�R)��>�O��2	� �����D�+.�WJ�l�0'L�w�?}U�R���|������nHh��w�	� ��̃ ���|}U�����]�Y���	����D:@�b�c��c1��WF��n+N�zK���{G���'.q�"��9�rqF-vv`D�":,[�7	ˤ-!i�qa��]���b���7m��l[O������2��1�������g�C�MV�-u�������nGϳ��f�	��(�[���,e��mGܢ�X�٧�O�{�ax���+���d�8��*m[u��۱�۩���ө5z�k$O$��dMƤ��wY�^���,G�1?�x��ʻuwQ�F]�	,�A���`n�A�U]X��ȌqE9�l��yb4�L�G�v�ύ��|h���c�X�$iHh����)�^����M���ȞFcȚ��8h�b4�&'陘������r�>4�S@��Ҹ�6�p6���M@I�mN����� LG�A�D�5ն�d�܎%"�����<��h�����A���"aK}���`��̃��40�W�h�u]��?�bk�~x����,F�G2����0�������@i�4{�9������{�O��լ�<� Yq��4��1�~�����{��.���������ҍ��z�h�Jh����;V���0�B��p+&X��qu[A1�ʐp��{mbm�l��-+������7��;u�γ*��I�ύ���<�j�/YM�cULdqb��!�^����Z�)�{�)�f~��+[�dO#1�7#e^��Z�����DA'�� l�"HBS��2Q�`���H�IF~ڭUp�!�<�eƘ�!rVV �"tϔ���H@T��ce0 �� 9�x&�2�14q	9����FH�$BA"!���rL%! �`T�Fd�D� @`ԉXE!�,Y`R??noC>�MlYX�B"Q�HaB#T� �����)bP��@�K�Xr0�/��,�s
?L�U,-(��A6E`0!��~8	1&�V\eH�IH7��X#R5'ƃjQ^ ��D���<�=@��Q7� 0����oH����E:7���=��;֎u�71�%$i;��,F���F��b4��ycu�^ό��c�~�cN�Қ��~�J���}�:�<�/"̷U�H�.s�E1�O�leי*�cm+]�#y����JfX�b�BG�6ܐ����@�֕h�!�D}31��|hO�>�fI,��Ԑ�<�j�/YM��M���=W�'F�,��ҍ���b4wb4q1T��hV�o�Tsg��ǋLC�)���3?f~]n�h<f���*�q1��h�]:�*�2̪��̪�4��8�b'���x￧�{�)�{�8��'��L]u̻��֗��\ѭ�?>�
�uU�q֎@��4=$���yR6' ���Z�)�{�)�^��z�7E���nF��V��b7阚���h<f���*����P���B//'.�����@䱚�)�y�ՠ^��z�LSIqyww����M=f��mր�b4{�4S+��"�9$49�Z���~��h�#@�1舤P
w�!���|E�w{��=�ww���f���X�'V��Ӻw���r����g��6:4��a��!N�#�S.w���:���mQ�vC���.�����'�[��g��rf�Z�8�{A��s����6���7��59[sBYk��ù2@]����|/;�] ;kr�O<�
�7�鱺\pG]�k��NFʺ�z;vح�df�u�"�Z��3 :C�������~?�Bn5΀�]���"%Q�:�PFu�^ݪEngcՊ�j��±]q�EK)����{��.X��LD���X��ϲ}2bɓ�D�4=���)�{�Jh����tj��O#"Q�e�^��h�b4s1T��h�ƁWu�,o$!0nG�8h�Ҍ�`{fA��d��(^	d�e��y��h��9���=g�9���<�j�ʫ��6D�N,I,Pj�J�&f8���N�^v��8�c�6$9zIg�f8��КƜ4{�4m��<�j�;�����խ�a	8�rC@��^��{* *[;����I����{�)�x��\fI('$����*�,F�ɉ���K�4��tn� �c�6ԋC�3��__��@�gƁz�hs�h�̋	�(�NC@��S@�e49ڴ�S���߳��<��' ��;����K�j����qsk.��W]�<OGTV�o�w�����v#"Q�N��|hs�h����߿fx���|��8����7"i�@�֕k�����x���h�#~����]+�VyfQW��������'>��7 m�
�I������;Ț[D^^N]Ywxh}3^��x���F��b4(.���<q�䆁z�h߳33�>�xO�{��}3��w�/ ��,��n.۳;h%��aN�q��B㖙��lk\e�-����0b�IV���_�������=��=�S@��F�b��̪��̭�b7蘊���h�3@�ޔ�=넳�d�8��9�l���}15]��$����ѐU\e�yY�Uxh8���f"��~��y�7$�}�M���L1 "�� �
�`�P�U�%4
�X�ƲA�cr<i�@�ޔ�>�I�?�x��b4��V���s���c%3�b�=��{#JӤ��jg�L��б��w��Ϸڦ�*K�������̃t�0=�K`v�,�̑��!�m�@��S@�e49ڴ�S@�pj��0��m�!�.X��ZU��1D������y�x��\fG%�iȴ9ڴ�S@��S@��Z�:7T�PR*��̭r�h"y-g���@�ֽw$�ʔҰ�0����������1[��Z�"��s�n�n�����&�3�9M�a@�J㖂Π36\�QQ�te�3t���3���I�rG	��-���sŴk\�Sc��v������c �7#�2�s�]�.����tm�&	���|��NSֹՁ��<�
pG�}[ \��6�LC@��ďL�t�t�<p���؃[qV�
�fp&$J�s��Ze,η^��3 �ݭ�bkmu�<�X��c\���L+��0�1b�1�(�NC�/��}g�/ ��@�e43�5T�'���̺��@]iV�"b*���x�����䊭��ƲA�cr67��(��2l�0')-�ڬ��,��Hh����S@�e4LEycu�.dP��̼��*�.�{�	� ��)-�:di+�P�9�K���|N��b��'6��^��������r��]�v��Z�eV��o���~�J���g�+N�Rd;���%�jHhs�og�~��f~g�l��:���=�S@��F�$b�6ԋ@���?�b]���@���Z�Ic)��D�4?��b�+���h�b4��?Gv]*�*�F�F��@��M�v���h�����"�#i��a�c��#����G�eM�KC5rM�M�#��w}u������p�k��wYM�}W��] �GX�72!8�u�o��%��=݈�T>dP�r�'2�,��4+n�%���@�ň0*$R��PCș�4�;�)�{pj�ҙH��ۼ��<�#@�֕h����O����r�����J	�Ԑ�<�j�/YM��Z�)�g�,�L16E���F��B��0�9:n��{Yz�H�kD@�L!���#�i��Z�)�w.���2ِ`l��`]^VR/++2�0�=�J��DU<f����)�y�Ѣ�I5��n-�rِ`wL�uIl�*��e��xT]�]���b���@I�4z��4T�P	��U�u�F�������ѐnd�q�$4�)�n�-��d� �+����+�;6J�S�6,�-�Q����cgqU<h�E�yٲn&b�����D&���]�@�X��X��b?P$�8���"�8�nE�{l���S@��M���� 8%���=��h������x���h��U H�9cns�h�e4m��=��h�ȬB�2cQH��@ݙɐ`ñ�Il�w�T��.ؖ4��>�l�m,����/|�7���<`��#����x����0+eSCD<�G���E�;��ƉX�,$1�^�b�I�RQ0h+��%�?y(?k"��"�ҐYh:AYE7�9�X@����ޛ��c��Jg'���5'����I��B��.��{�����|ޤ�� HF�n&���c�9����K�m���n�çs���΍�n�lF��b�JTvl���r�c���e���ۚ�'g[ [L���hE)!u�qۍ��������	)�YM/�il���&�*�����V�T�q�ܡ��ݻu�*�G*�!5R�۩:t�#���1�����;F��l[\R�vVB�Es��	N�s�%}���RߺY3��V���p1џU:%Z�V��5UGUT+,�ƞZ��l�]
�ԹZ�fduUV�$6���琭����ͱ���)�
����E9ݥ'���C6Ks�N�N�aeV��%Cr愺��b^�A�VYW�Z^].�%u��kY��$T�q�璭�@�Qy�ȳ�v"6�ge�K�]�5�Uy�����&C��M�P��X]��&�g�cZ:�@�F�St�im�tӷ<��֭��o>Y��c��n�䑈�����{l��*d��N�����M�p�����k����i�,+ֺ�A&���9n���a]nr�M���U��N�jf�N��� �VT19�D�:��S�1���[b���(u�u�w#j�@<�V볫y2�m�R������s���n�󕄼�4g`���+z�JO�`�s�61n�����C�![<k]U��ysu)��v^ѡ��K�9�Oo*L�!���|WTkm���0�cp#��[���bʽ�N尽��v�u�����6�$��f��e��;=�6�xN���ջK����4�x�\�j�T&���Ԑ���Q���\pl�/n����J�"���|�����t�/-g[��[$�=�)$�T���8u��`���jil�%�t�8w����d�(=F�E+Հp�
���^��ö��U�-��� �X)[��6���lP//C�+�WTpR�c� +b��n6i�M�u�b��5�b��u\��FR�^�,�z9Qv��S�{��w{��>��W� @<	����| b��~U�lQ"���{�������t+e��v5�]#��lt H�.�k8ܔ۞p�b����	:��E���uh���׳f콨�`�i��9T�u=���[��cIq�E��{^q"�3�����э�Ouv@lEv��y��`��sv�cJu�6�6N�æו^\�.����q�=�/�к���pb�m�u���A�X^�[�������:�TRӎN�����{����|�N͹&�ͭƗ3 P��+:t)sv)�G��s˺����������7ˀH������?w��ِ`w)-��%4kT�88,nFӆ��S�1T%mց����o�1T>�W�ә�rI���@��)��11U��4�����.�s,B����06L�vd>���~�l��w�|1̋$x�i�Ա�1=�Y����=��;���Hy�X�u���1�t�)n!�n�a�v݂��js�thk%Nf�2Z�T�}gd�K`ṽd�07��)u��hɚ�\�3SrN�=�u@h(�111�_<f���4.�o�Trq>p)��E$Z���{l���t����Z��׋�!�C�G����&~����_}��@M�Ɓ�iV��YM���ȱ��cr<i�@��A�ܤ��d&A�ճ*,Y�(�[;+[Og��F.6�kt��Mנ&#ؠ�!R��H�P�s�,��>�~�Y*�?yb4%�s33���c4̊m+�Y�fX�+Yll�06L�w�4�j�=��c�H��ے$��צ�}�zn/�'��F!�F"H�M]{5��'>��7$���0/
�2���4>��-'��@n��h{e4m��=��ؤS�i�w���iV��~���9V���3@�ޔ�=�W^
bJ	�b�Ȑ7���U�Q:M/c��v���g<>a�k����^�����df8��$��=���@��M�zS@�v����Y�!�,qH�'�b7阉��9,f���Z�X�.��ȱ��cr<i�@��S@�v�β���h���B6���/33Ic�y<f��L�P +� ~6�&��ksrOwо�b��2D1�2�e4m��=��4�Jhe����cs#rG;n�tS��#z�3�l%m�n�2=DDo`=��3"�8�rC@��M�zS@�t��2��%��YX�!f`����Bl�06L�e.S-A�1�F�ۆ���M�l��f~��3ﾟu�\|�,S#1�L���d&A���r�wGG14I�c�ǂp�/YM�{�.�#@���2&e�L�����cۿϝ����=1+Q6�n8��^ۗ��̫b�T�V�s1n�jW�$�e���lirN�����42���	��]��]���V����r�9��}�u4�y.�)�mC�n,�����À�0㦱�w�(�]�����Ops��|
[n���[���n�W��4��"
�� ���\��H��lƻb���ڵ��d���t��%ѭj�&k3Z�_��>DG�Pݿ?���ф�������H��o�[��}f96�ק^�'e���WU�9�c��N���Y��Jh{e4�S@�^.��?5n9$��yҚ��M���=��4:�W[Y�H��Fl�0'L�w�	�`{v���Q�$4�S@���h�����Y�u&E۳��e�y�07{ ����d�C@�ӫ�ذID<�D5*"U	�V�(����j�ѳ��v"���%��άI	,� ��̃t�07{!�Z����qE�)h{e7�?D�\��}11.6�����<��Z�y�j`�&%�'	�@�e4{�4Δ�<�)�{Z��ȱ��cr&�4{�4Δ�<�)�^��z�u������q�$4Δ�>�z��4����J�]FF��"G��]��:�0i[r:wcq6�f����g���`��oQ��u�m�?~�4��{���V�o隡9T� E#ƣjHh_�Ɓ�t��yҚ�e4WS���r&Ԑ�'��7$�s��s�>�����8�? l@��ߵ�nI��צ�{q����#lM�@��M�v����=��-bꅉ�f8���49ڴ�S@��S@��M����c�FƱ3Ly2zW�����M�,:G����H����I�W9k�[t�07� ����H�h�88,nDӆ��t��9Br���A�ڪ)�,K>X�n9$��yҚ��Z�)�{�)�y�b�����D&��CC����/V7ZO�{��� ��ْ"I�F!$$D�H�Tŷ!s1�\��Dz������;�t����KIf[t�07� ����Z��߳�fw|/��Q,pc��N;C����f�Wc�Q��Mf6H'��x]��'����r� �mI@�}?��49ڴ�S@��U��21�F؛��9Br���A���A_D,S#1�!!�v����=��/:S@�=��bX�q��'L�{�	�`{����:��E�#���M8h�Jh�)�';��ܓ���7$���|"E��w���x��ĥ�\6b����n<�)���3���bc�d�rmm���1��l�)������
@��XE��`ˤ��[�ֺK��Bݥ���Og�Ϯ�n�mr���s���$R����[����������7+:�5�\gbO)�jϫ�d���%P�7/m�Ӟ�V��gZ:ظ4<u�1��j2A˽���:̹�5���5u��-��������ܲ
���r\��6h.�U��GE�5���4���*9x�^���f�f�f4ڿ���R[t�07� ��R��7?H��6�hs�h����t��yқ�$_��""��*̭���=݈�Z�~�J�.�7\X�9jHh���b�w�@j���ZU��&i���9�Ӻq��i�(�ۆ�yҚ��}�����@��S@yו�E&G1���8��H%ŷ���L�5,�:�5��.AZ4º��-����E! �� �N4=|@;���zX�4I�c��7���^�ڡ������p�s�%����?u�Z�wM��FTf nDӆ��ύ�49ڴ�S@�^Wdn~���rI��%�6L�{�Be̱V+�̢����4�iV��9�g�9,f���M �r��ic$I�ɒ)Cڷm��a�͓�Ձltp���^Q��v��՝")8�nE�{l���t����M�v����� �c��Қ�#�Қ��Z��o��9}����I�E$�Z�>49ڴ�O,�I��x�$��|��+�n+�t�M1D��A	����ʟ���F-�P�|&]GA ���ͨ<P��0HA�`@�	)ؐ1@>BB֑"H���ۭ�B����3�|��>���6�D�aް� �·>������J�6��i���FF[S�Rt�Q�I��@���[|��e��¡
�'$�0#�cBB��F)ʟ<LF0aJ%����� UH$���L<h��>UJ�5C��^E()������L������D�D�,�~���|hٗl��#(���̬�11^X�h<f��t��yҚ��K1�MbX⼲�+@\�����[�~�j�OW\�d��Q0���X9LW:�qƜ�F�ء��5�Mqˤy-�^^	ӑD�{�)�^t���;W�fx�����/<�� �s!M�$��Z�~�J���{��"f'�����D<���!5��|����z�h�Jh�)�u�tuc�ԏ$�̶ɐ`ovA�ܡu	��(E� P�J�R	��G�@>���r�I����f��L֥�Yy�h��hffR�3�V�h�)�S��c�b��$a���N�q�r\"ܻ�%4�n��{fK��t�M]c�cThl�G�8hΔ�<�j�=�S@��S@��7RDDF8��HC@�*�CO�rX�u��DU�Y��148%�'�Z���{�)�^t���;V��j��ȲBLLr(�4{�4Δ�<�j������������?�����H8��F�q�$4	�`{����2��0?��S�E"�#T3ߧ�j]]a��Fj��#�f�WB��9�.������\�V:@�̕��0�w�[h١Zj�9;qk�y�-��Ws^��|��]�Om���MܣћG �V��#v۶�۬d���k�p���[q��y���SE v�s�m��V�Yn�̞#V�>����\��Z�\j浑ZqYڴg�6�յN�.��mU�z$]�����Θ��	�b�@kÛ��[�k.Y�]f��K#ѐ�a�)���!�N�⨱�,�e��u�1��!�n~�	�m�������S@��S@��M��JS$ƲG�6��+@\��&"�䱚V�h��Z����4�q6����t���Ѝ?�3U�mր��h�J�A�Q&�x���yҚ��Z�)����[�_���DDF8��HC@�)-�:dݐ`NP���_ZP���d�խƗ2[D�ۖ9.�.n
/=U��ywPΛw%\�&l�9k`N��d� ��)-�9�E�b��M8h�Jl��f~��������U?PND�Lǰ��4�n���~��$nd#M��$��z̦��;V�z�h�Jhu�,Oj~�	�i�4�iV��b4wb4�!ҜԷ�$ƲG�6ۑx���fg[���gƁ�;V�޵]�$iI�U�,��<��u��m�[�����k	����b&�Mc@��jHh�Jh��hs�h���\���#�$X��`��2���)-�:dݐp�f��̫eEa�U���W����m���� �A4
��sy�c4�!���bȼ��/
���cqhr��h�Jh��hs�h�lqdY!&,nDӆ��t���"{���Z��;��e��e�1��u�=.��fs�V4��[�A4ϱh�P"��S�u-֑XmV����*r���A�����M�S�MbmC@�@�e4{�4
��hs�yVI�d�m�"�'L�{�	}.r��}W-T�4�q6����t��WUM��z�M����y��5����r>_?�drd�<I�@��V��D�}3�~������=݈�>�f;y�$J��X�̓���s=uF�p3���n�g�9��V�v4�qhb*b߀l_�[d�07� ���p`{{&c������=�S@��S@�)�y�տ߳>����ȲAĆ�%kI��tʃܤ�ɐ`x���F��F�q8I�̦��ZU�y,F���k41��ȼ��̢�����ZU�}3<޳��3d��znI�T($;�K3a�.���M�k5e`3�Z���6#S��>�&���tz-4��/q�q����91ó���/�����7���a^n��Z��n#�M:� ��`�^qѳ�S;.q�)�O;�n��F��[wn�\���9Om[<r)ʐ�96 ������'g�t�Z��Hm��m�+���դ�C��<lr�t���6{	����|� ~Q5�P�ן^��n[�b4�ݷH	�����3`6�gh+�Z�rvےz:�:�eV��݌�=݈�;�B?�1���ۭ���&��r&9!�{�)�wY��?u�Z��o�3Tӷy�vfV^y�����O�&"f*��f��ύ��R���Y"����R[d�07� ��P���1�������m��?��u����3�@�@��u6B9"mLI�&�۞���D�T�ɾ>us�N�Gu�'��Am&7$yH�܍� �gƁ�fS@��������z�ߤ#r&ff�jkZ��w���8+fA@"� �!@-a�H�����;�Z��=݈�?!��*��ƙ�v��e4�����[�ύ�r�*�1��㍶�Z�dݐ`wL�0=�K`m��ı�r&9!�{�)�wY��<�j�=�S@�ӫ�16�bQ���a�H�
�LFDkp����{u2b.5l����%������G 6H�Ĝ<ߦ|hs�h�)�{�)�Z:�X�A,qE�'3�Il� ����eA���c&	c�ǃqh�)�{�)���<0c���+_�:��S��-�_�97$����w$�rw��SH�܍���M�Қ��Zٟ�w�oƁ��~����&6�p�r��%�6L�{�q����Z5;�a�e�#7&��E��+g�v1ƛf�UF��g�����wc8��N��ˤ���ؿ~�ɐ`ovA�ܡ�>o,�1��6ۑh�)�߿dLALU�3@J���ZU�z�iYƁ�8�䆁�t����M>���=mW��@ﾟr��,�ě$R���q33��ŷ�;���<�)�4���Gh�D�
T�d��@����$	c�,�9��<�j`l��d�`mwd332�k��+OOf��I����3�M�,�g<��&L�44]�6a��6��߸��؍�d#陙��b'���@��8�����7#i�@��S@�t���;V��������)�A���$��k���<�j�=�S@��S@�U��D���������{gδo�{���LRX�h	ū�y�uX^]��ehK�c����K�I=O�RM���ܓ�E�(*���"
���E�Q_�DEj �+����+� �	�� �+Q@_�Q_�

���E

��PU��*�����+�"����

���E�PU�dATW�ATW���e5�eob ^f� �s2}p��     z�(>� J *�         ��*��(    B��JH�U�)J  �� �@PQ�T�TP     )*    � P )  F ��\A������,p ,�\f�8�.�@}�N=���s� 9x�;�AӀN�}�G��D����7������G>����_V� �@    1 �>z��)���A� >�<J�@d����C�oy��p}xz9��i}��^ ��e����P\}���{.�׮��t=� �9�  �  `=�m���� x>�
 @  �Cw��{�=z8�>ޞ&����n 4�[�ޥ{�u���]m���{ʯ �}��;���}|��_ ��.���}Ϫ�x S�OW���[�Ww���ͽ���W��u{<����}�{/���ON� ��   @!�}})˾��[t����-ٯw�}������^C������� � AAE�     td@��  H��� �: �
 M� `D'@  �\ P Z   P   6 ( D )6  �t � ((.� Ro���K� �=)����μ  �����x���ӝUg۽��=�����x��>M;��.3݃��7�z_n>ԫ���)������@���R�  �'�UJ�T�S�F� 4 ��UI6�R�	� "��d��JT @DHjJJh���P�;����Oʋ��uP1�mC���B�
���(���

��(����Q�qDTV ����a��01_�B �B_����t���sP��hL�����q%�<��7������Cɤ�� 5pO�^m 0�2MT1I$$�uS�P�1S,)�sB75HcTԅ�ɰ�]HSFq�X�>	_S��BZ["�d�>N�Q�E�W��(J��״��g�	�ļ�H�/l-S!L!B�b_���"$iL�� �%�o�#r�9<�=8|&b��dJ�a��J���F�	�|���8ٜ�]%�l�5����Ā�*�,U��H%X�`0&�F��0�,@��Ev4"�"ōS�
�$�5�%Lk��70�� ���F���dP��"Q0�%R	A���p!�l��@�C�,<��Ϥ'�s��g����=�J���M7y�!sxOL���HĮ��"�$p�0H@�L��<�-|=U�0��h
��`P�k��>���32a��(�������5 p�al"a�@�"BF&0)�F�a����A��`D��I�ل ��B�@�B,r�5 G���ׅ49�cbIL$w��IdS6�<$a�fo)ZBT%.��4L7�� ��!䄒�2����x��a��}��ệ3�_xt�^���1��E#���)7�aJ�BANq��
0 E;�2z��cBE� ��� 0c�����!��R5#B\��{���J��Z4%����d2�-�ԉJ@+_a���d����|=�_ap���P̳3s%�	e�i��%HT�]!LaH%!L�XC+ը:,`�� @��
���`�I��a��B��x�.��'W**�ZT��+�^Wn��7���Jo��}�.�!���TpZ��8{g2d+
B��;4��~�R�� ��BRS!Ik� Fԁ�������� '����� �)�0L���B�h|^o�D�{�<�ʉ/�q&c
d)�
����=1">f��4�^��O!XB沄�ˇ\�B�������OR�M$E��=<H�&�SIL����}ӏ �H>V��^xK�	=HR�c�
���zJc�S7�q�9���%%��y�)���#\t1 P�J�p5��a���0��̦�s�s�bD��`Ѕ+f�|F�R��{�E�@�,!ﻸ�s��)��K�e�StCni
�HZdY��$<J�&���=�d���.�Z�2y�=�p��nl����0��x�l�%�|����3Y��=7ƅe�$���	�>)r���3>sW
K�5�ɏ8篈K��s5��Q1)Uטx��)�ω*�Eߩz'��0����ϼ������1	��y�׼9aJa>0��� ��k
|2�+�p><t8�<4�^x�p����ni�/�C�<=�kp5OOLHQ�t�i����
8h���Y�p�!wjJK��i
�+�"P����ԈT�K�mO�cS
*H���ձ	�sۧ=8�*1�ĸo!S��=��[�̛���!o��\0��|0��D�qʙ��d��#&Nh��0�r��*᤻
g�����
��9��3|��4%eO�����
�!
a�J��@(0(b˚P�.B.�g�[InƦG*������lO	MT��I
�0�~�ȳa!XR]�J��@��#�)������t�	/�y�7�sjy��*���i^jkjBuQ�yy
T
�a/�}Ἶ�>�$����<�|�_��T�v-@���!\6�þ��F)H��|���{�9ĈbEX1�E� `b����<繡hK�Ï���eY}�Ynj����E�����d&\�3�[��Z��
IhbT��!aR%T�M�aR�4J��T���\Y���8�)���=�j@��=�>���T�@���c�!R��I��a��=1�=�E,�=��z!�<!<0�i	i/!
eɊ`��)�bF���%�c��1
<�T�w�u�'a#�Bq���a�!9.c2�a/�ω�Hf��
D�!�����B�g$&^6����#��0糟i��3����i���5�¡
�$i
�+�CI	s�|�s�I�=���Xzm�>����zP�#R*R�o<߼��4=ebG�0|�ϒ�f���BHY���}�L��O�aP��(U1����,h@dH�<��%05x||C=���Ut!s�o4�� �x#b��f���7��
SK���Ʃ�E+"S����l ���?{��d�C!�D`��>�O3��"�)�E��@���� no�o��fy9P�Hs�t������>R��#�+��$J�N�!��ǩ.q�B���FBἾ{�B{M��OT<�g��5��$_~����B��$��<+�@�7y-۞�p�ƾ�+�&��9��nC�!H`B���Zc7�y˗�� �,�H������Ć�q����B� �t�x$Z�����̞�
c�hKy�HSS�����\5�����0�4�'��A��G� ���Ks����s�n�7���F�11 ī��Vk����~e�Lѐ���i>��c
!0#��B�<8�i��3�c�0�F����.BJk�(��B#FR����"P����d�L&)���J�F�rl�������ДͤB���q!+��l��S�PōdTͩ-�9��XR��Bs7� D�-�3���$����	$�0�n�%aB]�q���f�+#-��i�&s�%4�6�Ä̀�# B��,7f����P<�3'�O�� � ��H5�X����L&�D�f�)r�^!�L8y���p 3�$�M�L�J�(���
`X���B���"¸����O]}�Ma�m3��)��{�a����l)
i$�����|=wx�z@��b1�j$
����H0����P�fCB4q���B�hD��F�*1*�Z�"���Z��
�	�0bk����	� D��}7ɆO=X�H�Hu�t�� 2&U�h1��$��(&���ґ`a-�`�=xp	�sN �B��p��oxp�S�0#�N�C�� �1@�L�[���W5���,*��MmHb�C0��GZpɁ躐�ĽJ�4���br$ �HX�ug�{�z��X��E�~#C4_]<�LN�jB�����`�1�V D(���)�CZS�Id5x$i��)qՍC�d�$x::������ c�����7ܞ}0�y�IC�BIL>�/5�eq2�m���x��|tI����Y�hR@�$	&2[6�-Z|i'}����vC��}�Y 1_�D*D(�B
|��:�+#et��S�R$ ȵ��҇�K��4���f�+�*����4#@�@=4<,t�)����-���1L(D*k�S�
e7����p��9	w�&b�@(F*B0���B!~�ӂar��$q`똒Ɏ,)q�0S&�@��t2\�`l)�cGX0� �!� @�ӧ�N?��m�� 6�  � m��`L�n�[v���+;-�eT���8[@�Cm��5�ҥX6��;��UU{J��!����-�m���[�E���W@	�KU�H4N�X�� 6,s��^������й[��v���`ږ����˹6ڣ��v�p� ��)we�v�h�cPH���ӨTծ���T��-�u�����8�ʶ�R��Ue9�U���d8[x:@�i�-��N,�J -�.�lp�� �m��5mJ�$Cm��;�Jm�    ���X0[V�my��J�s����r�t�E��K��[m�jNu�u�-UP 8�5�6�m۴����! lp�   Am������m��6[�zԟ����j� mNJ���mI8��:�� �?�}��[G lm�`!t�om ����Ӳ  6�RC`    ��M�I6�  �v �m� �[A�u�m�V��� @ 6���]����[\[D����پ�m���   	6��$�l�[A"E���  ڶ� -��t� ��v�۫Z�6탂��m���l-�m� 6�-�m��H>��m���V�%ڶ�	   ��[x ���k���g�	˖P�q&$@ � ���#m��l6��  ڶ�kgN` �ۭ� 8m����K���	6�  ���$�Hݹ��  �� ��n�m'l  m6ۭ���C�;%�Y.��@5P6�$�[z�N �[�gm��m�  6� ]6�m��6� 8 h�mq�  ( �ٶ[Cm�H��k��-��u�m m� �8  @;k��P�s0[UucqU)l�ʷO*� J�`�m��� ���ŶG� p8	�ȓu��v�$km�'I�6��� ����V�n�v`j�̖�]R�)-U)3؇�.�N٤����a�uЦ
{�u���pW\*K�J��� M�-�l�OtQr�Uut��e��C� ���  6�HN8w ��)�K�%���uN���`���m��� ��	��at�f�G`H/-�,9�ձ�mp�y72��su������[�--�G��l U2AUT�+/U��@m�i 9��T�m�Z�x�*l|Z��p��a�� $�l�U�8���m6ؐ��_H�ėm�� q��p�,�6����Y6ms��N�N�����Iz� m�]"�p[% ��m��k� ��ۣ^��ey��ۖT�ѷU]���q��c*�VIj��\�r�V� mt�k��vCj���үKu��Ð2�셨M�
�����W=��8�',�	zkܱ+�D�4����kK�N�;dZ6��l�(<ԩR;V�u���P:��3b���R����m�3Uz�q�c�]r����h(���-;`#\��<6��:Y�G;6y��Z�q���N:�����2s�UC�^�0�OAHS�=��j���m�����ݱ��۴vĮ����l��ܖΖ�k�w`  5��ݦ��l��p5mU*�Zl�7E��մ��P���f]5��EM��w�i6�7m��6킔���&�l#W��Pl���*�6���)��	e� $|�uu�����l[!�藐U窪�,n���[B�(s�q��M�� ���':C� ��K�f��[m�rFN�j�ڍ�b�m���kp��$ � m&՜e'Kn�$H�pN[@�ɽl���dhx+UJ�-J���8ﾶK#�I��`m�m�Z�i�6����Ls�U{,lg�W\���{�<�턃�p:@ �06�� m��BEU�e�j���� .:P�N�� ��L�i Q5���m�[@ � I�lm�ͻ%u �����l����p �  �Vp�%���Ѳ4P � �[@�i�   �   rۤ�mmm��c  ��m[@  ��@]5M�m����ջmm�8  o$ �m-�e�-궹�rk�v��H��z� ��'J$�plX�{IL�װ>_����r\U]���� �m&�+��nCqg����C�8Mk�����i�]k�Wj6qmJ���pS��8  �Hj���J�UUl   ؛u�-�3 2pI����K��H��m5S�����c�"�� ���$�R�m�cm�ځ����]�'Dڗe��ګ�.�Am��IS�n��-ܚ�u�I�l���g���K%6 �i�J  �մ�'I9m,�j���m$[%kM�4�+E� ��	$h���    I��h86�m)dY4�,�T�  [xN�v� �o� H�{  -�[_}���d	����y@>)��UU@mWV�mn�6�S��m�U6�� �.�$9�� 	�#q�u�J    -�,��"�@m� m�6��d�K��  m&  8 m���l ����-� ����M��RL$��-�;!�l5��s��	m�H���m�I�H�qö�����d��U�V��kD�@K6BM��-���I[5��-���Ć� 8   ���m  [\m����$H 8m� -��-Mu:Fm�	���8�[s�d�f��8iI��p5*ԫU@�`��m ��i��l    	 @���� ��Ҥu��8�\p9Ͷ� ���Ggl�T�!�ضWnj�����	�� [r9� �`�6m�v�l  ;6텺m��ņ�,�	e��=JOm�5^��|�|V�YF�V��ͩW���jk�` ��V��ڃWV����[/Uն�J:�S6ԫ�Un��VU��[k/.�l�[nI��<ְ�m�۸۴�!� ��`	$-����WQ�:� �l�      m�r�I�  HK(�    m�8p�T���٨
c�R� 8ݷ!���{kƉT�=�<��<���n��� [KzΦ���I[[~���l���M�A���1���"�]9J����X� �Z�M�ݴmY �*��*RZ��P9�t|9�"��mGCZ[Ժ-r%�mTmv��H���V�;S[Tk�����*���c�@k����ݻ`妒5�գ����v�iy��vi� /Zj��K/R��1Vg����ݮ����m h��mۓh�+�@uUH������S`�b�I#  �6�m�m��A:8����@V.��n=��N���5N��l�O�)�:�w�}��-�e�L�L���;oj����d3i6-� ����h�$!��3���t]-ת l �v z��v���ۜ�n��H   m� � ���� �`rmqmkXqm  p����  ��   ����%� 7m�km�i��[v��\ m#�����  [\;Z�hsv��6�H ��[p s� ԛn� p  ;e�ݶ  $�m���-� ��h�&ְ 6�m:`H�       �n�j�mAmlp �      �bF���pm���J�khH s�ݩ4I� m��m��KGm  �H  m8p8  �Ӱ�n� ��  p��� ��[v�g$b@ $�,0� �m�H��	�k� ����@ $p ps��	l��ޠ 6۶� [d &�2 ��q��Zl F���_���m��[�m��ԅM[m�  	m2�R�<�����hE�@-�h�l�kn�x  �  6��m&�m[ ��d���	$�p  ����8  mi��`� @�`�a�k[@	n��@�l � l�m��v���8tr�ڻf ���&ʚҞƶf�-��ad��l�8�G9Ij��5�:vڪ������ l�  �$6� ~� ��� ���UlpUU���ڴ� ��h/^�v�m�v؝
�nl����]����A/,d"^TЄ4 S�
��m�����U�Zn�uP
�+C��%ZR���l-�}rv��\��  l��սڀڶ�ۅI6�m�m��kh  6�  &ݭ�j�� [@ ��L�@f��͝�Ŏ�7Z���8V�/{�����{��T��$@���#�z�������(�7�bH���z��T�"�A�"@9@��� *��=���:$P*)�|��E=Q�x���Ԃ|�P��h
����Q���O�TtB������q|R��^���z��\ �<5O�)��������bD` h*t@\�<U�
!���=U'Ȅ"�T"  H���P(# | tD1*}z"|� @�����'���EUO�H� H��$	�@#c!j.�� �/UE� �CDt��(!�8��QE��jT���� P>X xPTz�|��1����u�Q� ���1X$("�
H����E���D�F x*�ȇ�
#�8��P�x!�T��,<T>�_���:�Ƙ��P_T�G����H��)S�� tEL4}EM�A}U��M@qT�(��� �z�ER8��|�
"���e��@���P��ys����n��ͩ9�5\�s��K�lf�<�۪jI̔�WC-�=dΉ�$�Y^��e��m��gX� �@���wm�[�v�b}.�fB�v�[����s�p�[��+�a��X��>�s*`�3dg�SXv�B�j���^�=h�gv{r'h0d"_�Ԯ�FNZ��m"��( 7-ź��pMP6ʞ9l`��r2F�":m^�l��u�X`��ʛ5�v�g�Ó=gt��v��Q.��]k���Ze{b�����J����(���v��L�p'��rⲏ*sg�8FB�7j�ۮQi�$s�[���vx�R�k[b������v��m;�������'��<�����%����"9��kk\��I��[j���
���Ʒ;D[��]*�9�۶ӜLvP:q7 ����AAΨ�G ��vs�$�R�q�kqVl�z:'���$����J�ѵ�ڤ)��&HGX�5u�"����3��ЧN��1��P�%�������Ol�U�;u]>-���m�z�յ���9�9�Ik��1�˰ ��(W��cF�x�2���/���Nؗ��7 -��l��SI�%�ܔʣ�/I:&�����;C����UN�,q�]!��q�z
٩T{vʫ*ԫ�S��s����m�J���Ύn��1����i�a;N��nƺޚ��ݗa�݋.Ҫ��*��-U�l%֘�V�z���e){EO/Wg�m�M�X,��#�s�֚�p�5�2E�x�z� ۗ�G7����7$��	x��m���h:[j�c�=�%p�F��1Pڎ�v6[��esrʵ:(�\�3�]�b�BU�<��hj�mЅ��\��jm�JA"���b5/e�v�mڣ�mtnT��$�-��@� �'OZ�J�sQ�-Gh�+ꤑ�")9#�ٙ�5띢��N&��p28ȩ�pջv�.9���Ac�+ԬS��tB��u�0�3m��p$5۸��~�D7����$�T��<1]�?�bz
}�#��J#7��4����ٷg�nKa���z:n{n�<;�k[�e,���f����;vs��,@���ڐ۝p�ݲa^�kn�dH��z��B�6�Hbz�\�h (�9�=vY:Z�	�n���ۍ[&��9I�B���rû9�cC�}�z�H�	�NCjB�*GmXw9Z�� �K��1���J��;m��ݧ�1��ֻ3!���.i��:��S��O|�����r�����vn�;��nE��eݻ �π�T.�L�wd��wS/wc�&ffM�͞(�\<T�DL<@LK�̪ ���rd�;���f�fL�uO��n��w`ӻi7�r� �u� �ٕ�� �q��i�ն	5�w��n���vG��}Qŀr�^�[cH�N��f��+ 9� rH��\0��(�T�)޹��WjnK��!���':��퍮R�l��z����9����QwͶ��}�|�9$x{��̬J	+,��M�ɻ�3w�I�{���(B 1@ ,"	����
 �� u�}����rI�{��9����X�c�V�!ڶ�����+ 9� rH��լ�J�����n���vG��<���K�X�$ժTӰm� s�< ���`�2��@�zMc] �Yӭ�k�7��e��6��Q�낐k<�`n��..:n6�%��m���� �u� �ٕ�� �q��i���	7�w��n���vG��<���P��Wb�V�3 �ٕ�$���y1S� "�"11�#�;�p�;%;v��v�v�`;#�I����+ ��J�-1Sn��o 9$x{�fm* ���̙�A����	!L)ܳ���)��������p��
��b1]$vu:�
�*k�۵c�V�!�m��'�� �ٕ�� 9$xvEj�P%v����L�7ve`;#�I��͐�X�$ժTӰm� s�<�����ɕ�oT��V��WN�W4�����Ҁ�ݥA�:�
�Q�/�%D��U~  �Jy��.1;-Rlh���w�s���.�iP�6h{݊�qk��J!Eu��*V�*����g����A�MnW��n���n�l��qqZg����������@�٠.�u��d�p��‵����;V�&���wc�;�%��`�Xω+,Iڦݡ�$�ީ/ �u� �d��wc�9�>Xݫ�N�ē�_vg�w���wc�;�%��]��Wl��0��T3$�����3#��^N��hD�����P~S1�~���i��gY8��*:�&L�M���F�H��ǬI�,͑�Qc'�Z�ܳ]����!�����;��Ɲ��0[�w�ݝ��6\��=v˧G�j`/5�kk��6�#�=bx�#S<��f6�8�Ll+/��:�WF�p�ڭ�[�3#��ك�=��$�=����F՛m��)��n���[������۰!��76xxW��ٸ�{ :ܜ�*���TDSvz���j]G2�S��+n�	-p���m[*�`�j�*i�6�=�r� �u� ��z��ʷWV��5i&�\�g�����`G� 9��R���V��[`�X{����;#�9rE�r�j�n��ڱX�ݦ`�ǀ� ������`���bNպn�m���wc�9rE�s������+�!v%��}���vz�g��\6Э�Zo�-v�y�v��і�ur��������;������X;'�c�U�L��ws�O=�{9���d"��Q W�#��!�������f˒,UWf�W���7v��0�`��X.H�w\0l�Z�*"&)�w&$��I&{�ފ߻������*�]4���j""b����PɚU���og���_�m���qɻ�p�(�����9n:˫�\+�v�9KrQ���N�މ��a+7���5�s��n���ŀr� �h�P���4S��w\3�$ɓ�o��@[�tP��([��i;V�i��l�9}ذ\�`���S� =8"�~A�~��䓾�N@�J��ĝ�m���X.H�w\0�p�9}ذw`�n݃T��V��9�p�7u� ��b�9rE����������͜���^��GR�f�)6������sM�j��t�;�K��l�a��6��7��r�b�9rE�su� ��U��I&�R����0^�Y�fN�wE{�����s2I's29��[���]4���Xo���9��n��݋ �q��ګl`��74�̔�e��(��(=�� �����(�T�f��'��6P���V4;��w\0ul��}�<�� ��ݫ��c��i4���jkp<l�k�]��b(*6�ˣ�Z�ᦋ���t�4�ݶ`�Ȱ�G�w��n��J��ĝ�6���k 9$y�uI���'c�r�"�9�)ݻ�[�;v��;�p�7u� ��E�r� �ȭbv	]�n�i��`�Ȱ\�`�`�
���&А6�ƙ�r�"�9-��9��0���UBJ���>úwi�vw3�\ܛ���Q�θ��ϟ9�f5���ֺ#I̛����2�\m����[TmǞ��[�f9�zݎ݂z3p��y�3ʭt�ۀ�[��乇u�t4�SҴ�� ��	�X�͛��oh����=B�6kv���逧p#A�,gn��:\ZM�v����}�`�e��媋�j�Jn���P�&ݐP�l�&�s5�=��93%���n��f��*�ז,=�������(J�mt֠��n���N��MZI����w��ou� ��E�s�\buv��&�6��\0�`�Ȱ\ذV��C�lv�X�;L�7��r�"��D%3�׵�w���8�7D�U�M�n�vZf�� �͋ �u� ���HJ�$�SnИ�k �͋ �M��ǀ������P�*�l��ܷ.�uɞu�^(h�m���/t��v�۪؞Jq'Oma��C�s���������32t�<�������ot<TK�d�f�sg$�}��s��h(ۑ`�"�;�p�9�k)�MաSN�i�/�,�$X;��`�>.U��i��I�I5�r� �u� ���݋ �j|�$6HL�D�P��(dɛwk�o��@}-��5BP��u4V�])�E�*�0�l0���Ml�/+k��:_F
���[���v[c�jƇv��&�� ��b�9sb�9�p�;QIJĝ�t��ݖ��y�6+�ܷ��/vx�2�t�5�IX���m�M`��`�pô���{BlH'�H�fx46B1"܄��(Qc�	HfE3%IHK���WbQ&�40eHԌ�ɠ&h@�	3B		R�����Є�Vb��J�ס#27yPP*���@��Ufʣ
hF�c��EH`I�$'7@�rY! T�$F��/�#��.*�[C�?+�8�D1��
�E�U<>DA�@Q\  "����w��'�v,�U��T��YN�j�t�m��vG� ���݋ �͋ ��Ym6	]�n퍦`�p�9{�`&ǀsu� ��vz���5v�hI���O��[�P���O8<k�qnl�P�	�=Zzwb���ݫHmݻL��<��_}<�d~=��)�{~0>R��	�R��J������ 潼�K�Gwo�(��{~0K{[
ޅRuץz�j�QvX]�*��8�｟�l~0^�Xɱ���vZc�j�t�L�7��r�b�M��L:�_PO���� ��_e��0�/AX���ڴݖ��sQ�`�� ��ޭ�
�\K����˫��,%t�':���Tj�߿���o�\����g�,=P�Ù��;=�su� ���FŀrV�����$�m����\0j6, ���ݗ��t$[�l�f����� 96<��7gֱ�ST�;�i�/kb�M� �����S�厊i��ӻj�Xɱ��p�7��sQ�`U�{��w�w����({�'m�=r�[t#��q��G�u����3��[�5���l8�ԝp�����;�n0�t<��M�֧��N�6J��vϚ6	M��6����ͯ�X7T��7F,�k�͡�k	�ݳf7V�J����)t��uv�<N�nH�(�3s��8sK��A�n3����{`�.��������B�K�K.ٚؠ���NC��s$��j�8+\��Z������-��[�8R1;��t�'n�6�M���������`&ǀr�[)�i�+H�L��{�5 rlx7\0�[bNպT�j�l�9�ذ�c�9��ou� ���X���m�$Ą� rlx7\0�`�lX%mEv��[$�m����\0j6, �����n�(~��q�`Q��lj�ثnܮ���ɺ����X8�s�.�ěJ��!��'����0�G]`Ϯ���07�k%MҴ4�ݦ`�lX}U�}��S&I8{sf���Ҁ��ҹ's29��ӫ��wlM`}<�n�aﾻ���� �T��`�'n�6�M����\0j6, ���V�e�1�i�;N��`Q�`Ϯ���`����PE|
�6mC����f㱫vK�W`�r��n���f�@T:I1X��n�n�l��S� 96<vL�{��M�X���lbL�I� ���	�2��`��,����YN���t�6�;&V��og'��:���| �yxw���G�wv,���+�6���n��`��, ���	�2�nϭc��ISN��f/kb�=�W��O>��J���Ҁ�l�()�ԓ3(�|ηZ�Ѽ�*�.-d�s���"���Ɤv:جm�lMp��x�X�\0	�ذuK��;v�n���'d��7��MFŀ��5ʷV�Ҵ�lwi���j6, ���	ݙXj�%݉;V�1���u rlx�̬
���_+��0	P�+��M�I�	� ���	ݙX�\0	�lX�6�Qs�,���&��W��?>m�Q��w<L�i�kMN��5�ܮ���� �qg��f��m������`��`&ǀwv,����ګv�u�ou� �D� 96<n̬���X�*LISN��f:� rlxݙX�\0�|\��M�ڶ�lM`&ǀN���7��N�b�9�.��I۷Nۡ����T^N���@�٠1$2[���ݾ[[sM��aR�V{tj���{ ��`w�vGK"�G,�k!Q�`��2�Z�ˀ��v랅c;0��:q�lr=�󸺍�J.;V��^&�nu��6wW6OK,�Tl��6I�Ӯ!t�*J�DL�����-������ܬˢ�ј&x�t۶��.rqBn_�v����YLC���u�Q1��!\tl l�.�+2fnf�rz�(,�sx��-EBѕ�Gt3ۋ���Ǆ-���m�ۺ��g[..���6�]1w�m���x�6�͊ ���̙/8voR�1f�!	;V�Si�-� �FŞ���y���{���ܬbN�61&$&��c�'ve`�p�'Q�`�]��V�I:@�o��_�{��M��:�� 96<�"��`�����n��`�ذ�c�'v|�m��?w��qd��k��O9�e�."�B�.�oW-&t$t���[4φ�^�W�ݻL�%��, ���	ݙX�\0�>.U��n��i��M`&Ǚ+�XAO@0Lt'˿w� M���ŀs�]F1ؓ�n��D����J���ҎfI;��ފ ��<��r��LiZCNݤ� �� 狮���x�N��� �n�J����L��-� ��ذU��π{g���`��R݈��v��R�d�:ɘ�<�x!d��-7�:�]s�t��LIڦ�$�T��M� �ٕ�ou� ��ذM��S�b�� M��>u��P����Lg��`Ϯ�l�mؕ�Ӷ�7X�\0	}��E0�Ku�L33)�#jh^m*۳�X�*MZTۻv��K�lXɱ��2��`�|\��N�m67I� ���	ݙX�\0	}������M�n��Qخ�M�F��ϕ�ۮ*��Q����ŷ�����ub�l��CM��2��`�[ rlx7m�N�1�i;M;I���_kb�M� �ٕ�v��!+M+t�m�[f/��`&ǀN���7��n�w+m��)��t��M�	<�����~��I��L1X�FH�)P���%��$�{���C�R�lTӴ�x;��\0_kb�M� ��i*P.�.��/�6�4F�q�I�Q*������:	s$6����v՘,��1��{�/��`&����v?d�ֱ�T�$��v�3 ��͊���>呂����2�t�grj����-;��I�:M`��X;��z!yU?m��;-o� ���;,�*�ݺm4&������o��r�[�y*�~�`ݛ�SV]T����3RP�:P̮1oG����=y:PND0���<�`@$H1 р�<��T��(EIh|/"p �`�ߗ�| �V3>� 2|k�E�F�9
"��B@$x���? @�B�i��x�!d"3�`EH�a�"�u�.����1�j[mA��! '��"B&�^�|␅F1�@Y ���R.�
X�`BA�0��&V@�"@b_6�L�	�ZōKU�e!c#�Cû��`@���! ���A5`�b�"@"�8�!�@�߈�G�%�}��um���8M�C]Jv5��p�b�pZ����rk�fu�k���#��;�M���CYB��Zi���csCŹ]g��@���U� �-\n�IyJ}b�U�̭�N�Y�ģ�'�St;v��Z��8�r��Wk��mY��$�բh����vĖ	E��jjv��<j���K=p��۳�pU�[c�Ej|�/G�	V{Qj��˯���n�� rݞ,�ٻM8洝P[uv��1r�ڍ]�;B��7;�Sm#�$�;��������8�2d�D��9��c�0p��8�id�`i$G�����]9tC�	%���s���ؼsp�;l�S���[Q$��c�ָ��� �s�)�ԙ��:�f��-�=Q;l����2(Vi^;	]����
�k ����'���2][;�:���v�cEq�s+$Mu/�ۂgvx�ZUr�
��U�V�l�u1���)p�֕�P�f�QWiKn�=rv�^����zN���3�Ӟ7Ʒlu��O73���t��$�9�ɣ�u��	��]�V�e'��;���T�ٶ
��[u*��&^�S�v�U� ��qk��X��V�cvݸڌ�%(!�R�
�$���݆{ޭ�Wc�U�kk�q�'-,qU�V��3���P�v5�B{u�As;��4h�ں8ٵ@ �[���Ug`una�n�k4��;]��#���L�r�z���35��@��{T�vGO8̶�5����\�5�c�LD�k��qJ��^'����T����m@�AtG KDi�n�p۲w�t;Uקc�L�:��.T���V��/k�hj�[;&  TM�6�
��ʸ�,�tx�lq���;��rUa�tWs0� A��v�v34pS�n]`����8��S@���Q3V��Op�bȚ�f���\�I�N�m.�ۂ�,�hT[3���*�I;���=�u�HR�fHl��	�m�M��A|T�~_�T�A4S�D:!���!@5C�U�{'�=��sL�f�/TeIv��h�A��]*�l�zmҖ��0u;l]�7vwS�n�ۭ��p 쯇�i�F��=�f����q�vK�h�n��8�jy��V6�i����\�������su;2�͙d'T^fPY:�vu�:W4�:T�:v��g�}���ͣR�& w�� n�MK��k�����m�]�9]���=���� <��ԥw���w���)�̑H8Ju�ԷK8^g��*����h�APq�7���w���q%n�6���4����`}�`�`��H�b-�Se4�n�X���~32gs3g�;g��kv(nWk[4�[k �u� ��=��ok�X���ݓm;�m�$���\0\������F0T۫E&�v��r�H��Ȱ�p�;5� ��*WD
wbL�c-����9�IV�Йx���7O4*� �^��f��źh���M&��M�}�`�p�;5� 9+c�9�.�7nĝ�t�7&n�$�{��sD0L1b�Yg��z`�7xg��lD%'�Tښ�ꭶ&��}� 䭏 �� ���k��ҷJ�MYm��[/ ���;��06"'��L��Ք[b��i;�I� ����`�p�J���t��?���hHc��t���oQ� ���I�K�ۇnX	��I��ykS��ة�hv�ou� �� rV�ꪮX���6{��mݵv�զ��Py:P�f� {sf���ҹ�2Ogg�Z1���h��n�0����٣�2f^d�L���@z�t�.��M���m]�M�z���吏6?�\06��*&:��cZNպm:���;գ��� 9���&Ǜm�����}殪�k*�\2��j���l;�j8�Sbt�g%ԏ�n'U�ᴥt۲�0�`6�< ���n�`�[�[J�*m5e�`6�< ���n�`�p�&Ԉ�[b��i;�I� ���n�`�p�mlx&�Wie�M�C�m�}W�3���� {l�c3�I����W�v��_[�{=���n��-Zci��\0�[ rlx7\0o޾�x��==-�u-�(N�[v��{�uk.祭�J�ʶnV�8um�s�5�Y�����c�9��ou� �T��M�էm��I� ����U��]����&�� 9����Q�ui;V���o �������`&ǀsE��V�Ҷ���0�`��� 96<��zk��ҷI;��0^�ŀ{ﯾ�|�?$�߷��N ���*)z}<�w�z�
V��e͉3;��MY��ֱ�ǣ1)Ҙ�P6q��c�[i�x�l#Ĕ��������I�N5ҽ]�癟��]��
:8�O G[B�&�ۙ���^�cC�5�nV�Rr��p8�uX�$�C�Tm��J�:��˝I.N��u:!,�RC�t촅�٬��T+I�_�ӣn��4�3��Λ[YǌR�q���۳/#/-��޻����O��C�LF��mv�K� �"J۲,�Ť�'o�o�>|�C�
�äة��L�I� z~��nN�^N����}[�@_j�w��<�M��۶������W�d��`�S� 96<�&6�wlV��v�0�`�[�vw�� ���K�X���@���3��_W�y`}<��`{깳<`�}w�vZ�N�E�M`&ǀz�����&�� ��ذA�$S��ݻB��Lnݶ�&�qk������ꖷnv;:){v�뿾���s�p��n�N�����`�p�9r�/W����xb��n�vҶ��� ��҅��&K�I�Kz(;�hfL3��}�]��k�Bi[����i�nT��M� �����$�)[c��i2�&��c�9��ou�T$�����9�mL�b&�WwT�nnf���Ҁ�L�nmq�-�wE {sg����'�;������Y9%9�Kv���L�j�f���nt��s��f�io$�I��\0\� rlx�`�]��m�v�u�r�H��$�Cu���� o��Wbe�S4;V����5�lx�a�}�U^�U_%̬�*E�N�t�1ؓ�m��+M���I�+ �ʑ`z�꯮���v(�V�m+n�n�l�$ٕ�r�H�M� �����P�1�}m�B�XQ�����5� ��.-��3�j�k���[�d��bF�o��}��M� ��M�X�,�[c��i2�&�M� ��M�X.T� �j+�YWlT�J��m���I�+ �ʑ`��f�7��e�DL�D�������~]�@���I��]T-�|�rI�{�L�ݺ@�V&�`�R, �c�7vـ6�,a(�Q�� *�SR�n�[#���k[�p��yԮy��wE�n#���*k�͵�n�+C�hi�n�\ ���n�$�X.T� ���c�;v��ں����<�M��X'V�`m�y/U���WW7U7jn�Tݘ��b�>���<�/U��x�ߌ�;t�V�mZCN�I�˕"�	$x�`I��mm,�[c��iP����x{�f �x���� Ģ"�O>'!{Җ�.ɛ�ܙ�n�,��v���[��NwZִ�F�d
��5wn{v��2�^7nf��Ľ����l�v;$θ<�q�Z랓ն�R=��X�9�Wh8�[曝6�MJk}c��q����
��N�wk�ϰ;c��= �J��+�>�ےoEr��3��D�ڮL���D��t�f�k�m�m:N�8û1�g�>��:�����>a��k�N�4�64��=�u��n������Ky��aۤc]S��v��,u��e]�Sm*v��'���I&V˕"�	$xŲ�Lv˶�m$�I2�\� I#�7u� ���j� M��X.&� n�ٖ��n���;����h�Ӳ�&�I���e`*����,�z��c�'n�t�o ��I2�\� I#�=�W���~�����_K+P�MqEh��Qۧp�����z�i$�%���6�҉\���Ʃ�g ����*E�H�r�H�`�kԕ��V�Ӷ�u�r�H���Ԁ@�EX�$�H��.`�}x{�f �x�R�a�9b��M�mU�m`��<w\0��R���ŀrun� �L�+ʺWuT�nn� �;l�o���X
gwu��z�Lv˶�n�f$�X33\rޏ wwM��� {_!h���cp�=^X�Q���(謎�]�0�Q��+g�6�n�o�w���w�h�vi2W~`��{X �w�w��y%�\����X�����i�n�X$� �;l�o |�]�^JQ����P�I۶��6��=<��ea��]9u5F
Q������>�D|	!L�2N�'��13\�8F�#���S� �hR� �ecIR���8&�:�D3��R�p��@I�F���T1"͔�X$T���#���p�h+�ԈR�R�1LW�\G�WC���'�T|N����>DT�*�z
�!�/� �C�/@D
"��� <�@���7�߷ =���9����������Ԓ~��* �[�@��@e��@]�*RV�mZCN�I� rVǀ{�����>�� m�X�%�6Q�$�*��/E��F���f:�z�S�q7�i�ppR��7Tz"�d�7e��MԔ����xy�f �x�B_H����ZT��f���T��o ��$�X�R< �G���%�ަ���ě���n����n��Dɻ�xn��>ṃN�[j�m� N�< �G�n�j���L��[�q���iݴ6�I���e`�#ͷ����v�,�(�WG&��ً��,����-���xF��۬�Z����tӫi�w\0	$��	�G�H����m+��Cl�$�+ 'I I#�7u� �MjRV�mZCN�I� N�< �G�n�&�XA�1Tݖ��7SRU��)���I�M�X.T� �j
�e�5M��۶����ޞ�p߫��I'{�w�N�J����r��;��\�%��+�f�^�Ǝ�[wL�;t8�u���8�N�j��z#���O#���1;�[lV�7�m9d��6zy݋'bi�l�,4�p�����t掺�.�N�Ѿc�Jٞ1�H��K-&T1@����m�f�.��zW\��*�zp�F��I�M�ܶ���%� 㬱l�5�ҘΎrp�Ʒ��(=�y��D.s�궫'�{����|�ݰ�c��/\���Q�Ƶ����קm�%2F��:��:ݷM&;e�e�7i3�{���*E�lx�`��V v�hi	�X.T� $���p�$ٕ�w�~.0���鵀lx�`l��9r�X�eD!ؓ�m:m7�n�&̬�*E�lxw\blM4��T6�M�X.T� $���p�
�v�Zmb��*��47%�Sr��趜�h�ƫ����$pYT��f�tč�6߇���`���M�X~�%�J�4݅�.��$�~��?ʉ��WI��	�ԥ&d�lL�@ggR�<��,{ZK1�lT�J��m��p�$ٕ�r��X&ǀlRSi��v�bLi3U͙L^ԋ 7��*�w!�w�<�b�v����u�r�H�M� ��M�X�bE�Y���Jh�u�e��LL>�	��`zSt�B��\n4j��{���|��zwr=O���ޚ�'J/'No8[���d]V:���hi�i����\0^ԋ 96<�UٱO2�V�j�1���]�u7xT%��,!LE"�X�A���0R����f{�x�~0�m�M$�J�-��L�mH��c�7u��}sfx�7�^��J�6U�V�5���g�6?�R<�] .�]1S��"gGX;5Y�WN�Bq�PUv]�l�$�q�xnm�HV6]�Leӵm�w\0�`�7~�\�;�������ڻ�3v9$�I@e��\�;�����/������%�X�N�@�I;l�9z�� ����)��z`���9�pL�B4X��j�X������l��$�{��rM>R@<ʻ�aذle\�:�ݥn�t�o ��ənmq�-�wE {sf�/2���7Z����ٜ�c��g+��c\���Km8<.��N6u�ww|������vCH'�	���9{R, ����`��R�I�hH��-3 ��H��}v���3vx�2�t�I�����(y�TȞb�Rk ;��wu� ���ڑ`�*
��ݱ1�Jն�=U{&x�&�� ��H�=w�O<_�����]�X�L�7��~���. w��{����&�؁�Q�`Qn���ߑΝ�j�u��msm'F������>p�R]�t�Όܗu�nC�0�Ѻ�d ��J�ݎغ��˗;�޸u�LH���mnzyVE�I�:W�7��#���S���s���N@�-��p������%r,C���ui�;\���мU�I��J�.2�pq>����(���y�ء\�g�y��(Vu��5K[c�۸�{��ǟ�;���-F�:��ҷ<���������sz]�K[�R�if��_��K��ىvi����{�� rlxw\0�`�)Є��UV�i]� |��?bQ�UCݿ�����f�Dɽv)�E�����-�m��l������"�M� �R���M��ف꯮l�Ʒo >}w�舏BJ���>P��B��y��r��nL�we�6pA�6667ޟ�o �`�`�`�}����� � � � �������lll{�y�pA�666?���w����s�q��V�rWaE{�5Ū6��T9	�v,+��������o-����t�>�I��s&��� � � � ������A�666?w��8 ���~�Q|���������� � � � ������i��m��.��A�666?w��8 ���X��S�C��C� �6?���N>A��������� � � � �w��A��66?g�ߦ�黅���͛����A�A�A�A������ � � � �{��x �ň9������A�666?w�?� �`�`�`���K�&n�d�w-ۻ8 �����|������o �`�`�`������� � ؊� �������lll~�2�4�3f\˚L���� � � � �w��A�666("U�����}�����������lllo�w��A�666>��	�Ի�M����)�w6qE�\�h�b^3NWu�n��u2��U�|�wϏ���\ݹ����� � � � ��y�pA�666=���8 �����|������o �`�`�`�����f��2m��7vpA�666=���8 �[����|������o �`�`�`�������
� � � ���~ɹ��w&d��˛8 �����|������o �bS�b���b�`����' �`�`�`�߻�ӂ�A�A�A�A��v~���7e��7wx �[����>A���߻�ӂ�A�A�A�A������ � �(*@r9�o �`�`�`���O���n�ٶ�̗wx �~�?N>A���P������ � � � �~�����lllo���x ����w{��u��ku���W"���inݸ]j:�P�ƽ0�t��Fg4����~���7p�vY��s6pA�666=���8 �����|������o �`�`�`������� � � � ����3fdۻnI��3n����lllo�w��A�#��A�����x �*��y�0	���;�>.S�
�i�w�� �����Ҏd�g}͞(�y��ʹHui�I�ۦ�x������\P�<P�6h%2JY&Hd����:
���3{��Ͼ��M�m&�;ml�7��~��U��R����3��h^N��c��)Ӓ�)�y�7��&gs٭ع�v�	lS�ɻt�8uz�\N�44�VЩ4��l�wc�M���������p�����='y�T�75E�� |��<��(QTu���5���wc��}Wf����wlLwbH��y�����3332w/7��/�����Q���Wm�$Ɠ0?W�_U͙�/7��=��A�$�ɞ�k����ݫv��M� 9ݏ 96<�~��I>�������iG��� �B!'&�р?�Ĕ��'���l�T��VC�� B:b^։ÅHB �4����FU�T-JS��`qF5�$�VT��|�j���I�wqP���H�($b@��<�H0 E�%��V��3�����$N�ë
@*�p��
���fo#	D1��5#Ä=-2������	�`�"�`B#�%�w31�ݶ����hk��e-bM�a{c��NY�w<#F���j�^����x����#�7DW�˚X$#C�ix�:�U�:��khጇc4Ij�D�ʚtTNiYӝ�U�7-5J���6-^��6�Ģ�ӣ����W8۞�=�a�y�S��q���v��Ua;/PS��t�l:�3���h��[pby(1ة�%�{�r�UJ��i/C�� .;��1M�v�P��p]��V�դ��ӠNȻ$-�IZ�S�v���p�	]��)��4���k[�A&-l��H�Ɂ9�t�/ 9s�xе7S^��y��k�Cн�6{2n+���A�v�E�<ݺ7MC�ж��a3;�.�b�rB�y�A��$h�IJ��0F��$�f�qᮋIU ��cm�ٵ�d{M���"N�)VΝ]���U*��C`�L�G��l��U���yh 
�<HR�mR���LR��N@�
��9���7U�^�[���lpY��K�E���k����ӝ9�흶�F�:r�t�KJ�n+��L��[:�Fe�V���9�3�L�gn���vN�UR::�wen�-�]�V��,�ݔA��������[la�齳s�Ҷ�U�J��m�6jk4Yl�J�R��q���[!C�m�f�IѴ�v�ݻK.�T�;Y:�]x�.��6��YW�CM@ �[���j���Ѭ��׋��h\�rM'%����tT�N�<L��e�rjl9�}]cm ���v�.u����L��٫�n���c�XV�:�}��4� �3՗m�C���*��tU
��g�����u�=�b�A�8�����BՠZݥ�\J�Ud�$�PGchv��c�]���l;��-tCZs����)q�Vy6��ZazN��!��8+����j�6ʠ���(v1�V���t�[)*=6��Wm��:%�d���γ�z0��]��4g��9LP��PA�`)W���i�p�7a.�u�窙�x�F�)������~�Q:/�x(�M9�'�W�Xl.rR�b��[�s۞o"��Z��sn4���s��C��<��j��˝Y�]t�ݷ���V�5>,�j� l��#`6� ����͋�/B7��f�50��i���r���]&�b7Qkb�R��&�����e�<��mJ�j�c���-����ی$8�A�m��Їl��OkZŘ]��%�X�=!�o_���nNO�e9Y�<��Y�ku�j��fW)��t[�M˹��˗K&i�UGy�e᠆�Z�lWm��<�w\0�s&L�y��ޚ�dO�	O/0<�m��s��ou� 9ݏ 96<�_����䍞k��i؝�lf����wc�M� �u� ���j���xd��3;�oM _oM��f�P���� ��͜S7e��K���� rlx;��\0�����w�~��k�����>��&��g�}%�u�k�'CЌ9��Y��ں7����������E��	���`�p�wc�M� ;%D���]�X�L�7�ᑙ����%�$������� gwM�Ɇ+ꫳ��17jݷv��E�l�����]��3λ� }w��S�Zt!۫Jӥv�����]��� ��� ����<�le_��ݴ�m�M������� ��< �dxm��~��g汞_j����L:��'{N��ܼ���V�O]{l�Ls��"7igZ4�`�2Py:P�6h׻?3/�\�O� ��5��-�hT�l�vG��N�y�4���N��;��i�I�d�2912�34y�4�N�;JL���' ���#�!T�g�'��f�����;
���wt�6X�.��5B�7�x���q������R�Tګ��n�f���������� BmB��HJ�vH��X�W	GEdwKGX�E<k���'j:{��٪z(H�v)��m�?�~�0� �u� �u� �V�\�B���:Wm� �dy�v?�~0�n��
L��b�T\�w7Sjn�����<Py:Q�$��y�4y�4�Z�c��b�Cl�;�p�vG�I���MA��r(��G�����~��_���m[B��h�� �dx����\0�\0�_y��d��I\�'� 	���G<+�my[ȴ�v��,5�9���+�#�c�Đ��� �u� �u� 9��T%廻b��CM��g���RD�� ����M� $��6���v����ou� 9���吏����BƮ��H�i�� �dxɱ��`{�3���|_�Їn�$�V��M� �u� �� s�<�q~W ��"�T>�;��tx[l�u'4�H�_T�ƍ���p;����:�Xh�G�'�8�k�g�^�4�u��-͍�\kjnn:�s�����Y�kn�m�f��ۍ�n��9�]uTC\u�^6��<[ p1�ڬ7vxe,1��l��v�e��<��<���س]6��Q3��	��=��0;��`w5�\'MAQ��\��M��r{9���M6������y0�[n�˺e�+hə[���}�{u�.�|]�[n�'K�zuQv�t�Lvպ��m�;�~0�`;#�UUr�吏ݍyv6��SE	I@e��_$���@��@]��_3*��jG~��j�ҡ�h�� ��� 96<'�]��L�`�֎�!R���"$93&L��͚3g�/'J �dxaP�c.ة�đm���
�fdۛ\x�hۛ4=�g����b����&C��D�BwDSn���H�����7��y�r�+�6����~�����Ϯ��Q
#����:��+�wbm$ݴ�f s�<⯨��D(Qv�� �]� �;l�(^��QD����Є��I4����ߞ���� �dx;���Lvպ�����؈�
{ך`������&ǀs���c��wV�����ou�$��|}�4�N� �̃�185h�gtڮӥ(�Dӡ�r]�C�_j�n. �j.N.zqZ�={�@�٠.�t�ɒ���ԯz̥m��,i��� rly�����]�>�� >�w�	D%JU��~�v�M�$�m�y�0�`��<S@��~P=�����I<����	+e&��e�X�v�0?}��W6g� �� ���ɓ�mq@^r�(��H�i�� �dxﾪ�履 ݏ���uJJZJƂݶ���z����a��y^wF�Sqf�T*\���i;���V�������ӓ$��^wM vl��%��S�m��w�៪�� ��� 96<�"��"fO��r�6�ݴ�n�nl��� �dxɱ��`�[q<0<�R�1̔�2w�� �ޞI=����*���"'�x
��Ͻ�M	,�V��ƛ���M� ؄���>�ޘ���D:WV[r[4Jb�Y�pv��آv�\&��ݗn����עn��'��-��X�Q����~gJ/'J �n�2f�}�4|w(j�V[e�M�L�7��� ru���ٞIB�򈊣���arUՕAw3uuV`}�^ |��BP��n��&�� �uO���]+v	'm6�?}P��5���� �;l��J&x�� {b+�T���ݺi���9��{流�"��� ;����]��BP�[q�ݿ�~J�s���V8z�Z�e��N�Z�vny:n[.9��v#qԁ�l6^om�N�nɹF��ym�"�t�^�2��6���m�`��tFX{N�֤��=��/X��Ό�.��9mz���$uu�:e�N�;%\�vӡx���:ܼ��F�{J������8;(H�ʙ�ɃMƃs9!��˶��\\���җ��d�.����K/'���u�5գ]��l�A�۰"�蛕����J�M�۩n4�zvh8z��oݷ����� ��w�>��(��C�ޘS���x�&Dď2P�6k�fffw��/vx�2�t��&I���)C̒�Kn�o ;��su� �� sv<��e˺j�,i��9��m��@�٠�L�;�oM v��
f,���ؚf�� ��xɱ��p�9 㤮�`��5�i$��y	�knܾ�N/E��brid��':Us��{��|����$ݴ�g ;'� rlx7\?r�l~0�^��SE�N�Zci��O;�w��OD����N��4x���@v��@�ٯ�$�ó`�!S�C�m6�xd~0�a���$�^�M _oMw�1�02��Py:P�6hۛ4&L�̒Q�߼`mo�U5tM�����n� �f��&d��z|��^N����s��2T���(�C��q�Fδr��'ء�Q������Y���?}�{�萳�Ԏn�o��ߞ��{����´�x˶*n�E��n�g���D*�^ߌ �� >}w����Tڲ�v�bi��\0���߾��D�6��9�%"֧���S� �b�$j<�0�͸���r B!��$# @��x	��J�Ĉ0I������K���Ԋ.i*b�ʤ���LU0�Na(���R2�c ����.��"�J�cQM�&tpF�:�F4��N���Cj���� 	����
�<��D|�1O���t���7�O;��`삼��$ݴ�f����UT�7�� ϻ�=y:Py:P�5��tJ��
�������x��(J:������ǀrc.���hh�D>��F"��Ѹ�r#��.�Q[�6^��q��u��E4*uhv��o �u� ��Ҁ=y��ɓy��ޚs^c�`"eޭS`4�{���xɱ��g���ꫳj)�I&�&&�m�ݞxɱ��`�p�;(د)<�*drbe�fh9&d������<Q'�����p"�$#E"z%S��@�SCUE�����w��:^l������m���{���x���	F�[U53:v��7at�k�e�:s���m�]i;sZk�����$�4���{����fRj���i�-��tO?� s� s�<�����`�m1 n�% {3f�&I���hݞ(��0�O���t��V������̝(�L�;�l�@��@y}P��ݴ4ݶ�?UW�U}�<`���fl�|�&w��3^c�`"e��S DI@]��@|ɓ=����h^og$��Ѐ�3��������7nu�ɨ��j�y^�ö���6��!�"6����˲���m��UMu*��<�=5��mع�����'m���ݔ�ج9�l�b0V����k���DMZ!�e��^�n�L����bLE��=��-�0ܳ���[��%��s�N�W�s��B��c�+�[��+�+ckn#yQ�%�ݝ�=D�����ﻮડ��I�Y&�7v˚K�nL室�<r7;*��Yí�n#v�Ց���.?����|��ʧJ����-�@'��� �u� �u� �ѱ^R��M�4��o 9�� �;l�9��0�7y�	z��������퉌�I��$��`�p���gw�x�O< ��Rj���i�-������>��y�4�͚ד���X+�iwm4��� �fI﷧�fl�@e��@e�@�#诔c����Y�f��Au�2�A]�n[�c�����74�N9cdn�WͶ����h^N�^N�3/8��@�~Pirmۻ�737y$�߷���0�QC&o�&J����/;��=��@fc�>�Bn��`�p�wc���2w/�����‵��`�yP��
&$y����y�4}�4�N�3$�vg����YJ�V骶��m�&�@|�כ\x͞(כ49�Av�Ӹ���nH�B����|���:��t���v�Ʃe�e�]q�z逳k�*��?~�Py:P�6d��_oM w-�S�wm;E�4�{���xɛ4�'J䙙ܵ��D9/2�2�0�f wg� rlxr���}�K��M�z���h�I�+N�m�U}Uw}�4��^N���'{��;6J�%N��lm��x;��\0כ4�͚�Ifk����Ӵ��鉑ЎՕ�����Ni�v��Kq=u���v��g<�ޅ�Su�6���UE�Vp{~0����c�9�p�;Z��RV�[����d�^l�3'p�ޚ�g�/7��ʢ[=���L�w.���ܷwy$/������G�$ﹳ� ^oM{�ұ;���˦�m���{��wy'�����A��_�? ��C��<���{�ޙ�m�m��O$LI@e��@|̒{�����;����ޤSi�����6��+q\�)G%dam�ch��:���8sw�FnT��[v�7v�I� ��<�6,��R�(�Pk��7[�M�Uw2Tբ��h>��w����� z�f���I#�̫�UhV�I+V�ݏ�ޭsu���,{����	��T۰nJ/'J �����ؠ�f{ͮ(�����J��Ri�ـ�ǀr�ŀz�t�2�t��2jd�1'�N�2�k*��v׌몛�
�ڸ����4-�kec�l��+����r���� 88ܜ����=ٷQ�w0V@�Y���tH��-�&�[.��n�]U�=���i�U�M!�3��#��ݥxف�[	ۮ����c���R�4�sM�`�A��F��<��mr-Ã(&#��k�4�d]�y�t�s���cx�>��:����{���x:�zٺzCOk��]qm0����� �=ku���h��]]�b}ye+m[���j��6�y`�`�p�wc�;6��&��2�V��=y:Py:P�6h>��s3;�r���;wwm��&��M�� s��L�;���P�<PW�C��/s7WUf�DyB���^������f���S��[���ح�v��9sb�;�p�7��� �ċ��p#�1sZ3�r	Ѯ�=��m���[��;<.�t��~����s���ͭ�p��`�p�vG�r�ŀov�:�&n�a����9$�߷��C�ɦB3�h~ފ�'J�F9��7I�[f s�<�6,?]��� ����],�m�t�4�ݶ�=�}J=
*�������;��0�7xfu2���U�wx9�f�����tg�� 96<o�HR��.���އ����uћkA�'t-�m�log�׫����T��T[�ӫ���ou� 9� rlx{�+�
�iڰNƚL�vG���吏��{�z���[���ح�v��M� �og&����(�@h���Iv"7�n�= ���;btR�hv�6����\0�`;#�M� ��J|�	��M���f��f�
����}���� 8v��tH��]��uf�ms@�E�r&����
���,F8�\\���s6+| �v< ���w\=U\����],�m�t�4�ݦ��c��gv?���͚�fd��gk�Q�bI�E���~0�a����;�� ;��v)HR�������0�9$�{�w�I�~��N��xE@�)	2o&\�2���([���KÂv5m3 9ݏ 9$x;�m����NF-\��^�"̡Y��y^wF�Sqf�DX�S�L!�v#[%&Zv;M�$� �u� ��UW�}��<�o�^B�V�nҶ�Zo �vـw��`�n����P�G�t��t&��6ҫi����vG��<����j!+h��t�e�`|�$��y�4}�4�'J��I'�3��+�K)[j�5M'wm� ��4�N�^N��ݚObj�L�$J+Uw׾�@����V�>'���"�T1��*>i*�,hc(�+��TB	e���f��j6��������0a��H&�"E$Ɉr��["!���jE�T�$�X> (�E�E�,�>O��8$�>7���4�`2����m5&'��F�b�n12���j�N�:ً�'$�=���m���&xW:b�.zX�h����n0�vS#c�7Yf�ŐmͮI�W��iLEh�DUR��I[$@El���G��m�al�$h�w[lٜav�p�$��#���� ��u�V��:^ C��מ�+M9�ld�9�7�s4�k��g��ؓf��v���MI��ǰ;h�ˑ����B"���0<�Nu��7Gm��ⶣ7*�%o<N�Ά���5庺��7%�룫���16C�7kP�� <nKr(V�V�]r�6ææ�ˈkn����^1��qV�$3�U^mZsw::6��!�:(r���Ў5�Lg�Z^9;�O;d�s�'8����sv`f���Q,�ۣGA	�ݲI��p@r��t0;6��s��l�݀(��b�y:Z�hX� ���`�n��U	�^r2�9ݭbN�!:6��H�]��Wcs��p%\u�xƶ���l�DX�@���1\^Ts�f����=�jr�+n���+*��j��9��\�Y�Z)Bl��
�T�b���*�����ɮ,;a B��;d�G*���ưll4HH�ҍ�\��R�s:%���`��FQ��n��˞^
}㊙�q�g���{aƦHx�4���4��b�U���j�ӝ4�T�<�D��n�8�>�na�-c����9���׵��a���w�) �vɚ�>sù�j���^8z͹���`��3��ӀBn1��ө�����ᇩ@Z��T�=��
]�3�$��ݖ�N9�9�(�4*�\m���U@`�������C�	�7`�h���/\�1L9�X+n��:]j�.�Tu����p�Pk{0Y��c�W5�\�y{ j�@�Ӈ�^���t�Fr�Is�f �:%�d�F�{f�u�#�J�{��<p�vWͨ��s��.�	/b=,�@�V)����@p* b�� B���P�QbUM�Q>@F�>��������s.i�vnL�$��Y{b��q�V�q����/g��^�S��p�ZN�n���	l68��j�Y�pT����=���z}�]�a�;N;Yd����L��%�·n�8
���[���˭�,�.y��^ŵ��"�O��N��{Ir���Nx�L�Xs��[T:V�\c�aq;���c$��q9�}��^����
Z��O��;�K�n�6��.��n]z��k�j���\������E�=�$���p�4����4�v4�m�$��� >�w䗒J.P�����B_���I�;M3 �� s�< ���w��rI$��k����������0��< ����\0�`�0Vڱ4�v������U�}:h͞(��(>d�$����@vl��uhv�+l���\0�`;#�M� 9��PJ��I��c�L\k��Ҭvux2�D�[�z�y;==q��u��{�_|cĳ��Mݡ��[L�G� 9�� >mߔ(�C�w��-�SUWD�n�����I'���Ρ��%R!kVi�X��?�k�4�N�fN��I�+���.�R�պi�������}�>r��\W�ww��r���̧�ww�ҧ��4�v4�m�w}Z⼻����s����Қw~d̔D_wO����S(wbl�M^]����9˻��2�]���H�˻��q^]������󤮒���u�<�$�k�������%��[���q{TJ����}_UQXݘ+m��i��ۻ�{�S˻��M����������w!�]���v>�)31��� �~ߟ����zww|��=�wr�iMrI4D;�m�uiݴ��]��˻�Q�^]���r��4�m�Y�%A<��!�Y�ܧ�ww|�9ww��S��Mݧm�cM^]���r���ݙO.���6>r��(!� oy��켶��?~?�����&�m����ݙO.���6>r��\W�ww�܇9ww��We��*�V��BT�I��۝a��gWe���ZK���b^��_�w�(��0�~ ����~~ ��|ww|��>d������i���x��u)�춮�|���V��.��{�r���<��������|����)e7E�`4�j�������]ݝ�����I_}<�����O��}��o̚��X�2���m�����m������m�>����uAk3k%�vY�;���zrBf��C������&��]��k��������.���˻����[Lv�7b^/Q��r��a9�Q�6|�[���U�Qn����~ ��~ ���>�����g�����}�>r��D���Л�I�0�D�N����d���%;���wo�[o����~E�wvޙ���\�ܗ]t�wm�����~�e���$����T�ۏ�˻��g�r���2�m[��n�n^�ߒh���y�g����҃���J���� ���~�5wM1ݖ��o ����=	BM���;�z`ͻ�-DBL��@ ��@��}'}'�_��s�ך^�&.��v��]*S�;:of�JAf�p\m���t,un���-�v�vy�5��^���ʖd����ZB����գ��Iɦt���c�s��d�ȫB��H�pwf�Q`W.H��t�4YگN��N�������������A�� �1��ɋ��Jn�m��ϑ{An�4b���nh�Z�����y���-�[��+nf�Zw%ګ��.�9b��`ތ�ĝj�iq�b:�[`4�j=� �u� 9$Ͼ���������+LUi�[L�;�p�I�� ��{!E厄6�m4;l�I��}�}w$~0��v2�R�V��HM��L�{݊3'J�6�3$�ﻧ �^K�'Bn�7m�-5�n���Y��^ ���{�@rL���9�`.y�Q����<��k�n�� =��Mm3�ѷ*FG�s��=q,���`������X�n���ג��n��Ӫ�񹻗M���.i�$������P�U���w'J�6��`���WM1�V�m�����{꫽����y`6DRlul-�M5�n�����9rE�r�"�9]؊!�y��.������ͥ@s35�w� �Ｐ�p��"�J]�X�.8��ehx�K�3/�㡷���q��\�����Qn�BV6��X�#�9}�`��w�2�	�ʈT�ӻj�l.�x/�,��UvI�v{+ �����:wi�m�i�w\0��~�D4�O��@��o�߳ ����;f�i5v�n�N��UϾ��x�D�,K���59ı,O3��8�D�,K��6D�Kı?~ߢz�n���������n����ND�,K����'�,K��{͑9ı,O}��q<�bX�'�:�?P��F�/E�n.r�[�۾O��n�qV\���n�Pm��[W\���|���6���ݸ�ı,K����q<�bX�'{�l�Ȗ%�b{����Kı;3����bX�%���!��K�]�M˹���%�bX��y�'! �5�$��ޖT&@�p���3 e^̖T2�@ TȖ'�a92ͻ�ݥܻ�"r%�bX�}��q<�bX�'fw��,K��=�s��Kı;��dND�,K�{�K��䛲��ɷw��K�ʯ�6'������Kı>��gȖ%�bw��Ȝ�bX*A@����`��o"}�y���%�bX���:ffm��f�-ݸ��bX�'��{�O"X�%����"r%�bX���;8�D�,K�;ۉȖ%�b#��gMW��|�v��]ڴ9u��[t�<��k�m�k���x����f�=��O�~y�4�ss��%�bX������,K��߹���%�bX����ND�,K����'�,K��'{�]�ܷ]�w6���,K��߻���%�bX����ND�,K����'�,K��{͑9�eL�b~ϯ�����f�3wv]���%�bX��~�q9ı,O3��8�D�,K��6D�Kı=��vq<�bX�'݅��n[��͔ܓ7n'"X�%��{��Ȗ%�bw��Ȝ�bX�'����'�,K� ̉�o���,Kľ�����.�wa7.��Ȗ%�bw��Ȝ�bX�'����'�,K�����r%�bX�g��q<�bX�*���d.}�I�X�]ts��������sɱn#�v�M�=�y'��-9Ү���%���q����G[�m<(�Q��yz㛈Z��f�]��ۂnCX�����m�x->�L*WaY�����ݖ�{df��`=�n5��jx�5����`S���Q��r�f8�
�:�Ar�{n:z㘁5٧9�:ֈ�ɰ$��g�ܢ-���ow~�y#��wS)����RxV��R�J�K,���8�Kt����;g�p����zx��&�����{��<���8�D�,K���"X�%��{�����Ȗ%����Ȝ�bX�'~���&�$ݗn�M����Kİo��jr%�bX�g��q<�bX�'�w�"r%�bX���;8�D��oq��w�w�^�`�ȳ{�oqı<�{��yı,O��6D�K�W��bw���8�D�,K���59ı,O3���Lٷ6f��ws��Kı>����,K��߹���%�bX7��59ı,O3��>{�7���{���;��,����['"X�%��s���Kİ��ho��Sؖ%�b}����'�,K����dND�,K�>�)��.�\۸��gF�x�hi���������ZW������v�d.�[��b��w���oq�����ND�,K����'�,K����dND�,K�~�gȖ%�b}��3�-�sf�n���Ȗ%�by������O�"�T�Z�D��F�B�j>TODL�?�,O�~�Ȝ�bX�'��É�Kİo��jr'�*9S"X������ۥ�.�&廹��%�bX����"r%�bX�{�|8�D���2&A���59ı,Os�gȖ%�bt�p�6��.�.��l�Ȗ%���ȝ��~�O"X�%�{��jr%�bX�g~�q<�bX�'��6D�Kı=����K��3n�M����Kİo��jr%�bX�g~�q<�bX�'��6D�Kı>��vq<�bX��~��.�v�㛠�gVk����c�\;!�@źX#��ۍy�j��������r��\ݙs75<�bX�'������Kı>�y�'"X�%���s���Kİo��jr%�bX�{���4��l͛�ff�Ȗ%�b}��dND�,K�~�gȖ%�`߻���Kı<����y�2%��N��.�n[�l�͗vD�Kı;�y�q<�bX����ND��f �j�@ >��,JC� qH��H	,Z)��N����$P�x��ƚH��o�C1�eeX�X�%aB#B�#4��n9��
-BR%aB%ee-��kJBR�ٍ�-��Xa�YIB� ��FYx/O5_qT�)�ۤe`�+/��B>�F�*��/���g�J.d���<��#H�'�rWX�VNЌIYP�/�zB3�R���U���%؁u�)ڗǚD�C���9�X�1@��bD�C�
	 �Uċ$�<A]DO �����D��=_AQ��!��\��|#���O3��q<�bX�'�w�"r%�bX�w�[�����6ٻ�.��yı,�{���bX�'�߻�O"X�%��{͑9İ?ȝ���xd�'8�8]2�I�GODnjr%�bX�g~�q<�bX�'��6D�Kı>��vq<�bX����ND�,K���|0����sM;џN���XM���t�h�d�k�ч>og��U�w!��K�\�n[��'�,K������,K��߹���%�bX7��4??�}��,K�����O"X�%��aNmݹ�n۹w6D�Kı>��vq<�bX����ND�,K����'�,K����dND�,K�{�[�L&i�wrm͜O"X�%�}�sS�,K��;�s��K�C"dN��6D�Kı;�y�q<�c����}�}2\�I�г{�oq���D�w�q<�bX�'{��"r%�bX�{�;8�D�,�P�;�{���bX�'�onu�&d���ܲ��Ȗ%�b}�y�'"X�%���R�����%�`��f�"X�%��{��Ȗ%�bS���ٻ�w6�\n�֜�A#������[�jL]��AQ�e[��
�X$���E����{��,O}���O"X�%�~�sS�,K��=�s��Kı>�y�'"X�%��{9s:n���e7weݜO"X�%�~�sS�����,Os�߳��Kı;��6D�Kı=��vq<���L�b}���m3f��K�3759ı,Os�߳��Kı>�y�'"X�B"}�y�q<�bX���٩Ȗ%�b_>�뻷K�]6M˹���%�g�@ȝ��͑9ı,O��?N'�,K��w��Ȗ%�by�����%�bX�;�)���2M�w73dND�,K�~�gȖ%�a��@�����D�,K������%�bX�w���,KĢ| �D�PT|���)�N���r�ں6ۍ1K�8�i#is���m�k�Q��;�St!�]���Rw]cp�=��j{s��]�����A�Yf���[*�l�ձF�V7`
Uٜ�����`��5�M�.Ƙ�\a8�1�M��a��p��v�ER�K�+��J�1r�G��s��y��b���Ew6��d���l&�;���=��Κ��v���3������eɛ���͙:�"�GbsI�t���=)��K"-���e4�ݓI��3n�M����Kİo~����bX�'�߻�O"X�%��{͐?ŞDȖ%�߻�É�Kı?o����`�LJ�������ow�߻�O"X�%��{͑9ı,O���O"X�%�~�sS�,K�����]�fM.雒fnq<�bX�'��6D�Kı>���q<�c�a�2��٩Ȗ%�b{���8�D�,K�;��;TX���7������'~��N'�,K����59ı,O3�w8�D�,K���"r%�bX�t��3����6ٛ�.i��%�bX7��59ı,?�#�����{ı,N��͑9ı,O���O"X����=��}��@�3�/=������K�V�7Z�9��Róv�U��7T�ĝ-&�e7����Kı<����yı,O��l�Ȗ%�b}����yı,�{���bX�%���0�ۥ�.�n[��O"X�%��{͑9
 j�D�0@����]�Ȗ'y��O"X�%�~��59ı,O3�w8�D�,K��'2�&���'"X�%���wÉ�Kİo��jr%��)��=����O"X�%��߹�'"X�%���-�M&4ͻ�6�O"X�~�Q
f�"X�%��~��'�,K����Ȝ�bX�'���'�,K���a�r�&kB�������ow������%�bX�w���,K��߻���%�bX7��59ı,N��ϟ�6xk=��NnlGiV9:�u���wCt�G�=��u��������~z�.�a��7<ObX�%��߹�'"X�%���wÉ�Kİo��h 3ș�q��oE2���N2q�q=$�;�<��ے�Ȝ�bX�'���'��� G"dK�����Kı=����O"X�%��{͑9�2�D�=�w�3�sM��ݗ4�yı,�߳S�,K��;�s��K@���#Ȝ��}�Ȝ�bX�'{��q<�bX�'����L�n��M�3759ı,O3�w8�D�,K���"r%�bX�{�;8�D�,K���"X�%�|���.���]7-��'�,K����Ȝ�bX�������{ı,�߳S�,K��;�s��Kı?�T�N~��a�e�V�a�nӬ�knܼ�A��N�؞��M�U��ͧ��qlƆ��ߛ�oq���w����yı,�{���bX�'�߻�O"X�%��{�S�,K�����&�	�f�ܛwN'�,K��w��� r&D�=����O"X�%����Ȗ%�b}����yı�{��］r�&kB������,O3�w8�D�,K��S�,K��߹���%�bX7��59ı,O=���K�4��7$����%�g�!���?�zjr%�bX����Ӊ�Kİo��jr%�`|��HDj�@��Q�R�¨
��A�"n��gȖ%�b}���ۖ�]Ʉ��s3MND�,K�~�gȖ%�a��>��5<�bX�'������Kİ~��59ı,O�����w��m9�l��Kۍa��gZ9�hF;�s��f�r\���G������m���fn컳��%�bX7��٩Ȗ%�by�����%�bX?}���bX�'���'�,K�����s.��6Sp���ND�,K����'�,K����dND�,K�~�gȖ%�`�{���Kı/��ofnM.�u�r���yı,O��6D�Kı>���q<�c�
#���bl�����Kı>������%�bX���8i�%�7mܻ�"r%�bX�{�|8�D�,K���"X�%��w��Ȗ%�b}�y�'"X�%���%��&L�M��6�O"X�%�}�sS�,K���+�?�g�%�b~��͑9ı,O���O"X�%���("0dZ�
`>��?nW:�9�l����q�q��8݀:�/-�B�X���&��]8Ń�.�Kd��]X{�wf�p�����z�Q�Hq�݃����:��+�t����j�<e`,֌Vf���>����n��v�Yz�Wnx��̩c�
�

�ƹ�	]ظ��Z��r�-�S[�ќs0w&�a���=�H�&F�����U�ݗmÍtl7Glt��M�t��)�h��rrI<�6�ɹ�r���$�x+��(;�֧z$��n�5��n��9�D�7������ow�����yı,O��6D�Kı>���q<�bX����ND�,K�w�:d��M.l��378�D�,K�͑9�#�2%�߻�É�Kİo߿f�"X�%��w��Ȗ%��{��u��I'=����7���%���wÉ�Kİo��jr%�bX�g~�q<�bX�'�w�"r%�bX�tߌΛ�74�fn칧Ȗ%�`�{���Kı<����yı,O��6D�K���L�߻�Ӊ�Kı;��Ùt�ٲ��fnjr%�bX�g~�q<�bX�'�w�"r%�bX�{�|8�D�,K���"X���~���=���V�u��,��ܗjz���e�R �sT�sn
��Y�qiu�r���yı,O��6D�Kı>���q<�bX�����Ȑ2q���;z)��N2q�������"�vK�n]͑9ı,O���O!�!\��,{�jr%�bX��{��yı,O��6D�Kı=����K�.�n�M��Ȗ%�`���S�,K��;�s��K�ș��͑9ı,N���O"X�%�ٝ{�.M�K�7.�"X��!"{���8�D�,K��͑9ı,O���O"X�%��{�ND�,K�w�:d��m�a�	sw��Kı>����,K��߻���%�bX>����Kı/�����%�b]���w~���o��/;�1ufey���8�g�����8S[�vwc�-�i������aY������Ȟı,K�xq<�bX���59ı,K�~��<B�H�}��H'������6S7v]��$A��6'bX�%�wx�D�,K�͑9ı,O����O"~\��,N����sn��6Sp�wS�,Kľ����yı,O��6D�K�A"3��qa"r'����O"X�%�}�sS�,Kľ{>�rivK��2��Ȗ%�b}�y�'"X�%���s���Kİo��jr%�`*�bo�߿���Kı?����9�Ze�.ٹw6D�Kı>��vq<�bX��3�߳SȖ%�b{���8�D�,K�͑9Ǎ�7�����q�
�[����&�d�^�+n3/b���.�ݺ㝤��k���v..��Mݳnl�yı,�{���bX�'�߻�O"X�%����Ȝ�bX�'����'�,K���öe�2m�fn͹����bX�'�߻�O!����,N��6D�Kı;�y�q<�bX����ND�,K���:d��m��vIws��Kı>����,K��߹���%�bX7��59ı,O3�w8�D�,K���칙�w&ws-ݑ9ĳ�02'~Ȗ%�`߿~�ND�,K����'�,K�5@��.	��؝��6D�Kı<���/�wv�)��.��yı,�{���bX�'�߻�O"X�%����Ȝ�bX�&^o�2���N2q���A�� �+b�}p��
�T��{6�,��@u�bd�u���n�G]%j�9yY��7���{���~���yı,O��6D�Kı>���p?���Ȗ%�~��59ı,K�ӿ���K�]tܷw8�D�,K�͑9ı,O����O"X�%�}�sS�,K��;�s��Kı;��fsd�%�3lܻ�"r%�bX�{�;8�D�,K���"X� !�2'������Kı;����,K�����inM̲n�sgȖ%�`�{���Kı<����yı,O��6D�Kı>��vq<�bX��w�w�%ʓ�V����{��2X�g~�q<�bX�'�w�"r%�bX�{�|8�D�,K���"X�%��(���ՀQ0� E`"� @"b��@Z����V�ަ!���8f2�H���ie��d-�jJ��P�J	u��=��� ��E7��(� 1�k# �"�"\���6q�"B���� �8��P���,	ġJ�'P=C�`15aX��H� � �,`����J��u��\�Q�Kv�����:]�=P�Y���N�7Movݮ[k��"�w�nS3��MkP�X ��n7�S�v���݌�u�vҭW�ЃoT�<i�n_Acm�2�7���U����:ѩ^�ʥ�N�E��9��c����'E�iޓ����+�a�f�k%Vq`G��q�[VW�T���v�m̭I��Em͕N������V�p[�mix�W���Vl��\H�h����b���p<х�
Ԃ�`n�n�T��-u���m9.��sӎ^C{	\�B���ώZ�'�[��,��H�@�^�b�t�6��>p;#����@�ѓNO�>�eq��b�pt�6���ǰ��u����Vy�{i��<vx��$���c�ض�<t\�%��6���=�U汰iɤ�WX�6]nݑ G.jR2[��-�h� �V�*⣇'5u{:"�p[m���"���+�mK���c�'c(�����x�G]�k���m�;��8�W]��mخȀ�[F�xjʭG*e���֍m�:��js�mg=giTq�
�%%�ۗ��rE���!5T�������s5�@x���!*�b��m��gK��>k��/���"Bg<�vjez{瘺�)�UiH��0��x���t��2�5��8T3������Udm�ն���ͨL-,�V�J��
ʒ�ZM���Th�!��2�gl��������W-"��UҞ�v����^ζ�Y���;h> !Ӈ.��o��ꜻ3�gk�%�Yzq�\1�G^x<�t��	��j�j�jtU lU��G`݊��-�˻9��R$�\�ڜ�1�t��^g��N��6�ݔ�H�iB�n�N�����Ӡy���t2˹yU�G[��%U��9xW��GCM���f!s/'d�gT���)�W]��v\�5q�
��l�'���0
�3z�wl��8E�ç�\qncV�六�k�|��.P�mi�Ks* �_΀�
��*�P*�x�( z�?	�����@<R�OY&���m��.3I�h��t���]�e6���ԡ��L퓭rִ\�<�2a�K��Λ��l�h��3��s����7��83j��e���u��P�<u��n��6�t$��g4��p\8去k�tFlT"�I�\Rn��Lk����f�����많���j����knWn��C��m�y�zx��p�5�׭����sǲ3��u�J�7;�}ߏώ97����(
�R��U�t��\#ûte[vuu��	���W������9�ۜ2is6�3f�.n~O�%�b}���"r%�bX�{�|8�D�,K���"X�%��w��Ȗ%�b>��`X'=�[{�oq������wÉ�Kİo��jr%�bX�g~�q<�bX�'�w�"r'���"��lK���\�����6]��.���%�bX7��٩Ȗ%�by�����%����;����,K�������%�bX�vv�l��6l�a�����bX�'�߻�O"X�%����Ȝ�bX�'���'�,K�E�>��59ı,O~����&�f5��ws��Kı>����,K��X�����{ı,��٩Ȗ%�by�����%�bX�}~���̖�e�k�/�kbq�3�[)e���5G�mE�� =\�$��ųI��|��{��'���'�,K�����Ȗ%�by�����%�bX�}�l�Ȗ%�by����6Krne�wlۺq<�bX����NC�@*#�W�TǑ6%�����8�D�,K���l�Ȗ%�b}����y���,O�����t�˹%��n��"X�%��~���yı,O��6D�Kı>���q<�bX����ND�,K�w�:d��m�dݒ]��yĳ��"�����"r%�bX����É�Kİo��jr%�bX�g~�q<�bX��>��`X'=�[{�oq���X�{�|8�D�,K���"X�%��w��Ȗ%�b}�y�'"X�%���~���\�1Ɩz�]!�RRq�P���f��H�3Y�N�d3��î����.���%�bX7��59ı,O3�w8�D�,K�͐?�O"dK�������%�bX��?[�se�sf�n���Ȗ%�by������ș��sdND�,K�w��Ȗ%�`�{���Kı<�}{/�4�0��n[��O"X�%����Ȝ�bX�'���'�,x�Vx�
?�R�1`C�8`$O ���jr%�bX��w8�D�,K����%�vM�w.�Ȝ�bY��U
�|q<�bX����jr%�bX�g~�q<�bX�'�w�"r%�bX�w��3͒ܛ�d��6�O"X�%�}�sS�,K��T�������Kı;����,K��߻���%�bX�϶fK{m$ܙu�,����N���p�n�}�Кi�.����k�ݵ�Y���y~[�.T��Zow���D�=����O"X�%����Ȝ�bX�'���'�,K�����Ȗ%�by���L�\Ͱ̛�K��O"X�%����Ȝ��(ș�������%�bX7�߳S�,K��;�s����oq����}�2�9�
���%�bX�{�;8�D�,K���"X�	��=����O"X�%����Ȝ�bX�'�ߋ����f�7Mݗ6q<�bY���2}��jr%�bX�����'�,K����dND�,��>=ؙ�y���%�bX�vvܜ�n���ᙛ���bX�'�߻�O"X�%��G���ȞD�,K�w��Ȗ%�`�{���Kı?�~s۾�ݷ6m�֋ZtȐ]ks�zņ��M���bw�Zk]��<7:r��Ȗ%�b}�y�'"X�%���s���Kİo��jr%�bX�g~�q<�bX�'z^��L�M7mܻ�"r%�bX�{�;8�C�F9"X7�߳S�,K��?w�q<�bX�e�� ʆ_C�������x���n�sgȖ%�`߿~�ND�,K����'�,��Dȝ��l�Ȗ%�bw����yı,N��;f]32�I76�����Kı<����yı,O��6D�Kı>��vq<�bX�%����Ȗ%�by���L�\ͳ3s7$����%�bX�}�l�Ȗ%�a�ǿw�Ӊ�Kı,�����Kı<����yı,MT�������,��wrK����0����M���]h�"�+�	�ܫܜ�m�]����9�~|q�E']=�;��s���zε�\[���3g��v�3��g)����kvQ��hx��䫲�AƐm:�&�(=�bx�t���.�<oa��\�+ҕ�Y�_Z2Gj�)`xn6�vlJ6�Z�f�f1�;�+�W��E���H�ri�5�f�M�c3p�����8səy������Ru6��>����i��7mu6&�&��!��<�Nz)B�ND�,K�����yı,K=�wS�,K��;�s��Kı>����,K���:f��n͚n乳��Kı,���ND�,K����'�,K����dND�,K�~�gȖ%�b}��rr�n���37u9ı,O3�w8�D�,K�͑9ı,O���O"X�%�g���r%�bX��;/�4�0��M̻���%�bX�}�l�Ȗ%�b}����yı,K=�wS�,K�	�=����O"X�%���e�M�M7mܻ�"r%�bX�{�|8�D�,K���"X�%��w��Ȗ%�b}�y�'"X�%���9�̲��eə��1ْ�6�xWF����g�7i�*\"Λ��&fnIi���sK�t�yı,�{���bX�'�߻�O"X�%����Ȝ�bX�'���'�,K�����d�YM�г{�oq������������cȜ�b~��6D�Kı=���8�D�,K���"X�%��۝2is6�2n�.�q<�bX�'�w�"r%�bX�{�|8�D�,K���"X�%��w��Ȗ%�ow���\�Nz)B��|��{��>���q<�bX����ND�,K����'�,K����dND�,K��r�電��6i���O"X�%�}�sS�,K��;�s��Kı>����,K��߻���%�bY��������I�1�Ϫ��.�В&�ӤkC:4�\I�v+"���Հֈ.����3759ı,O3�w8�D�,K�͑9ı,O�����L�bX7�߳S�,K������d����72��Ȗ%�b}�y�'"X�%���wÉ�Kİo��jr%�bX�g~�q<�bX�'z^��M�M7mܻ�"r%�bX�{�|8�D�,K���"X� �
0�}o� �Q�P���D����K���3��Kı=���"r%�bX�u��<0���d��ۺq<�bY� �߿f�"X�%��~���yı,O��6D�Kı>���q<�g���{���+��,���D�,O3�w8�D�,K�͑9ı,O���O"X�%�}�sC�N��?_�:6i=�t�k��r�-{`|j.&�.��<t$Jw&m��}_]�h���J��y��7�2�_dX.lX4[Йm
����f�ٕ�r�"�9sb�;�p�96��Rm���M�۬��˛���v?��`%��ۦ黺j�M`~�ﯫ�� �����ҀhfBa�̙���n���/,ulUi�V��;�p�7��`O��}u�l(�	�d�*���À�+��'4hӺ�ۧm�0��T��/���k���ӿ�������u�o������r�"�9sb�;�p�9>�K)RJ�V	�v��r�"�9sb�;�p�7��N���v��j�4��M`�͊�'J9�;�l�@[�tP�׍Hui;-[j�����ٕ�r�"�9sb�9����hT��0��T��b���lPy:P�ͩ $Q?�����4��4��#Y3�]�lH5�f3�g{ۇu�)�Pn8(�e �۔^��X��ۜ4����1� �Ѵm��uЌ�#U��d����?8mtn7z���E8���u����:��bPx�؍q�H�f����.R�Z����J�9Z��0c��LpqR&-��4�şWeܽf6΍ �g�5�&�6Hw-�ܹqiѧ}�ww�������2xC��ͲnK��f����I��f�:����b�[
���?9�}�:-��]��61�h�������9sb�;�p�7�2��쁔��t��5I&�\ث񓹙����J����W�w-f���4�Ӥ4���n�� ����9}�`��`�!k)�j�'cV�0?U>���o��@y�6(9�$�3k����YN�TҰ��ݷX/�,�6,��{�+ ��a���ڶ]�+���u���nZ�r<�D.�9���fuq���S�B�v���ͷ���[o�����w]02���u�V��ն����I=����S�H�NÈ�(�}wJ���lP}͊��w-lo"$��N�J� �=��r�"�9sb�;�p�96��!��c6�n�_dX.lX{��fV6Y)ۦ鴕7I&�\ذUV��l�V s�<jɷv�������M�M�Ź.���p��3D=�Y�I-s�N�B���N5��*��M+m`�`ݙX���\ذڐ���wN���i��6� z�f���lPy:W32w/��)�J�V�[�� ��� �͋�q�0"�e$���π�c@G7����a������ԏ�B�*�B,���b1#�ԣ��8F����'���!	!��FB$dx#
q��G1))[�4W`2v%$�J��V6K���;��q"||����B!sG>�O0�9Ģ�4i^/}�LN!���t���	�T�`�#�P��S��
�sGŋԝ$V�H)�#O�ԏ�*�@�>HS�Bhą,��A�S�)J *	���*��D�E� �0(q"b���A8*���4P`��}�����:���۫nݪv�M�~��ﾫ����7c�ou� 9�ΩjRZCbv��i�����W�6g� w}�r�ŀokl�c�.�6�-]4�[t����{kq�kv���������\[`�L��M��� �� s�<�6/�U���`�M#�m��t�-3 9�˛�����(��(QG��x1\ڻWuT�誻�1���Ҁ��Ҁ={�@y^jݎ�Zt�$���`����?�v(D ЂH���-K����aH��X�B6 X�VА?%J�;���=�������wm[L�/rt�>d�3�wO�܎�.�t����s�,prb�,u0V��/2�mƥ�S�G��7n�{i�Y5��n�7\�Jl�hL�vG�oT��w��vk�:��E���ڦ�E���R^z����ݏ���� s�<�_]���^�:����mݧx�~0�p�vG�oT��sE�	�ШM�� �� ����Ss����T��� ��K�R۴�:m��� ީ/ �u� �� K�D		D$$BIq0�ZK���>h����:v�`�K�@��N��n+th��j�8.j3ѹ�T�>����v��^�m��ˣ��ذ�/&.4�h{q��\��	uv��Z��[�C@��'b��38ќp�27\3�E�W덩z�v��6�] ^ʹ7R�m�M՛�Ʉ��� 4�]��P�1�,�E�n�v�.����؉�]�nmf�f���D:����g��Bd�$���t�.ԯ�|��|�=�^�p۴��Zn9�c�\t�r���ӷM�i*m	7�7W��x{�f�`;#�9Э�wn�j�:C����9��3�
�w� s���}-ŀnԅ��E��t��V�0�p�������Jg����w���>i���i%M+N�i����\�`�`zQ-�� ���:���SqwWD�]��"�;�p�7u� 9� s���}�c�\��a��uu��ą�\"��i�[�������T7Jr���:�ZIs|{��`;#�9rE�r��QJnɺ)vT�ـw��cI�	�" �~U^�����Ns�o$��{� �u� �Ҩ���Sm��� �dx.H��\0�p�&�*V2�5M���$�˒,��w\0���Э�X�v�Ӥ4���s��`�Co4��ݼ�m���ߧ��;�� r4�[��:�'9���Rm�GRx�,�t�LW%�)��i3�I=���˒,��$!k)�J��t��l� ��ؠ/2t�33iW̓'s�5������C�L����N�y3/	�a4��L@��;�=��$����j��!դ67v�Zk ����+ 9�<�$X5^�[e� We�v`�^,ޅ	Ww޾���Xw\0��v�Z�ҷuj�LN�!�&sR�6h5˛$��c	A:��3�$];W=)U�m��v�`6G�r� �����ʕ��MSj��o ��"���Ҁ��Ҁ=��\ɓ'r�����c�V�!�m�d~0�p�l� ���R�����i���� >�w�}-���QP�$Đ�P�@�W�>z�'ys�NI;�Ӳ�+UU%�݁uf }�� �(K�%���E����@fd�@e䐡�wtDD#s5ӮR+�-ۣ�И��.���@�T1�ظ�u'C"��m�}���w\0�p�l� �jRvZCcwm����`���˒,��_]���z�V�m�6�G���xz)�N����L���դ�ۦ�Wm� sdx.H��m�	(����{2�b��v��h��&�\�`���3� �{+ 9�<�|8� w��K9��v]ۙ�R�:�oa�b�]��u��S�������g���$���9]�LkL��c��T��O�	��Nsx�.U���Ӻ�Oqol�g��rto^���M٭t7+]Y�����ZP��/f��xy@]��+<�۲��up��ƚ�v�R`�vȺ�����Rr��Nk�[;�0���pMX�dg���܀t�W&o/w󻻿�US��C��{�za�a!K3d�b�v^�]�l��룘��t�v3�X��u��5��ڷb�ګN�Ҷ�@��wfV {7g�y�߻���]��HHK�i��wfV sdx.H��W�$�_q��)Q��2̪ ���m�P�%3��L�����*�ZE;MZI��$Xw\0ݙX͑��.1;-!�����9��0$�ߗ�{��}-����?G}tt$F-9Q�f�y��E�r�3���\͙��B�Î	�y��qX�&��f��+ 9�<�$_���a�?�SëI۷LN�wm� sdyϪ�����F*T��"F�PB�J#!0�m� �m�{�+ �K�YJ�7M���$�˒,��~���{+ ;=�st��!X�U�Hi[k ����+ 9�<�$X�%�Y@�����0ݙX͑��"�;��se8Ь��\���+I=��Z�ۥ��]].��=�B��9Z�d���:���Yb��w���x.H��`�2�	տ*�]$�i�I7�r� �u� �ٕ�� �q��i�ն	5�]��@ffҢ[)�-a��&�I��	k2I%	�3.e�z�����<���ZcJ��:N�0ݙX���\�`~�ꪽٞ0�bn�t����u�� ������+ ��}�}:��Ά4=[[)ۈ�tv$�έ:Fn����@�-��غ�7���rV���Г|��y`�`�2�����>W�V;T��6���w�៪���%26� s���}-��9Ѳj���	�մ�wfV s�<=_U}w������`�P��MZ@Ӱm��D(���� ��ެ��"$�x�ꦜ��8rI���/K�3vݶ���x.H��\0ݙX���m�>�w��'n�9�)�����\�װFޢ�����l��G6+��=u���Vn)���'J36� z�g�I���2�~���//�n���Z�V�3 �ٕ�2N�y�4�wEw��s2I��#xv&�'M�7wm� w}�r� �u� �ٕ�IA%e�ة�hm	7�y�v(��(��T���t���%�V;T��6���w��g����M�V�� S�dP��2fd���3&Lȯ��*+���*+EQ_�EE�Q��Q����@T�AP!PP$E b�E `�E `�E�A���Q@�@B
���� ����������
"���QZ(���(����
"���(���Ȣ*+�∨��
"���(�����*+�*+���
�2��w[����@���9�>�a|    =                   4*PB      PJ�
 ""���)JJ$*���@ �  $HRIJ    F   � P  
b ) �(()6�AJv ��� $  
R!�-��
� :S']=�� ��ܞ\\w�PV�zruN�Ͻݼs�b�X �����}���;�)��
� � �(  ��P� ��}���M\w+�&��y{�-� ���w��<��d������ 7OK��^�彼 ��zi�ӫ� Εf{���5�e�Ó��]� ��J��ut�w>�^=�  �    `   (( h0  �=���x�v׼mu��<�����z�ū�->ڸ�.�&�w  �Je��N=�x5y=]���U�C��+����Ԫǻ��Z�{��}i��K�>Z���޻ǹټ�   A@ �&�z}i�}�uy�yy�}�J�sq��v� ]�S���8ջe�[��}��r�n >�r��;|�u{���  >ξ]ٽx��w� �ҙ=W.N�7���۽�r��� }>�g��zi�ק�^���{��� �   ((�}�}��m�=�/����j�&�ۀ>�G�)b�����׼x(�� `�fJD

$
  �D� )@ 	A@�@�"  ���V� ٠ R @ 4�Sm%J�@ ?�L�)T�Ǫ�$(  D�*�I*�� EO�	L�*J�2�"$&RRH@2x�B��o�O���b����_L�̧O�ڇ�ǋ��DTW���Q\UTAS������QQ_�DEEb��
���	!3�J,����Y��0����-
Y�r8�[
�6�Q�1�F1b��(q~T�M��k߸|6�\7�M.�$XH�l�X101�-RS#�i	�"D�CK�|���~>�-	��>[�##Ņ3/HR%��1K!��u������o�
�c�!�s�:��6�d�J��F��R4�$:B0E��-�S
�Ӏi���E"�0Ѿ6iL0t�\1��9�h��`|�k��Đ��0���@���H�	��&kE�D�C4�f]��|sl���z6B�K�*J`F��i�١�\v0�B�3}9�WZ��,)�
��M�!o~	�a�v�[&:�
K�P�1��P6P�"PZh6t�D�:� �����g?|�	L4�0�@�D�Z$��)b�#<��K�� �J�hA����DƁ�������%�$	�4��,X�}͜�/��mXҫ����I �Ƙt8tN� ��V��	F!A��h�4x$J	8iSp�O�7:	�|��RBl�b���c�o�҆�}�����0��.RT��4�k���DH�����jc��@�nHM�hѤ�IBSP���+@"B�jB5"^o}�X͋�s�Sݰ�9������מ�������C�P)"�$k��I�s0ᡆk9��s����33���11��(�[&)���!\M!$"6XC3[�y��&HM��!�ũ���.Jdk�(JF"E"�(gy���~4����\5�#BjL��5�"S4��+�P���T&���nہ�%��l5u�k|6�	ԁ���º6��|��j~/#L+�l��*l��.��ٯ#!
Ʊ����h�+;�!��ӛ�kl�J|������\�u�#u�Gj�1!HQ�)�r��;��U�B�- R���ChӐn���
��:	sS��G��*}s[�����0�3�	�UM��t��jfM�Å�xN\&�h�H1�4�0�7�.Ͼ�8����
�d�K�HCA
9�K����]h�ܳ}%1��e�Me�vY�l�9����Di�.h�.Z�k3R�.r�O��h! �a&%F���i"^h���}ɲ��<h,hU�*B�`1�:b��u���8�9�_����k�}�L�+
ߵ���|X�XH���obs�aP�$!�<��+�[ �  �B@���qaC;i!�$�,i�s������L����O���xi���'�Hl��kp��t��:EH5ֆSBT���3W|ap��D��.��	&k|��cJ�@���&�� P�9�9���4b�0`�:��|3\�796}�!\��k[�|uۤ��{(��� Ս-��rI���x��
d���	)	7�#u�$ F��1�V��J@��0��5�لf�h��L�ߞɰ℄*B��NJȌ�$"@�E�$\M������j,�N~ߋ+�BD�`��PbP�F�0�����`f@�!��Ct"ԍ �H>IH�J�|h�h��H^&���MQ��2�ŀ�j�!f䉁0���D �MM��"0�L���0jˆ�sG� @ԉ�
D�5���i�8r�.��t2}���� ��n	��h�b�$�a(� 1b�
�� &&���J��*Uq]?�:��t�IH�)pѤ�Z7����`M�H�P�Յ1!F$qb@t-1`��kSZ5�o\]��ɣ��3C;��C
B���B��	d	h҆�!
�,a���kV�m�m ��+�%�s鯾�|���+0�4�F�*E�>e1%�a�N�?M�a�3P�.vݦ�sk���M�Cz�>!�����I��2t�DRG�����Wn+��!�!H{��Ag�2��#���-��:tM����>M��i۴�E#�7������������*1#��0u�(W	sY���V�4�1 �a��3y���p$�Z�2�B0��bB��$�K��g�4n4"@��`F D���%S!��_����\���K�.]��t������B�J8� �|xm�D��$�D1Ѳđ*Wn�0�	yÁ�f��ec
搅� A
�:B504��h�.:�S�0�B����v�0�	e٦�@�\t���)��/�5�8R0���K;5M�a��)��wg�; Ł��D�`� !@��i߷����ph#���į�h$v��5pB�^ϳ��2�#�!B��%��!p���ih�"Fˣf�P�asZ��ޜ����,)�M�!q��.�p&h��D�A �٨S4hۿ��e+����͆�Lt�7��l���0��Dh��"h" i��\ɘt�$i
!-0X2%q�
f�B�pc��#*Bf����ۡx����@���&��ZĴ�}���ɸ� Ł��[�kBJ�Sp��%�8��["dX�P�[��6d�IÌ�o@n���!N?o��GbKg��5����`� сaN�k���0hi6�>ԅ�4���\�C�͍k���1S4l"U�I�h��V��H]t�
CR�˲�F�۬��Ï��}R���v!�_��r$�J�j1���o�-d��vF��0=V�I�!L.�����h޻2�n/�H�D��Ltlб�����q4l!\
���@���A.��rb��q<oaoam���;z#s[߼]�@޴mBA���bT�G��n!h6Ѕ����r﷝\f@��ߋ��!@�_��!r뮔�$���%�h�@���aL!T������H��!1�3��Ԅ�`X�� Ȅ!O���}��a�G1�)��l���,A��@��~X�q#N�-! �Ӂ"@������D�!$���]�kT�)�toQja�L�WLCH� S㥅5��W��SW��Tƺ�.k��4l V�	�I��I!��:PL$i�F4��4�>�y|H��@�>B*�6��I�8��:�Bu�s^@`}�Ɓ&'��H�␊�6|ˋ&0+��|ɚO�08i B P B�`�#V$L�D�Ł �A�Qp+�#\�N��y�!xЁ�}���0��2aD#H�Ō��$6�� B�����}u$aH�a� ���\��Bfb\	L%������ L�BD�1�Ip�-�
kt��ѥ��^{�s�	��$�.�N��ː�� �a
�&�	!H�4� �N����х��p&2�(�a�4!XЍ6�`@�)��V�Z��B�9&��Q,ܛ/ٿ��W5��c�fq!y�D�Gpjb�~;͕�.��3���96o����E�p�ĢD(A*�q*D�\^	��`���v�	p�1��l>C��4�:A�R����@�<�}��\���F1ۨ�
0bm�
�y˾sy��77�q���(A����}�x�iփWD,�9�:��Q�Pk��٭wE\8W���\�LsZ!�HCxnm��)��y�˓a�2���NE�S�3)��!��0��),�).Ss�K�>jJB�jf[ h�L�jQ�u����_�   � �   :G�R���oM���l��RR[ô��` l��d�� m�e��Ap �km�H��h�� m��[mћ��k�X�nllHS˥f� ke�[d���-�9U*��xbIz���l]R�nS>��q�ڮ���W������5m5�ʭt��e$�O�|6��b���m�#P�q�2��mtU�,(u���v��E���ဪ� ����3W�����W0P�>���B��K&��޿߹��np k��m m�   -l�鴂@[x-���#�I��t��-[�����ꪀr�."Z����ʻ �g��Z�U�V�W�	�I�HH -��`h�K����m�@  I �'l�I��Ͷ-���;i��,j���� �-��[#u���6� �ĀpR�m�Ht2�mx� Hpm�kZ�oP  [@ ��[@ [E�Km�� �M�rmrBK,p[@dٻ{��jӦM�  $ݵ���ޮ�ۤ� -�N � -�m�	 $�$� h6ٶ��� q��  �J $X`$փ��m ��h[d�۶�f�8 ����\���h5^[p� �Č6ͤ�I� �"� ��-� �f�	   n۰  � $��f�69d�G���� w$��kn� [E���     ��i6 8�$m����Cm� �9z���[BB� 8��K5[�A�Hh�m6ݎh�!'�m� 	6ݸ ��-6�l����m�-�R�  i0l�  ��m� $ �prޢYx �h�#��`�[y�Å� [Am 8[@[V� �����k���U�� In�	�[�m�h @ }v���q� �[Bu�-�ht�l�āV��+J�veX@j�xp8�i6��am	��K��v�m��j�@	�	��m��[�]��h ݶHr�m#m�cl�9"޲H�յW[*�Um.���c:@rxz�0K���pH�d �٧��>@�WYX������v�fN��Krײ�<�m��;l��L��-�[@ $ِ�i-亶�m� BKM����l� ;m���֍{g0p�`�m{6���   6�[ �5�Ʉ�Δ�� ���>�k~�m� p	 ��H  '8�7$�k��<\8n�5n�m*�uR��  � Hpu�۶Ƶ�q�86��g�  ���n�=�B��m� ��E -���  �h  [d!4�m6Z ��dβ�A�[��gCdi�f���>��q $ޓ��K[i ��6�`l�  m,�n�]�U]uVһt�!� �UJF@آ7Y�;sUKc�T��g窥ej	e   -��� �n�e5� H6��  s�m�-k;d��+�R�l*��1m]]w/5��P�;@R�p	�S��UU[q�k��lR�[@V1 ���φ�>VI��[j�ۭ��M�p��u�� m�M�m-�l�v��	�M�t�4ت��#a����Dy��u�,� @m�[v+0�5�ݤ�%@�+���T���g��>|��Z�X�0�C`��ٶ-��ɦ�Y��Yl���WX
�1�b����7n�v*	�+�/n�۶��I -�m��)��SL���圞�kӪ���9�l�l�n���lW��Tx
�99Z�Zॡ˄e�[@��%�k�t��hemR��>��&�*�6�Z�X$�v�Y�й`�M$���v�m�����U
g�2�]mP�P�	*�EѮ n���m�$�"�I�-UUm] �C�ں��ݕ@tU�R}�FH; 	,�m�M�n@  ����m��_i�L�Ad��Yc`����-�$$m@ l �m:]$vAn�pm�,sF��L .��@���
���Y]#UUR�rv�&bܫ�/Pp  6܎��p  �m�p-���Hiˢl��$Il��l�)��඀�cm�۷le�`:���C`|�<|����]'lm��;WT�dګ�\�p*�W��z��鑀,k[l���� .هm��`h�og ��!m��h6ێ�[d���V�m�rG�m��cvͶ�޸ $H�8 $  �H�ӭ��6��	l�F���1��p�+��lLm�*V�[].�H��3��v 6�$ �m�Mz�6�V@%����jq�X2ۭ� ��8ݴ����� m��Jl�$	6�m��-� �K�^��6� p��� _�ϝ|U����]��c�Jk��9"ޠm�U�}u��[@�����lkY%�֒8I�������f݀ڶ4R��ޒ�ٰ�� ڶJJ\-�Ӄk� (=,[Zk�gDN�L���[+pM���>\S�L��Y��k&kSkq� N��y,�uն8$in�0$��lv��ӧR��%8�Y�� H�];a8�V۶DX  m6cj������N�v��`-�6� m  
Y^��8-�m���K��$6�m���Ŵ�l�گ� ���u��l�# ,U�^�-��� m8 �mA��l���@6�m  m� � �	o  �$�-�����@EΌ�^@eP9�t���UU  	   �  m�]�i��-��5닦���  �[e�b� ��Ʃ:��$-����V��mm���uH��n���:@ KV��l��6���Nc��SY-�u��2��l���P@W]*�� ��mЪ�b��*�P �f�h	o�!l��K����9n�\č �Nm�Sm�z�6�ݮ[Cm� �d���i� �YWj�L�kh�\����!I��@m�p�m��¦��p=#�N�u�٥� p s8^�o������_����`6�,���� �D� �m,�     Ø 8&�Lp�������H��M�� ��H���  	 	���h�Gkr���H�p��@      }:� v�Lq 6[oP�gXnH r@ 4U�  ���2-�k-�ݶ6��   ��%��-��e��� Ͷ��� �m5���vj�Z����
�US���zj$෬�#pt�t�� 
��z��������y�j��ۀiV���6�
U���� 8 �n���`    ��>I6�i�h��0�`��;A[ AͶݫi���2@ H   �v��!QKr�T3��lN����.����yUZU��(6ְ݀��%ӺN�Y+[K��; ձǊ�(����V�`�H��j�Bl��[p� -�[n�t�%�lP��	 5�l$Z�|� �]m�ޮK&�7m�mV/l\�V�VS=!N�z�hĻI�.��,0 ��R� �-���UJ���ʽU�UR�]]K�R�]n���T [���&ŵm 9�[�]��`�`���UU�/n��I�r�V�S(n����HL�e-�K"ȍԋ����Y�lù�-k1m�8	;H�i8l��[@;i�[ջl���hH�K^��m�f�m�m�m���4U����v�������� 4=R���U-����`��k   !�^�	6�u ����[j��U*қ:�6�-�l�� m�A�Ŷ��A��m� ���V���i&Ŭh��6�@ �  m��6�;E0�n�6� m�@Y@��m��۶���| �����	i6�k��lj+$�H  �Wl�6�  o  �Z��      -�ݬ�7`�`l�-2   �����m�� 8  �ȥi�n-�mn� #Z��� Vm�Zl۶��  �I����;E�m� �    "�H� d
�� m�:q������$i;f��y��v�l�9k�   �]�� l��@���  � �m��ﵙ73���   &ն���J�X�*�U@GTkim�6���U�e���Z�U\�de��X3	eJ�I�H  [N �k���~��m��� ��9�Im  ��  [@�L[@ �Ŵ!%�Hj��Z$m���ݰI�Ul8 u�@ r@� m���� �9;v�q&۲�P@UJ��#�V�j����uͳ[M��5��&n��b��ܣR��<��Zֵ�����UT�
'�� �?���
��S�qS��ڇ�?(�@N(�UJ�"Az>Q.�}H#�� �+��P���	@^��&�'��Z�kc�C`��pA�M����`�C�N�tC�\6���m�O�Q��A_�MU�p�.��� ���N4��¡�צ��~T4��$|l_#���� �� �A���L@j
S���D>�"� :��| ���
b�q� X |
tB �}�bjH� Db��"1d� �+��PT�@����#�Si��'ʠ�1��*ï��p8�PG��P+�4*=�x^�-H�0��`��,"�<ET�A�� |�u���>>6�E"�bPh�"!"�j������ >GjńF�)�4^�'�E:�����(@T�A���SA�@H�)�� ګ@�
@~�"b�_�""���������;�wu���ߦ~� p]Z�)���qN]R*�<��iZ݃b�����2鵴8�f�^R�6ز��=-�Ơq$�Z�>������=����ԃ`��*���i���u�m�I/]�4�U���6�+g]�vCvQڡݭ�z�3�ڠ��&���S;[gUr�Z�#� x� �U+��:�a�V�G��i�L�A��y�nUg8$LvfI5�ڦ�3�n��,�դ\�QT��ٻ)0vr.@9]*`����4�U#��9�Wu��X���;R0��S����8�-Y�Ѻ{Y�\;���Z�w#lA�<�|�V뫃ғP�E�.�k�C�ˎ-��ˋv2X��U� ��T��T��yע�x��e-
�T�`�qs�
2Z�N[�<�gx�g6N�'Q����v�Q�i�ge����Ȭ�J��À�1l���ԍ�q7m[b�-dR�3�m{ch86F��aA1�49r�{[����n�9%�;î������N�7k
@HOJ��_elL/<��X�Sh�-�	��k�Y�ݰU�u�4۲�I�u
�3V���]���E��ܪfiׇ�m���;!���Us��]oA��Gv��v�L�FM��۔�c�2c�:��-U*�ɐ��3�9�){�mø7b�m�#�,�m�%�`)�+�T�\�5wgv[��ld�����ۣ�
��D)v�c��ܹ�U�Ùjڬ����/P�t]:��$�7n86+e�'n��O
YѲ� �ƚ,�i/�-+,XS/�B�m�Xړr�d.�Y�E3�A�Z�)���{k�����3����u�),��%1v��{�jIl��dT��Q+��նd%�GI4���:L�6�l�ն�z���Ā�s�U��,�qv�=�yc�V���\�р���mr"==-:AꔙX}�9����ZJ�Վ=*퍻g9��i���gi��,7�Z{B=�i�eYvf5n�,��I��f��AO�U��$p�$�^��E�9��	�=����j�\��5�jY��^
�M:��Q4휍��g64�� �%��6�=��%������7�v�n<��B;:ݺ���si�m�fvq�7��8�9�9hθ�<�v۫��l�ۉ���[va薻r�,ت]��T�=��T���D���Ʈ���vkL�f�� 4��&t���\U�qFL�nә�]�n�svuI�5�f]d��EQH��\���<w�nɱ�l�Oa�v�^�p���S�g�eܼ�L)�eʟF�A'����$D��ؚ�H$�>������L�bX���7q,KĽ����Y�D�kV�5�kZ�r%�bX��粦��?WQ5Ľ��kiȖ%�bw���Mı,K���[ND�,K�^�f��٣Z����ֵ�7ı,Ng��m9ı,O���Mı,K���[ND�,K���T�Kı9��ѫ�\��j�%�k6��bX�'��n&�X�%�y�}��"X�%���{*n%�bX�ϻ��r%�bX�����In��4au�D�Kı/>ﵴ�Kı;��eMı,K��}�ND�,K�{7q,K��w<�5d�&h^д��(s�����$���[s��Dے�V����ZK\0����W�w�{��7���w=�7ı,Ng��m9ı,O���Mı,K���[ND�,K��w�����C������oq��'3��6��Z� "S��dq*DDb � EA�A\��J���"r%��w6D�Kı/=�kiȖ%�bw;�ʛ�bX�'�-�>܋/�V~{���oq���}�fț�bX�%������bX�'s�쩸�%�bs>�iȖ%�bXw�z�ɫ0֌�e��q,Kļ���ӑ,K��w�ț�bX�'3��6��bX�'��l���%�b�����V�5�W�w�{��7����}����%�a����y��Kı>��dMı,K���[ND�,K=�;�����m!@���P�dzב�B:7%π|��:uv��t�\i���Yc��Y��D�Kı9�wٴ�Kı>��dMı,K���[ND�,K��k"n%�bX����jMh˔ѭ]d��fӑ,K���͑7ı,Kϻ�m9ı,N�}����%�br����-��B�
H[��]HJ)p����h���%�b^wߵ��Kı;���&�X�X�HbA
H$�; �Wf�dO���m9ı,O���q,K��{���\�h�n��ֶ��bX�'s��D�Kı9��iȖ%�b}�fț�bX�%�{�m9ı,ON���\�urh�h�nk"n%�bX��ﵴ�Kı>��dMı,K�����bX�'{�j��Kı?'�~���>˴�T�N�l\��7JCk���Z�������&�]%wV�V��m�k����%�bw���q,Kļ�}��"X�%���ڱ7ı,K����r%�bX��.d՚5�.Ys4D�Kı/;�kiȖ%�bw���Mı,K�����bX�'��l������~~o�}�m�PM5|�7�ı;�{V&�X�%�y��[ND���i����߳dMı,K���������oq�ߝ�~��έS7ı,K����r%�bX�{ٲ&�X�%�y��[ND�,�>W�j��)�R�A�(p�(���A< ��LϿj��Kı>����h�r�5���5�m9ı,O���q,Kļ�}��"X�%���ڱ7ı,Ng{��r%��ow���O��cvڠq�Wv��t���.�;�`Ŷ�i8�i�t�$���+�$�1�[�Z��Z"r%�bX��ﵴ�Kı;�{V&�X�%���}��)>��,K��fț�bX�'���	��r�-�n�Z�r%�bX�q,K��w�ͧ"X�%����"n%�bX��ﵴ�Kı=;�/�sE�ɭL�d�թ��%�bs;�fӑ,K���͑7ı,K����r%�bX��֦�X�%��jN�\+H�1�g������۹������q,KĿ{ߵ��Kı;�{V&�X�%�y��[ND�,Kþ3��շF�e�.f���bX�%�{�m9ı,?*G���X��bX�%�����"X�%����"n%�bX�|#��D�b�X0`��#	�"0Dh0	=��?7�6�1Ә����cR�h��5x��^1��m����6{u`-y�d�^��pí�v�G����^�p:��{Gc7�ێ���Ʈ۲UIԌ�M�)Dl��7ZٔLl�q�S��[vj݃�F�z,��Hu@:+8�..nK��$�f�n��`��Μlq�]v�1v�L�:.�ߏ��kzh��h��dv�T���ٕՄ��SV�@�\�-��J�t775�=�{&y�b����<%��)iI3�a�Ѩ&��=�w���{�O~��X��bX�%�{�m9ı,O���q,Kļ�}��"X�!�ߝ�~��έS��{��7�ļ�}��!�#��,N���"n%�bX��{����bX�'{�j��Kı9�n��Y��ѭ]e��kiȖ%�b}�fț�bX�%�{�m9ı,N�^Չ��%�b^w��ӑ,K�����d��kV�֤�ֈ��bX�%�{�m9ı,N�^Չ��%�b^w��ӑ,K���͑7ı,N���5r�ɣ2�7Y�m9ı,N�^Չ��%�b^w��ӑ,K���͑7ı,K����r%�bX��=�~%���͸�Bfe��4�ۧ\�b�{\j����yu��v�5�6W�غ�r]��ɓY3E��ND�,K��~�ӑ,K���͑7ı,K����r%�bX�q,K���'}5s0�d�5fff���Kı>��dM��=͍4��B�^D�K�{�[ND�,K�׵bn%�bX��ﵴ�Kı,;�<\ɫ4kY.d��"n%�bX��ﵴ�Kı;�{V&�X�%�y��[ND�,K�{6D�Kı/{<_j�։�kV�5�ֵ��K�2'��ڱ7ı,K���[ND�,K�{6D�Kı/;�kiȖ%�bt�{�5r�EѓZ�ֳV&�X�%�y��[ND�,K�${��p�Ȗ%�b_����r%�bX�q,K�秥��Hl�Ҝ6��/O�7F�q�۬����fBgN]:qL���C��A��D�,K�{6D�Kı/;�kiȖ%�bw���Mı,K�����bX�'�'�v�I��nMjK�h���%�b^w��Ӑ���ș����V&�X�%�~��kiȖ%�b}�fț�bX�'~�L�f�L�3-�u��ӑ,K��u�X��bX�%�{�m9���ALTM��Oky�&�X�%�y��[ND�,K�����7P������{��7�������r%�bX�{ٲ&�X�%�y��[ND�,K�׵bn%�bX�~�~}Я3��2�|�7���{���{6D�Kı/;�kiȖ%�bw���Mı,K�����bX�=�����q۳�,b �v��J7%᧝q]��^Rlw<:�O[.�<�y�=�z\.34D�Kı/���m9ı,N�^Չ��%�b^w��ӑ,K���͑7ı,K��ڗ5�j�j�f��ֶ��bX�'{�j��?�c�2$����.�L��v����Ԓ�����{É�&F8��8���h��h��Wmz�V�I�1d�iW9���sw~V���N7V
q$u��s[�x��n�)0֒d���w�h������[�s��h;�H_���~QƓB��{=:�\J��i���,�b��\�5���[*��ʻK?,�������07�t�=�٠^X5q7X�1	8�����Go�����@��@��io���Cmɠs��h��mz�{f�}�㨏"F��ۙ�w��K`��ޑ� �%)���"$J9�@��@>�l�9�w4$�{�nIG������K��[3Y�.h�z�L:�8�ѳi�7B�q�ݶ;3�R=]��+Js�/5grg��ݸ�RW���
���T9z-lN�O:Iq�*q�\�!�ov�e�S� ������xs�g�m.h{s��..7�ї�N��ܽɓe�Hz.���8n�%�!:Z�3p�+�ۉ����!������cY���6]�M�'	]�����JgW��}��ϻ������&��9^��:]�
;V�N9�qɸ��ֹ7W[-.�k��aFLS!#�8�}��s��h.�������:	1d�i9&��#��t�.����0%J���$ɓ�4�{^�޻V�߳�$r�M���4�A��1���=�Il��$t������Z�m̃$�$����4[w4�{^�޻V�^.Մ�D��I�$��͎�uͨ��V	�ً<���fN�p��R����1�N!���9m��>]�zz�^�߾A�o��r���G�#blY�7$��}��P~�E֧w��ܓ��נr۹��qR'(ےG�r�-���-��#��t��� �hɊd$q����k�9�w4�{^�λV�՜����L�F'#�;�ڰ5%
;M�|:ݛ��u`o���������w�NB������t�\��+���4\l�=hyՈx!��q�g�J̬����5I��;�D�����n��v��m�c&6)�zz�[�+|�����>]�z�`�Cnd(�
␚��Nc���V|��GB?ب��(���SCEi�6Dpa1j�03B\6���d�����)�(���p���H0�A!�D�My ���4�:��J,,60*�*�bq�@?AP��7�;�K���D&R��t�E��������a��ȣC0	�m�C̔�*T�J70WM-�.0#m`Fb�E1 R�� �F ���P"���|(qAR m0�	�A��jUAX�u7{�?��;_��y�}�㌐N!6�Xl�����{[�u�6|�{-�X2���D<�A���ɹ�V��~���n͟L�oy`f�ڰ=��'��9�;!�z��nn�%Q�c�o��T_��o����#��뚫F�g�j%j�������������˺[���+Ee)���Z˽��#����8���;�j�f$U���&$œ$Q����|���-��r&�t���5WJ��Ĭ��W�L.�lۑ0<���)�!�z+"�W���y Js{����|l���C&�ɪ�/-��r&��gGLw�o����k%�3�ۖ2s{xz�ړU'n�:�ӷ���86�/�0+ӴCNH��gVn0�˺[gGL.�lۑ0%xv�b��N!6��9{w4�{^��;W��V��|�2���D<��q�9��{���-����;����A�x����ErH��g����=<�}}��q[�w;��m,��BGqh.����s߾A�o���K�ǹ���4�n}¹�c�'����ɝ����)�2Tq�ҼN��թbi��)�;:R�8v� ���-��Sg��m\:ť��T�`�g���O�M��W�ܸ���Wlk����ϩ�(���<v�c��rb0��]a�g���$m���]9Gs���'������n�f�˜�����n��]m\k>��;L�4��[+�]+n/�~\��g[$u\	���w�{�z�|��Ƿ^�Cb���mF�]"I,ܞYC���9�d�aD-����v�8u�F+���=��+��֯�V��|���ց�����`�D�2brf�8���V��_Hv[ڰ�'5���x�Z��r��1�L��~H�~��8���9{w4�{^�zv	T71�ps'�������˺[��L	-�j1FH'�q����˽�@��@�w��w�;���,Px�j��&�k�(�8ٻ��u��_��Ϗ�$�;h*:����y$��I��+|��ڴ�{_�3�~�}}���B=	&�m�9Vv�����I(���{V��V˽�}��.\wأid�28�@췵`u�f�S=�����6�-�&$œQ	��^����נw�ՠ|�����j`�y"N"by������˺[gGLH[��ʖ�%eCW]�yͬv�n� �3h1�%�����+Y��[�7 \i��v܉���-�����t��:��d#Q�b��>]�z-��˽�@�]�@��v�F(��nf�{�ٹ'/{���!�t>P��뽛'1Հ|���\��9��J�)���-��r&�t��0h"�D�6���h�]���7vՁ��:�6!-kfoy�(kj�GW�,��f=��xcpN�a�լ鋌\ۑ�:a�q�q([N�11��O�m��GL.�l�0
��Yj�YW��2�$t���t�uȘ.����Z�,H������|��l�0<���6H��х��XY�v�R2���"`ywK`l�����8wv����~��B5� N&�t��'��ywK`w\�����>:E�����g��LJ6U����P���n�
����#�7D�N�6��6H���-��r&�t��댸�D<rB6�s4�{^�޻V���k�9m��h"�,��Erf[��L.�lIl��˺[���qFҁ�&��>]�z-���{f�޻V�g{��M4�&8��[d����0;�D�����������ߛ�O����v�1��+۴�x(8��6)�	 ;���c͠���NNٮM�\�������6B������R�vV�Q*�G��֍�m�n�h�'\d\n����m��8l(��w�9$;s�&�m��Z6����v���"��kG��y�)���i��+;;,>�;��H{1º�1�������/b7��v��q�g�An���wn�w�w̧�\����E�an�p@�g��6��u��g;u"�	;�%6h�{��1�*�Ͷ����0;�D���SA�GLwF�xȠ�J~Qɠuv׿߿bG�z}�nh���b��B5�!'���-��GL���K`l�B�4FFG���n�}�٠uvסW��
����y�� �M�`����[˺[d��R��[�l�;k�k=X��iۡ����$�!�rL1�6�O��;cq�]��/.Э�`r�-���-��GL��[W�-�K�5�Yu���f䜽�|b,B+���Ԃ'�MP�*P� �`���"���^�f�sf�w�h]��H2ۭ��4��(��-��GL���W�J)����'���itx,B'�I3@>�l�:��XNc�IDNn����=��Ur�r�]���^c�Il.�l�:`�٠w�\X�TA��a�a3�v��h0s�7fӷ����:E����?;�s���8��@�s@>�l�:�k�9l�;�&���&&�z-��TL�[�X^�XNc��S���R4�� ���@��M��X�@�(U٬u`g[�`%�'��-�(ܒI�uvנ|���[w4�v���w.(�25mǠ|���$t�=�1�ˤ��*R����ɤ(���S�_5#j��j�۳���6u�fZu�,M���i��1�r=��� ���.��[���#�
���^#)fe0oL`r�-��-�����v��m�X�J~JI�uvנyoK`l�� �����W(Y��-e����-��-��GL��Jq@�Ԫ���$0-$�g�ٹ�O��^�I܉DFF914��6H���ޘ���[�z[�������TtQ%�K@r7;Z�sr<n^R�;�%�n�Eg�ʝ��z3�VD[��Ǽ�2q��>��(P����V���$��$Q��@��}��bGo���{ۚ�;f���.VF(���n=��נr۹���ػ}4
����+��M��������X���'����=�V�R%C�����s�h���y�o�rO��lܓg���C�H�!��8i4����Ra�!00��@H�C�6�����$�
B
?Y s��M��Hb�h��B!��ZUBEbE��`� ��T�yV@�"W	xd]�FC0# �H� �$c���D���A$�hw#)DLF��S�X�1B �c`n�S@�@�8����E�=@��I�&����F
R�с����]	�*ɨ�H���*� D�����-5J̥�T�M��/��������t�ߟ��p ]Q��*�Y�/T���]��3uۮ:ع.�ɞ��������om��D��(�q$�Z�ͷ5��ݸ�H\[��M������΄�M<���N ��=�!J�H'��!�ϓ����V�`.ƫ�ѹz�)�۪��c�պ!w;]�e��pMXpԭ�,� �%�^W�Ipڶ$��7n��9/B:��e�jۀ�Y�	q�u�Yƙ�ܖ���.ҭ< s��ڔ3��{s�</i���H�,���Z(�f.s&p�w&;X�M��MQ&�#.��їi�9�
��^�x-�g�d�y�r�&���΋c.�����;?6�4�KÂu�����n��]�rFe8ecYѭ��OY�c'F��TjJ�loE����(�G`��^�/d�ێZ�٘�o5��Q�a<�>ɥL\u<v}3�Ggs���m���%ͧ�����³�6C�l�ֶB˜�I�8	Y�<��W)f��hM��=��d�ۍ����7a��57;n��t�Z �4Xn�q�8�]��/�22�lQ�MRvi�<g5]�\�:�n�>�����5�;d���/k�ݝ.CG`5�{��\G@����ו�˔���W���t-2�ڷgknQ�{J��*�#[���4�ӻ�]�u-�1��ʁ���ږ�����]"f֬m'�W6�n5s� 1tP@f�vۢ�v� �WS�(6i�R����t��vͶrE�F�*Ɠ&�\��k˛8-a��]�U��UR�ju��cP66�7ns[��u�&Kqts��sP��;hS���FwOY�e���*�|����]s
\�D�`�X��΅�2���c��ř吐��͓��ȽX��F��g(�6kvVUW�p����mRJÆɕ��Ij��FN�V!������7�M�%��ܭ��Av�.���`/U6�Z�\���a%ٷL:�e���qU*�NZNsA�7����S�"`^p��.*qG�c��!�z � ��tt��	� �x�
���{������)�q�]�6W+=���;�<nr����n8�k%��'��qD �.:���׳q�<�;q��Ҟ���0����^{���J�
���t�=��[t�/��u�{r��
67p�����X*����E�+��E�ݶG�|c���ջ;����n��Z���委x+�m���S��RH�4�ė^�T�$�����Uj��ݝq���4vdGU<:u�s֗���'���.v+�[<]:N#�S&Fۙ!���Ĥ���=�-��GL���*씯,���W�5ʰ>���%QTf�ڰ��,����1'B��d��z,����3�J)������`E�.�M�C���M����4�ڴ�;^��n�^�:��&�#m��uȘ��e�6H�{zcӒ�o�[�ƨ�g�O60��q�^[;��jޮ]����[&�k�=:qv.�ac�[��$t�=�1��r&�.�5M"~rr=��������w�rB�_|oy`wi��>��Ԓ��=����!�LRL�v�h�iq..�z9n��;sr6��m�j����Ș[��$t���Ioo���f6{���c��N-����ޑ� ����Ș�"�+Hq�5g�R�9��t;�z��`�Jwk1���%��v]J�6�2�������}��`�{���7;	j�K۫�-�57�8�bm��˝�@�]�@�s����o�?~�����ԐM%#m�\�X���v�͝X�R�!QO�Ձ��k�;��r��S1�D�Z�Ž�������z[	JL� n˹M�"~rr-������:��ڴ��V�|U����I�$�i'\�����۳�'G�E��5rg���0�:�Ʌ���&)&h��:�Z�}�@�m��>�nnHۙ!���Ĥ��Ș��$t�=�1��u�JN3#Q�b�8���V��n�~H\�k�h�!:H��Ҙ��7���V�q���M͇U�D����dZB�0 �o=��I�qy���'�bs���s�h�V��j�-�s@��po#��>z|M�=������Z�4x��>k�7����Fz��皉����b�6�r?�������SI{��%�-�)muK˴e+1r�5\���9�BP�L�����=��j�r�q�1�O�@NE�[n��z[K�0=��0%HGhW����,�`ޘ��r&��&[w4�ۛӘ���mbRM�ڴK�ǳ�wmX����LDBى]����}�e�5�V3n9�;�ej��۲�����f,.#��d���\_m�X��Ů���ʙ3<�]��<�;��\OR;�؜�͡\ ��Eu�v]r ������V�n�ѡ{�`qq��7K�On�;���ϟ��+���nu�'F�h��ζvCH8��gK�k�m&�$Ȭ�eI�pðN�s��K]�,��غz��������|�~|(�x����)�vs�۬*�]��g��c,pm�8͵р��yu�'Y�F�c����s�`cnՀ}�|��kvl��&���rD�91Šv۹����?bA��M���@���h\�Z��D<s�5w��=�1���Lm�L�:`�uLI�H�q9&���Z�}�@�s@>�l�..R�"`�8�%W&����l���/�;�y`c������q������ka�*G�ۤ�n8�պ�Ms���m�W�����p����5������0:\�����$���I�j�՚��ѹ$�����Snх�鹰3��l۵{
!L�Ǫ�R�1�͸�B�������j�-�s@�s���f6\N3 �F	Š}��6mڰ>��P���vl��I�k$�528qh۹�{����=��-�>ՠ}֒:�8�5)v6rf�hy�ppG��/�~{>=���wm�q_�ًZ�n	<s�4���}��]�@���{��=�{s@-��'	�Ȧ��s�`7M��B�U�}6��Z���7߿${|{Q1�MŠs����j�Q��P�T#�q�,�o��s����1�Ld�܋C߱{���`Ǽ�����	yV;�M�����@��I�I��{f����Oy|+�Z��hZ�L�xԍ��eK6w��/<��u�^3Gm�8l�nMuۂ��)�~m�~#�@�v��ՠv۹�߳>A�o��z�\�$�A�cQ���`}��oaL�wmX�{V:nofK�LI�k$�8��Š_{ۚ˝�Of%|��s��h\�Z��D<qMq5\VP��8��`o�ޛ��9�p�";_��s�~�M�'>�ڙ���d�=�ڴ��V��n���k�=���ff\�[��n!HIW8��ܫ��+�n�bs�p�i:c^�[l��R��q��c���L�FF�����@�s@�s���ՠ���"D�H	�l�:`ywK`t�˺[�B��@��I�I��{f���Z~�*���U����X�ssS3<U��T��yl�"`ywK`t��˺[��w.$�A�1Dqh.����7$��}��w��]�6�1�/;�����������]v�=��m���\@�ژ��V@��`C�A�vH�7m�u�v�	���Ս��vۤT�mXӶF�"\o���IϷ��Z���*�$����Ǘn^���Cm؝h^Scv�zŋ��զ�FP��On��{g��N�j����.�J�ݧ1u�ٝ�Ճ�(�쫹��m�s�qY�.��]�]�����[����~�����>���;gX ��J�l�s�J`�$��mgVP���n��(��Ο�wpOD�$n288���ۚ˺[�Ș]�����)Y�����73@�w��/���+|��w4��e�#c�M����j�>��VlD���Ve���x����qJ�$mF���~�ˎ�=����>]�z���~����U���2H$�&2@NG�cnՁ�����=�ٰ>��V�B���7��Ƹ���kW��0��$�5�r��݋�v�U���Л4t��cg�uq�,���}l�"`yoK����t��Z��1�ѱL#�;]�f~�� �
�X��V ?;����{ۚ˝�|�z�\�$�A�cR�����{V6�Y��IUd��X������f$��I$q��iǠv۪��{��t��j���=���;S�2!��nf���k�=�3�_Oy|�zm��2��!0O1��1����stu�7��q#�96]0�\�z�P�5ҟ����9�nHdM��m�H����@���X۵��	.�d���/V�Q�MWYY�,˼Lu�L�:`ywK`uv��fbGW���I�Lc�7"�/�߶nI���7)C���88+��@�`�RϦЂP	H�F�-@�k{ki��%��0�ȇ�!BYS�.��;�����9�TiI�!3J14�a���# |@���p �~C�$	����.�c,�� ��R$H$()�c�����hZr� �pu��J�u���44��Ch/��`�)��=�x�m`|��� T� �"�*#�|��!l(�7�ߦ��Of����HU2LP�L����\v��������k�-�s@�{Q�Ц9�6)�N-�nl�K����n�ڰ>��6�-տ{�����a�$��ή�S�]�j��pu-�����v�Dr���o�%�����'7$������U��v���ϔ(�Cv��@�1'�ǒF�#�ӏ@����}K�0<���%-�-J��E��nf��_j�-v�=��%�o���{ۚ��2�D�n6ؤ�@��6Ә��m�V(K�S��6��r㑷1)�(�n-��נ[n��_j�-v��R.jC�!A����v◶
��X=�d�s�����vi���q�3�&�C�9�m���}�@�ڴ�{^�r���@ٓ$��S�}K�0<���$��w�n4)�~��dIŠZ�Z����w4����x����c�8���j��ֽ�wvՁ��s`7Ḿ�ى:F�q��iǠ[n��>������^:�)B�9	
,_��������5���_;:���:Lل�8:ȝ�.{m����z͒.ʮ�{YCE��X61�;��c.�\��ӱ��e=u���n�c=��G.�ٛ{+��ʹ�4ri؞9�n͹�@���$�r����=�d��;�"׫X��q8.׆Ò���Wmn����nע��̥�M�ӸsD�t�qٵ�[��
vt�p�����n�������R�.��%TZ:�������˷�Λ���`k�ಧ�jbdC��4������]�@�^נ[n�w���"n7m)��\���:[I0;o�`J��q�ۘ��H�-�{^�m��x�V�k�hV���M��0O2�H��}K�0=/�`J�G�0L�""�L�:���]�@����$��:�$�����+2�8W��u6盋�miz�U���Y�ٮy���G��ҐIG?F�2	ǠZ�Z����w4����x��s �1��j�I�g}w��6�T�`�B
T8�8�;m�v�f�n���f$��I�G�n-�w4����j�>��h1V�&D��s��JS��"`r�Xws���2�D�n6�RE�Z�Z����:`rޖ���D�����?*�1��!�ª/e[;��k�k�Qزa�8�C\�����O�@�Š}_j�;m��:��������u{���ID6�&�&�:`rޖ���LK�ԑ��K�Li�d�1B)3@9o��k�l��T����!�*�I(��s��l����uUV�Q�ѱO�rh�V��_j�-�sCىr�M�-�bRE�pj 7��V9�6��� �{�76 ������v�vƢr.մt=g��V�X'wk1�����v7H�6*�)�,|�cnՁ��:�1�s��h3k}6�h��L�x�s���|���߿bE������n�w���܎4��G�v�V��_j�٘�����q[�\��q�ۘ���"�-~���_-�~�����9{�f���*`��� $1��u�]�;��뫣X�Q����m���g�;|��~��>��Z�V�T��O�	1�z�N�c���۬�H��ۃurg�GV��O����_	�0L�&(E&|�z�ՠ}�ڴm��9mi�Ē��LS8�鹿z!U������XNc���Yn{�,c��0n-��-�w4����j�9lĝp�H��HUrl6D������,鹰Գ���@�.���&)�'0i���c��76�X��m�VqBDE�@:���]~�.j��՚̉L05Z^�� cUl(�N|�T�l�E=������.y7@�|��&9M�w�*j�=�#��H�-���'6TGH��c��mO.K��y��k�ʻZf��v�}��@wl���PO�a�\n\�Z닩s��]9��PN��^k�Xk��r��u�K�
�m]�`��N� к�u��V��\"�E�������mv����gPy��,X��-ۋ8�c�x��;�|�o��^c����}����}ӾE踦��I<�?���>��Z��h����\r&�8�H�-�տ�ّ�G��Z���,鹽�2f��Rd�$�Sr-���4�������ՠv�WI�1&�H���V3����{6�X��Д/$������/���m�4���b�Ǡv����ӣ��t���_|�.��B�O�nEon5��V�nNc����Oܓ�m�ɒ�#���|:��8�yͳf���mo��ǎՁ��:�G�%��o�������RAH������?s�n�%
,s˺�>u�l����$�K����I���4����=��&��&N��t��Ytb�Ŗ������+�r��[۹���ؗ-��=���$m�q���)��_\���u������1���S8ݸ�ss�w%av���=v1�n�<gp�-�ڳnӗ���fr���|�b���8Z<�O�0"�-���K`N���6)�LI�52
93@�v��~ċ毞��on��?$w��M�$���bі�WrO~��ٹ'�����U:!D��X%�v����J�MO+��C�����z��{�ۚ�h~W�_=����dpN$7��;V�(����ڗ�`u�9�;���w�ݬ��n��k���m
�hD㎱�k�����Ϗmm����8��{��F��9z3�X������K]-���&�h-�ˊ'���#q��v��g�d������K����6 �666?���f�A�����۟�j�3F�����WZ͈<�����k߮�A�����~��A�,lg~͈<�����j��lA�lll~���]hֲ�ue�d��j�A�llU߽���A����u��؃� � � � ����ٱ�A�A�P��6V �(@�~<��D>pA�w��A����O~�-�n]�Ժ�h؃� � � � �����A�lllP�E�	��w��lA�666>�����A�A�A�A��߸lA�lll�w{�����z�����3q��N�I�iHN$6�ᵎ6蜳h�\c���\7d+��-֮�A���ߵ}�6 �666=��~�y߽����A�A�A�A�u��؃� � � � ���~.�Z�&jLՒeֳb �`�`�`�������"�������y����؃� � � � ����f�@S�FA �`��߶K��솲�5.j�3Wb �`�`�`�����yg~͈<��*6=���ٱ�A�A�A�A��{�؃� � � � ��5����f��֌��6 �66/� 1D� ������A��������؃� � � � �����A�llP,~��y�ߋ��u5n�\�.�Wb �`�`�`��ھ��y�׿]�<��������b �`�`�`������A�A�A�A�|�!��LRI	��$�~ ФO%�،T��+Ah�!As ����hP����e"i,a)��\T��2�@ ��^�R!�5T:}� �aN�|� qCB��)�F,q�� ���bA��:�ld>n0 zT3[u ���@8m��7q�H` V��o�H��LG�M�PC��4�)A1�1 @��)� �H�D�!�vE j�\Ɲӧ~ץ����I����8p;���������\��)s�6�`��Bnnwj�c��N��)���.^����+�^֥�7�ms�.�E��0FZL���Wem[r-k��Z�U��;F٦��q�mB���讥�y�)��!����c�k�t崢B�m���z�a�R�F�9n� +P��s*��mnV]����{TB�B�K#HM�Xu��b�b�]�HGK��On�n{kK!�N��r�KQs<
٩L[�fn����=�2�\�-��Y����-Q1S��yml�Y�$�w6'`�޵�3���Ѻ�����+,x��Hy�-�,�5�N����3�qKϠ�؊���*���XÑm��8��XV�UB�qѝ�»�B�wI����(���m'����i����	�i;D`�����m����N��X{'l�T��
���*+7��y��V�4}��yVA݈��mgĒ9Ĕif]�m�E�rp��[b����'<�<l�`8M�-pk%s��b^�2�@�;lgnܤ��5�A�l-��e7f��ӻ�:���t��q5��ڻlqŸqx'�����&���M(��J����(ZGk)ݖƈ�Fٴ���v��$p]"ls[X������GfC�v����l\M�u�;x:�C 	�sh��M��[��i�'m)՛f�X+t;��9��j���8�1Z���*�#Q��ui����L��'v�`������;'7KQq�+l��f��ت�ܽ2�]p��Ƶ�
\���氘9�9\�Oe��`2D��;j\�t�Kё��	�(�G6�Г�ڨ��\�R��i����aL�M�8�VEd��rHml�D��� �5�N2���$K�]p',�Y#N�Ӷ�ڶ s�+jUR�̏�+���:5MT�N�x�j��
�;zjCk��nW�D��d}���ޣ5���<6H\��UPG�� -���*�5N�a��Nt�<�>�{���(�Z�>S�8�����@�x`�x6j���\~?,�=S��һ=9ݲ�Q�zj:�.L\o[n@G9Cg�/lVu{m�\;��p뵻5��S��9��Y\�'X��J�6{vR_=�:P�򗳋�[���*[�K�vw 1&nC�ru�1֐��X�x��o:wd� FvQ. kuؗ��+c%r����������+�v�N��Z�Փ�,K��m�FN�OEr]8?���ǑV;VE�c�Z�^��ѥ6�ΝGTkҗ<��T����D�ssy5��њ�\�u��muN�����u��؃� � � � ����6 �666>�~�AD9~���؃� � � � ��{��ѫ�-՗5��kWb �`�`�`����p؃� � � � �����A�lll{�W߳b �`�`�`����������������Z��.�L�n��b �`�`�`������y����؃� � � � �����A�lllw��y���&g	2�N\�F[�]�<���*� ����f�A�������b �`�`�`����p؃� � ب���߮�A����;��u����欓.��y����'�ݵ`d���:�qՁ�c&gk�R�:Ѷy�+7n=��`��Ş���έ˯g�ۮ n�W�25?�ffb��� ���X���O��Lۑ06Z�l��0$."�x�j噫�s4nI߳޻��Tx ��-�Q���M���=��v��D�f�=�LC��i�8�毞�z�V�Q;�mX��6O8:9ʪ�.P�����r�=�u����mX���y%}��9]�Ȣ�N1�"�-���=��y|�W�@�}�@�:�q��ס,^�F̵쭗bۮ�����ݧP�Ԫv�����f�Å.�q5�6��߳`c��V��>P�z;A�o�X�x�pƘ�4�Zk]�@�}�@��s@��|��K��PqLN �*�ͧ�`7�Ւ�D)I#� P�@m1G
R�b�1
��������@�jנ}��W ���Y5\�B�*���V�����S���ʴ����5��73@��@�k��6_D������%b˵��\�I�qF!�]Uۤл$�P��N�����y�T��.(3��c����~}~m�_j�-���;�j�.^²A�d�]�,řl��0$���r&K]��f~�H�=�x8�n1�"�=�mX�nl�ID�ڗ�`f�ٰq��!16�BLQɚx�Zk]�I>�w�r~C�`@��8I%�w޿+���)U5�T�<U3�&K]-���&�0;nD���߽��߽��q���1G�ٞݍDT+��5����3�6��{�+�B7��o��18�jG�?����{w4�j�;Z�z���0J�!�Š[۪��!L���6ڗ�`<�s`59#�pq&��1���h�v�?�/W|�z�s@9ځ� D�H�b������}N��|�������a�H'�$1��E#�/_j�-�ܰi��1���>Q��Jz!Vx� S����f���;��g��T�eC�.+m������"����0/n��Ks)�z��]�1�CXE4I,gvݼx.ӽp����4��k�@g!���tk��æ��� �{4��[�=v�n��捳Cg�$KȽ2���v�u�1[G��s4��.�݁�y���gu�6���AF�� 蘃TPp�۩,=[�H�6����i���}�����󿂗Wk$N�Q�x��
��)P�Z�C{=	D�#��[�\��N��$�$��U�K��Z�i��1��//ٜa����{��\�M4�BLQɚ�77�I)��Kڰ5�ٰ�j�	,ċ�x6LXӆ4�1�"�/��z��Zs�䭳 �ՠ9����4M@�fff+�ڴo�4�j�;Z�z�����y�#�@��aDD-�n��=�{V��6������ی���ֱ�͕���b��=�Y�o.nYmG<�8ʞ�^n�������[�`c��V��?��~DD%���s@/��@�$��(��;Z�{T.$�J���s`6ݫ���؄�!${=a�9���nb�H���-Ύ��"`t�����Yuk�EW(��rl5(���u���ܭٰ1��z��Z�k�"jd$���>�s`j��I�%�|�{6x�X����oϻ���¬����.5�R�ͧ[����l�<�x����a5'%y\��`c��V��6x�j�
�CW}�qR��S��z���D%2n��`l��X�q�ꄔ%�J!*�v�t
�«�s���������=~��s��@pD��;��+�w��hr�P�I��&ne��D%.�v��/j�yX���"w^��뇗�c�$Cj9���k�=	(������V���������<BMї.��셺˸==�k�k�Qػ=���<jb�:u��ۖ�~m��\s`>�j�s�u�B��3j^Ձ�[�92!�!��܋@��s�g�.�=�KڰkިJ"#�(�=��_+�,M���rf��������k�/j�-���9ڪ65�9��)�N=f$��%�X��l�ڰ�
!r����3h�o�׹w$��t�֮����S�U��X�����ߗ�nSٰ;Z�z�]1)��`(O�H���uv�k/��X���Y����ᱻ^�n��l��7�ɂQŠ[۹�^>ՠv����3�|��w�@�+�o�P���73@}�s`c��V�c��v��BI/~�ٍ����La$�m)"�=�׿���X��%
���V�=�3���Nd�71H�z��3��e��=����������W�@�ɑ�D�s�`7�Ձ���(Qw���������{����b#&*D���w�;���Ѻ��P�4A�M�k@�&s�q�D�v2��XԴ'���qmcn4�f�w:h����O�Pbv�j�cq8�cQ�]�M�s��&��0��%\9�.4���՗ƻېcq���5q������p�#���{t����%�i[�	n�u�b�8��e�u��NwQ�s]�r-�N�:�m�ip�����߾�w�|;c�&�)�a 7H�[�ɷn���V^���3�)�v맡��l8R�W]����~� �S����>�����{j�{�d�R���JciŠv����?g��ؑ��`n��`>�9�B����ƵW9��ʞ&�����[n�x�V��կ@�.�N<�pr�@�����́����ԔB��=�e����l�R`��h��h�Z��ڴ{w4AዹpY�~h��f��Tn�"q��h�pw��|>y7��
؆� ������CV�~�l�bm�"��k��@�}�`7���B��7)��P�\��qr�3E֮���{���D�0$HT�S�'� �����ٹ'��~����k�����#�~�'&D4D7��X�mX��l�J���/j�ܧ�`^۲8
	�2b�L�/j�;jqՀ�X���(K�
!%Y�{���{?����O�iLm8�u�נ~�߽�|����4�ڴ�Z���7��.��F�Zݸ� �7n݇v�c]<r\ⶌ��e5o������|��=%�d�����gɁ�#���ֺ[��\Ç	���\��ݫ��(�Ty��t�����Z]��ęD��	��+;X���T�>���!A! bö�'/P�D 5 A��GR B��X�E*�#.)AŁH����'5�1�4��A��	AH�Î�h XD_f�<1;�b��ѵM�  �l@����Q�2�+ $��i\x�h# F	�{��t�*b��L�	� 4)�1J(k���>,��VՌtqQ�Rr�������y$��JT�s��=��^[��w��h�gar5Ȍnd��U���2��Dy(�=�utu���k���v'b�!
~��yl���s�6�:�l�7;�v[��j�O&39(ak""�'$4���x�V�ε���3�g�9�<h����
	�2E1,̦m�L�]-�������_��G���65�I�lSN-���zvA��#�m�L-%J���Yk*��O9V
"{���;����c�#U��{�:�ARw�N��x*E'&N�ݦm�L�]-����U~�J��~�qg��hsv덜��f�wM�T㎎r������[xw^,v�M�{�������]�n�=��ɰ;�8��}�2���j�:�+'���JH�u�׾��1#ݳƁ�{ۚ�o�1#�
�ƌu�<��`k|����j�D%3�[�`ej��.Z��""�7$4?��f$����7+vl�N:���zX��ĔI52`���w�ՠg���%�|k�ͻV�J%�����͙�Dt��g�(s�Тb����آ�.\G(Gc]l�9}�n�c�d��Qڰ�99�mb�.z��]��&���<��s��1=V�ign�'�H��X��:�d��y׮��(��:��鳆�T(�l�y���v�v^���6w,G�k�Yu�Ob�3u�h�kԵ����m	�b.�m�/*�ckLr�X��g?����^�w���:���h�%�r�Q�^�b^�k�gh_�q�D�6�hJ���ٻ���0LȆ��ԋ�s�{���"`zH遻r&���]��K*��Y��ݹ�GLۑ07�q��B�I*�v�:�9<&�Up��`g��Vz��=3���X��6]��ĜJ2AI�i������b�}�4֯���;V���s@9ܪ�~�l��5U3�r�X
g7g�;���r�h�U,�m��11A�=(-m���܉]�;r�N��҅���S��f�S1��E#�9�j�>��h�����|����s�瓏""�(���'=�l�W�"��U
�9^�h�_=�v����(�ɑ��I3@��@�Z�z{333�]�����{ۚ�ʍ�`��S�r�X�76ͻV	%9�zX]=���"S&R=�v�����ߗ�fo4�;�8����2��J�RFuJ�ݮ�).&��,u�qv�syu��v�E�r�1E#�(��p�����z���S���D(�C2�f��zU{�)�A8�ә�s�ՠs�v�������j����ƶv�G8U�MM����^Ձ��sg�"���k@��ՠs�w�s1��E#��Ng7f���ڰ;�nl<�Jq�^ց�;�MH�h�R4��h[w4%����u/j��i��5%�`�j���7S%�l��M{ŷ]qg������;u(�.�л�������|�0뤸*��_��`oZ�lۑ0=$t��*#cX/�Ɣ�@�Z�{����#�~���������Q	L��rm�r��T�O9Veǹ�ݫ=
L�V�h�W�@�^�e���'��ݫ������V��Iz�%1"�Pb�@���s?|K<�.u��jD��	 �N+�����P�y/k�2sv���Xo����H.�Nѹ�r���;�=���3���z�5�3�Đv�>��aM?�R���[���Z�<�v����@��{�KbM�h��)�@��@}nՁ��s`u���F��3kI�D�B� �}���} u�u�\��^ؓI&A�JI�8�Z�]-��d��0'J�yj�W�bʴ�e���ղ[l���^��% �N���L�5d2�JSN������X�r�J���5�͔5��7\\��8W)�a�s���n�ݮ7X棟=ن8э=���z�$k�m�ۮM��Ռ$��G��x�s�;WvW���`�rG�D0X8���O&xŵ۴�;v�=�sͶ�f���P��*,�v��WW��lp�]s9��s��H�pl֨�;.]7Eq��ޭ�`e�	�����{�޺�8���o�ݒ�{tYgFdv�`��ㅳ�9ش��ئ9^:�1�7I$�d��9l���#���06Z�l�w����'�yn��YM��נqr׾H�i��)�B8*��+3y���S���(��g'7j���ۚ��J��26I�rE���˾�}l]����#���L�u�$�ƌNa"��.Z����9�M�k���*�Hr$(5f9 ���,Ls����緱Ж��WIڊwb����"�qȴ���9�M�k��qڴ
�lI�����s$���2�}
!�P�B^��n��V:{6����ˋbX/�Jcm�@�k��ۑ3�/��:`wO�0<���^VZ�FҘ	H�=�3�.v{�@��������;Z����w��xG���GLގ�-IlmȘj����9�̘��ZE܍l��2��6]����Z�w�[�[T��F��@��AsZl8r�t����-��I0�\�6I�m��;Z���#�~��=�{s@�j�;p�qli9����u�ܓ�g�w$��훂� DH��GzV�$D�iI�GHt��ο��s���=���7&	�#���L	$t�ݹ��-��r&W�$�D�Ɉ�rf��;V���߽���W@n��nՀt�*fI�1�����a��a�c��k�v�u�X���f���Gb$q���`�8)����կ@�܉�$���"`j�IJ�.��%��-��}I0=�"`t�_���27H���rJG+�9ɰ7wmXv��<�e�N�X8��9-Y�'�B8&'3@��ՠv�k�O���nO�qUO��%ACO��ޟs4���dɄh�1��@�jK`jޖ��GLmȘДV�k���i�gZv�W�nv��������ֹ5v<�y�+3v��n]fu��O�:�nՁ�i����{S�Vu��m�Ms�=�w4��ZkV����}����/_D��bd��Ǘ�L�����jK`n�D��GL�jh�&+�S<US�M��BJ^�wj�̧�`6ݫ(Q
{�ݛ%����6���H�q���w4����_{7$���=�F����l�SЉ�#��9���L��#	��5��p���B��� A$@�.��/"�mf�N� Π}� �����l��>D��ObYj�u"	@ �:�@�T��l��ЕZ�y�7/������$�o����A��k-n22�J�A�V}��8����l�L��Nzڸs��L���v��1ezE-QY���Ō!���UvQ6�6U^ݪ�"�
�ΓOOt�U@d
�8Ւ�vWg�Le"�3r��j5�h3t��9���@AKUU�hө�� ��=B�WA`ւ�ȴ�WG!r@uT�k�)���NveU��7X���X��b3�=�0�;,���-�M���#�$��'<�s76nݝ����
�9:�P��u]uc�D�g<�7���I�f�g+v��웈����ee�L�NKf��ˎd�P@
��w
�*�kH��Pqh�a�s�q��cp�X���an��j���X")�RCCq�"�a5۴���qӡ���f^���k��W[cr�j��ڽl���i����`�u5�(U�Z�V��h��қ`u���6�+s���E�%m�WL<�T��������3�*�E�)�8�]pFե����э:���y���U��
�:��8��8���M+ԭ�}f��7L;nk��݌��t��H���=�s�8���:�U;\u�m�q��5n�sh�u*�����vĂf5m� �m%�`��G	��:�\�Զ���;Dd,���֫y�ۄ�3=�� f�5�`$�@k�m	����T�{E[�M�z�H�\X^p�H&�ɣ��m�9�I���v:E��պRX	�"Ү]��Ӻ�U(r:ʺ퇎����������9` s'I��g���b�*���^c�z<�_
�V���R�[��2s�d����>M���Br�
d]��c-��79�+	\�VՒ7V�r���sT�2��8�Z��F#����lq�]`U���5UWNF�I�nv����cQ+J��:#��U�v:���V�W@Jэm�^m!i�wTN��d��-�2�H).=��se,�m��8���y)<�U�ʝi{���|�3�"7I�m<��J@~@(�P�b�&����>A� �"CA����!�ϡ���ͮ�ฎ�A���[\ZB�tkh�*�a�����7����v��؛�:7%�wb�r��Zg�]���[��6T�cZSxǈKOc��ݻ+�s�LP砕U��n�n�F7���֒�N�+�q/cg'b��p�m�f��v��"�T�F����#��m���z�;3�f��U=8H3]چ�H�::vn5{�wwu�/���q�e��;VSf��mj���X������/��"简����X�i��pm��>�h�[�BKВ���}6�g��rg�����19��v���^��>ՠ[n��33�bA̾3�1�$�M9"�'־����0$���r&J%\[Ncdd�G����{=�{�����sa�P��{�ݫ�Ml�R⚓�d��E�[n���@�jנs��h
�Z�@�X� �
4I+�GW��m���-��]��nף����w{�_>|� LL��1G&|:��v�k�9��>�CwvՁ�������L�MO96{/��x��(|�rw���-���>�o����ؑ�jK� ڃ�K(-f[��Ɂ'GLmȘ-uz�Ļ��j4�`G�on��i��1��J"�q��.vv�$�<r
D����;V���k�9ǎl�ڰ<��!KZ�'(���C�ռ���lc�ey��x����|�<�v�u��1����f�����H�ے.���k���q�&�0=�"`t��Ryi^U�J�řl��tt��܉���K~���9]4�'�$�-޾�ܓ�g�w6Ԅ_�#�ˊ���# H`Ep 9��/>z��ZW�$4&"LRI�ݦ���S����͇�P���{}�`{�<���b�<�k����S����L	::`ñ �R"�1!���X��H t�[Ӡ�b^�(2�u&�ܗ8��s�'�H{3TԖ�q�J`5#����@o��|g��_H=�{V�S.M�5Y�"�-���~Ď��Ɓ|���9�ڷ�?$yU��sD� �I9�+�����T�=	B�̧�`wwo4�o��$�M�!�s�v���s`|۵`�Q��+�����~��������6!�#R=�}�@���������]��*�Eb��uv��^\����;-��+s��]���frE�@d��E�}m��9��Vr�lD}!ܭٰ6^�4��hⓜU\����~P�L�[ڰ;��6ͻW�	B�QT{���W"&+�S�*�2�/�����LI07z:`yr��B5��?%#�����yhyu{�f�����9m����_�f�m���-�w��d:Z�,?���ߜ� ?��{��>��I!I��I%7�=���(��U	AR
�@3߭����\�њ�z�Ug�U�8�,!�كiX�'m�sͩ��4(- ��gŹ�X�짫�a�M��;F^�,U2� r�ڧbes�4<�\��n��6v6
�)�ܻ71�
�u��ɭڱ�n�D����!#���i+�����9�T���n�����/�5%�vm�q]��s���Gh�8k�W,�p��Af�E�:I�g���qy4u>zq�ׁ���-�����G	9O��g��}m���A�:m$\��k[�4g-��~��Ü��{�f�m��w~��8�]^��ԒK�nx�xA�bm�3�I!wKƒK۝��Z�um$�����K��ű��6F���椒���{�%�GV����ޟz���^4�[�ܩ��,���"���q�I/�����H]�񤾯�W{�|��O��]�Ɉ�$�bԒ_s�����~O��|�K����J��ũ$����܇|���P�u�r��̧H�KϵƌY|�dݺ'*��װ�SF(;m��J����[v�y����[o�}�?�Nf[~�p�-���F�B4���?%#��K�N���f~�Ψ|��G﾿���wm��~�Ü��}�9�$�&%�\Q��Dq�_|�W��M$�����_�_�U݋���I%����$�����8��AH�&�-I%�;~ϾI!N��$��:/y$�\t�I%�%C���Ci9�|�B��jI/~��3����$����Ԓ_s���䒹\vAdx/���J�JG�g7#]�;p�i�^���9�����r�&Zo���t^�IN��4�^ޞ�y$�:^4�[����<u�CT?��8�����Չt����$�����i$���{�$��+�a�&(�H�ũ$��o���$+�楳oMD$�L_"u?l ��'ݞ��$����4�RtI{��Zʴԙ��/�߱���5$�;/��$�뻋RI}�߳�K�Ԗ�i4��sRI{s���Ju�I�����0N��ݭ��_�Ũ����:�vq�4��/$�WH�g���!'X,k�Ch�n��gm����}��� ��m�Lv�qLq�q��@����s��u�p�=���O<�P��u6��).�"�+�`�>���&m�Ls�s@2�*,I9����rMg���脕c����}6��j��%�	.��["A
�E�sf͚;Sm�I�Ɍs�-�������X�,�X���B��>a���su�q�Nq3�Z���[bǜ�����kZAs�V�����wa��\�鬽��Θ�L`{o�`rޖ�� ���51��� ����>ՠus��s�s}��~Ď��Zژ�r(Ƴ���`o\�09oK`{z:`�1�x�.��Ɩ(�8��v��uڰ�>Xl%
{�{6�jvN*䔯0W����`{z:`�1����}�@�̥Ĭ��H� �3��(�h|���d���^p��0�mu�f����W��nk��<=nn��/�U5i�K�ctq�� U� 8k��tn��<ps��FӜG��JÑ�7mn0I�5e��y�F,q�k��-��8�gF�ķ -�[��V���`	�۷�x�oa�!��@^�]Ey�6N܎����,�v�'��:;:[{��߻�����~e�<�:r�00�q	��:�]���,X�\��=�o8��Hs֍v��B8n��ߟ��k��9�3��?(��c�Z�=(��?�I�l�G�hq���}�@������8�W��Ǔ�qȴ�c���g�B^Q
��o�`c���w��L26���$�-�v�hצ0=��0;o�`M�I�$��kMO8�珖�Q������l��s@2�!bŖ�~�9RO���'�����ca�`ye;�����<t�v�R�Z'^YV�1����}��� ���ĺ���"X��Z˝�^~�	�� ��
	�� hԀR ��ҁ��'{=��ٰ��Xv���DDB�kkC����r	�&�z;}��s�i��Ĺ�|�.�= �.R"a�(�bs4?����IoO���s���ޖ���t��\�+�cDj8ܓ@���h.v����{zc�%�/1#.�Wx�+��D�&��z�D[<���"Y8���Vz���ww����I�ɍ�8�_���}�����m�L	��*V��*�eZ��`{z:`ޘ���D��ޖ��_�=�xKr$��SjL�v�hs;빣�P�1!i*	+�=�KY)+J@%��F��(Ƭh$5�0b� z+@��@%�!	D� �G� @��*¡���P*��0�2�"l!�C�}��1R$R�H�!Ki�N�H�F֡M�W4���#117� �t*m��K�����*ʒ��(@ B�Km`�R��X���VP�c�r�����οi�!��)�&�,�Z���
�j���D4H�!Ve3j`qS�!�H`� ��p��aU"%�`l!��Q�(@��BL(P��>y��JJc
�Ƥ�(�kbs���In	��G�@��
$ �P#F^qH�[��Y@!y���>G G�>\;�_�`���E@���T����
�J�%���r�X��Xܩk&(�$b�Ƥ��}�@�s��s�sC߿~K�����*�dmȖ)2�Yx�[��ގ���0=��0?��g�^����܆�,�#O����f����	v��ka�ynY-3�v�ʝ��0<��M��o��4�v��>�����~(��d��X����8������5��=�1����-���遪������rM�>ՠ|����f%��nh;}4r̸�ı�ɍ�9\��zJ"{X����V�q����@�}��w$���3k2���nk�`}�v��$�c�s�c���Oq���~q�`����7Kqb����c��
��:鷝���l�=A�u���ڰV0nm��V�)�{zc�}�z[�����Zژ��$b�Ƥ��}�}���}l����	�Ir%e��%K2�-^`��ޖ����?�~����0=�<h�WBd�x��M��?�~_t���7����������C��T�����5�`w,(�Kqޟ}{�ٹ'��nIM� �F �R��0w��5�d��WK0]���917l�Q'm���۰���@�rX^N��]�iQ8�\;3����7l6ʾ:.*tt=:�<�r�d=0v�<�m�j���v]���K=�W����XC��S�ۜ����N�F���V;V�`��9�g���sX]Z�xz��X��}1 s�Vj��vy�K<I��Dv6���n��:���p�4��Pبy���o5�%$ɩ�f��)�ik
����u;�g�{.��MGb��<�s��4]���,Ȇ�q�'�[��@�s������߾@s��@�}3؜ı�ɍ�c��z[oGL��{ ��}��26��)�9�y۹�s�i���{�x�8�|��D�H���5&h�䷧����|0<���&�t���jdm�ƣk�h���?�~����v�s@>�l�U�
cS�X<$��G����讹��YP��m)���ᱵ�W��8�r%�Lq�!�|������ ���@�즀^�w	�"c�N!6�qڹ��RI%�	B�|�y`o�<h.v� ��E"&D$Q������q�yB���ڰ7ڰ:���,$s"Q����?�������9O���7����ٕ)^QJ��+/,�����-�7����	���/F�[��18��$�BAG>��b7[�Ծ����ٜ�nӸ�r~���_��KD�I�r?��o�4�v������8�|��xK`��p��Rf�}�|�P�(Jd�|����ڰqڿB�ċ�孩����JI�{�x�>����rT(X�+�����{���]E�ۑ,�c�9��נ^v�h���e4�+�L���	��U���Ձ�J"{�y���XOqՁ�Q�È[B�I�*UJ��Qȭ��f�9/�������[>_H�&��Iޢ�"ɑ���ng ;}�4��h.v��s@��;p��̈mG�h���~����}l����ٙq9�'�&G�h.v��v�h���}�@�v��#h�	0Nr�?%J"+���1�`}��6PV 
��T����׵��T=�$c��ƚ�4�v���;'����`{z:`zE���aE���U�I��	5[��y�r'Rlm�y��T�������ڦ�mL��8�mbRO��]��oL`{z:`yoK`M�K�0�Y�V^U��0oL`{z:`yoK`{o�h�Wp�"&9�nM�v�hOq՞I$��(QU���`�ܰڊDL�H�6�s4�;^��j`ޘ���t��Et�ayyX����\�Xv�́�%
q﫠c�Z�>��ٹ'��"��B�
��ߍ��C��ۉ�R<]g�y�:�9]����J� �l.нظ���f~����l��q�sk`�v��ms���V�P��)s̜�8�j�ƽa㓮^�9�v����jI@��E���d;78v�7/4����v.g���p�};<[t9�I��ґ�=n �ntG9/WX��!�+�gcg��T\�g�V���g��:�l��*cC2@�qD�ʷ37?~��ϵ=�6*�wk��Я,rn.tv�=4v|9��N��r�ع��n�n�<��9�?�o��Xw���:��C�Of��OfU<26��)�rM�v�o�331#���@�]��>\�zoUC�`�81��)��-����-�����*���ۃ�F��@���h.v��v�h{�~����_X��H1��G�t,���ޖ���t��ޖ���D�������'���m8.�r���-\ٶ�Gk	9B�?�s�IgM�^�t�̍����b[�+�����L-�lm�_�_��Wo��w�G����m1��˝���"�%�Of���ڰ>�;Ve(X(�DF�Q����V���k���\������s�PN�<�c�D�����m�����L-�lm�LWҬ�Q��I�r=�v�h���}�@�s���߸Ξk����㭘Q3�O���^Ѻ��N(�n����؜X��Ǥ�z����5&p���@��D��ޗ���+ ��h��W�f]�����������=�:`�پ��}b�ȓ���c�H�����s��f�Ӣ��'PNrw9�nI���h�Wp�"#$�6ܚ�������ݬsa䗢*��`ޓ�$�Hy"�m73@>�l�?�����v�hs�s@�+�\F7�mDim]1�ǅ�Cf�5�Q㰙�����I��utL�[�
8��rM�>ՠ|����۹�s�h��bx�dq�9���_�L�Ƕ����ݬs~S&k��E�(�d$�9���nh����&���@������j�V�S=Ǽ�;��l����В�@ �H@I�w���f������E$dn6�)&��j�oL`{z:`ޘ�ݢP�Y-�p�`�ۮ@��y�ټF�)���]vͫn���l�$&G�"#Q���x)�}�٠}�v����D}!ܧ�`�֣���,�ewy�oGL�������\�Dȁ�1�Nf�}�|�k٩(S'q�,Ƕ�ȱ�`��7$�/j���4��� ���@��A9�'�&G�0oL`M��{zcm�L���@�	`��2 Ek\`̤���р��D�X��d�Qq��U�������B�HF��Ј�p��@�R,)���ڎГ(X �h�B0S8�H���s�!�P0\�G��BB{�I�[5�|���i!pŦ`��$�!��ֵ��T%��Mn0�	t�@N�Ձ��bs��У�G'n��X�qýu�nɽ��\����>[.��۝��Zq��V����C��L���n������ʱ�e^�v��d	IL�n��Z�jJܦ˶R�G�q�.���Lh�;
�k8eC�-U��mt�֓�a����C�	����F�l+��$�s�κU�����]�y��Bt*�h�/������v�W$�[��..�N�Wi�9�4��d�-�W�Þ�0kh�\]^���k��٨b5m��WU�8�u���"[��ڱ�C3[Z�6�9�	bU�m[Ky��K+$H@��M���c�C���N�w6�Uv�Ǳ�l�`p�����6� ��u�����X%\���:)�w:Rx�I�Ό[���G9+�I��/nڷQ��G^WdЖ��ѓ)�93ɺ9�i:�;Ng[�H.UV�N��s�W#�p��z�k�.����k(Ӯ�����s��`m�����9�llll,���Z�r�Z���g�9|�9�s�A���- @���굕���ם��6���>.�����0kl�n��ܐ���ֶ���ض�UUSx�s�v�wV��&�T��m��/�o>+�NMQ��g$��UUL�쨻��5�5��Y�ۉD2]��>'�v�~e�ڦ�@���� 3�f(]Ű'�UM�Z�6�Tڌ����a��Z���6%�j��@J�<m�U���cA)]q�[�:8|��٧-�[�fbt k�ҏnm��c��A�< ����A��l�J]c��:�Ѧ�GU���ܧJ�F׉���vEc���T`��hU��m�`d�1PJ�`�[D�0��U�[��tJ�;nV��C��YGr��r#Z�ӧnm��2Ԗ�À�ٵMK!�o��t�[�����$n��i�J ������r�rՉ7
�]�Z:��"A]5�,��mR����y���%���d�\C��l�f�ZЧ�>���]��(莜J_�N��A�. Q�E*��x6�x��f�̓�Zp��\�E�'gn,ɧ�;O�e�P���mTƶ�<�"�	�+���lvl�9�hfxM�b@87V����]��s�c��FR�e�w�]&ӑm�MC����]7]�9�w W�"��XS����n_!���R{.�3��v��f��[r��bg��y�a�J-d5�8ç�0�'&g�6���|�����n�֞g\���;�7�|��K��n�Ӹ5>H���9�)�N���RgH&�͒,���{����"�a2bNI�������4�ڴ�v���z���Ʀ8㙠w/�(�7)��q�,�v�RI{���r�����|�jt��|��������yBI)�Ƕ����q�I�&A��G1�Z�;f�y۹�w,=
�S�ǳ`k[�.rJ��'�E��coGL��o�`ޘ�ߜO�Rx���,+�S��&���uvB�s69�6��ޭμ�)zѮ���sʼ���	��0oL`M�遨�P�(�#Q����[����qg��!/(J"#�y~��~�`w/��39�O�����r- �o��7����	��06]t+�Ë�8�k���$�DW����1�`>�j���4�݉�ğ�Ʀ8㙠ޘ��} ���ގ�mD 8��u�;hR*�p��m�h�-&6*��S�k�<!���\���6�h�A��̀}�|�q��
!%��{�����dmds)�}�ٿٙ��ۚ��M��V�{�P�"$*�%UW9`gqڰ���TDD%�(Q�;�S�	DNb����$����t�H���m9�����g�X�ܰ3վ� ���`gqڰ;&Jx��L�G�hWڴ����.v�|�����@���V]���j��.t)�HN�Sk�H�Ǳڣ����-����-���6l7���&7#�|��M���{zc��&ˮ���+qL�9�;���D�w����ٰ��4Kv'���jc�9��;f��sg�DL�Ǽ�=�`cmZ��$cn6�)&�����\��Z]�zw�T��D�vD\������I-R�F�K#��H��v��?~���> 篦��}�@/�)��,�HF���-��m�Qk˛"n�2l;�-�3�e�y��r�]HO$���zy۹�^٠}_j�:����.R"dC��!�3@>x�~�	L��{6�{Vw��L�%�I�JH#Q��<��ק����x�Հw^�����p$�K��,̼���-���� ��K�r̯�	��#r=����<��^��;��l���Iy���ߛ�?O�7G�����=���73�*�6.��$��]-����Ӎ��q�<z�:�uL�v9�{pZ��	V��XN�;{Yۋhͧq��S\��".����gj�!ЂRG!\���u;�g�A�MY\�P�c�����5�yH�z��5��g]Ԙ(����#q���;[<����wE)�wc���w`�u:we���뛄#f�3V�4Rg��)�.��T��s3��tn��$��WN.�E/8�k�wq��f���}�E���a�d����m���o���09oK`v�t�ޒ�]�]�e��mbRM��V��*���/o�4��7��o����F�G1��hv��;z:`�1��}uL�����A��mǠw��������g�ث������"dC��!�3@=:c��&-�lގ��t~�Y�ݝƞ��q[R]*Q�V��>����Q��7���n���\l��-_6�ϯ�L���0oL`ytR�0J�9ʮr�ɰ���Do�yW{�V}��}_j�8�Ux8�m��I�<�`v�t�=�1��} �������y���f�}�٠}_j���4�s@�7�ܑ���ĳ1��} ���oGL��q����n�n�
-�v�0��'@�Jݩ�q�^*�y�\\�I!�s�����0;z:`ޙ�y�s���㧔����'�rh�n�}�������{zc �%C���Y��[�7$������;� 3���T� Z�B*"Ȃ��%A�h��h�n���RVbN@y���?��}�>Lz}�	�0oL`|�U� &��$���Z�;f�y�j�>�>X���܅D)!IU4��x�tlL��%އGm�zތѺn6z�e -�����wC?��]j�j�x�%�bX�߯�ʛ�bX�%������bX�'������%�b^}�kiȖ%�bw��z�&jeњ�f���bX�%������bX�'������%�b^}�kiȖ%�b{��*|��{��7���߽��j���|�r%�bX��֦�X�%�y�}��"X�!�2'�_�*n%�bX�������bX�'g����I���Mf�%֭Mı,K���[ND�,Kݾ�Sq,Kļ���ӑ,K�� "�� ��[�z��Kĳ���_�����V�{���oq��Ov�eMı,K���[ND�,K��z��Kı/>ﵴ�Kĳ��w{�߻]��;~��%2�$�1���E��O&�������!���R�5鹤D�fY5����S�,Kľ���kiȖ%�b{��Z��bX�%������bX�'�}���X�%��v����&��ֳZ�ӑ,K��u��7ı,Kϻ�m9ı,Ov�eMı,K���[ND�,K�����I�.5�e�f�jn%�bX��w��r%�bX���ʛ�c�"_����r%�bX����jn%�bX�Ͻ}�kE�SFL�nkZ�r%�bX���ʛ�bX�%������bX�'������%�b^}�kiȖ%�bw��7tJ\55r�˗Z17ı,Kϻ�m9ı,O������%�b^}�kiȖ%�b};혛�bX�%Cȇ�"� �$X�{S?�����f��Ӷ�zt���Nv�B�Gm�<vPS�F*5��]9��8y˷-:w\@�Ap�l��D�ձ�����r�n��nc���[�Wg�v�)ũ�(�&'{���c.q���*[cZ��Om����6�N+o@�^������N�#XZ�U�i9���`�]�"rn�m�q���iO<n9�ܜ�vW��it��d{7[����&֜5�9.�)���e���MI2\!�5s��(s��M�RONtE�i}��cnI�=u�7/b��FnZ�RS������oq�ߟ�����X�%�ϻ�m9ı,O�}�q,Kļ���ӑ,K���_�5�Yi�ф�թ��%�bs���NC��L�bv{��Mı,K��~�ӑ,K����Z����2%��ƽ?hˬ�љ�-��ӑ,K���혛�bX�%������bX�'��z��Kı9�}ͧ"X�%�g���5ў*4�n}�7�������s�}�[ND�,K��~�7ı,N}�siȖ%��&D�����bY�7���p~�l���������d�>�֦�X�%�����m>�bX�'g�l��Kı/>ﵴ�K��{����w߃�1�P��u���qס�N�Ѣ�rj�i��NmV@g%Y����ֲ�Z�I�9�}��A9>�D$���7�,K��=jn%�bX�����]�M3D�f���bX�'Ӿى�p0�$T��P�M�'"X����m9ı,N�Y�Sq,Kļ���ӑ.��ow�߫���%ȕϻ��,K���[ND�,K��=jn%�bX��w��r%�bX�N�f&�X�%������5�5�u�Ku�m9ı,O������%�b^}�kiȖ%�b}��7ı,Kϻ�m9�q���}ߓ���I!�sؠ�|��%�b^}�kiȖ%�a��}p�Ȗ%�b_����r%�bX�wY�Sq,K��亮�\/.CZњ�k$�#vz�����bx7XI���|�׾qۇ�۷=%]:�,�љ�335�'�,K���7ı,Kϻ�m9ı,O������%�b^}�kiȖ%�bY���Vh�0�֋t\�7ı,Kϻ�m9ı,O������%�b^}�kiȖ%�b}��7�C*dK�ߥ?g,�u�W�w�{��7���ϳ�T�Kı/>ﵴ�K�҄:IƈQZ����)��8@*>�j� ^(O�2��MkZC�l�m�n��x���\6پ,a�mNRf �_y��#+��0"/���϶xE�t~�7�`��;¬I4PIJD <G��I�Po~X2�Є�Ay�G��S�<�(ٿ �9"Մ���BݟB$Pa�*�b��O"tND�;LÉ�S5������fSY�0>� ��oi���*��z#��@<�	�(+�T]�Q1@�/�z�b��	@N���;޻�Sq,Kľ���ӑ,x��{���v���]3���|��x��Q��3������bX�'}l���%�b^}�kiȖ%��&D﷟�Mı,K����F��L���Է5�m9ı,O�}���X�%��������,K�ﵟ�Mı,K���[ND�,K�{/�5)l�ԛ�鲋ى�`a�X����A�L9ۣNN��]��*i�<>��&k�w��7��,Kϻ�m9ı,N�Y�Sq,Kļ�����}"X�'_�*n%�w���{�jF��'pU�����{��'{�����%�b^}�kiȖ%�b}��7ı,Kϻ�m9������[�ow�~�?��I!�sصjn%�bX������"X�%��}�"n%�bX��w��r%�bX�wY�Sq,K��u'}tfk-�4fj���kiȖ%�b}�fț�bX�%������bX�'{�����%��X1H��!�K`$R�H�P+J$W�7�k�~�ӑ,K����MY�h�Z�r���q,Kļ���ӑ,K��E#�o?Z��bX�%�����"X�%����"n%�bX���P����%�)[Kj�n7KuͰ�i^N˳QG=]y���utL%�Mu�:�Y�������owY�Sq,Kļ���ӑ,K���͑7ı,Ng��m9ı,{��Ϸi����9�w��7���x����Ӑ���"dK���"n%�bX�������bX�'��z��O�/���{������]�N�������,K���"n%�bX��w��r%�bX�wY�Sq,Kļ���ӑ,K�ｙ�kD��L�2�kDMı,K���[ND�,K��=jn%�bX��w��r%�`~�.�{��|D�Kı?~��8]jܚ��e�M�ֶ��bX�'��z��Kı/>ﵴ�Kı>�dMı,K���[ND�,K�T��j"X ��n�~��s\FҐ(��`u�etcc8�==�m����(:�����t���-�'����v�Y��#��h��w]�<�_�_���!Ě�Kr��]y�m6d+=ѭ%on�dR;S�{���vrB�q�v�L�Z���{y�\竁�\=y�Խ���Ks�5Yk0c7�8�d��.��WA�"�9��vc)�%�m[�\"��,Mj�{������;60?�6`G�[%��[[�-�{u�`�ì^]vͫn3[��ݻjՙ��t�7;���7��,KϽ���"X�%����"n%�bX��w��r%�bX��֦�X�<ow��oϥ� �r�U������d�>��dM��#�2%�~�kiȖ%�b{��֦�X�%�y�}��"X�%�g|zj�F�[�33DMı,K���[ND�,K��z��K�A�Dȗ������bX�'~͛��{��7������M����KM[ND�,K��z��Kı/>ﵴ�Kı>��dMı,��3������bX�'���d�a���dֳZ�7ı,Kϻ�m9ı,O���q,Kļ���ӑ,K��u��7ı,Nzv_ˬ&j��e�m��N���D]4��n��'��,�ΐHե���VG����똀j���oq�������"n%�bX��w��r%�bX��֦�X�%�y�}��"X�%�����Wg�Ւ��v�|��{��7�������U|��ȸ�S����i�&D�9�g֦�X�%�{�~�ӑ,K���͑7ı,N��8]MfWW-�mֵ��Kı;�g�Mı,K���[ND�,K�{6D�Kı/>ﵴ�K�q��w����.:n{��oqļ���ӑ,K���͑7ı,Kϻ�m9ı,O������%��{��[~}.Y��2�|�7������͑7ı,?1ϻ���}ı,N�Y���Kı/>ﵴ�K������w}����$E�j�b�
m1��\�:K�\;p�ι��}lm��xSYz�dц�&d���'"X�%�~�kiȖ%�b}�g�Mı,K���[ND�,K��6D�Kı/�=g��5$��u��f���"X�%��u��7ı,Kϻ�m9ı,O���q,Kļ���ӑ,K�����,��ɚ�j��Kı/>ﵴ�Kı>�dMıN�D�#�"��EB�n&�^�|�ӑ,K�ﵞ�7ı,N|{g����h֮��ֵ��Kı>�dMı,K���[ND�,K��=jn%�bX��w��r%�bX���7�h�\55r��5�7ı,Kϻ�m9ı,? Ǿ�~�9ı,K�}�[ND�,K��6D�Kı/���c���ŸrL��I��nn�lv�Hܜ���Y��sև���N�n��-/��u�m9ı,O������%�b^}�kiȖ%�b}�fț�bX�%������bX�'�u��%�5�f�f�%֭Mı,K���[ND�,K��6D�Kı/>ﵴ�Kı>�֦�eL�b~����3Yn����ֶ��bX�'}�6D�Kı/>ﵴ�Kı>�֦�X�%�y�}��"X�%�a�ոa�jL�33DMı,K���[ND�,K��=jn%�bX��w��r%�`A�S@TH 2��o�\�;�gH��bX�%�N��n�I)�[�ֵ�kiȖ%�b}�g�Mı,K�S���kiؖ%�b{��l���%�b^}�kiȖ%�`���ɻu����6ڬl�B�HN<z��r�=��j��㨖�\�h�y��j���{��7����[ND�,K��6D�Kı/>ﵴ�Kı;�g�Mı,K���jk$̦�j�-�k[ND�,K�{6D�Kı/>ﵴ�Kı;��eMı,K���[ND��2{�����>TvxzЗ&������d�/���m9ı,N�s�Sq,�"_����r%�bX���6D�Kı;�x�u5�a�2�d-ֵ��Kı;��eMı,K���[ND�,K�{6D�K��#2&}�~�������ow��8�q:�]78)<n%�bX��w��r%�bX1����'"X�%�~�kiȖ%�bw;�ʛ�bX�'�CPQM��ڷVkS声�^9�{5�k��pl2�#9y�9���5��z��3Wv�v9RY��۔�٨��j筘�M����z�
���.����Wu�\uq���=L.wm�sv;n.��R8wo*\��5��J-5�d��#Ebu����魤�iʉ�ST��hN��M�5��l�9d�����N������\\@? � �]��t9����\��c݆�nK2灶�i�������1g�q��6lg��)�r�g��2�}�w�ı,N��l���%�b^}�kiȖ%�bw;���NDȖ%�~�kiȖ%�bX{��kF\��h���%�b^}�kiȖ%�bw;�ʛ�bX�%������bX�'��o������w�����~�����U�m9ı,Og��T�Kı/>ﵴ�K�AHdL��߳dMı,K��~�ӑ,K�����-�f����kZʛ�bX�%������bX�'��l���%�b^}�kiȖ%�bw;�ʛ�bX�'>=�٢虔ѭ]e��kiȖ%�b}�fț�bX��ϻ���}ı,Og��T�Kı/>ﵴ�Kı,'�%�������X�#]�kFm�qƋ���3�5�E�n�xzЗ&������D�/>ﵴ�Kı;��eMı,K���[�DȖ%��߳dMı,K�����k2�4e�M�ֶ��bX�'s�쩸!�!��@ �D� �H��Z�@  �+1�5Ĺ�}��"X�%��{6D�Kı/>ﵴ�Kı=;���.�ֲ��-ֲ��X�%�y�}��"X�%����"n%����/���m9ı,Og��T�Kı=�I�h��՘f���33Z�r%�bX�{ٲ&�X�%�y��[ND�,K���T�Kı/;�kiȖ%�bXw�z�0ц�e�.f���bX�%�{�m9ı,N�s�Sq,Kļ�}��"X�%����"n%�bX���#�h�����]^�2�B��e�m�h�A�Ө�Q��6!��X�����ϭ�I/����<X�%�}�����bX�%�{�m9ı,O���q,K��w�ͧ#���ow�<~o��3��AU�ŉbX��ﵴ�Kı>��dMı,K���6��bX�%�}�D�Kı9��=�WD�M��[�ֶ��bX�'��l���%�bs;�fӑ,|�k��J�)�L5蟳��D�Kı/������bX�'��ѩ0�jj��5�7ı,Ng{��r%�bX���Yq,Kļ�}��"X��"w���q,K����p����f���Y��r%�bX���Yq,Kļ�}��"X�%����"n%�bX���ٴ�KǍ�>�ߦ�b�Nv����9.ݭ��b�����nB�عU㫵����q��h�h�nk"r%�bX��{����bX�'��l���%�bs;�fӑ,K��w�ț�bX�'��;�����sRffk[ND�,K�{6D�?�c�2%��{߳iȖ%�b{=����X�%�y��[ND�,Kþ3�a��5�.Ys4D�Kı9��iȖ%�bw;�ʛ�c�U�Dȗ�{����bX�'~͑7ı,K��Y�n�ɭ[��f��ND�,���5��g�T�Kı/~��ӑ,K���͑7İ(�� �O��<�Ok���ND�,K��g�����������oq��}��"X�%�������%�bs;�fӑ,K��w=�7ı,O���p]v����umڼn�G`9�y5���ۦ�lں[�ɷWE�N�����Kı>��q7ı,Ng{��r%�bX��粇�D�Q�D�KĽ���[ND�,K����4jL�jj拄ֵq,K��}�fӐ�@�DȖ'���*n%�bX�������bX�'��n&�~ʙ����p����f���Z�ӑ,K��{��&�X�%�y�}��"X�%�������%�b^}�kiȖ%�bzwF_�S5rh�h�nk"n%�g�02&}�~�ӑ,K���ٸ��bX�'3��6��bX�"{^�����%�b~����r,�7-��|�7���{������&�X�%��+\����� �'�D�A&��u�$D�Q_�Q_�AQ_�QZ�����"*+������Q_��Ƞ�B
AP"��Q@�PP �E��@�"AP*E `�$Q@�E b"EQX�*�����DTW�"*+QQ^�����"��򈊊��"*+������"��숊�������b��L��Q-E�<�� � ���fO� ���                      ��$(   �
 @  ��
J
Q  (�!ETJ    P(@T���  �    �E N��N[���<G�`���������d�e��k���P8� �AAc)��@ F�
b0 ���J0 �r�@� � �
 Ҁ14  �(     � (�)J14A��� i�4Xt�� ͂��6JY�}q�N� 8�����]�Z� [ם�K�.��>��/��+ͯy��{��y�����>U�t.,��ۭ���cռ >�(     �J�����  41  � �k�7��� ==�mnn�m9��w{�ż��� �y�9��qe�׋yon�ޱ� w�{w��g���\�;�y�:� �-�7mŗ����7�����|�@(    ( 2 �U�ݗ�6��˼۶�.ꗞ yKܻ��{���3���3��v���3���� ���m\�.�� >�J�uu��UӖ�}�;/k� ]�k�Ӷ�[�ux��\��mx� � 

 d� �ﵦ���w]��p�>���zO��Û�yO/v��ŗ�q5/p �r�9�;�/&�  ��[�y����^� ���nO/K�{������l���y+����v�w��yz{/ ��J��T�T�F���6��)P  "��U*UL��b'�T�i�� ���)����   DSD�JE��N�x�����g�9�_��'�=�׳��g�EE|/���������ATTW������QQX"������P���5��h�i��!� ��&&������'~)t0p�SD+,������]�F`GB�����{��F�k���N�5:sFؐa#L,����
=�T�M1�}�7�|ƚ"@����
�0(�bсJF��š��iR���SX|��m	�"��������O����|4`P�$���
�"�p�Ct�
0*đk���o�]|o�^4ֳa�#�� 0�] B�0)��6}�u����s�����ٹ�t����Z��@Ƈ�"D��0	CJa�0�	bk4m�@�
��c����F�u&[����`�f�֫D�ſt��e7�@�XE"�t1&B��0�@���`�b�(��SG &�d�t��r֑Z1�ā]!�
�0i��~5߷��D��z' 0H�,R&�8#�H4tq,��(�X����d B1��Pb���#MSi@�R�)��4Ӆv1������>�_�$��2n[~w�P��91��l�4ٜ�r��ƈiH� VD�i��H��˛f���Ԁ�!�H�T���a#@�`I)]8oc+�lv��#KB�4����N!��H,p~6|�)   �P�@Е8�ĀS\�t��p!LS%R)P�`ˆsf���_h���:C�-
�~B	T#Xi���CK����Y|sYf��B|��7�ɽ���G)F��>!]I�ۮq'-	!vFJ�&��uLxk5��N�������#��M�P�n�,�TڼW���� P�c���qv5�J�b��HA��쓖酲�h������c�hX���#���F�P�Wbc��#$ @Ɔ(h(`����E�ˬ�ȕ��^F��p�/X�0�Cz�'# B�i
�>ь��.��Sf�"`�+�06�i1M��I�b�1$�цm6B�����C���7��77���B���o2k���g��!
0+�C�,h��cP"##!$X���J��t�R^���xb0cCK�t��ƤM:�N��l��
�&>�uXҮ�C���#u�>�Q���� <�����p�ҝP�F�J�T�bbtx}�ā�:A���GF��4)a�0a�����!D�+]HH@)��F���uv:H�Yk��P�!M\6b�pI%I��Ʌ�c�B¬B��q�ƺV�jI��I��) ���b�rM�X�H����������h�!�8t��H���l$w|B�fI��L:�4j6@�H�FF��۷d1����3[H�h�N'���c��Ia���[�y��9L1Iuu~ɼ�H�_o�g9�R��`��<���x	���0��>�Ǉ��lٲ5 �R�@��F�J}��F]�d%��ٽf����Fs{�q��#Rx� ���.� Co ѱ�Mf���������[�]V��_sGЇ�
�Zi�t�S�.����H]`����X�5�P�bAHƑ����H`l�0"�  �
�+D��F����@ A�*F�d��&M�P�:N5�ti��:&�2SHIip���+�#Y���oF�CA��֓|>z��ُ�F���p��u�&އ��~tSQ'�Ʃ���	�8aM��
�mĠE��������Fd�Β�$g��čt�;8��P��c]8K�y;�l"¡�jhB�	��	�kdH0��s��%ц�<B�ʒ�k����M0Jh.��M���1 b�P�@��lJhЁ>~�gĒ��]x�Y�	M,�'�!~8����C���б�F� ��`���*®!� ���E�ia��>v�m1�CdJ��{�n�v�Ё]nfG�\���+½Vé�� PцȜ��Q&�6�k�P�CN$���$��X�hh�6�$x�y�i��u�E,R� �@���1��H���+�CA�%t��J�L�)M��b�$��r]��5��"n���޶��0�$��xˬ�z�l��� �v<����&�(čHFe �b���#���$+�ٔ8��R�!�4�hB���$��J@����A
���V���YB��6I$*j��Tt��(� h1X,@�5�H#6D#�"�z0���t�>�>���j�$�4t�0NĴ3-���&���i�2k�|f���A���5ћy�}aHӉ�i��Fo
w�<!�>d��H��D
��Z�F8F1�X�cF@bSf.��SQ��8�C{)!!��Md�"l�5�l�F�� U�!5�s�Q�6L���y���\�4R	�ڸ��K:��r��_��)h:p�gh@�0ٱᄏ�]8F�����º�1J�pͤ)�	�j5�C�"4`F ]��䌺.S��}"��

�6}��`p��%�CG�I�
�:p1�A U�@�@���<#�w9t@����u�1����J�V @qBCg�W�P�rҲ���B%4� ,�� c�'���FJƔF Q�ƌD�$��D�*�jF�En��C��0�Q! �D'����D ��Rd ��"	,���7�� ЋSdj�]Ed#"����,!����yx��@�ѩ:f��2���!+���#�F7f�isykR��ai�fЉCK�\�)�vF8x!Ml#YS8oٹ�4��#�%$�}���2�Z�s{������)��U�L#͛��!u����#(Mѻ�[���"�٢�ā"]d5˚8l�ٲ��7t`H�s7�w�m&��4�XR_�Xr� �޺}(h�u�a�� 0_��2��j���c���ԇɴ��6J�!�8謖e �Q�"8#@41aH���	�,��D�p�� 9���� 1�%�c�D��)���Ы"� �x;�qb�4#	���d�	���U��3h��,�4K�]a��H��5�Ást����q75��ߞ�����8 qG�°�A����`qi�+
:(lx, ����cc�|y��MJ�)�iͰdhF'�M8 @hs�M�}�>~�(J"Y��6kXj��A^���~���`��]!s�}����|
�iu��kWAg}�.�Zt�1#�,���xH	
�{��1x@��)A󏃢5а+,
�ƞ����@�H�	�ƃ�:WJh0w�$�T��t�۸Bv蔗줴�#t�R4���`(@bH���E���D�a0����arn��p��.�l:7�`R!"Bt������K}�ߣ��  �R�� �� $  �`�  � [Cm��  ����x @�m6� p���V�UUIj��V���H[Cmj�[-�mt� 6�  	,%� �kh�  [@$�Bڶ� ��8/F���ڶ -��)ԩ��c��՚��m� @ �SE �9b��(L]��P�C����v�v%{@<�դ;�}m���Y��9�R�ʶ��K�\���
eLi�)��QR�0;�`�8�]6�� ]�Ia�  m��-���i0   8�  ,�� 5����6�cm&۶ΐ$��m�m&ăZҸ�0�Z���;2��19BBuU@Um*�0���e6�h�v:������ m��@�@-����v �RkR` 8%K��h86�	�� $�I�]��U����|��v V��5�\ #n� ��$� �$��m� ���ͮ�g5�0 � ���@R�UU.�R�*�� ��6�H  9m�����%���׭H�I#Esm�����	f�-�U�� m��i� �v  ���m��b��y�@  �t��4�D��  K(�l�[pڶ�t�  �aqÿ'����[@ 8 �m���a�A���p�  q�'�0��[@�/��� m��	� Б�m�$ �mm�ݰ9m� I��$[vؓm�� ���  	 hŴm�     &��mm�`t�D����$ ���A�l-�e���AŲW  �d�[%�Q�출p��t�����@?��H   �����eɭ�[V���6�m�m����� m�   hl�қkin����۶��d�-� 6�z���BI�  	�lM�$��5U�)ԫU �VҠcmUUPR����lؐ�� ��m��i p    �Ҁ�`�m�-� 5��H  [[m�l��B�t�E6�E�Y �Jm%��%��d��n���Hp8m� m��\�!�k����l��i0�6�u�ſ�� i��` ��n��H������p�C:i
�5�	�)����sm6�l �-�ڶ�  �` ��$g@  $� ��   @��R�Y@�h   ����� -��am[@$Hp[%$6�	�sm� m�s��k�I��Ӗյ���3 ����{����d������V ��J�J�+��4@�9��u�z��d�iwKϖԄS�-v`0�s��Q!�   nܽ��:Cm�E�Nm��Г��RgӜ[@ �ٵ�Kf;m�� �'G�h��Ku�'`� �I$m�N��L��l�M� $>H�l��K��J6��v H   8ᴛ6�� 8 s�e���Hp���LK(��I�$6���l��v����6�A��[sm�m��` ���`]� �mp� x<  �$��,0���2�! �	eBA m�π	۲mE�[T��m� k�6�7n�pi����鷻ӠI� -�ʱp[N'BKl۹���-� [M��� 7m�� �ȱ"�56���� [��M��޺M�By�I�l��  �X6�	m��n�-�I�F�d��e�5��jj�6��Fvk,�ݮ	 �@� Ӷ� 7$R�R�6P�j*�zH���a���[k(t�t�gYO�Nkɜ�P�y�2�0��T�n���@�I-UK�e����[*�mJ�N��pf��2 U{��T�G��v�4�zL�̻-<�m�9�mU[l�ppj��mm�m����� ����6�դ[���2`2�,2G�x���e��kH϶�]\�N�4.Yp�0���0 m��if
-�l$��� 6�t��}�vY�����rA���Cm��mÒ��lj�U�hZ�X��5����mu�[���) ܄����k���ΖݻkvZ��m�p �6ض��I�m͵�6%[kkݺ�X �8��f��m�� �j��T�AVyj��� �[K:ȶ� 6�.�`H� ۝< *�Uҭ�Uդⓛl�<����[pj�8  -��sm�   $H 8  H[CE۴���e��m�\.����-Ԩu]T�=@W*ރ  pH�hk[l�	�skz��q  �8�k��-��Ӷ ��[O��5֕����m�   p̈��-[��� �NJ5�K�v�K(�m��������ɪ����*C�YxbBK�rYg@�nKd���-P9��H�F�%�6�O���n%��)25K��9iIj����n�`�� րh$�h� �� H�mmŴ�iH �i\��m[�� 8V��s�ж��� H$m�88����~{�y�m�� 8�e�9�����'�ݒ�   �z� @m�m�H��` ==�{�9��4P �   $� m-�m� ��$�������  �-�9�8�lZl�ͤ$��t�   ��m��C]z묷D�[xz�Jං�v���m�E�pW]]@UYI��oPti�mmv�1�����{���M�i!���h���.�	9@iV�<*�U]+�*�6�۴�n;IEx��ĺL>&�Xݻ=�����UP��ml�ܢ6� [! t�K��]�5uUAH�^j�݊�e����7��7nݰ�GTʵ]@ GXXk�l� �    �΂@�n�;m#�ڝ�n�� ��` :�U8��k��g,V��g6���B۷lm�s�q������{޶��&ٍ��޹��6%YV��� ���F�f�`[�̽Z} ��P*�%^�U�� n��m$ � kX ���mUV�9��K-V��ҭ�+��q��V6�*ƅ����S}��m�s��f�H6� -4�`  U����j��j�$�]"Q"YVж�m�6�� mp���   [BG-6 ��5�6l� �D�� 	  hh  H�7�[�  	     �l$@ sj�� ��[p�fܴ����6݀  �` �   h � -���� ��    �ۊR�*�J�WU*g��F�ޠ8�  �<  $��� �`� H    8 m n�	\�-�	  ��l       ��[�� �@�� [F�ۃ�m ����Cn�͸ ��� $�AƊ��Kh  � $ l6Z��`v�@6�m� 	 m���A�V6[a��l�sm�[h�     I�p� �lᴛ�  ����i����J-$8l�m��I���m��kX��@�I  �[��    �iխ��miW-�5���k�� ���l�k�[�NHlm����0�]-,�,�n��P�^���l m��n��l��mn��6��   H6[�6�jU��
Z�
U	    6زu����`m�$kuIv��ml@m�fF�5�l0 h  �  @�[D�5��h��@U+;-T*Ҩqm  -� 5����	������ӎ�mY�  ��[@[���[R 6��mz�m[@�-�  d�`�h��I��6�6m�koc��@ 6�Ͷmv� m�tK%�\����6R���)UJ�J�uJ�N�m���[́�` ٶ�� �#��m� 4턄��V۰6�].  mm  �I���79�ڪ�հ�L�r�M~���Ai&�h� m���$N��� m cZm&˒���  �o�[F�9QʁUUT�̇ �V�R�neН�U�h�U�mGJم���6�b��� c7���*��R��imR��p�vm��U/=+@W b��@P"�am��5�n��n8�hN�� �K�f��j�
�m��pm���8HR��UU[OK6պ !�mm 	6UP�rԫ/����;���   �m����  �m�M�"Cm�6ͳ��� -�kz����;���PT�/� "�X�W�/��mp�zQ<+��`)"��x�������X�/�:*'��D:���
;TY��F�> ��6'||<�*|��`�=�@�PШ��Q�D(�l6���6� qE*�|�� �6���� �E`�AH�<��>D8@]E!,�Pv�&��B �RET|�Tpi*�T>�� �H��A����"����G>p�c �@	�|(���H|ET�ȣ�Nx6|�o�!�U�>���xR(�< ���t�D��@�T(��F���@ �A�"�  ������ ���q
S��$D�T�4�	τB�Th&��hx
���":>CB*& �� �X
� Q �C�N���� !�� ��S�¨������PH %¤�*)o���r7�Iwv�]P9����Cv���T�T��hQ��t�d;h�6�I�L[:�흋\qZBӺ��U�OW۵���d䮡�ınM�jx��u�r��X��`��.i��L5v�eG��痌k��j��i]��{eWkkv��y uk&�Iem���V����,�dh67H�[;�S.���A9U�S�V�`�5pV��C(4J��]D;C�-����MO0se'�e�U��FG��B�v���8v3�lm��ǯM��$M�mp��c�8j����p,���#�7"��s��.:��.�n�9�4-dV�U��(�X��e��S�i6Q�րFV�N���e�W���4���9` i��Դ����v�֦�
!7�ڀw]:�4��x��]��0v�j:�m������xc8�rg�H#mt<$L۔�M#��u��l솮�E����=��H��Ψ����&��\@sx��V�
��Ʃ�nL[.�[#�p{ce�[����2���ԑ>����y��VK��5����1�;Q�SՄ�L̑�oh
ۥs �Ψj���ܑJ�¦�$�6�;dr ���ˌ�7�V��{]a��äŉD���kV�wIÒ�v+2�����^�i3�$7J��{7f�%�*�.�c�p�z^6	|akd�Mά�a	���:�D�䄎pH�B�l̙F 
�j�ܕ�]V)��0Rյ T��T��l�*�i����+�å�Cj�F�hj���6��Hgki��rމCG6���\ݪ��6n]���A�ש����m��ɨә��;��m�@U��R�ю���F\�H��Nb�j��=35ʵ&���Z��v�(*�sE��L�Km��k;�H܅�nC��ٱU��}�J7l�����o9֩�Jl�s�]�MN�i��븕V51�u��V��jf���(�ʣC-!"0`�@S`G QDУ�� ���~��me���c�����N'Vd��Dͷgqi����^9��;���m:�i�w&�+��p=�P-a��O;���΄`�P�����r���Ǔ���[�����JН�p:��4�r� ۓg�E�x6�m�H�vԳq�u�6��v W�[�`<��e���.��P������ݐ^{c�&�e�� AqD6 `���ٕ��#T��o=�v��C�=��ʼ&�������W��/G�w*��ـ?�������%IU0�_����L���$kQ�&��}V�K�B�8�]&�0&Mi�^IL���@�72'��Š�f��빠�f��}V�m�;���Ɯ��=UL��0�)���N�K�.�@��TY'��mD9�4�l�>���u�@�u��R��$cɏqʱn�x�5�O[�썽dxsE��rog�e2���<X)�<qE����$�@���@/$�^F������� Q\�u3Y�\˹$���o�hX �T`�X�P ! U| �PC�;D�*%�{lܒ}��7$���@�{�&�I�H�M��&��빠�f��}V�{��ع�IH�S���f��}V�{��{���|��#x�#@(ӓ@���`	.^IL��0�)�w�����-�:�t3qSK7&���si:L��v�%��:�����C�[s��yy�>��S/#L�J`}=��	�W�<&�s1H�$�;�w4�l�>���u�L�߀��ʲLb�QE$7$�｛�s���F	�1@����F�
�Ul	@X�P*��'u�f���ٹ%�wx�1cr6�qI4���٠w��hu�@�T(B~I��#qh��@�u���f��}V��O�ޏ��N��Վ�6�L�A����dn���%�Om�^x��s�c	2ϻݱ<%��IDؚr|��s@;���ڴ�٠}�����JDژ"9��l�>�ՠ������|��yH�
ɠ}]�@=m�~����s@;��׮j�1��E1�q8���`fdi�fIL3~\p�I��\�Ъ�v��!��Y�@���;�����LR!�4�%0>������sqG��.�؃���s3�%�5�޶�c�9����m�L�ذ��w=���'��55�m��ݦ��u�\��.s��Z`L��8�n)&��v� ��h�l�.V�P����H�]`$�^F�d���{'Xv�ӷ�ErF����ҭ�������}_U������ڭ
�0�;� =�ـrI}�y� {���훒uh��FH�.�)(a 0�5+ g���R̺�ֵ�#�v���-tȜ��C�˩�\�6���`bd�sZ�m�L���u!q[�Jm�ck=6䂶�j�۩]=m������9���v��w;��{��!M�q�xun4)[K
v�"��mI�Y;ęy�Y�-l����1;t������u�h���t��Ft;��"K@2�ur�d�9�6�/k�W[|i�w��}ޱ�7����i$�b�5���Y�3�%w&Ɯ��x��m<<�a
)zz������n��\��yiq fIL����1�������[f��빠������,w�m��L��h�w4�٠}]�@=m��W�d��6��H�� �hWj�[f������h�P�a�8Ĕ�M��Z�l�;��hu�@�������@��DK#M�� �qq]�ÍՖ�uxko<�즩#	���y^ԎI"�[f���s@;���ڴ�����1���4��;��m�?�"�Db/�D���R�i,��W����oX�)��A�s�����26���hu�@��V�z�4y�VG��C�������okw�7v��`�S� �q
�܃�ڸ�< �wf�T��[��� 7{��������-Q�6»�7^�X�wnG��[�����h��ܩ;X�'�<Q��M��%2(8��;��h����Zm�@=���Qch��"��ٜ�UM�u�< ��w]��G���q�$��hW}w$������O��P� ?�)b�K��3 wwLW��hBUݢH�- �٠w��h�������Dҹ�%b�@�u��m���Zm�@��h��D�v��9�\��)�gս��:Ny�4^w/vģ�J�e�B��E.�"X�, �ݘ��Zm�@�u��/�J��Py �9n��?��� =��>L��L��?l���%�b^��ͧ"~PCU5�^��;�Wn�N��q�XRe&Qb_~��6��bX�'{}���X�%�{�{6��bX�'��z��K�2��L�Pwwwp�[�&R�)2�9@M -	�߸i7ı,K�߿fӑ,K��ٯZ��bX+#@|�k"{^��"X�%�g���i�L��f��fMı,K���m9ı,?G���֧"X�%�����6��bX�'g}�I��%�w�����wߝs���:�Ļ�����;s����]�+�:F5q�͗a{rH/g���2E�Y��ND�,K�f�jn%�bX����iȖ%�bvw�4��bX�%����r%�bX�=�RzL��Z&e���Z��bX�'��p�r��bX����&�X�%�}�{6��bX�'��z��Kı9��n�_u���֤��6��bX�'{}���X�%�}�{6��bX�'��z��Kı;�{�ӑ,K��]��WY�Lњ�f���Mı,K���m9ı,O������%�b{���"X�T�'{}���X�%�߳��3Y��Fd1���ͧ"X�%���^�7ı,O{���Kı;��7ı,K�{ٴ�Kı?"w5���8��pD�0�����g�0�6�q�V�-�mY5�cXc��ݰ���1u!֔1t���t�O�W[�F��)m�����]�\@nR�nwa�nrK�؝����h�n0k\��m!1V[����f�ǡ+y��EnҸd9u����An��vb��ѐkCjȼ܃���	�2�{\NX���g�n;����V�ٙ�"RnCe�َ���]��z����;=sp�2s�j�Ҏ[d�%��o�6N3����7E��0{�7���%��w��8m9ı,N��eMı,K���m9ı,O������%��K}�^�;���q�wR�)2���}��7ı,K�{ٴ�Kı>�k֦�X�%��{�6��T�%�g�ץ4�L��f̹�T�Kı/��fӑ,K��ٯZ��c�	D�O߿~��Kı=��eL)2�)2����{#B�r���&QȖ%�b}�׭Mı,K���m9ı,N���q,Kľ���ND�,KǳZ'�Ɏ��f\��e���%�b{���"X�%���["n%�bX����iȖ%�b}�׭L)2�)2����k�˅��2�[�D����3��ؚ�aj��b���m;�Ѳlv�w���^.�cB��߭�7���{����7ı,K�{ٴ�Kı>�kև�g"j%�b~����"X�%����o�VLu%�N�w��oq��K�{ٴ�6<�DȖ'��z��Kı>����Kı;��0��L��[���[��)�w&R��bX�'��z��Kı;�{�ӑ,`$,K���Sq,KĽ���ND�,K�_M�aj��kF��-Mı,K���m9ı,N��eMı,K���m9ı,O����aI��I���eꃻ���.�6��bX�'{}���X�%��P�߿~ͧ�,K�����Sq,K���ND�,K�(���~6S6��#]�Ɍ��If���
�[�|t�pIygm՛����4��գ��4Uǻ���KĿ�~��ND�,K�f�jn%�bX����a��bX�'{}���I��K��Zw�4+�,m�$�9ı,O������%�b{���"X�%���l���%�b_{�ͧ"X�%��٭�d�Z�3.���Sq,K����ND�,K���D�K�6�����b����X�!�� Pp�6�"���A�(h�Ŕ�H�	�"I&�Ə��+:���4+�(WK
Ƭ5��u�0��H�@��T�����6>K Х� �B_�O��?H�Y ���~����	���A
+���	D � �����pޕ^u�TM( i@OhG�: ��AG�(uڪhҾz�����H�
Dh�C"z%�ﻛ�*>���%��ٯ֦�qRJ�Ҳ�)}~|���ˌ��EȲ�D�,�Q j'��\"n%�bX�߿~ͧ�O�j%�bw�k����qF�Bj'�~��iȖ%�bw^��ֵ���rᆿ"e���,Kľ���m9��Q5�����Sq,x!D�O~���ӑ,K���kd?D�K��Ǧ��Ն��KJ]I�.h�]R�\��ԄeD7��hy��q���R
'TUId̆7&����=P��j%��������%�a�H�������%�b{ߵ�&�Y��j%�����r%�c�VR�u���+�qA�j��,)2��b~����!�D��j%��~�ț�c���j%�����r%�bX����i�cȟ˕5����o_�K�kZ�.5���iȖ%� j'����q,KÊ���߿f��%�bw�k����~ j&�~����"X�%�go�i̙Mj�����7�'"X�%�~��6���H�&�X����jn%�bY� ~������%�P�`�4�B
D4�P���TO�4�>�����q?�T�K���E��hW-�仙K���L��^��Mı,K
�}�{�I�}� �	"w��&��	ϻs&k3Z�i�΄:�"$��ɠ�����#��g�4	T��ι��'��
����{P���{��7���{�6��bX�'{�l���%�b{��6��bX�'��z��Kı9�����]f�̺�&��"X�%���["n%�bX���ͧ"X�%���^�7ı,O{���Kı>W�iwr��q����XRe&Re/{��ӑ,K��ٯZ��bX�'��p�r%�bX�ﵲ&�X�%�ｻ���\�3!�-�m9ı,O������%�b{���"X�%���["n%�bX���ͧ"X�%������+�qA�j��,)2�)2�����Kı;�kdMı,K�����Kı>�k֦�X�%���~|a�H�o"gq���mx�� ���n�N�x\TYJ{r�G�2.��l��[��c]R��ʑ�r����-�NL��6Iq���e��4W��c��c�=�ݟ�Ş�v{,�:{v�c�m��#z�W�Q�i�gٚ�<������c�2����j�ތ��OU���.�Kr�P$��6�\�M�;�^�g5�HMq��8�\z{n���2�ێ�绻��䭾��1U�����s�Ԗ^�v��1�\������u�f��u�V1t4W}���q������s����%�b^��ͧ"X�%���jn%�bX����iȖ%�bY��W2e5��[��Sq,KĽ���ND�,K��z��Kı;�{�ӑ,K���=*n%�bX��wE�u��CY���336��bX�'{�����%�bw���"X�%���zT�Kı/}�fӑ,K��l�F�%]�$ww#t���L��^�{�ӑ,K���=*n%�bX����iȖ%�bw��Z��bX�'5�ۻF��\dw`\�)�I��K��Sq,KĽ���ND�,K��z��Kı;�{�ӑ,K���s�.�5�Gh�yqZ�v��d����gm=Kd5Ӯ�'����J����tE�%̕7ı,K�{ٴ�Kı/{�eMı,K���l?�}Q,S){��t���L��[�ƺH��Q�5�ͧ"X�%�{�{*n��2"�@k�2%��߿p�r%�bX�~�~�7ı,K�{ٴ�OΪjRe.��|�v�(8�XK��)1,O~���ӑ,K��ٯZ��c�!���}����r%�bX���쩸�Re&R����wwq�(�G"�_�&%�b}�׭Mı,K���m9ı,K���Sq,K���ND�,K��G��L��\��ne���%�b^��ͧ"X�%�{�{*n%�bX����iȖ%�b}�׭MıL��\�U.�:�Y,��a�	�c�����"֢�wNLᵧ����)�v7i�����fR�\-�����%�bX���쩸�%�bw���"X�%���^�7ı,K�{ٴ�Kİ~=��<L��Z&e��fT�Kı/}�fӑ,K��ٯZ��bX�%���r%�bX��ײ��X�%�y��֋�.�Yf]j[u���Kı>�k֦�X�%�{�{6��cEb� x�q7�/;�eMı,K���m9ı,O�v���kRS.\0��e���%�b^��ͧ"X�%�{�{*n%�bX����iȖ%�b}�׭Mı,K�d=�fe���Z��r%�bX��ײ��X�%�{�{6��bX�'��z��Kı/}�fӑ,K��,񞐥?fLɒMjkB��k���噻p��I<���{�]�'�ZɅ�܂Z��w �v�%���I��I�wfӑ,K��ٯZ��bX�%���r%�bX��ײ��X�%���n�F���c�;$�2��I��I���{jn%�bX����iȖ%�b^�^ʛ�bX�%���r%�bX�w�<�2e֩3S-��Sq,KĽ���ND�,K���T�Kı/}�fӑ,K��ٯZ��bX�'���/�3D5��[s33iȖ%�bw��*n%�bX����iȖ%�b}�׭Mı,b�r&w��6��bX�ǳZ'��kF\��k
��bX�%���r%�bX�{5�Sq,KĽ���ND�,K���Sq,K7��߼1����2�h8�5V;v|ی�Q���#��<Wc�1�DifM���h֥�Y�ND�,K�\����%�b^��ͧ"X�%���l���%�b^��ͧ"X�%���{Y�Ԛ2��[�*n%�bX����iȖ%�bw��*n%�bX����iȖ%�b}랕7ı,N����噖�nMk3iȖ%�bw��*n%�bX����iȖ%�b}랕7ı,K�{ٴ�Kı=�rh�5���\�4f�
��bX�'}�p�r%�bX�z�Mı,K���m9ı,Oy�'K
L��L��i�����Q�e�6��bX�'޹�Sq,KĽ���ND�,K���Sq,K���ND�,K��찞˚�,�2\Q�k���ԏe����G9�oBk���-�dù��'k��a�3�K@�}Weѳ5���v[�]���U1��8l�nټ�=�wv���sчv��խ�}��J� 봽�Qn�6��P�c�:�h�Xl�O �;�%�6}�Ŵ��ZMV��W�b�"��l\���� J�J��(� hΝc=c=��6WY�O[���w������<�l��8�/]�.���82�6��O6�&@�X
�z�)�52�k%O�X�%�}��m9ı,N��eMı,K���l?�}QI���p�aI��I���,-$��\�����r%�bX���ʛ���&�X�����"X�%��~�ț�bX�%���r%�bX��٭�ˎ��f]k5�Mı,K���m9ı,N���q,KĽ���ND�,K�_l���%�b^}=��=��3,˭I5�m9ı,N���q,KĽ���ND�,K�_l���%�b^��ͧ"X�%���_f]I�.\0�ְ���%�b^��ͧ"X�%����T�Kı;�{�ӑ,K��}��7ı,O{ۅ�������z*���;1dsV�����;&V[y�dx��#Z�Z�����{��>��ʛ�bX�'}�p�r%�bX�ﵲ&�X�%�{�{6��bX�'}nM&�u��F��aSq,K���NC8F�@i@�|� �t��'���D�Kı/>�iȖ%�b}��7Ĳ�){�eꃻ���vIre/�)1,N���q,KĽ���ND��5Q;���Sq,Kľ���m9ı,K;{<�2e��[�fkY�Mı,K���m9ı,O�}���X�%��{�6��bX�A&�{ߵ�R)2�)wnXZ:Ih�]�2I���Kı>��ʛ�bX�'}�p�r%�bX�ﵲ&�X�%�{�{6��bX�;=�^2ɦ�f��sZ���n*��\A���f9������J۞^MNK�a�E�e�Z�3.��¦�X�%��{�6��bX�'{�l���%�b^��ͧ"X�%����T�Kı/>�հ�9$�;�.E���L��L��m�p�uQ,K�߿fӑ,K����eMı,K���m9ı,O�v�{YrJeˆZ�7ı,K�{ٴ�Kı>��J��c�8����4n&�g��ND�,K���R)2�){�X���+��ͧ"X�%����T�Kı;�{�ӑ,K��}��7ı,K�{ٴ�Kı;�rh�55��]]3Y�Mı,K���m9ı,N���q,KĽ���ND�,K�_l���%�b}�I^�2ےJf�L����kn��k�*�sma،*��a�0I�Bi�«�+��~����{���?5�&�X�%�{�{6��bX�'޹�Sq,K���ND�,K����L��2��u�Mı,K���m9ı,O�sҦ�X�%��{�6��bX�'{�l���%�b{ݸ�F�-K��rI2��I��I��מ�7ı,N����Kı;�kdMı,K���m9ı,OI�Zz��]�!.���)2�){w=6��bX�'{�l���%�b^��ͧ"X�h�"_��46�P�XV2RB` �E�X!�H0�!	(A�"Ί~Q�D֮~�7ı,K�Ӻ���.ff�]jI��iȖ%�bw��ț�bX�%���r%�bX�z�Mı,K���6��bX�'}}���tSb4.ܬv��9(�9�m�Q�u+�r��&9x�brܠrű�\+v�}��KĽ���ND�,K�\����%�bw�ߦ��>���%��~��K
L��L���a�FB;����L�Ȗ%�b}랕7ʋD�K�~��iȖ%�b{ߵ�&�X�%�~�}�ND�,K��&�ֵ���ѣ5��7ı,Nw���Kı>��J��c���Dȗ߿fӑ,K�]�~,)2�)2���^�;��#�����ND�,K�\����%�b_��fӑ,K��nzT�K��Q>���ND�,K�{��\ɔ֌��k2T�Kı/��iȖ%�a�#�]��9ı,O����"X�%���zT�Kı"t����1D��)
/w�}@�1���4�,�5��0>G��0-N�A?l��꟩�' �4��((�.�[W�ő� 6��tie�� �c��b�Y��m�]u���a w�9͵O�1#��3I/�`2D�tђ|!A#���J���jD��b��a#�����H�q~Vx��Hc>�i�Z��S:Cy�ֵK���AL�ЁU��D�h�9�?,P��o�c�"2��"�	��)�	�|��P�>�a�#!�1�I
%P��$������]ܻ��$�� .J,3m���[ݪ�i�֤�rD1�撷f�R�wf��js'JNݹ�m����)*ݲ�p�y��n�q���-б��eZڣ`�@-���vi"ki#K�3q6�jd�\EV�67[[-Pqsİs�rcZ5ń`]l�܁��kt�P;�B���#iy�]��n$67H�[s�*Y��1��[u�v%m�8yz��6j�mm�Ѵ��6����c�FEJ�iP jR�ɀd�9��� <�.¹��=�|9�ʏfش�Z;Um�PvMa�8���Y@Qɩڕޤ�[�z@�^�0���Yx��5�*���T-R��aX.��{��5n6Ɠ7k:���aF����z;g�][�a�6���%n�]!�'��:�ˌ�M�3i��UNX�\v�ΰ��L��u�k\ˮ��W����<i6P<��h��ۮ�[���ӵ��`p����<u�@�.Bm �=��Hguΐ��/D[-v�ݔ.z�vr�C\qJ���Q�h�Xþ~�;�x8�Sv�qkc�M��s���d���\$g�/�J@ t��]�{]�흨� 3��4Y)M�[t4���ժV(�v۪jT2Z�5�@F��l��۰ݱcۧ�s	��vm��s���y��K�<jF��q�6�P���ɛl�����Y��]+䕓�X������{p�V^��wY3����l�A��s�* �<va�ڶ�H���Y��޻޳1mm� �����L���I4E�A���㍴�t�/8īU W�nr�̸�OE2�[U*�scJ����Hd ۄ�7M�\�M$�v�h����J�vݻ ��J�mΓ�h�OW*��[mng�g��pE��Bm�ݙGF8'�M�؝���V˴lp]t����(v�c8)�qJ�[5͛֞*!7)�2 $������$���v���svڎ���o��m͗���p&�7j�:o:6�nQ�Q� L�a� �:CGWj*UOq@O!���ȃ�W�8z�2xͮ5���uڸ<���Z2�%u#.6
�����S�cmΓu`�p�Iű�;�w��n��]<��w��t�oJ�,�{wu��.͙6�5rY'�8���b�g��6���\�n����*� �A����t�a�FL�Z��i�pl�9���䬠n;m��V�6�N������Pv#ڽ�*�[U6\Q�m��Ѣ�]LQ�Vh�76aL���FD�Ɋ[��1�ݒ綢�]�t�j�K�g6���w�.�o�{:[��������d�?\��7ı,Nw���Kı>��J�'"j%�b^�߳iȌ��L���->Dr���r��aIı,Nw���?�Q�
�L�b{������%�b_~���ND�,K��GK
]n���K��Ôr\�;���a��Kı;���Sq,KĿw�ͧ"X�CQ5޹�T�Kı>��唿�L��L��6��pHEkV�J��bX�%�{��r%�bX���J��bX�'=�p�r%�bX�k�:XRe&Re/l�ٲF\e�)ɭfm9ı,N��Mı,K���m9ı,O�sҦ�X�%�~�}�ND�,K��2Ka�ΚkY�Χ��*��t�&���9룫�d�g��mFۘ�=v�gp����}����ow����ND�,K�\����%�b_��fӑ,K��nzT�Kı;�z����'-�.,��Re&Re/��M�|�����b\�}�ND�,K���Sq,K��}�ND��j��X�{�?5̙dֲ]j�fJ��bX�%��6��bX�'{sҦ�X�%��{�6��bX�'�掖�I��K�k���Ijܷr�5����Kı;۞�7ı,N{���Kı>��J��bX�f�k����r%�bX�����2�h�3Z�d���%�bs���"X�%���zT�Kı/{�fӑ,K��nzT�Kı/=�fY�5,��d�X-(e�K3���*��ѧ�8�ӻ-sɡ���5��8���w�{��2X�z�Mı,K���6��bX�'{sҦ�X�%����6��bX�'ƻm=��%�r�V�J��bX�%���m9ı,N��Mı,K�����"X�%���zT�O�[�e&Rޜ�:H�"��8]ɔ��V%�b{�?J��bX�'5�{[ND��x@>tj&D��zT�Kı/}�fӑ,K��eˣ�5��R��Fk2��X�%�}�{6��bX�'޹�Sq,Kľ���ND�,	I��=)B�
��������'-˗Y�A$Nv�&A$w��m=ı,N��u7ı,K�{ٴ�K)2�)n�V����w-
�li鞦:xr�)���O��E���Vn���We��z�l�%֬�d���%�b_{�ͧ"X�%���n��X�%�{�{6��bX�'޹�Sq,K���w&���ѫ���K5����Kı;����Kı/}�fӑ,K���=*n%�bX����iȖ%�b}'�h�&\5�&kY�Sq,KĽ���ND�,K���D�Kı/}�fӑ,K���۩��%�bs���I�.]f�\ԥ���r%�bX�ﵲ&�X�%�{�{6��bX�'޾�Mı,��� .D�~��6��bX�'Mz��〜 �n��)aI��I���w6��bX�'޾�Sq,KĽ���ND�,K���D�Kı9�H��&���`�ٷA��c[T��N�őT7��tݳ��s��`��S:n�U��ٲ��Ȗ%�b}��7ı,K�{ٴ�Kı;�kdMı,K���m9ı,N�Y�<B�3T��њ�*n%�bX����i�~:���'��["n%�bX�����"X�%��^�t���L��_i7T�ݑ�.̳5���Kı;�kdMı,K���m9ı,O�}���X�%�{�{6��bX��i湓,��MkV�aq,K���ND�,K�_l���%�b^��ͧ"X�%��m�)aI��I���^Z-=�Z��e�fND�,K�_l���%�b^��ͧ"X�%���["n%�bX����iȖ%�b~B	��5(ĚUK��?�˻��(
4W!�������j?�[}�68�A�ژ�6�<pOF'I�
���:�V���Sp���(:��o�li�@���}����ҷ��t��a����Y��ݰT��n�鳱�c!��]���#��[[������r�%�<�H�g�9����R�[���=�P��u��t���땸5˩�<�X�{<�!����5	5�ՐS�1D0Rj�i�]�]�t�D!l���������٠H�CprFy��*�����/kKWT�ı,K߿�fӑ,K��}��7ı,N����Kı>���K
L��L����5G�q�w"�r%�bX�ﵲ&��*��MD�=���ND�,K���7ı,N����Kı>�m��e��%��kXD�Kı;�{�ӑ,K����*n%�bX����iȖ%�bw��ț�bX�'~����5�W2CE��iȖ%�b}��7ı,N����Kı;�kdMı,K���m9ı,Ox�4x��f���њ�*n%�bX����iȖ%�bw��ț�bX�'}�p�r%�bX�z�eMı,K���F���i��йⴽ/N�{N�ŮCu�}�>K��1�s�8�Yb����8��r,��Re&Re/{o��bX�'}�p�r%�bX�z�eMı,K���m9ı,K'{|�2e-�j椹�&�X�%��{�6���:���'}}���X�%��{�6��bX�'}�䉸��T��)}���i��ո��r�YK���,K߯�7ı,N����Kı;�o$Mı,K���m9�2�)hy�O`�ݧ	w$N��E�bw���"X�%��{y"n%�bX����iȖ%��Fj'�_�*l��L��_/s�g(�dwcn�YK�%�bX����&�X�%��>������%�b{�����X�%��{�6��bX�'}!
f�
{R�-��� �qPnӠΡ���M��l�������ҧh�\ �m܁K
L��L����X��bX�'}}���X�%��{�6��bX�'}�䉸�%�bw����2۬�s$4[�6��bX�'}}����c���b{���6��bX�'�~�H��bX�'}�p�r%�bX��m��Y��Ժ3Y�Mı,K���m9ı,N���q,t	��"w���"X�%��\����#)2��M�wwq���(�YK���V%��{y"n%�bX����iȖ%�bw��*n%�`~j'�~���S)2�)0�}N�#N�\��q���bX�%���r%�bX���ʛ�bX�'}�p�r%�bX��{,M�e&Re-�6ǰZ��ې��t��5��6�l��j,�,e�O	��U�W.k
\�fӑ,K��zT�Kı;�{�ӑ,K��^�7ı,K�{ٴ�Kı='nh��r�Z�rf���Sq,K���ND�,K��z��Kı/}�fӑ,K�ﯶT�Kı8}�Y�5��s,պ�6��bX�'}�����%�b^��ͧ"X�%��_l���%�bw���"X�%���m=��,3�nk-Mı,�"�M{����&���#L-qs��)��\Iq���@��K,�$�@���/���2H�w2y�d���\��W{�Zu��<X,T4�Mu8�z���;����r�����&�;�K�d9^����������]��[f�}n���,Țm�H6D7&�y�Z�٠_[���ٜ�a�=:��#eܒZ�q��t�7��Xr�ٽ�0��x�떋J�5s(��/���������@>乬+F	�	73@2IL	����J`K���s�)������n]�r�fqË�$��$��Ki;�U��v���}�������M��r�`2�f���\$�=�.��L:#�Mu@��c=v;/�y�8)�>uN��;�ƭ�m��jU��r�v"s/2nGg��)Ƃ#��md۶��y�(Nڲ�X<[%�q!v�8��vn5�z�H��`Uu6z�2+�X��	��B�^�;p��Yy;�����}�����mMN����g͸ܕ��/;��C���]�8Ln9����8�ي8�H�Mܟ����� {wf�n�������[i��vԊ&G��ٜ�g{��݋ ������N(�pnM�֘I)���{�kLn�0.��k�	܅���I"��T���n�, ����O�����q}v�ԑ9n2�T�����M���֘�)��T�*�v[Z�`��r�Zw.I�<���Io[C��ۋo.�&�\=�;O �0Z���e�������n�\�0.H��}��;�s��O����.&��`��,�R	�"T"٩��~ٹ'�{���;���%�aq��i�	73@���̍3��%���S�����	^�r)xF���4�w4�٠_]Łԩ�������9t�Ԋ&t�d���ssw����0&di�??-�������l.!â��'&b�F�Pk����v,6�=�b�����郾�"��;�����̍0&dk���������Lt�����@��ڒE�}��X̍0�)�.F��s��{iW}۹W#�9۽� =�لMR��75��"�϶5�� �H�#����pgF�����8�j�ት0Eؙ�Y*�$�1�� �lc��I��}P:��5�z"i����lJ qG��qblU͇�$ҥ�p6hqH��Wq Ax�\Aۤ:0��@H
0Uv(`��h|P� O��Q���|��S�Q���O�%�f���7{�`�5�dl��8_}I����7i�����0&di���<+$x�Q�X��@��s@��s7w��&��3$�u�"��w,�����RG�s`č��s@qg��wf]�*���h�nX���۸���wb�%�i�fI_�8�%~�4�ŧ����
ID�������u�h�w4��h\�E�#Y&A��� �%0%�i��F��4���:�TI8��1��4[w4�.����WNA�oG&h$i�/#L$�������;�#���5=��ײ�7C��9��õ�ʍ��yg��;sbs]�\�tW}�^F�I)�/#L�4�>����"CrE�� �l�/��hm��/��hZ���G�EŊ94	y`d����0�S���{���X���۸�?RO{��`��X�٠_u��>�6X)$y����4�2IL	y`d��_9[C���&��n��k��r۽�VJ zJ
�wZ�4�Ẻ,v��4 �|�[s$��:�`0'lj���p�l�a�-uCt|r/T������o-�7���7��{<o: �fx��sٻe.��cG4���օȯU�bv
0���㲴[����ַ�O>;3uP1c��^�uI��zP³�ܵ����Qm r�;V4-��T�k�A�d�s���{���t���<�
�&�������0vU���w�;J�e���>4���N����, �ݦ��02H�^F��E�H��G c�rh�w4��h�w4��@��J+�' 5�cU���#L	y`$���0�GfD�r(�Ȝ����u�h�w4��h�Y����q{ޤ�2IL	y`d����0'��k~u�[��%�M&��fc��S���$�vǤ�ε.z]��{p�A=�T��7<ת��4��#L	y`$����l5]��w��Ŗ�-IUD"���""D���<���i�}�i�/#L�����Uw�Q�i93@�빠m��]�����bˎ��J�$�b]k�_u��=�2�{�4g�$Y"Jz�
�ު`K��I`K�� �Y�vp0H������9����m9A:�T�sp��s�cS�F+ɻf���&��hR��[{�:�����n�����$����s@>���&��&(���_u��	$���0$���W���*���\��wq`���7�n,.�I*WIe	� @���j��#4�b�_�����}��7$�}sDj�ơŎ94�S@�빠�4���,n3b�M�`I*	�`IL	r4�>���:s���Q�uFÎW1H��Vn\����v$8���`PN�g��������$���#Z��n�h��[g.�ڸA�A� n��~�ŀ[e4�w4�T��%	�c��T��#L	%A�3#LI)�vr�\1�kI&h�V�{���'��f���(F*�/w��=����"pjb�d�-�]� �%0%��'��\]^�u�a+۬�Ls�6r��-�s�C�>�۫ٝ��@s��Ro#Qc�A7�m���������h��hZ����O�s8��/���:�V�{��u�hs��0X�f4����uv��]� �l�/���>�J,N�Ǒ�i'�{��u�h��h]�@���r��8A ���m��`d��`L����W8��8�R�X���V w��5�w-2a	5�zi�jۧDB�>�nA�1�)�4���4�f6R=lt�nft�1ӠbLsm]��xC������t�p`|!��&:.L=�Z'�=n���f���������Ū��L�ɳ���
�Ә-��wD�9oV3$�u���'-��[;m�v.+���֌�ݮ�^���3���\��뱷gq	�v�꿻��{�@���s��n��q��ɜ�3�(oA7h�]�+� �OdI�UjK���TnkL���	�`$��y�ޡ]�"ݵjI�ן�R��۽� 7���n��ﴻ�2�����Z�٠_[��uv��/*��� ��Q6�h[f�n��=���:����}���9��Ŏ94�w4�ՠ�� �����_�Kr�Z�[�b�&g�%���8z�{��cf�6�CprFy�)��8j�X���۸��޾���`�l�/��hz�'qH�`�N- ���s�w��qs�K��T�������h�\v7�$L�)&�u�h�w4�S@/���ʕ�$�#SpnM�����h�Y�m���]m���ly$��u��q.�M��&��^F�����4�C��v�pVg��<r�܆�����z���L�Ze�h��.&�����4�2IL	r4��*K���$$�lnf�u�h�w4�S@�빠Z����Os�M^F�%A���8�=��F��J`}�X�X�f4����u��ۻ09R��{��`{��;����$���{��u�h��hl����ǗkF�,$�X�#�YݧA�GWDp�i�n��q�{`��=5���~�?J�H5�w"� ����� ��� ��s@�0��P����@����\K�&�h��5��J`]�{�19&��93@��Zg�ߛ7����ŀ�iw�e���N\Rz��RK�&����`K���8p�+ ��D�*r�{wrC;����	����m�����������<}�ŀn댽�uj+f�,�'l
�箍E�۲�rk�)q�:2����i��D�qG18��/���;ou��n.IR�`owL�؟[CQ���� �����~��U����, �߿L~�ŀo����r[��m���&di��F��s�\�w7Z`M��p}m��eڵj'܋�R�����`nn����:��Is�]�7�����_�Ĕ$s���/���:�V�{�lܒw��nI��)!��B��eH��B�#aY=�N@G��� |�8h�hV�V0��b�!��6.� H��� 0����(�J�A�'�`c�,`��Oi�<`�BCqA�I! ��"�)�	!T�UzȿV.�q7�F(��
 �@Wݪ'���PdڐB(r$�j)�B @qXmLR�b$��;P�b	��K�-���@�n�*%ZWv��ݪ�a`) ��u�fڕ�M�˓`m���A��㗌<ֶ�{b�F�s� 0 ޫ�x��.�N�R���K0\��U��),���f��aze��+v����F�ݽ�zs�Vy�j��K�V�X6�mH/d.���h�[ �$牕��,;��j��VN�vW*���]z���c�˧MA�k�4���e�� U����T��6,�'��(��\����<V��I��\BL.��T��V u�	���ӢL3�L�Cw5`�j��i
�/nN��v:��6�vj��$R�`!8U��\��k�@V�P�B��l�9��t��z��V]ld���Wb�zB�p4�lzzޠ�*���[ rgn|�S]�gu�� ah�����ke*uW,ad����v��/�M�`�$[<�c�����Sse�����r8����Zp�14\`�ͷ!���/3ց̝��� 6�p"�2�\�}S7]��BP�*��n�b��n�6�x�7�6��]��PlR�ҡ�a��=	�L�3�EĳsYs�ѭ��ڔ6k�R�Gt���U��n]Mq����c̩�<�ᢸ^g� �*����s�&��9��ؔ�n�Aظ딂����&l�(i�vMڶ(
����jw>6Tz��Md�����ZM�[��9ݐ �:o0͛�Vܮ�T�$˴۱��΅�U��PYt�Ζ-��D[ ,$j���i^�Cm�q�U�52����]��l�]�am�eB)��U�Uy`x��Cd�H5�b���̓@5U[Q�Ӧ�+�ev�PM�Y�h��.��*��[m׃�m�)�l�*����wnr�9�8���UWaՔey�<�����6(�[��j�UI�WTm�'Wj�u��v^��	1 �ì� �[e����Qׁ��m��71����"�e;u]�/ne���52�-l�CT ݗ�}�w�w��w��rq-H
?#�b�(�C���:��ATM�b*=��g=�߹n.��v��\��n8�O����I��=v�ӡۗ�M�!��S������u�T�u�p�J;z�cr��;�z�Қ�zuN�\3͹��
ɸ^��E�ֈ8fؐ:v�u�3�Yk˺1i9m"�;��g\����6̥I�Z����9Nt�W`I�{*Gtr�'�$4�n�d�]a�P��n�̛�v4u�۞q�y�v}�\q�U9�r�zؔ��2�^sv��Mҏ]l�..+!�s�O�w{����˻�N��R�_�w_s���`�vr��*�a��ŀ{��#.����LnE�����������^~��*���{�X��� ��.G*�����i���u�L�L	ۃ�[�#�\nEqȰ9R���w,z�� o���J����X��>���,M����XI&*J��s�IW�����y~����A����~��A�A�A�A�߬�?�.<mn�<���2'G����!q�t7�+�8�V�?{�ܮ���sl��b �`�`�`�{߳b �`�`�`��߿p؃� � � � ����6 �666>����A�����g�_��h�)���Y�y�߿f�D�>F+ ��yCb�A�6?ٿ�y����b �`�`�`�{߳b )�PA�l}���f�ۓ3Xi�Mk3b �`�`�`�������A�����߮�A������ٱ�A�A�A�A����lA�lll{�[��֡u�iu�M3�<�������]�<������߳b �`�`�`�{���؃� � ؂� ����6 �66
T�IS��]�wq�r)r<T�	������ٱ�A�A�A�����lA�lll~��y{?~�y����?��c��vɚS��n{5�7���r�-�=�4�A쁡��,�;�V�	9�������n�s`�`�`�{���؃� � � � ����6 �666>�~�v  AO��� � � ��߿�b �`�`�`���~�D����D�\̗Y�͈<��������b �`�`�`��g��b �`�`�`�{߳b �`�`�`�{���؃Ƞ� � � ���j��3P�R�Z�b �`�`�`��g��b �`�`�`�{߳b �b�Q��
F�%jt����yA����lA�lll��~��A�A�A�A��Kw���s5u.In���A�ll_�B"����~�͈<��������lA�lllw��y{?~�yw%?j~�jh�)���Y�y�߿f�A����o�؃� � � � ����؃� � � � ����؃� �!LT�1RU���Z��e�[-�,,]����b�J�6胹5�����<�s�x\Y��b\���N�kY�~��������6 �666>�~�v �6667���6 �6667��~͈<����{�sZ�.�-.���5��y{?~�y����y�߿f�A����gJ���R�V�����F]�E���\� ?w~����:��M��q�n�s����	�1�2)&�z�4�=7$�u�]��~�V�À��~�������<�N'�"p$rh�S@���`2S �%05q)坋Ut��g��l���²ok�Z�@���s@q�˲�퇱q'cj7�[������@/u��l�/����8J<OS�c�n�ǀ�l�I%M���`�`���+kY��j'���.IL	r������ �6�~E,q
)����4�)�w;V�{��z�4{��[1�I�<�����:����rJ`K����<�
$V�hT@���.j�&�N�t;0`�c���/Vnl�h�b���.�
�Ѷ��2d��֞\�v�6+9�+;"�r��.��K��=; �F6tsڇ��<���@N�vzv�����Dkm���g\��M���o&Y2�i5�Y����e�/W�W�$'�<SI���:�\6-�*��60gE�s(�aʃO`}
+ql�hn<y� �X�q�����X�[n1�(���T�����\�����nѕW\=������lNZ$�s���^����z�4zi�����< �ܬ����W.G$XrJ�K�7eh��۽`I�����g=�h���2;�rI0�`��ӿ~J�� =m����m��}�W9�����5�rJ`I�M�p�x����&�4z�hIRI�����8�=�`}�fH^x1܊�B�\��]�8��B�&�w=�S�X���&F�)Ȳb��3@=m��P`fJ��../��9�_����y���r\WW�0�f��U����0�S�s���L���_�/zD�6Ǒ�h�O�@��s@=m���L ��m��n��.X�RH`uUR]�7��3wi�.T���2���`Aݸ�\�H��ݘ%J�{���7zq�o����ix�D��I���M&��t�]��F��YQ{q�v�:�k�6�28����OD�H��/����e0��UR����`m��DX\bwi����=�g����X����L�IR���v{��rӿ��1�7~�ۿ�`$�~���K�s�+�8�����zq�{�{i��e�6����L?$�{��Lͭ�������h[��ڐ�]8]ɀo�4�9%��O��5�rJ`b��w����<�h���S�¸9��Ɍ���ƫgN�]��$�������4cr%��<���-��Ɓ{�����U�÷{ }��}m����c�I!�o۸���M���`�ذ{f�ԩ%T�R����_�(�\��� ��~�̍03%A�.F���[�q���$�I>���n���rO}�lܞFh�Ө s��M �I���PBs4� ����ߗ�������&�ޯ*n��c[tO���d��˂�Fr65����C�a�	�qð+o�ߗ#L�������&֌�k����2%�ܙ����]���`��,��RK�٫m���mHH���ɀ~��� ��i��J��wb�wt�=�H��7"X�c�$���h�4��#L7�%�ݓ~L�o���{�\E��I~�ŀrI������nI��=7$�'�$@{�'�y���c����Q�}j�e�uu%.N:�"X�dԚ��t.�Z1��#�H��e�Ix��n��W*�o<ݑ���̻�7omzώ7]v�����#���,�[���U`Yλ�냞��T��3nq&���e�;vR�ې�a,�X.���bl�[���:���"�'g�z�;KWm]����p�Usa�+�	��ɓ�뿾�-�����g۝LE�.+���]���>8�^z׆v�78.� t��n�.j��V/v�24�����s���L~�h���i�9rI0��~J�RM��`��X��ٟ��M��>�0x8�M���^���/���>�w4��hS�QbwIb`��c$�0�J`fH��fG��A/�&D�AI3@>�f��n���M�����<�я�x�����:&�e�ӛ*�����.�_a-u<�����Y�K��!B�w'��ذ}� }���I/�ݽ0{['X+�e�ֵ5us�;�}�~GH�����}�ذ{w~�l�˥����"�H�"�wt�?�ۋ�J��{�ذ��, ��?2��ܲ�rL鑦d�02�4��9����^��ߦ���/�d�����X���`~IL���I���di��������ܑ����O*FËp���=��ù=���;S��{�����������[�Ԭ������L�0>�4��m8;�q���rH�����K�T�U�����߿b�=�������W{AH滛L�0>�4��<s��P�"���^{0R�'�8�Q.`l��[�&�K��2@r�|�(H��y8R�P��� �s�.+J��y Cj�"���!
n!`���`CB���$]z$K�B�<�K�Rc�D��`�A��ЈT�P0E9��� �>J(��\�q.N]�[LfJ`|��RWk��*����Ԙ~��]���0&Mi�fd�׮���"V܉bm��L�;�Z`~����s����`g����#L��~y��hGm"=ɫ3e�D��r� ob�/IW�3m���Z�&@V��:�U�3%0�J`}$kW8��L�� ������2&�s"rh׬�>���=����{fuU$���v�d����$��݋ ���X�{f ^�@>�����~M�x�������&$�`L��w�!p�BI\"@>D�:z���ύ�9��K�;�$�0JI3@;�� �����X����?U$���Ó��Ki�ӹC�����63�����m=v6���퍏5\U�wr�"co#�E��O�=��L�ww4�]� ��4��lQ%�0U�z������s�&JрI6��$�>�$]h��Đ����Қ�{f�l����wb�?��;�ww��ے`~J�&�w� }�� ���X�S{��k8�D��˷$-܌钘��8�{���d�`�)��T�W���7 �*h`��V�ƹ���I=El�[��N!��sr��y�����%q�:�Z۰nz��y���<��Sw/Oo6\Cَ=t�����5fs�jlmenxbݝ��!{2�nȃF�q��B;V�ؘ�g;U<�\<���8鳞r`Mc�ʛ�a���f���|^�-v��!�r�sM�-�M���
�rm�����GX;x�k���X��]rt�K'<pm��V&�sn�=ɮ���X��vQ��<?综|˶~Ξ�U~���߿4�2�S ��L钘ׄ���������73@;�f���s@>�f���������=�����M�ZrI�ww�X��ه����X�ޘ�#coc�E�r,ʒI��z���02���̍0>Y�)���z�$�R���?�wʒU���������Y�u�C,�F8����bR7;v5tq����YMּX��[8��r����1��bHLrf��}V���s@>���$�����������Ʈ̻�w������j�O�Q���ޘ��,�_����׮�R��U��I�}2S�#L�qs��fzoX����V�yZ��rI�_[��/�:������{�6�d��֋E�)�%��,~�k�?R������ޘ��� +��N�t�
��� `���˺;��T)�N�!��x��m�(40 $�8�I��)�{��_u���/ʕR�a޽�o�tm�N�XY�U&/%0%��_��fF��R��嶅��[jBKܘ{�|�Z����h�@�ܫZ���X�cWr,J��zw<�{ o���$���� ��G|��\cW�u�3#L�vM����i�/�u�ʩ>�c�]bnX��@�$L�t`��k�+u���qm���B����ك�����q���zP�I,����L~�ŀo׺����WW����!�17$����Ԓl�_s�;w�`��3�URM�������SvKe�Xz�������Sgn��;�ذ}���\c��}�u�3#LfJ`K�����U� �F!$EO��&*o���� �lm�N�XX�E��l�?%��ߗ�nzoX24��e���|��_�-���٦�� %��u<n��&V(�v	ܖڐ��9n���݋ ߯�����U/������`����w,Đ��3@�}V�{��}z�����ߒ=�H�	<Mڀ^빠{�����/�U�\UU���hS%W�U&��L	r4���N�&di�}T��x�H<�ɠ_[��w��`L�� ����I�q	\K�x���;Yیu��#<;�錧7L7r���Tpt�'=��Ʊ�l�Ւ��0�ۙ\�Oa�}����S+��Gk��1:"G=G(9���k3s[E�v��N�=�u�v;W*���lpl�� �9͈Z��Kn�ݎpZM���� [V���w�c+m\V3Q�˛��묕��Ň(<ӌ*���"�k^�ݸ���	��9�a>�{�G��\s�q�T�8�c��
�{Am]��tm�;���\���$M�r��hng�����]� ��4�w4�I+X�F��u�3#L�J`K��_��,�ĕ��&'&h�Y�_[��䒪M�y��ذ�Z޹m�9,�ܘO������< �{f oY�}�TٌcN3B������ ����%0%��a�w���;�qz�y���湲��c;qۗ�p��Uu��<�7��21�6�8��"�h�@>�f�}n��}V�}qUW�db�$rh^���~��?6Y.��}V�^�4�(�ưrdrI3@�#L�d� ���L�0����0������w*�J��M���@����>��hܒ"V$�0���]`�)������`g�ߚ`e�'Xo���>�3��v��Q�'T`8X����	k���Aٜ��;��-�f1\�]�G}T��di����_�u�fd�����(E#HNf���s@�}V�wu��]��r��cq��N��R`K�N�̔�ϱs��į���: ��8(�D��w�ŀ~�݋ �_x�����ƭG#`�)�/#L��0%�'X�M�E�%�B�ɀo��X��W�~����}������Z��7%���ɍ�m��u��6�h�A{q�v�:�Ƹ'7n+�X�Aǃ&F�4�������Υ�ý�� =��v[�
�	k��&�d� ��L	y`}$i��*�6o�c��.X���ۑ����7�n,?$����`��x�#cob�	�`�NM�]��n�|�Z*b6~ ���~��;����4�"� ����n�|�Z��h��h��ɉ��,ln!ș�]E��i�\N:&2=t��e��κN�S�}�I���q���������wu�*I0���`/i�;��q�Z��3%0&di�����I׫�K����>tE�%�B�ɀv�b�?����ڴ���/ yI&�]�"��UR������޾���`~J�$�w�� {���$unӻ����:�32SfF�I`W>�(�#�(:8렦��ܑ9� Ί�%e+�(M;S'�H��􄑟}�M1�',�X/8�a�tjFti1ЄP��ʊ�G��1N�,^�F�Љ�#u�|�w=������J�UmR��T�R����Z뙀��$�:2d���Mԑss!�i�k!��s��k+�6�J�l� ܯ\�]���m�T��F�.��	�	NG��:uF�'.չX��q�;��x���e�Y��5ۃ�w'c[�Y$�;6��0�#�6��gLM���meM0d��觬v��+ڮ��-�1
��E����	�0MیҨ҄��g���LŊ��)�օ�i���m��^u�)�۱�[Б�	���m쵳8��ʶ�ca��X$�uu@ۑr��U��@��V86�x6f�Bg�R�n�esu���%�nۗ���&��v��m�y@����Vp���lU[w.�tm���g��d�J��y%�n�s��!�t��:��Nu�2�����m�*��0��r��2��u�R�&8�b
��l�N-��6�\ex���Ԅ-���c\�<�rV�t�nys�n' (��n�X牵5m����ԯ3�*��	Ӭj9h�:ឤ6�'�U����v��'\t6ʰ�m����.���nIc��`� &��y��ɶ^C5�t�m�쭲����u�NԪ���W�.:�e��-u�<�4���v�g���S�u��d��5��Bol�l<7
�f0۶�PX�NC�L���c%�52��]�(cVq9%�Z��lyL�.�s�Q�L�.�SgY�˶RT30`\[7 ��]���艣z0�` ��\�6��Ol�f��f�ճJ��]V�u,�r�;`�kg�`I��m7YY:��[�e���,��)�]@��[]���y�W�MU\��wU�ۜp�"ziP�4�]ʵ)�J�����2���R��q�α�^m��.�sR��P�*�:��%���Q`
�ġ	;ks�n\�nM�Tpݔ 7i^^{j�;�ݩ�-���>�0vzk�8w��k<<eO<��d�1�S�É��U�#�`Ԝ�}���ݡG9��1�P> � z�6��QLD:!���������߭�����
�B��+m]r�v�ή[����*pޞ1��na�C��3u�E�RV��G=�����|���oBNͳ��(k���e�`S)ȩ`�m����yw�f�(n��[�o)u�RZ54�
��az)����gD����n�\3�zbRۖ���x��ٴ��[[.k���̕d���&"�7�=v;A��4[��w���U�����ɧ�T9�n+9�{.��X5���Z�64�q�L�jA���~�J`L���#Z�\���M�pG��"e��ܘ��ŀn�,~�k�{�3��I6}����[p�8zv�`^����`�)�/*��Ee��X�Ӳ�X�U*}��$�`Kʃˉqs���&��u�m�q$<�E��f�}Қ�����ZS��0f=��?�G\R�p��k��n	^8��Y��-� ݳ�7c{���M��W�dy$r|�Y�h[w4��hwY�_ t�&�MffM�9�{f�"G�J�-F |�M��7��m0%�A�\\�]�f_���7!��G����;�����/�S@�۹�w�B��f$�F�WX�`}2���H�I%�̩��9��u�Ew�`E�o���H�/�:�����\SIާ���< z�����Zz��I�̀�����.냝�s*ۿԩ)�/��p���w��02���̍~K����/i�bHLrf��}V��빠}zS ���,���g��G|��We��{�w���rN{�鹤���F)�'A�s��w�d�0$��`go����J��REw"���ݹ���b�=��^UR_��^�~�`��_�Ii�]�]Uz��#L�d��#L�T��r@�3�#m�l$`��#��/\��p8;4r�OnP��G�w���y6Z�KW�}�_3�z������#L
��bb�f$�"H�w]���L�۸�}~םJ�9����"���&�d�3�{��`d�ۚ����QE!Hhu���d��#LK�f��$��bs�Ibc�4�j�=�w4�)�}��h��,� �F�A��^�K6[%/�� �v:��y�6َ\�����Ɏ$��8�w]��Jhu����ý}� ����)mڐ�+�3*�8��zL7Z`n{w�̍=�9ʦ�����RZvw�w|wb�%�N�x��&���+Fy��[��q`s�N�n�b�7ޚ`~}��`�۴�|��v���=�`~���9�=>p�i�/�u���Ă�E�F�b�����R���ML!!�[�K�M�ø-�6�Z�i�S3�#R�����S1�db�.%�P��t��5�ېٞ_]r�D���v8iQ�hq��-��#{r��s�nݢ������z������n��,��d�󥆣;`�e�ed��E�ţu�D��c�g���j6�!nR����@]�p�/� �-u2�ܹ�T�[ˣ"��$u1�;����{݌���:N������ݮ�wQk�@l����][<q���s5����\���ݻT���h��H�_��3#L�WR���)�$)��s@�v�����Қ��*���s�Ib��L�I�fF�2���H���"to&2 y�@�빠z���|[��w��@��O���y!=^望�T����	���3#X*�ۦ3�:�X��eʶ	��vv��h��Z�{9S�n�=�`y@�.��E����r/�;�v,�^��=�n,�]� ��^4�~j���h�νI|�q#9ʢzkL�֘�`w�7���q�����;��h��hŻ��h�`��!{�j�fF��`K��`fdi���oGq�&�q`� �w�s�w{����=����[#�ʒvƲ�i2�cn�����O0qbx��Ry�q�F�1�"���s�Ib�93@�v�3#L	�`K$i��2����JȚ��<�����6v�b�;�v,�ڴ^H��L�O$�93@��M�=���nc���F��H!��/����<���X�~6'n8KWawqK��?>������<����7�w4��,(܇��h�ՠwu��/u���%x���$�����oǈzz�87��6kx���!�d����a�Uj������C�݄Ѧ?����Q�$�u�>�$�t5$���}�IU�Zx��.�写s,ݶ�w���y�!${�m�ޝ������FO�R�����q�%�lw��m�ӳm參�K�]F����������M+�Ь�|�U~T�I��~�ͷ�?�f����r��1G�UQ��@`�(��B"��H��A(�U�%M���7�5$���|��Ɍ&'�$�t��I%{����%x���$����K��W��1翮ثe��V����sf���e�[y�܂�p�Iy6:Ϳ�{����k��t���r��ϛm�������oW�01���7_��I^�Q�$��l��	&	ȣ�g�$�λ��$�����$^���Kׯ���ԩUUݱ�����
���M�m%z/�I"��Ԓ^�~ϾI+�wCRI_Nm+��`�"#��H�)5[o��p�-��}�ɻo�DMk�w���-�]�����8�j�p��o}��_�͵s��jI+�j�䒽%KRI}��Z){:��`���rv0V�����'������뇵\�z�<h��a{h��Y.ۣn���t�ٸ�#'�nmT%p<]��oE�-Z��B�O��n;d��	�(�<�Od��c�8��2��5����v&�ɂ���˷//>�خ����q]6�6ۤZ'1��������;���s���VA�*�{v�+8]�Ƿ��뭺��~>>ӿ�<�m�ɖ�L=fճs��
եa�opGhx2�G�w���ۖĈ��6;�u��-���o~�������k�J�W��o�{�6߯_c��m܇�cr������I+�T�$��g�$�λ��$��S��&�LdŎ+��������o}��������J����ف���l���6ٶ3ڑ��#��\��$�v��K���ԒW����%����D��h�)>�$�-�m�ԩR�gs��������{�f������:�����9S��[;u�j�v�UN�q@q�Y�ݍ�a���{-o&5$�jI+�j���wCRI^��$�e���$�ӓ���&�������{{�{4�iB	�iD�GKTj �#D֊�T`P>���������9�m����&0߯u��J�M��i�|�q�+Pw�g����������`zѥ�q�%�lr�$�wg�?��u����*�j���r�Y��h�ՠu����;-��;����q�Fӟ�Lnpd&OyL<<=v%8�/V���ggv`�������o��m��C�������;-��/��@��s	�������{*RT�'X%A�Iw�禧n5%�`�(ܗWt� ߯u�f��A�������¢9`���}��� P�D�"�(mBh��q�BB�$��ςQ�!t|���cC|g	V!C�6��S�!�#���Q��Œ�����+�]�Lc�!F2`��pbr��c�H��H#_�c
��XB&��)
),���%�90+��g#!��b?����=�"l���Q�uP�|�P@�kh����/�޹���}�Jh�S��/�cR9�8h�ՠ{vi�}��0:�'��8�9���}���MZ[)�{�S@�S ���x䪩�pu˖�.�F⻻эjLc����d�Y��A�@��a���֡�s�������;���N0-٦�׺���������`֏���c�K������M�v����=�w4
�Z�14���cr��ZIPf����n���v�`}fA���ڊ���<�RT��8�=��X���~��zZ�\iu�&Fӌ�˗!�}��,��U\�~��|����[)�_uՏ@�,��1��n�u��]r�=��ێ�u�5�5ҍ\�q^F��GS��s$���;-��=�j�:�M޲��#��/�cR9�8h�y�ޓv�`fn���%A�;3�|+�F`�&"8��S@�����l���;V��k
�v	2@ǐN�;��F[����u��T��/nX�K@��0-٦��%ř[��	�Z0.�A��Is��$q8� �H�DM@�c���n�������&�Y�m��G�v�Ֆ��f[E6�@q��V��)�,�=���<���ӧ���K;
V.#e.0��g���#�ݫQl��&=c�4�f����t�GJg��N��c��H�:���"��v4�u���ܘ�}�]<v`��	=��N � 9d���Qn�Y.�nq���z�a5��&T�&�t;3�-����<&weW��ݽ���A�pnz�)7b�nA�8���W�="���"k�u�t�*?��v�[���ݰX=��X%A�w*�.}ЋwZ`{��j��Ɏ!c�Šu���e4�n��;V�|4��"�M˗!�}��0-�ŇRo޾�ot�@�x�&E�1�����h����v����=�)�z�0x;"�ڷ%�I�׺�T��8����Էs@=yY���~����AƉ6N���g�<&:Sc� ��+^^	wK����;iD"8�l���YM�n��;V�|�V�;������YG��hG8%įW8�d��L���l���xeuF(���,�����ߤ�?�%���h���i�;��qX��:��,Ԫ�?zw<��i�w#L�#L��>�#���*��8�Z�S@����:��h�hF���R�<�&`ȒF���U�p��k��8�ֺ}�-�fq�������{�9��t۹d�v��{�ذi�� ����W��`z��dj��wrI�����s����ް7v�`]����UI��İ�_H�ڷ%�I {�� �T$���8��F�	`c�K��,V��n���J���� �O�@�[����@�k*bw""Pw�i�~J�V�����=��n�� �I$��9����j���C۸x+x:��zsv��qk\��u�>�����e$dN8�C�� }���-���e4��T�&���b�7I�]�O�9ėzn�h���с����MR`�s	�8��>��h���=�]� �������L��^�z�I��s����`d&��.�>�>��� ���5�Eo7�=���ȡ�JB)#���:�h�l�>��h���<��I�Fnz�H���v3�3���/\��p ���˽�m��r�}���:vv~���Mj����ݦ�F�r���24���=�\�3iDF������e4S��{���,���&L�N�P`d$i��9�s���'�������`zзbq���`�w {���)�{�S@��uLbi9
V]ŀ}�0������=�d������?�4%#H�{�'Ocn��ק���Kk�Q� �.���cwZ�����,�Վ�f��h�ݼ.�v�6φt��]:�c\vڇ��Y�A��v���m�n��
�^����iH�un_j���F��vx��F
�g3'h켅)�]�8����)�0������ܯl�kb������<��tp�/<�s�Pc����5X�ݢ�.�vv�R�˺"���T�y�	��Ym�Zb��[JL9l���v͉S{�zu�=�����&CEĤr"���G+�'���� ��`Kw4޶hgcK�a26�b�k�0.�A�8�zM7Z`����T]Pʙ�E�p�:��h�l�-���e4Z)�T_��گUT�ܔ��Tr��Wf��� ����\�[����Lwf�܍024�.���t"�|w��cOV���NK�=b�8��Q�.�x�g��2� �YS��&�'޷s@�����g0����.�E�I0	��:��mă�Y�[e4z�����1���@�nf�]�L	%A�w#L��0>�J�[���cWǁ���wg�݋ ���h�hgcK�a26�b�i��w#L��0.�'XJ�g���=qvō����S;Iu��m��뇳�9��ݖG�Ĉ�I�'c�hmR`d$i�w�:��T-}й)P`���Ƥ��4y� ��Ɓ�n��=��,��5��i�,V�q9�˹'����rO���nqA T>�J�UoI����׀k��v�\E�P/*����F��0.�'X~�8���� ��_�I4;� �OF�~��	r4����׊�ޮ�9�������m���Zy�O'kӃ�)���q�ʝe(����9�w�o�퓬	r4�����#L��>�"��"K��<~�ş�6{�ذq�� ���y�����J2Yw�\Xf�L�F�2���#L	܋���v��e�p�,�?q���ݜ0%����I#�K����ݴ��`����R9	&h�S@��s@�#L�F��a�(�O%�*��rq�bnv��������gN��������-.L�3b�%!�u빠_[��Z{q~���v�� ����qE]I�L	r4����fT24��в�G�$$�bs4N���ÕRo{{��ŀy���&;nB�B��R`Lʃ&F��i�!�s@��ST�4��6,p�:���%��C#L	�P`E��u$s���Mv{��C�Ċ��0P��C��T.�|*b�hM1	�y�H���?}�B�4� D���D	�aX�#ÈxSqĈ6�@� b8�!G�l	N;���Ω6<IR	v�Q��C���@�1���!)��
� E#J����f�C������T@
:��̳3Y�-�ڥy�A`��i���	.�6pmtY���FJ�B̡��7�W�|F�m��8{uIٰ�;<ϣ<m����n���Fܩ20�m�5����w+	�7�@��Q̳�#.^ݻ�7\����yV�ۘ�ݜkd���}�M��e]جm;<�s}���	�0m�Ӭ6[�1���ɰ����Egq*�qtW�q�*�`�qY�A����ش��s��^�j�) Z'�#O/^5<���i�.0�ʹD�7ټ�s8���i{V!�vA��>���G�9�>�m��j�v�:��N��N�Q=Iǉ\틐փ��;\�+pJ�Y�F��v�i��D������"�K\�$��1��@-�v��zJ�ۖ3'����*g4+`ua�ک�����[�� k�h�q�7v��9˘v�u�<�&8s�����ug��ݻGkm����/��%�.ss5��Gk��)	b�1V����:ۏn��'vUV 	��:)�N�Yё���K4���D�o������Җz����P�^�;Ak��"�A�j c�xڷˆ��p�c��7+�=m���S��q�J�n���V-g�/8�@n�-g6ݱ�jR4����LjG*+.��q��E��,-��d��f,m��O\�p���g�$N.nC�@Y<T�ʇe�Ƿ'����m����[�v`�'��W;�Q���ki�=�x-I��ۦ�m
��f��z�+ K(@]]P
�F�kt�n�ʬ�T���ev����u{	.ʀV�ƀ�
��2R��	�.�L"�k5 L�a��"��k�@չ�ʛ0��Im�vU��F�a}�7]�f��
�Ȗ��c�Q�u�����{kE�*��4,����j��������OZmC�咶ή����&��W����.-�$ÇXF�8n�5�1�ZM������N��Ѭ�,u�]��eU`*�t�@5r�  �	��S��!����@�w��L̲Om�N���A��i޻9#��u�Y��2�N�#r�49#,�:SGY\�t��͹1��9^��^����s�q�՛[�D�������s��k�Щ�\����2�$j�v.�@kX8��5��q���8�� �G���ы3���R���i	�ܕ�lT�8�s��0W�C��4I�:�Ѥ���e�k����=��'����s����w��_�Ҙ�߮M8����^H��e��u��]Ͷ�r�d2���Y����ܢk�I�,��r�ˋ@��ذ��s@�Қ^��V���MbXLt���L	�?��;�d�f��߷qg�U6}�8�:v��rD���ް2��ˉ.w���07	�09z���Q��I���M�H�Y���Is��7��u�W�)P/s���F�̍0.���}��yǤW�v�:0#r�"ތ3j��.c�j�\���N#�9m�S{
X1�i�⨪A�G�nZ`]�'XyP`}�)�|�������Xc��{Ͼ��<��O/��
s�{�M�?{����oǷ~T�6w����w-[WǀM��/#L	�0>������ԥ�˸�.ܸ�9~�T�����,����s@���@��s@���U8��dQI��]�����]���s@����1�ė�yj0ą�&��;��ƥ�J��n
�.�&��\���:��/v��Uڤ��{'X24�����W��}� ����r�n��G�\���Ļ�d֘�����`N��v\�D�s4�]��WsN���<,�%l+4�:WJ�Ic���f}�����׮��4,���e�5��X��T�v��X�{� �z�h/.�diĤ ��sOd��F�y`I��0>�+��ιۥoAv�4��,�{&rk�)��z��]��]��&�F�����w���v�E�﫿�5�^F�3����:���[�¥�]�c���ｸ��T�=���^��7�n,�o[��㶆F\Q�"�>�=ŀm�^�U7��ŀo��`�k�V��Uڷ#��`~��ojoX�Z`e�i�������ė�U)�ذ>��5G,Wv�I]`K���ɿ/�֘͝Od� ���~W7]�Zl�lG3�.�S�`h��L����4�n�zt�N5�\�M���&^F�3����:�����в�$LNf����o�����x{{ｸ��g���8�w��h�w�^��7�n,?RT����,ݯ�`�ȋwq�j��y`e�i�w;`}=����vJ?FLm�I����빠wr����Z޲��~�u��m�b�x���g�pk���]���ܼ?��?{�b���euc��d�V��;OsĮh%U\\upP�O3�����D�Nz#��[k��ltv�z^ڧ=����/�M���R�p����´j�N�iu�פ�Mqәű�ܻ������cZ�-�քP�N�WVe�nB�]���y�k[vf��l[Ђ��v8Y���q�6��'9i�2B�fa��0����=�:���Sʃ�&�k�:1]uc��m9��m6�(�x�縰�k�>���;�w4�L1�,1�jL�ݪL��u�;��kFɭ03�?�M�}ör�X��5$� �zq�{�w4�빠}_U�w>@�Lp���@�u��;;���}V�����в�9�ә�ww4����h��V1���Itɷ ��Kȹ:�[*'��ㅡ�\���h�ؤd2���nH���q�^��.�4����쑦�D�T�w��f�)���rO��oʌ`�`2A|�żM�5���$i��*�/vX~S&6�	��f���s@��w4���=���8��D'2&�L�F�r������F�\��2�Ƥ��E&h�)�{��h�w4g�����EM����A)ק$l<�%���xLt=�6A��� �y���F&��)���`����[��z���>_n��0�t� ݽ`�Ep�jN���F��F�r�����\���O'0ɂi��=���޲��X(�X"��* �qqZ��\K9�w�������糾���8��a����e4�w4^�����h[sT�na8hr4�������\�0%��y�*{tl����ZKu���G[��y�]>ܖ�s8;Z{p5�]r�aڛ��\�����.Tr4���MbY1���&h�[��w����[��z���>�Sx�o��r&\�0.�4��sf��ś�0/�Gl�8�wl������?{��`�0-\�0��$�\�/������p`^|�\��c�y"s4^����i��*�`j��@ާ��'�`�ٮ���$���zsv�	�����u�'�zZ�*�r���v밍߭����L�P`]���F�=���*���ڢ�w���02�A�w#L�`{=n���5I����X�p�=�`\��?w��u�ͭ(�IGɍ��4H�h�w4g���;�S@����-tL��Ŋs#jL�-\�02�A�w#L�`E�8��X)H�DX ���7o�D�ZBчn9�0\���iyf�cچ�-��;���ʇ4�:�&�;N�ȥF3�W��[�15��n.zceR�a;1l�.9x5�m���`�Hv�c/��6�8���.7)v��i�u�ݘ@��]���n��;%�F�Z۞ȱ�ێ:`�Vi^�cW;����3��f�	yvq��$v�	��W]co"h��K�\���d<+��mT��I�������[��=�����K[��J�<�6�ێxݞm�+ͻ!v�[�#cԫ�K@���F܍0.di�j�i��u	���o#�4z��׮�������Zs傹1�s$Kʫ�����������`]�����6��Ww,pŁ�J�����{�`]����]�7����ﷴ�;#��N��X�ߵ���������X���X���	��+�آ��Ƀ��+0�������M�[��b���n�k /�C�I����c�E��d�{�4����Z{���ɍ��8ғ7$���ͣ�1�� �H�"�$U�j�� ss�Owf���^����UT��_�w�8���&����`]�i����ުa�a��8ӐNf��}V��ti�����#L�@�J:W=�.��U]`]�i����L����u���Z�.H��ŐpX��Řit�0j�%m68�q���u���<v0�6kn�u�L�y"s4�]��-��>���=ː��^6�D�h�n���:����/#OW9�ޙ����.XG%�&�w�^��>�ۋRqRy_]�~� �ӳ���P�*=C^F�|�uRuX��d%X�cH����������t��K�� �IF,�4T�l�e��XS��81f��D�E��M��hmbt>y˴f�3GXB7���Ec,�"X��H`! �@���,(�0	��|�lSi*�A�5���`&��B E��`D���P�$$�[)+�T_.���Hҕ�B_!M���D�2������v`A���A7C�R��"4�ccU� �Z�	����g���t��[_<Na�������`H!@ J�!���=�G��E�����0*��@j"qh�����5��u=�Q��3�[۹�}����nj���#b�]���qqs��~L	�Z`]�4��>�@�����cnbN�4�]��K�qf�/���ް.�4������\^ذf�N�q����7�&G�v�ͷX]��l��bL=��mBp[-ҕ�l]�4��{'Xy���L��6R1�?���8�p��}_U�{�w4}�ŀ}��,��U$��7��?(ܮ�ȥҪ�����y`]����@���ɓ#�"O$Nf��빤�}�lܓ��}w'|2#����^O�ύ�;�[g�k�F��V��}I�w#L�s�\W�7����/����%�/�rD�C���Fi��X�)D=��z�cNP)�9����]Rh�t��ԘOd��F��`]ɋ ��j�".�%�j����ŝK���zL��3u���:�.%ޓ4��S���!�	q`��X�n��?��z����t�5�@ndmH�r4��{'Xr4�y�./���Kݽ��o�V��5v\�wq`�~�`]��3#L�`u�ˋ�LX�B
�vt�f�5�Zm�k�N^�7]�����6�Z�Z�F\lk'="�nW��8�u�s��N�]-�h�<��j]v�ip�v��� Q{T��e�u�����{6��x�	�8��zy�on�g=wKt`˅I�l�k	0s��-�b�^���e�t;rQ/C�qq��2cF���S��V��.��o�{7|�iR�U��9N�8)�g<��p��Ơ�Gm�����O!��s�M|eՔ)e��e&ZPݱ7;l=��qt��mՕ�+���<.
���Mt^}�]:UWX��i����܍0>�ՠw>U&9���y"s4�.s�険��۽`]����zM�i���`㸰��ŀ{�a��IS~�v,ݽ� �o��)%�9-����02�A�3#L�a�$���ߖ�o,r ��"]�.�ۋ ���hz�h���>���ˍ
$�+`կf�y�Uٓ\Q9��P�գ�=cdǧ ���O&&�	ȓ��z���:���;�S@��s@��X�"k���\�rN��ٿ"�X�'��	��"�O��sy�ܓ����p=z�h��2�68�dNf�ޕL�0.�i��#L2��"Fco"�4�w4z���]�޲���Rd��� �H��ޑ��&��3kF�`~\��uo�3��/��5��qrh:J�GW8�I�sɖGs�{��K�d�2����ۿ�`]ʃ\�0.�i�s��J�#DR4cs4z�h��h��X�ۋ?�&ϻyc��q�h�y7$��߶nI�����Em��hQ��s=��f���rO��l�����4��4z���]�޲����jʱ�D�%���̍05,�z|��L�`}���뎀�ù���ɅS�՝ggq�WmKځr�ۂ���.���콹�#�\�=wԘOI�.J`fdi�3#L�PM	������f��[��o����ל�9��vt"�q��;U��Z`L����:�%�L�rkPI�����/u��>�۹$���nKUBD @A!��T����n���7��{�ӄ��v_�0>����\�?sߧ��`n��25�{��6-[WR�r�qE!$ds�Y2'&��@�9��9U�z�ɶJ��m�WEv�[��X�qh��@�빠^빠}]�@��#��OƜ��rf���s@�����u�.F��w�{ս^��{��ܖ\� �׀n�0�J�}��X��s@��<uE�i<qǠ}%A�.F��a�%���03Ow����Qܸ;� ߷q`�������^�����R
���T��ٶ��:gm��������I�i�7=��;��g�O}8^�<��U#>�
�)�X�z[��n]�۲�j����ϵ�.Kš�eۛ5�;ӿ��>Z�K�v�0�b
qص��(��ѭ<z{D�<j�D ���`ஂ	�U�^����.j��9d�8�Cw'A��^��`҅]S9��d���������.�>�*=�S� ��T��k:�ֱ���mb��Kpu�EAʰ�z!�a�m�*�(K	ur�����ߗ��w2y�����s��/���0-F����@nF�f�Wuz�ڴ�w�{qg�6{�_H��N[�r^�_s�7��X~T�J���ŀs���^��L72'��Š_[��wu��*�@��V��pG4�&]�E���{q`�������_[��Z�ˋ `!�x�1��Ae���˘��r�ώ� �^IݣZ�`��N�t�҈q�ɚ]��Wj�/���;��h�0ǎ��cc�'�8����ڪb�Q	
�H�FD�P"�B#X(UHE#�8�.�K��f���ٹ'/{�n��
���N8'��u��;��ÒI���^�_s�5��ݚ�����c��wu��>]��Wj�>ع%����SG3@�wW�}='XfF��`Z��Q{��;8`��h�<�W:嗑ru8�TC9�;-��y{h6o���$��$R]�	-��rO��������0324���y��ȟj�xndO��@�����s@�����Z��&��s�㙠w��ܓ����?� �)*�� T�xG�A���s��I���훒Nz����ƔC�5&h[^��}V�m�������� �lB�|�M]�-�w$���`I#L��0'd�`d����|z�l�^���l��&g���y�Ƈ�4����ι��&���{��t;}��e"ڮ���L��0'd�`}2�����ݚ����5vX�X�����J�T�n�L�������?���^�$Wn!���{v`۳L:�U*o�݋ ��ŀ{����l�B�9n����.s�9��{?~������L̍0k�H"@�@�����\���7��T��ndO��@�[��wu��u�@��V���<X�mŋ!����˥����.�{]�4�8���ל:� ����������q��;��h�ـm�I*_�*I}a���, ��5�Q&6�prf�{���ڴu��w]���x�68�l�M��:����fF���̅w���v9R������`�ذ�n��?�w<����-]�8��;T�y`=K�^ɻVvoh�1��������QQ_�PP ?��*#���*+�TTW�EQQ_�EEE�*����
 ��"��1"�1��1b(��0 � Ȣ�0��EQ��U��U��TTW�*+EQQ^(����QQ_�EE�U�h���������U�U���d�Mg�Ѩ�f�A@��̟\��� �         P          �� 
P��H�*�     (
  ���   �@ 
  � )(��  h (   DɥO=}m���Ҿ�������ϯ���\ z��&��z���z���}{}��yU����{��z����WϾ���zӁ�@�R������2�]n��J��^۽o}�S��}����U> {� P  � 	(d w�V��zV���;������W� �*ͪS&���r��xکT�O���R�n�=i޻�@
{�k�j�Ǡ�N���T�(w;�
��(0 z�B�q�����b�ZJP � T   $����)�EU15AVZ�    7X =   �����  � @\�J�^�ԥU� 'w�� �=۽i\Z�j�R��g� w��ͽi\�U�璘�|��k���{U޽�ڻ׻�m޷*��u*�  �  (PQT� z��O����UL��k�t�� �z��vsO{:��-O��/*{� ��^�q��!��;� D{� �O�'�^^N�35=����[� ��������ɹ��nW�{��=� P  P)C4	窖}����ڽ�w�v�rj��
;)b�4�׭\�=��R� ��ϕ�t�������,��}n���=_l��S\����}�_}��>��e{n �=��ӛ}��}�z|��}/n��J� 4�Om)J���!O�P��R��  S��R��6��@dhتT4R�  S�	))P  !HI��"D 4f������O�K��ޱ������w	]��gr=���g��
��NF_� 
��PAS�Q_� 
��� Ee><=�_����n�)
6�y�6�om�����0DFh�|Hpf4�Ä�b��i	<M�hՖV�f�mj�~�m3���6"�k�����&vY�i��vh�Y�%&"H&!a�q�I �JJR�����^{��B�'-x�*�k������x~��0��Ƶ���,�c9"i	[�Fh��e��<�`��8�!��	���I�s[3��f��/0�=4i�K��@c�`IJc�6����^h�4捜ld��g Ѵ�=� @
H�>����ѷ����� �A�7���`�>�f��	##��w`F�o�����9���k9����1���g�y�7���Q<pRO��燕�9^Fy�����s���o��s8h��D��FA[�����#p'l��y��<�þk�#5����F:�cj7�x��s�������<�<�p#�`D�'C�	�h��LC,3��l�Q!Ν�H�[����}�F��#g�~ ���y�ƽ�����~xe���)$�$Æ�c1$��I�0��I��ۀp�0�o���៿~S&�8~�x��,��_�w羟�"<'c$.�)��:`K��6!�k� � �cI�F��b�x!!��u�)`�4��Lt��Jb�K)�#�(C	#N�q���G��ⓆQ�0~4�o��~֐���Ȱ�Nl�'�l�?~�q�u�'4���:�kcf�B;I�	��,��0��i8�p�Y�w{��o|��u�O�h!m%$�~$Y�uS��z8�kdof�F��DNBF9,�$��`BK`l�G��4��W�1ש`��.##@���#sF�ڲ��e8h60���,��"ʒb�b�[Rj4��%qM)�ė�fI 4)8����A�xlBV�dŀ�%�$F�� �Hlx�����ËN!&	.*��I��ڐ.) BH$.�Rt��ɏ(�T�CH����!
`�5*D8&�f�L]�58RpӴ��&��sH���x㭛�$�;B2�0�m&C��a�g����<��	 Ã8a�<���ͯh�a����\cG��tU�$h�����$f�a������a�`�t�b���᱌ѽ� �4�83���#)YXӰ�o�M��Hlx$8:v�����C�Ӂ��d�NÉ�
|,8l8��KfaD$�b�B�;X0��,c8�`�$��,b���ma��b6�y���������/�1,��� �F4��.�K!�2H�08���I���q4� cQF)�ɃfW5��p���c��ɑ��Ieq4��1H���6�F�'\1��I�Ӳ�`Y��5�! %�d&�A��3��<I�41�C�8��X�5:d#��6Hc�a�m1�#4a�͞�&���e���N,�K��m�X��H��	�;3#@I}�or�ĄB�R�
��V+�mp�N���K�B������.��.ϧ�[��;RÜ��ōPe��s���ʝ}��v���w�}:V,�&Wm��o��e��������	.*:�(�Z�.9��E
�v_Թ|�W+�Q�pn�r�Q�\�.ߩ���[�w�T�u˧VR���о%�ۮ�X�������Ԥw�u�z���\[��J�.D*�P��V��r͝�}+.�K{]v�c��er"R�uUK��;��<]ַ�M�Jbm'��٘������j��r�c��4h�sla�?F%�ȳ|y�s����NX~����^��B�$�5Q�SK�L���Ѿ�8���Qk�w�p����'�+�J�0`m��f��e���$�fg�a�cf��a�6��m�8h��:p�F:B��4�#bG�$�Uk�о�� "���~֯B9��|�L��A����I��@�IHW�]*@%�b�8��ɊA���ǚ1��@����<g�����NE��,(����3��x�a�|ef0M;��p8p�M��:��x��#��4�fX�zI�fF��f���86c�`q�Fs0���+��aa���k5�G�����<��4�oQ������q��A�j-���fNQD`鷳���ef��-�Da��N쭜$���F��l����u��I�ǁD`F&�;�����-T`i�tm�4�x����$�xo�ov�;��G���0��1лN"Fos���dɣ	���a�07&K�B"b����:���1 ă,��FH&bD� ���H�K8��f��N�d���9A1Q�͟��g��K/ۭl���OCs�l����w5�0�s'F�ѭkm�4;c#I��"	��	B!�bLq	��0*2pY&\5�����r��5kC�-a�a8�<�,�F�bA�g�f���+yf:�pߙ�D�(��Hǁ���N��1k?b! 
�_�!v3n�+�f���9�a�
�[4m�e��h��6h��F Y��)��a���#99���΃3�p���I68���a�<R0l'a�����l&�"o�7����<v_��	&���=�-���x~<`Ĝ1l��Ć���s���7�H������%�n+Ă ���5�d�N3�>N����L9���%5D/��A8��O�cI�%�~~���pӰ�20�HLt�p<x���o	�<"������p���"�����Df�t`F`�l֧5���Bj��`h��Y��Ff���ћK�WI�$�qăq�H�N	&8�BFhd�5��8qb	t�����w�l��LC�Ȋ,|%�[�h��/u�Fk{Č�Lf�A��0��h�	���e���VCF-������Z&6Y�H*��٧�ٚ��M�0`�L)M8�dq�6��|�a��Y�R����$�����%�<P��1p0���A�FqӇ�$H&'3����l�/�<���m'A!�)�x0�h1X0IaC��$�dӴ!�&L	�14�HLEpT��R�0G@�XG�0RFC�p�~:z�k�o~9������°��8xF� ��h�!#�1�h�lm�Zָ\�4y|�8aa�٥��G�5���ѳ�L4�A��ky�9�Z�~�}o�㭞z�N�+�$?:Y�4d�C��1�:M��#��%�A�3��h�xXmǌ'�A�-��٣��hg#Y�HÁf������޼5��<d�uc���6ج��*�HM�8�`C%��4B;U�V���"wt��ߟ����� [@ �$p6�       � �/�  �������q�G>4*��T8��KR`      � 5�:� m��cjݷ��8�� [F�[l9$���6��H�������&�۸��� �l 	� �	BE�A��7i6  � �   6�   ��j�  �6�@ � )i�����[��vV�0q��U�� ^����k�Ft�*�dZ�ڕm�Z��  -���l��[�w�Mg�]^�<i.���~Ā	  @ H6�@�i�Q�U�Md� �m\�n9�l���ԍ�a�i0� �^v�`-M\m�m $� $HmU���ձTUu@r�r�:5��s�m�F��P�  	e�b�d-��̎�A�m�b�)��`k;S�Y�i]�s��v)PBvX
�ڶ�W [%��s]�5id��e�j�ZU��ۅe\�U^��ڌ�� V�T�M�k{g<�z�K��Q� 6���%Y�۶����A˜����v�.�]���:.N���%Fƶ7��>�"�p�j����:9�U���m<Y8%`��-tWnڻnNsJ�V+�g�4��;�S��]�����ݶ���(��V�ضB��Q��8%UR^�6V9���hu�ƥ��aKsq	��ĈHL��Vթ
�WH���m��ڐ㍶rt��@  �^��m� �n�,;�l� �`�$H�������4���ᮝ�� Nk��Ͷ�&�ͳL[�K7lI�
��u�(˷2�U/,�UT��A�jC�6�mnf�@s�P��}��+� ��P  6��m���0�`  e��m����$��$�m  ��x6ͤ�l���]���d� $   H-6Ӎ���Z�^������v��  -���ר  !����$�#m��Kz��h��ݶ 	�I�fgT��\�u�����v�p@uj��۲} $	:5�&E���F��� ��x�ڗM50I��pls�$��]�;s+e�l��*=TG$8'6�v�kv���Y% �P����=� -��K�E�Sm�u�K�l]�0��%��Ͷŵ���� �a�Im���@ m������{6� Zi0� Um\���r�U�*��@ ӌ[�\� $F� 8   ��m�i;d� �  H8  �` h H-h��  	&��5�	 �$)@�l ���m�m�$�8$�` $�`    ����8l   ����:msm���� -�m& m��m� �� �m� ��m����  6�	��`   �m��o`��N�ǽ���x �i    �@m� �  � ��� H��,�%�l �� tQ�� �m�    �˦�  -�B��  �Hm�     � ��      �  �   ����.��h km���m�� [@�l6���   ��Y�  �i�N�.���Yx[J$$���v�6�	[@ H Mf�`  m��   �.�v��(j݀�; m 8�v�kn��v� �`�'F�� �I�8�*��[�V�ҮQ�iV@[Kh �� [$�  � ���m�$m��=d���7[jے�ٶ� 4W p�&�ٶ��.�� l]��p ��6�$6؛\�]oeUU�X�� �\ksr��e���km� ��  p��[` ր�G  v�I��d(�%�h��u���o%%ڠ�+²�x�V [e�6 ��i%f��.�b5��z�h�����&ٶ��`�BI�m�X�SH�:	�YnC � F� ��K*C�-�M� j�$�K��� Нr�$m&� `m��`�m���a�nۛl ඀#m�m&l�Ƶ�٤������9OǼ��� *�mr��	��@jeFA�� ���XAWl��n� ���m�K�V��ph �H�%��@ m�� 6ٶ�a��` m[:S]3���� � ���P$-� m��qm Ӏ	lm[�L�݂@8��9m�I���l��m� m�M���T�
�jڈ�\��m��0෵:l z�����-@J�v�2�Gl0�)�UP��1�+�5T�vg�i3��p�_�}}ĸf�;l�]�$ 퍨8�jI6rڳ����vi�H�6�l� �l� [�]6դ�M�>��6�`h8 �n�&��y��j�`��[���_F۰ �-��wh���rBM�S`���$���}�ٶ[�m Hpk�l�z��Y�%�@m� H�n�Sf=$��p�,[JP�*tI��mU�ӂDݮ87m���@�N;m�A6�! h6�8  �d��I�I�E��'������� Fհ�յ��[sm� N� $�H  ��$p��ݑԶ�M�� ��6� � �8   iV1!'-� ���m6u�P�9!��$�6ؽio$�\ �6�`H� kV�o^[N �o [@M*ۤ&մ��[F�7A�v�pM�  ������-�:��  Vגs� 
�$�9L�Mp�E b�EK��!���5+YI�bX8�lf���Cx,�U��p�V�=�-�ln����EH��8  [G�m��jժm�����@m���$��� δ��%\�m  m��=����k -���݇[��npm���Mm��[m� ���M�8ȵF`zz� ݵk��ym�2\t���5�[MU�H1���nb9MS3i�b@c�4��i*M��kd�@	7m��e�H 6�;�ox�ho�[m�I�C�Am�6�Ո��h� �f��I���Vy�kk���)̷+[v�L��H m@p�ְ -�� �gm  ݶ��lAm  ll-�&���%�  �'@�rXn���\ 	    H t�HHΛ]&�c� ]6 kn   	  -�   �  8� `� ��[j�UWi]V��l]UJ���j���@���d��7m��[%����oPӂM�$p���Ͷ  � �` $�� B�ؐ$-��m��$ �[M� j�Ç�� �� ���t�m��%��6� �I�  �  ��ְ��Io]8l �z�   @H $ -�  m� i�      �  	 	   8� #� mm��m��ێ$ )���UI@�U��E�9�`  @$ց�ŷ� ���p t����ְH��H�5��� @ m�ڤ�6�5��@	���ѶŽR  ���J ��8��.�$ l����  kX�ci�D�mڻ`���� �  �  8 �ͫ`m  �       m��$  ��6ض��h h ��� @ H -�l�x    8 8 m���e��Ԁp-�`�lӮ �M� �dmn�� p�g �`���l�»4���-UԹfZS`�`�mY���-�T۰   8  �@  �  �m 	      [`�@��p ��  �m� m��` p     �`�H    l "�  -����6�ݶ�l!�i;1�i��m�6�d-�,` �  q��u����!m[A� v��� hlհඒI�  ��KM����
��6NZ�v����Y�h,���mm[�lB�u�V� ��@UU*�V��[!���c�\,m]�P   -,���{nҭUUJ�V��4�h��;Si�n��گ99������l�ӡ]����m��o-�����yR mm�66KN� >��  ����l	n�N��u��	�m�2��2�-�
vk�n�)v�����@EM"*}�����O�`'������? � �mA8���Tt"�P�sj�`@�!�z�:�PS�(x��A���C�"'�.���ѵ�S�+���3b�>���p҉��8���G������â>����ԚO:�A.�=}WϘ����? x��ʃ+�/�w�/��Ӛ�CH��VP}U8�����}�+@�@ ~�ht~Q�U����E��z!q��b*�D�4�D�P'PM"	
)�>�( �I`���aaw�4	�8 �2B^!�LW m� l:�u��I^��TCb�����W�� �Wc\_ǡ�!�����=�z���=O���� �!W� _U_Ϣ'���\ 6�<i LW�P�C��#������*�t�t"��H�JN"��T�����' 4 �� h4�~{�⇠*�@�<���_��E� &�������
���}��S�eBI=Ͼַ��kZ��j���F%�s�pUUV�-�N�@�6�vP	]��� �����j֣���[!�д7�j�vv���ks��.8�(�+��Iѐ68��x֛�v�.w;����+ry�E�u�5;��k��icOU;��j�}T:]t��-g<2��b9�`	:����i�ʫ���\E؁�1,���Ї����q�
���`�ns�q�ٶA��.�Xrvv��f�n��[,��ru���gX�EqՊNb�<;�϶�
�]ʯf�����[dH[]-Kaƺ2 �mN�س;I��Q{X�\�+շm�Z4��R�R/)*�VҭUհ��8@;%�J�:5R�s�n� HK-��Su��v�W�1O��Y�j�j�9K�������Y�Ô]HU�lMU�Κ�ݶ�]<��U-2�ײ��rg7��#t� ������Qƶ{WK�R����흶U0�����!ً���K#��n95c����4�YҚ�6&[�X��R��JlR���q�7keM��3��C��W�k�Rt���<�٭�h*��L��W���;a�mO2���*�xv`'K�&�l4�SWDiM�̹�Z���kD��K�i6�5,b��w0�mM�Cq���@�������ͷn�Ar`���b^�I[n���}��[�83Չq��mc�E]�i���D�bA��)KQD��^RV�ݶG�*P�ہ�f��0�sk4ǔ��ٱ;7g^�AG�*�%���/+�-P�Z�[�vV��	U�0�0�j��4n�V�W5$�w�ḱ>��!6R�	b���*�u�m���|��l��t��:vg�2C�= �dz.v��Ӵ�;PJ�����
IU�l@2[@pk��$Ini�k.���X$9-�C:s�[	j&���䤍mrU��U+f�+<8�v&s�kh��m�X�9�&ow���=����(�(�4 ���x*��|]��o�@�����&�����ǻ��^�{8��v,u�c���閷����[NՖ�#�$�n���b�c�U��oCf{u�nPy���+)���
�5�Aډ�֑%G�ݎ��%���$��Sj�vݴE�o.�����Ѣ]M�Ko).]��ZG����nv��HA86�3�
T�.� p 6+���Jv"k�蠦X{fݠ:#��hPB N(� � pS�>s��ʻ�����\e��\���	��v�쏜��dT�I:C�7��U�&�{������~�����c�����j騢$N��M�f�tB��.Q	D+������`f�4�7v�6�N"����ݤG =q�@8͂�܊����	$�U��{����ـy�Ł�D(�n�`��;�,Yk)i�X�~}�@tqR���׺���MѿI$i��Ԥ�A�v��W%�n���[j�(\�ۇF�nP�h;.�3o0�۽�4@tqR����K@f�4���iGQ���(NU������)�(H�S�HbP��@��:��/��D-^w_��U�}�ۀwsn�c�ͨₔ�	(Rv���KfL�>ŀv��~���Z�d�:�&�7�M/�U$g��V��Ł�{���M���QDH�'�V`z�`	BI��0�78�������&�8�0q�s�����^$��>/]�Ӛ����(;Nl�:��m�ݬ�ͽ�@tqR�Ih�@tsK��V���$HI$r���V�-���X��YԔDEQ�ιL�د2�YV�*��2�0=x����;@�$PS�_t ﾮrn�Ձ�{���֨l��M�m�� :=��EH�%�:3a`j��iGJ&�$�HX��Ձ��Z�6�`�l�U���Zf�]�Fu�'S�����4��+����v���И����cLX�.�w�o��$��$�G�@6���2�H2P�H�qX����F{g�3�Ł�{���f�WME"t�J��X��0y�0�J*���8����3v�6�RPH��)��`s�4�9����]��ܯ���~/@تU��> 	��|��_��j�D�� �*HӅ�Ź����4�3��V�f��6�B�"i�1�I����u��>niZ�/jpqY+v�`��3��'󾯾$����Իur(�N8���~,�M,��?��:��v��5Dd���6��p��T��6\s��YT]�Q����(NU����9�q�Z�2fJ���JRR����|��5���;�u`gsn�u�tN�(N�Cr;��s�rP���� ��,��u�b�
�.�U�Ug(���I�M��$M��#�
;r��F�];��ī�.G�g�]M��gj�k��Gjz!�M�;Hk��v2��bP��mrB����s��i�_ ��:�P�u�7�ڧ��*&:�V�'���t��<܏J<��}��{to�o����k���p�:�o1�9��:�g8��kb��B�ӲSls��Ah�vΎA`lR�;m���>������{��oy6�d����3v���扳�t��h��(�;fm��@v��Bu�N�pIrD��$J	ŀ{��;�u`qnk���ǚ���-�Ԕ))�q8X�T���18�- ��H<��RR��q'�`qnk�7��V�@{�� Nr���Z�V-6̬���̟Z��@z㘀�{�P�Jn&ȉH��M,wf�w]�Ώ5X��<���U :R4E�]p��܌qP:�ZN+"\���b�6�6[��$�"8��4�IBr�s�Ł���`s��V{�u`w^����Ҕ��,��U�~�uηOG�&bB	��ਏ�b|�?�� k�i�uX�<X�۫�xֱ:�d��l��@N1�@z=�����Vf�t�Q�*H������3W�����������=�r��($RS��p�3��V�����|�=�3�4�1i��u"�$ND�����è-�u���fz�.��1��<u�K�	��JT�n"D�r�-�vnK�� :8� Nr���V��x�p��˯�>e�%�G���7�b�?K�X�״6Jn'RQ)D8XܚX��˩�@����@U|@�W�;7	���y�DGJ6�R� :8��b�l���x�Ҏ7JR��D��`qnk�;�M���"�U�^��nf���Lv�U5�ڤ"�rX��Tv��Lgf�X	���A��r���vw	���ɥ��٥�Ź����tԌDqʒMU�f��ft%'o_���I��ꪯ�H��-���')8�,����}�Zs6�*@z=��s3j��5awWuk�"!BR��� v��*��{Õ��I���.���W�S���`w1I_�j�u#cR. ������?����� ץ�{t�Lv��	Sg2��څR�H�8��*F�C���ˣs��[����F�T�����3`����m���T�r��m��諭����+}��`wsn�c���q�R��n�y��}�Z�lT�������Z��A��r�DqX�M,�*@zM��Ihre������R6��`wsn�}�}���7�����G%
"u�QWuS!Jn�y�u�=K�,�a���N���Ä	�8���m������`7Lۇ���{b^]���q��c�����T���b� vœc������:u秙�q�xe5���]����s�et�vI�T���{�4c�l͹�:I����l`��@ݐ��ŴR����U�q7U.;�t6��Px�C6G]P�m����ϫ#����������ww~���y�ì8v�S-f�b�;,v,3���b�Zݍmvv�c&�8��t�'Q�n7+@��X׺��K��u`sr*�R�H'(�D��}�Zs6�`��6	ói+�Իj�FƤ\٤�`wsn��U_|���Ł���`s���Sq:����f��*@tqR�Ih%\�n�u��Q(�HH'��u`r������|`{l�6W�K��NcC�D�����3.��H��(`�6kL�7�c��՛uuis�$�Ss�k�ـy�!/�ϱ`/W��"d�ܩVnKu]����D+����{l��� �Ss�7�r���'��H���K{�K:�U���i`f��8��r���:l�K@Nf���܊�D��R	����Xך�f�f�� ��ŀr�ސR�e*���+�k15i]Dv�=S��vd�.D�۱BjFD)���ں��n.���S�`z=������@G�%��f��]��f�G�@sqR�9h9SK��֢8�Q�HRs6������r���3��F���ݦ�ʄ*�'3B���2�ѼP��N
9G��8��$$q�:�����ٻ�vC�c�I�7�s�v3���q���Wa��B��3 D4 @hy�x���@4��h0G6��F�4���ۚP�E�Ex�iH�D?Ҡo\��~�

y��~��<Q̿w��9J8�)m�'*Õ_U}�-ɾV��o��<���w���U�A�{߼9Vj=JB&J�ʓ�_W�5.� �����B�%BK����
"g[�X�}=
?H|�$��U)�Qj�樻*ɢ��і��3[���֮����c��+v_߽���r�b��"��Jp�>������3w�V������Q���`��L��U`\l�R�������~����~V��?w&�����f~�_�R�H��Gp�9��N �����w���� �S��)�uwm]H�9 �|��M,/?w}�Z?(��Gj�:��ρ���V{�z�y��%6��Ȭ�`���q|x���w�+�t~��e���=v�̋�D��Y�Cs�m�C��ruk8��nҲF��Z'X���`�}�Z�c������n��6��`g^�${�V{g�;�u`qw��"d��$EU����O�7�b�7��`�np��騢��"�Ƅ�;��V;6�%�=�9h�J2�@��#����wf����.��X�۫�V��B�I��qJi��s�}3�����Xr&H�9�E�{uV�6���Bss�츙�r�2<��Q"V%�cd1neN7K͠���'T���S,)N���e�!�Z����=/K��a�,�p�t�l~�w�{U��<B��6]�ȳ���6���H��Zt�s-�$�j��tЩ�P#�l�@z*L�G@����vݷ>5��6�&�ǻ���]�����7Y�&���vu�q�������,���y�]��~�>7���!u�6��6����1�@t{�l��6����m]E�\�=�;�4�9ݚX׺���h���l����m���@>�-�1�@u��GJ9 �AHX��,��V:<�`wri`w�69J8�)m�f�}�Z�c����t� ?��ô��S�R�u=<��Z�٦J;N�mƛp��sh��]V-��:��\Mh0��@{�r�� ��_ʯ��XG�yX�x�%(��)hN+��K��PS� .�w}��*��}�r���j�34��"	#��p�3��H�%�~U]�1�@>{�{r��J�#r5�ʰ3�uX�M,�M,�mՁ�x��J~��m]$�\�/��m���X���脣c�������Z���eۣuN-�t5G2�V���[nyB7;;�֨�N�eգ����?�� :8� �$��� =_Wٓ[�#�%�R��8��Ł�bs6�`���76�ss*��n檭`��^��<�D+!!T-IDF%Q��=�vـo�ŀݩjj�*FI))��Y4�3�4�3sn�.� ��%�NI#�4HX��0��������^���������s�Y�����S�7��n�oI��yE�+��A��F�,�ͫ��<�|���1 �6�4�5f:��R�H�C��r�.��l�`����r���V��v�����o���T����8�5J%9MI*'>hp�;��X��X��u��U	BJ�֘��5�DqD�p�T�`wsn�.��� ;�T��K"�M�ۭ3j��f���3h��t�%�\:$ikD��Ђ��t$�"9(D��G*����3p� ;�T�����ʼ����3v����� ;�T����9���GVm�C���H�Mw6�����9�)����ͻ�w3s6�o6�8��b�{��nm����FԩR7�9������`�q�HU?#��F��ٝ4�e�OOe15\p'{��t�l��
�y����Kl�w�Tג��l���z���б1�{�m�p�c.Gw9��z�e�-ِr�
�ۧ:ы����Ǳ���<��^�%�Z�U[���K�<�k�0�t�=��m��L@�,f%�Y�N��-k�U�h{�ݟ���e�-�����!{9�笖_�����}�	��!����c����:�Y�7G%u�VJݳJvр�\��*���]]ۺu$n?������ν�� =q�@z㗴mf�^���o�Y� =������ f���d��#�%�R	�����X�� ��@>{�l�ڽ�̫�.�mUլ�"���`��0��0�۫ �c[Iԃ%H�%
G`f�� =�� =q�@J��D����7i�@	V�;ba�-���&�-�Ѥ���v��U٣����|�T���1 �=����"��wUuV����5�ŕ��!A~P����5�*�"���6�`�<�M��ͭ����Ӆ�Ź����M,�R[�<X͞,R՛D�uwn�JBD��ʛ���{�@>�- y˔mf�Qȣ�%'��K{�K:�U����X��U S�#D��%J�-��U�XV#��Yf�V[v6\�����v᪂8�Q�B8X���~8��+{Y4�9�4�9ݛ$�n�qG���s��)��;� �;� ~�f w1�cR��#����M,=�a0�CQR��D%w5��}M���C����$q�JB�����q�H�%���@t��r�Ͳ�w3s6�ot@N{����ۓK ·tIFH�I#��r��'*�]
�Hs��2f�C�1��<u�K���n�#qTi��ν�`ori`wri`ori`r���'뫻jȤ$�.���?�L����;]�o��Ι>�E�)�%H��,���&�}_���ߕ��}?{��E��Q�G�m�����m�p�|�G�jaB��N!%)DDo���~��7~���7WUJ8��B�ν�`z���~8{g�{�K�5�TN�r4Ƞ�P�M�gX$�֤�Yr+p��ɇ^n[r$ �^��{,�����#��{6x�;�4�7�l�"GнAξ�p���Uڙ��������0=�gЗ�Q�wذu�Ӏf���UI�FרnRU$q�N)��X���9B�|�y��]l��*T����#�a���nOyX�0=�`r��|���<���/�fVP]�Uws����>�J7�q�ϱe^��{���&S���е��%LSN�@�D`z�Bo���!0��`I3�=�o :7 
� ڰdP�E�'���� e�LSnC�?c�p8)	*���&H�HBI�K+F2�0"i�0@�~Q��f |#IHOV�S�F ��!$B �v��oww;������?łeZ��B��U^�l  t�\��&qΨ��>YVڠ*VVR�@e�66LCl��e�"tR��k8c��kI�_:3�+��r�[l�Y .�J�+q�9$�y�	A�䷬�P-��m'Oig�B�Ӗn7bٝnq����]<��ZM��OB흓P)л�7�٦���r�^X-�^w�L�]�X�n��K�q��;�� :
$s++J�>%���ˮ@�.����c�"c.��5�;Ɯ��[e2fX5�}�|:����iA�'R�\;�[@��m�Q+j���]���������TDh�^g�����ڤ�sR���jQ����vm�XuM �tST����j��,`�����Ry ���^1�U�@�f~_��c�[k�KnT�r̭[u�5U[�t��#�=�+���6v�(�P��C3ԛ�z8�s۷t�%ݶ6�z@�/Kq� ��G2�G\��.�TA��z�n�n�@Gm�E65d.�e�	��*���ў�^%�]��������*=v�P��g&v�u�x�P��8��P�'HⅶjtM��f��!��u�٩v�nl�Σ��6����٪W�EY\�V	��]�)C#OA �;�����%ъ�
A����/d5(v�s��.�z��v�e�[l*Vç���N���$�w�ݒ/�uY��ڹÎ^ ���E|�/=w\n�h*�*
��J�}�Py6v�����&M��N��,�٭����eZ��i�uѠ�<��l����ee`�C�Uvz�V�+V������񀥵 c���I�t�=RN�aܖ�b��G����1a���gn��`m�ܒG5�7��At�ݓd90W =UL�jK�秪�4�;}|������A�lc��[x%�A��6�{��J�vʵ�Uԩ�k��[�9�G>����k[�V�b��I`22�a��6)n��v�=&�h�͂u� /C���z
� �OȾ��>�;�{���߅��Wh��YS���qd�zb�1�c)�v�X���L��Ssjn	�6�*L�n��WY�;,��V�<��1O����}�v����d�n���͉�B/,-�Ƴћ��9��/[O�oi��W2C�=�G"���8v��!�g��b�N#y���d�t�x�o0PERt $V���j�m�6Z�D05v�:��Mk���SFܟ�����s�}���wj�V�eXҴˬ�Y��23Ȧ��g�9�s�ww�����Z��F8��� ׯ���G����1{����@�Ĝ,�۫����ԒJ��_}8}��y�9B��=��q�9(�q7�����`orig����7��?���X;��5#U*)RJ*�p:!Ok�0s�0�`rJ^��5{}%JJ7$�Fڐ�9�4�:|����}8��`;::`+���Hz�Y��U1
'B\�%N�%�$N�$t[x[I���)�e�:�[����>�*@>�- �� =� yʛ��*T�ԧ)��Xך��N�US�VDDB��a�ߌ��0z�g�
"d�/-�����ӄ�q��=���`sri`f��Xך�sV���r�5f�� ׯ��s��(J%�W��:�(�rG��7�4�c����G�@u�fV`eJ����z	t������n�m�(�#�LJY9W����vR�5R�fk}��~���?m� ����	~��w� ku=EL�T��I�V�&�w&��&�u��U}������"NHIj��7��?m�&�(^�����X;�K��5�7)*m6�8�,=�/d_��؀��:����>�731ʕ#d�*4�`w�s���K{�K������F�����i�)'GMG�{t\�8H�l'K%��G�%��M��wo�|�� :=�s�Xך���h�Rn5 ��,G�@N{�r�����7L�qD��B��ͺ�8���ܚX�M,u���$��m9N�r�?}I(�V�V ������G(�"UG���*���Հfk<Ƥj�E ���@8�����O�ʐ����~tE�Rn]Act��̃�n��g��[(ؕ	Ѷu�+n�ʸ��n��{�*@z�L@8�t����IT�F�8�,�۫�}���|�՞�7�<X�M,;���ܩR^Vᵛ�����1 �� =�vM,-U�D�uwn��A���ǾV�@8��9�	nd�sj�7���Vw&������7��u�p	X�t%	"$�_D��U�lj�mL���%����e�#�<su�[��|��}eW�{r�2�u�3�۶	��Ns���Ӳ��[T�C�.z��mˣ�WLp�����6��A�!6��J�v�,n�V�j�%�9��i[��'C3mT��a᎖Bm�����fV��*]��s�����牉RXI5�m��Glsb0�C����O[[74Gw�޽��w�y�=��\,sӞ�D�����J�Sՠ��Xԫ:���p�����:�(�j@�r�]X�npu��T��X?��0u��u$�6F۔�G*�ν������7�|��|`��ϔ$�ON�:�f��Z��8��X�V7&�z�ꤽ�<X�|�[�Ѳ!D�$Q�a���O��k�0�k�����ӀwZ���J�R5*AHX��V�����O�S��?=�`��j��]��d��Gg�]a9���[c�T[��p�W�ԟ��ӡY?UU}iն�wR�N�%:���u�N������ ��,�ҟ�
�G!*AH���W>�u_���=���7�b�7�������{��V���T� m�`o�OŁ��ug�-��+|����ɭ���%r�!a��|��}�s���^�0>�P�T������F�$l��Q��X׺��M,�M,�M,�TF���	��G��g-nl�����8�n\l�wl���Z5�s�[��4���E �M��=�<XܚXܚX׺����P�B��7��0=�g�L�����t��lϒ3Z���J�R���,f�z��-d�*��`]� ?5�UU[R�N�%8܅��{�����������R�m��;�������%H7��|�� :=�� d����o�]���֙��k�eۣpҧl��{6I�&��y$i8�l�Qn�p�:kdl���T�}�_���y-���F���976��ν�`f����������6f�ߤh�F�ە�H�~��ǰ@t{�*@�n����E#�qXy}[���
R{�u�<��=���)А1D��d.s��F"�w]"�䛛�������"D ���D �Z���)JOg{��JS����R������{������0�Y�3m���p7��F+�\�n��W�k�J�{�`��uo�-��6��]���x�A�}�!/9nG���{��R�����k�JR񭪪�j��Һ-U�]��!/9nS��C%>���┥'{��^JR��lȅ򈉘���)��ŕuvZ���kx>JR�����)=����R���wۊR�����%)O3���o.J��*��*j̈A�%$&��#�J}�w��)JO������{��T{M������.�����"D���qJR��s���)����)=����R��2o����;j�^C0"��Ik�&�F'=�ZY��1.V�m���&��ft�����
r8(���D�+FE��Vs���AV��pQڮ�s�����z��v��g��2]��D�\H���:��x�]rbcV���U]�]q��K��g��u�ԑ�!8�O4lA�탈+Mf�l4�1���&��`U��R�8��������(��B~�/I�ʪ��Ң�"J�Xݳ&��,�N�cP�۵�Ol��l@Y�۫��cX�9����'�t�w��>���)����)=�����J�!v��"D �����n�U�����ַ��JS���n)JR{�{��<�)O�����)I����<��=���r!E$���R��}A�wq�_\�)�����$���<��>�|dB�������ʻ�Sv�I����'���\R�����<��O�lȄ!y�1F"�i�T�l٭��ټ�n┥'�����R�����>��)I����y)J{�{Ì �A�
:[�)Z�W2]]MW5�p��ž�Mbd����^��[�v�Md�����f;_���YWUj��U�\��!B����2!B���u�y)Jw����)JOg{��!B��f����Uݪ��U5fD �D���#?(G�s#��T� ���y)�<���);���JS	�m��(��@�X�K������*K����)�����)=���$?�����?����)JRw��C�JS�{�4G#Dmʌ�B����>���C�JS���n)JR~��<����H��y�D �@�G�S7w*���VIk[��)����(��~�JS�{��)JR{�;�JR�~��qg9&n�b��J�7I+�b��Ł����ػi�9B������﫳F3UwWtTݟ�D ���D �Z���)JOg{���� ~��>���!/���W$���.�sv(�JS���R����w�<��=���)JO��]���ȉ��KߗUT�|�U�+��+���"B�?})�)�}�n)L��7O��A��8�,x)shn1�1!��چ����gm8Fp�X������
���JL�"7WЄH%zĄ�Gx��o����E�� @�D6�:�@��P��*�� z('b� �/�#������?~�A�����<��=��p��粇�3���jի����Q��A�Ea>�����)=���JR����┥'�����)���٬ލ���Y��R����u�y)@|�3߻���);�}�%�2S�w�!&wt�I%�*WWT]Ң�ɚ�y�U�XV#�����dc&���'bRw��{���DqD�ND����}��V�}u}@�'�����)�}�n����H����Q�B�����亻�.��]"�g�)=���%)O{��qJR��}�a�)�}�)�9�P�w�j��xl�o5�j,��y)Jw���R����$?�c%;�~��)JN���_Y��}]U��bۑ��5!%)I����R������)=���%(3h���;qJR���֦�����jJ���a�!k׋"BR{�;�JR����┥'���Ǿ��m�v�n�~~X�yi�zV�n%�u�H��5,�tE;�.��\�,d�_7}(��ky�f�ֵ��)JN��}��JS����R����u�y)J{�{ÊR��~���[�淚ٽ�5��o�JS�w\R�����k�JS���R�^rܨ�!Bs�BsjmT�+���u��R�����y)J{�{ÊR��[�D �Z�ّ"B�K���oY��3,޵���	߻���)=�>������}��)I��הB����K������.�dB�	�����R�����)=����R������)8��G����ޖ��5�I�W#���Wsch8�]0 �5Ҏ���˂i����Ԉ�:$5�&��^��if+.![h� Bq?�͔�x\$��SZm!�3��1I��2ɠ�z�:ɻז8$.�`��"c'\W;zwNdr�m1m�H�w�X;2�#Դ�وw۲ěL.��4c�v�pP!P)-;���T���u�lw�n�����O| �I��A=��n)�ױ�n�=X�NZ�F�=�hں�x;;⣮�I;w�7��{����ߛ�%)I��ג�����8�)I��ܨ�!B��n�w$�UwWtTݙR�����y)J{�{ÊR�����%)O{�{�R��ｵ���o3-�5��fo[^JR����┥'��{��JS�����)=����R���;�j�B�iZ�5Uk"D ��-�y)J{�{�┥'���^JR��׋"D �Ǵ��3U�Z�u7ur���)ߵ߳�R�����y)J{�{ÊR�����%)O=�[��Z6fl�Hj�ա�&�����4���8C���ܼ!N�rON�e������'���^JR����┥'��{�Ʉ]k��A���r]\�������o[^JR�������~!|G�%)7���<��>��qJP>�fl��>���{�[��A�$Q�┥'����)�u�s�R���]�a�!kי�!�s�蛻�f�fkz5��%*��ݨ���/��j!2�r����]]��䒵��Zݛ��R��{�v���=���)<�=�%)O{�{�R������q�?�:N�u+���2���V�@vPckt��5��mux4hH�.�,�xfok�)߻�8�)I��py)J{�{�┥'��ݯ%)K��;�Y�o+[�6f���JR��s���R������)JO=��^JR����S!nˤ}�^,���vQwW*?"�]�8�)I��k�	�B�:	�B���"�"WP4 >�J{����);�:�F"���WEMҺ
�*�r!��{�v���=���)JO=�{��J�%�����)JOn�~3z�k3z���Q��ג�����8�)G�?����JS�k�g�)<���y(_iT|W�c�I�#�H��V-��<��-;%
��M����F��^���Uc]]ԗWw7@]ZȄ!~��*0�@��׽�)JRy�������)O����"(匿�&����M�5wJ0�T��׽��NJR{��my)Jw��Á���'��~��)�{��[�kv̵�oz�����R����{��)�}�)O�@d�������~�~�)JRw����ַ��k5��3{^JW�	�����)?w;�%)N�׽�)B~PM4��:�'u�^JDB7�;�j�B�iZ�S7fD �A����)�����)JO=��^JS	�m��!&{i�蛻Wsw6U�vkê�$RN!�$�����*�n[�Ȝ�;��]�U�Z�)ur��B���r �)<��vJR����p?ė%*쾕D �^�u+���St��W%U��)<���y�!�O����R������<��;�^�8��b�?�w�7��7���df���)߻�)JRy�w�<��=��qJR����k�!B��ڧ%��Iuwstլ�A�2O�����JS�k�g�)<���y)A�K߻���({�w_j��ݳy�5��o����׽�)JRy���R������)<�=�%)M���@����%pD6ण��w��[E��+U�en��Ӹ��%؃q'lY��sk@�sR=����$�c���H�a���ԝ�.u���U�]��cf�Un�\�Yْ��=�Ӟ.m���f�[�u�t�>��n�Y�,\�����_Jq���-u]e�հl܄:���c���m����#i� �"�#�G�H���r��(�6V�8ێ�kt6���q���﮺u��[4ܺ1A�����`���=����R9�m�q�)]۾����,�-���'�I������=���)JO����]k��A���4U\���Y�޵���R���wۀ�����);����<��?�����R�����y'��~>ެַ��捛5���R������JR���{�R�����k�B���̈A���M�ʹ�Wv���[��R��������)JRw�}��)����?��Lԝ����#�	���ں*n��5rU\�B���{ݯ%)N��}��)I������A��\�B�����Sjfn՞�s�v�Z�Ȕ+Es�z���gAmΗqo���G�H�X���[�������qJR��s���)�������b(�A��#�]uW�]]ԗ5wkn���R�����py��t��;�w�┥'{�v���;����/���߿��\Tu�p�#﷽�y=���┥'���^H 1�����qJR�߳�y)J{���ou�����[�kzַ��R�)I���ג��}�\R�����py)A����|dB�����*�L��&�ꪦ�#JS���n)JQ�Ͽg�`�)J{�w��)JO}�v���:#���f���u�5��^glv�W��;h*<G8+��#<b�;@�7_���1]����v�JO~Ͼ��)��n)JR{�{��!B��ő"Bg�l�|��n�ݢ���%)O��\�rR����ג�����8�)I���py'�90�c�mU���-M�Lՙ�!'�ּ��?{�xqJx(�)�� �@h�߳��<��=���qJa/�];SusS7SVM�\F>�A�{���)=�;�%)O=��qJP��HO{�#�ӳ�%��IsV��ռ��)JR~�{�JR����qJR����ג������R����r���:���v����i�Yڴ�b�\l�q��[X͒�ٿ�o���G]�ox>JR����qJR����ג��ۯD �A�uʌ"D/J���E]���������"D ��n�0_G�0�Jw￸qJR�����%)O=��s����������VU��{�J~���┥'�����)��_�!'���B�{ڝ�5W![��f���R��`�=�;�%)O��\R����{��������<~OA�mk�8�)I��=����s[��ٽ��x>JR������)G����mJR����R�����p�����������a��3k��t�F�Y��U��]��un�8���2�������6f�fkw�)=����R�����)JO����[�JS�~��������������WC{�o{�������D�������JR������)I��גJ~�s�޷�F�[7���޶qJR�߳�y)Jy�wۊS�(�I���ג����bȄ?NӢn�U��UWJf�T`����>��)I���ג���}�)B�d���}��JS�;ߪ�U�&nj�����"D ����a�O���R�����py)Jy�wۊR��� x�*�⁤�@h�����1����Ycz �hD���h};p_BLK(�%�ql��I@�BH �&�  �*��8�d��Ӡ�1D�L�F!����,2��XǉhU�(�X�H�*�q�-a�Pd6beCff{�F���0ɳ�{���x2L~6H��I��h �$�,��,+`��f�!�$���Fd��"!�&H$��Y$4/��H��z*����I$�@�,%��������v?_�~����M*�*���6M� �fѳ���5�5�3 ��Q̥��T�R���A6.�e1���m ֮ݖYWj����GkH�����g3X*�.4�����1�7ZVxz^s�=
�q�[�{ۮ�����m��`(�ͥ��ݸ�eV���	�s�Gm�mh�*�ۇF���M˸�4�3V�/d�RT�K�'��P�
���9T���V�η�/3��4IV�X�t���Jj�ڹU�H�I��Fu�-vy0 �d����Q��	ͣj��,KN� !ĪV����B���e�m��㍫�Y��Y��m2� ۳�c��v����u]CU��Ԓ[s��(ڒ�m���G*���a����K��Y�d&���n�����<P:6]�I}m��lb��������Q��GFu��vy�Xc���(鋸2��}-�f�2۷o;J�'^�zь�D�k��/I��uEwF��\gq��;�r��@G*-�ՆR��A����8�6���h�E����hLt�p��+hu�q��\[)��{�\����7At�:2�*����c��qZ�Jaz	^c�J��`Ƶ�=h�
��
I����jq���l�踲�ΐhꭳ�k����T�����)m�n���ҩ�֚��0�@N�A��[M��Y����']/Sѫ&0eݣn\�P�UF��H�2i��RP�粋���nJ���1��.��@NZ{iG&7,n\�cD��c��K=v�"743e�R�>uO6TUۍ�*��k�ul�j�Ӗ��(�E���45+lhM��\�=R��sR�0k�
 F݈���EJ� J�T-��Ԅ�����u�,A�ӣh�]�ƭ����{g�)��J�Q,�	n��o[R ƻ m�w^m�깶A���:�CC�l8��T�o`9�k��N���֎�v-�n3uǌ�>��QԒ�W(E�][���y�Eҡ�C���W��^ʏ㊊~AG���
�x����^��˺�k#5k3��VYԎݮ��I������c*)w;5�շ@8�`L<�E�B�]q��5r����������z�S�����뚕$��ژ�&��n֋�)N���\u-b-��]j^�Ix�W.C:B� ����Yj��=�a�ƽzf�6���b�]�Y��yS��;G*��Z�&G���';B�բMm��F�8!� �c^��n��mg$��:3iٺ��AVֹ��t�o1�*G=��D'����wf#��pu]��5��R���}ÊR�����y)J{�{��|�	.JRw�}��(y��j�B�n�V��dB��۱�)�u�s�R�����y)J{�{Ê�*�Ҕ��p�_����ѽ�o5��)�����)JR{�{��)�}�)JR~�{��)�u�k�l��f�n�{�ַ�R��Q2N�ﶼ��;�~��)JO��v<���I(DC�}9�!/�t��&�����my)J{�{ÊR�����R������)JN���y)Jz��uΪ�y2�g���fMV(r�Y�0u]�L�#������{���|Y躛����)JO���JR��^�8�)P��qD �Z��Ȅ?NӢn��͚��f���)�u�s�x�J�H@�z�~]>JR}��my)J{�~��)JO��v<��R��w*�]�&nj�����Ȅ!7�q��=���)�H�߾�c�JT��ND �A�KrV�.�W3u5��)�}�)JR~�{��)�s�.�I	���!B<�u�5��k{����oz��)JO��v<��>'�o�g�);߾��R��������ow�����n�����v���ş7#ty*���\Mwd��A��A˳uD����[JR��^�8�)I���k�JS�����R�����c�H�[�t��ګU6U����\�B����ב�!!����p┥'�w�(�	ϵ�D/��B[��WJn��nj�of�[^JR�{߸qJR��{ݏ$0�R��(��8l�O{���)JRy�{��)�{��-�{�o7��ff���R�)���;�����)�����)JR{�{��)�}�)L ��R��ܫW6����ڌ"D-z���)JO}�v���=���)H��ݨ�!B���S�U��WUsh�˵��)u��5�,TsL������nm��gkV��wh���WWSWs�"B�n�0��=���)JO��v�^JR��]�r!BZ��Iwh��n��#JS���R���}�ǒ���׽�)JRw��i�%	�`�%	BP*8BP�%	Bk0J��(H��(J��~�?��5�e��[3[5��g�	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP���p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bw�����(J��"��(J3�)?�r��J��(Mf	BP�%	����	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'��xy��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%(^���Ww3e�ʲn�(@��	(O3�(J��J��(L���(J!(J��;���y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�����(J��0J��(H��(J���(J��"��(J�w�<��(J!(J��30J��(H��(J�<�������P��%	BP�'��p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bw��f��٭����f���o<�J��(H��(J���(J��"��(J3�(J����ǂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	߻���	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP�{��8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP��}�<�J��(H��(J���(J��"��(J3�(J���������e�L��uv��-��mk���݅���ԓf�y�-�?\�-���-k���{�J��?f	BP�%	�%	BP��%	BP�$BP�%	B}�����	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP��߸pJ��(O3�(J��J��(L���(J!(J��;���y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�~���(J��0J��(H��(J���(J��"���
�����[�G �
AJI7+����(J!(J��30J��(H��(J���(J��=��p��%	BP�f	O�,�	BP�	BP�%	��(J��"��(J�����x%	BP�$BP�%	Bf`�%'�d�J!(J��5�%	BP�'�����(J��<���(J!(J��30J��(H��(J�����<��(J!(J��30J��(H��(J���(J��>�n�>3{�7�5�跽���(J��(J��"��(J3�(J��J��(N����x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	Bw߾��(J��<���(J!(J��30J��(H��(J�������(J��J��(L���(J!(J��30J��(O~��8%	BP�'��P�%	BD%	BP�&f	BP�%	���
([\w)�]�&nf�����y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�~���(J��0J��(H��(J���(J��"��(J�w�<��(J!(J��30J��(H��(J���(J��=��p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bw�����(J��"��(J3�(J��J��(L�� P�B̮�
�D�v��&�j�P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	߻���	BP�%	�%	BP��%	BP�$BP�%	Bf`�����%	�￸pJ��(OقP�%	BD%	BP�&f	BP�%	�%	BP�o����(J��"��(J3�(J��J��(L���(J���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�$�z���n����=�w���S*#,���z���o&�a/\h�;wm�n�+j5E��z���&�p���V�`1M1ƹz\��d�j�5F�Iѳ^Cb��cga�Ӝ�g,�=;��nu<ta��f�w4Y��B�N��v=��Bb�7uSn��c������sp�c[&r[��v�&�2p�R�Q ��M�l��cEr�VY�[L���T=���ƺ�vw�}���߭�_�ցu�.%�A����g`X��U��WBS���*ێcKa�zC��GLm��������P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B{�~��(J��0J��(J��(J3�(J��(J��;���y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP���pJ�����OقP�%	BP�%	BP��%	BP�%	BP�%	����x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'�G�V���v[5���k|��(J��(J��(J��(L���(J��(J������P�%	BP��K��%	��(J��(J��(L���(J��p��%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�'��xy��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP��߹�(J��<���(JT�(J��30J��(J��"��������)�jpM��W��P�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	�~���(J��0J��(J��(J3�(J��(J��;�~���(J��(J��(L����Q�~��y�~�~��>~�3�f�՚լ��؃�h���(J��(J�w�<��(J��(J���(J��(J��(L���(J߻�8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	߷߳��(J��(J��30J��(J��(J3�(J��}ÂP�%	By�%	BP�%	BP�%	��P�%	BP�$W��}]z�ȎTu �$���W�BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	��}�	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bw�����(J��(J��(L������!(N��]]}A_P}\�N�M�AGBvz����\�ub�i�)�g����FZ�6"�ټ٭eY��!(O{�{������c�J�������%'����(@�9_}�Eݢf�i]]M]�(@�����cȰU �������)?w���R������?�?�WZP!>'�*�&n�VM���a�!w��ÊR�����y)J{�{�┥B�n�0�A��ӻ&��U��*�]՜R��A �=��<��;���qJR��{ݯ%)O{�xqJR��n�5ws*��sV��]k��A	G�#=��m|��;�~��)JO6�F"���"��jT���P[.����k�ѫ�юU9��7ll��w&�[	6��M�auu55s�"B�n�0�T����8�)I��������;��r!B[��M�tM�U�r\��rR������)?w���R������)JO}�v���O�R��O}%ի�eZ.�T�ZȄ!?���d�)�u�s�S���z�< �
xI�~���)���ÊR�>_��]ܫW6��QWV��%���ND�'�w�%)O{�xqJ�,�����!B�M�V��D��Օs5w8�)I��ݯ%(��߼8�)���F"��9�!-r�ŒQ�.�Et�Nn�[� m�A�kM�S�[!z��N^��=�F�lvk���{�)�}�)JRw��c�JS�����\�������)~�����j�k{����oz��)JN���yb)ߵ߳�R��}߶���=���>D�iJO�}���{�f��5f�<��>�����)JN���y)J{�{ÊR�����y)J]�ܻf�l�n��{ٚ��R��d���my)Jw��ÊR�����y)A�M��<6�������)<��|f�oVo5���o,�ג�����8�)G�Ͽ}���JS�k�g�)=�����a�l����+EM���<��$��ՒX��b�+l��
�ָ�m�)c9�3�k�w�y����8�x�#��ذƝ�$��E)�N�%���U���u`f�ŀy���(�䒊������n����YW3Ws�w}�,^�X|�I)���7��Vq���JICpQ�*��DDK��� ���]78D���`�]vMQh���U���X�y�r��G}����ŀk׋ �(I����<��4"��{澋Y��Z���Xf�o!����۬�qi�l�����h������j�\6��!uF�`nޏ[�ܘO=���jx,���ۅQ(i뗹g8n��n��jN0ļ���$����l<Us^�Ɔ�b-Ga	�X�ca�����Һ��c!�A�a��ʐ6��P�)���;Nh�0�Pq��4�5����Q�%����������N��,�$�
H�������=�U�a����:�2��&��n.��7�u�p��`���%�C{�0����V�l���WUs�n��>IDDD���,{�0u�s舉�v�W)�#Mʐ"r�������݁��U���u`s^���Tu	lr��y�k�s�7�DD)|���w"H�TR����3^j�7sn��۫w6��M�Q���N7)2'Q�A����Ŋn����Ύ2Q���k�h������7c�RTJ$��NE�=��Ձ��u`7�>�	/�����_PUXL�ڙ����kg*����8����)���|�$�;�v`��p��Ϣd���cmJRP�I*��{�`b��gꪈ����`�b��V�SWw2�]��j������`����B����}O~�� ��#�M�8
8��x��>}�~{�0���P�%v��s��� P��.zrE�ٳcZR��Uѭ��9�b�;�Hj�{����4��-�j�x��ŀ7�0������9�^�G*:��6�V�m�ꪪ��J�������_%�A��XN�~�IJr1�,[���۫9���h���ڶ�ĊiWD���ĸ�~X3c��`��M(��h�`eqݭ��l�kT�ma����V	%$��d��V	%��h� �"pQ=x(c��ZP��<�50*JL)�!$ۢ�,�N�D �)�<=�� z�	�D%G���$�@?8�����y��]X[���3E ���I®j���%�$�Ew}���wذKz�[���[����	ȣNU��^,I;���t��V��,�~���6�-��Y���v�i���;h�#��r' �'4�I?Y'�=l��WL���&�n���׀l�u�7���~�}���aZ�%?UȔ	
Q98�o��޼X�x�Kn��J�srq3u)�'�G���]X��VV��s&�J��Q7*J�ʰ��	K�ߖ��Հl�u��~���Q	bEU}���6]XY�Z#�u	$hr�rL@;�b� qR�������Sۨn:��i��IM<�v�0����.���[8��t'����}��ک�6��np_�߸�nEHT��b��4�%%D�N&�vf����#}���1{�v-�vq���JIU7j���`�ŀz[u�(�s�Հ7݋ l�u5Uh��V��5sv�>��D�wu`{����`|������Z�����J�7|W��`V���]��r����\��|*vA�O���gda��,�ոJ��:�=����!ø��g�.�[`:�vqv׷/%'gO63����w��knÑ�b�K��nt=N����5����5�����q�
�N�jv%sz6u3�#`g]z�D�S��s[�e�����R't�i:�`�\�+Ҏ�\�C(�9��v�6�͒�'��4�l�s�w.Ƶ��d��;x�w{���?mv�4�p1/S�W�Iq�7E5�&�u�%u;u�e�4���bR�7u)AI����5�X��_$�H9���9�꫒�&�3k4�ͤ�*@u�1 �I���_��Sf�ߟ��h���cnU���}X�n��Lʇ�ߗ�wb��t�D�:	)��)�ꥯ��7=�;�u`unk�8��I��Q'��7���>P�K���/ ������`����(rP�1�ォD��p.�{\ئ5�n��RP �!*�&ֻn 3�3��
�U]��լ[x�K�X��_(J#��u`{ǧ�m�N�"�J�:��u�l���A3��k˙�ߵ�=�z���ͺ�8���OUȔ�B��u�<���x��L�}� ��Հ���)��""Q�a��|�=�U���]X[��?U-~�;1��J2AH��m5k ׯ�F�wW��u`��VV��A�i�(H�Ө��<f��9�T0Q5�Cu.�����L�Jɦ�А�BnU�ջ��Ż���ݺ��o�����GA%8�$�1n��7[ŀko�m�t)�eo\L�i��T܎������۫9����V��������tܕu5k�)}��`=�X�n�>�-�ܫ�6xm�'R��8���w^�۬u�X��`	B|����zy��Jk�����������_��Y\��̊�Ȫ'ȯ��|��Jr�D� �q������b� �R�I�ї�R��t�D����ݺ��UI�z����y��u���}U�${vyȔd��8U�MZ�wb�=-���\�u`�]X[�Z#���6&�X[��/s��W���9_�i������a
#�Iz���}� ���Ȼ��\ګ�����6[u�|�s�����`��`~����yS<�����:%B29nr+�Hfa��0j�3\�3=n� �2��b���n�M]��;�b�5�ŀ�I}�_����׿0n	)�$�9V�*@9�q�@H���˰��I4	�M��P��vVb�w��Vsv��7��䧪�� 	� ����7[ŀk׋蝮���k��[Y�fmf����nEHT��be��(X�ۍ�(���d.ʪ&��m�^m�r\u�òqve���К��똴���3ѝ��Bd.����,���й�P�Nv�2vU�6������ڶn�W��͍2)�ǲRG+՛#t��vݭb\�U�:�sn�"�E��hAs1ԍ�8L=�ۭ<á��6Gj����Vk��y��.l�m�S:M��WWk5�����i l�nw���{�/}�F䮡�'V��6�e�.g1Gh��2h�A�5�R9�-�_�_4�)���+ �o����v-�vf�Ձź��8�P���7*���րw�r*@8��U]�[!�ѻuH��Wt�j� sϫ �o��)[��Ձ���:��'�9Q����wX�J+�Ｐ��ŀz[u�l�n��؞�n	)�#Qʰ7��V��X�k�u�X�B�W*W*4�x�*��ufs!I��Dׇ.�I̍5C8�2a���wk�����\�%w/�����@7"�� 	���f�e�ڥv�w?���Հ�B_BJd�݋ �}� ��s�{�sL&���'+k4���9 #qR�Ih	}5��5Ȕd��ȜQ9V�W������}�>���Ӻ��D��,gΛDqD�#i�*��=�`~������([}�W�}�ذ��,���GA%]��ڬI�Y-�Jb�14�6�73j��t�Z��E]Wg&�n��\�yX�m��?- �� #�R�r��Ṧ�����WU5s�k�ftBP�N}ذ�|�Ǻ��#��% ��"p��� �Z����E
��~K�	���8ϯ� �w#������WY�����s�y%�{r*�}����\�S� C�pk����Q��P���ǀ������ �ǔ�ƺ㈩v��#lQ��3b掁�;j>��HM�@��2v*��z���>��m���`�\�B��Hs���;�<�J2AI$jA�X��Vk�V��VnM/�U}��^��DqD�(������>�Ӏ=�s�СB�|���]XL7h�*u�%:m�`nSs�k�f ��X
!D/ZI$�%�}�������凼G�F�lN6���`��EH1�@G�Z�ٿ=�E�C���,���Hn��Zm���	��Ř¸��ge��5�� z�,]k��7=
?H>w���G�m�'R���`~��}7ˀs�Ӏk�f ��,�DL�����d�S� C�p�~��ܚX�۫5�1�6��R�NE�������0}ذu�p?�DD�Ӏo�z8��#$q�B����X��k\��ـbk��"#�!&������S��٠�Z�%��`D;!1(f/�JD@ �P3�T��{��r6f���)tF~����>�\F��ο�(�"ʇ�P�)�C�Bv)�2�QD.J�fF!cb�c+���8?SJ�J�1�ԇ
�UWQKy�ɶ-�m$ur��^K2�,O$�aW������q�H	mnl�N<�U�tO \X��6y�R�&��ۅ�Yx�gi���78!�9"T�U��l�nl�n�L��mA����#Jۢ�Ɯ\�0�h��`�C��ɵ��Um�V�vZ���*J�񹺒[c����>�e��B��ƻl$m)��y���9rm���<<��Z�V���t۱�k�p]j�۱�|q%jŴ;UA8$T#+�14C��i�k۲ZYKE: ��x�RT�U���@A��nS5u�۴�L�hZ�U�s���V�*�P Pn�j&.U�Q��u�1������m��9m��W���%Q@{d�f�β;Un4��@�V��ʉ��^�U�1Tp]Wll���*�[-��E^��`�kE�m�==v	�;��;����lu��+���k��neKW�r��GI��d��W6�j)�/$����X��n�����O8h��`� [c�JjK�7cDX��m����#;21�u�=������t)�݀-9��	-(kl.Y�[����'qK���jڲ@3m�7�YK<\����UG(���u"F�t6���3���T��!7��ە�sʪ��N���g@-;[p##I��d�s� �wk����v�7N81��r�A8�t��b��m�A4��"�]恪���͂&]�
��Rv	ɔ4Vͧ<�.ݙ��6��2UT��t!49f�R��j�pj6	U,ul��k+NZ���l���V��,��$�t#h�ڱ�q����dE�ZO9h�:���kkm��r�jBC[̐�5mPl[]In�P��:]���������+�v�MU�s\�z�`��պX�m�K�Jd���(hvl��"MQ$�c����[r�blsj��[�<��b�����j2*��r�nR���{��{���wp8���Pg�
���
y��GB
��p1O�<_ww���w{����Xt��4�jk; v���=��+�krS�mq��`'��k���ƞ�'�����ǊW���\�cS�&5F��1ۃT.��ӄ�z��bM0V�Vr�h�bR�s�؇�i��m�\�/./N�n���ש�M7���;�y��`8`4�U-�h��*MʓF;%�-�t+0)-^m����c�j�^(�����p�G+p-M;N�{��K��&�L�45�l)g��WfZܴɦ ��Q[�{�Z� {Z� ׶Ϣ#��>}� 4���E#�QJrS��V��VnF`[ŀk�s��IL���ueի�q�'R+}�Ł�ݺ�3^j�7j�7�`�R4ې��,��]k��k���"V��,g��n@qIQEr���V�������Ձ�ݺ�9��j�)I*E rB��tc���^�<S�f�x_,ltn{BsɃ�ު������Uȥ:�ґt����;���7��BK���rr&���'"���`w7n�>��}_!w6���=�`sri�_W�$o�z8��$��m��9�<���`��"��cֈ�B2F�nU��{����� ����Q/_~X��wwJ���n�Vfm�=��EH�*@sɪ������*T�Ϥ���A�r)$�����4IK����l�-�ݲ��tg_�{�ܯ�n�G#�8��i��7߿]X��Vq��UU\A�~�=���i��"m��]Z��ŀ{i�����=��Ϣ�����q��J�"7%X��V�78/�)J�J1D$�O��ŀ6�U��f%~��Ju �"�U/�?~V��X�x�:���S����9�I���R�NE���n�X��Vq�z�U�V�h��#i�H�T�9�1��^͛pX�Jh�k���J���T��)��-�d�*AI"$QI\۾��;�uX׺���Ձ�z�"8�P����m 9䖀��Z�����}_�g�=*G	)I%H�=��Vsv�DL�}� �]Ӏl��we��]]Z��ܼ�@s�R7 9䖃�N��|��k�G5X���4�ґ6H���@F�<���� 9ȩ��;��̶��-k'(���K��R�L���F�(�mh޼[o�?o���Yي�9�^���@N�-�EH�T��{��%.�AJRr.�~��U_}�F��X7ذm79ДB�ӓ�4���pjEvo�u`s3n���W�If�yX[�v�Ml��H)$�B')��<���� ��?*���Rc��DqD�#i�*��=�`{���kʽ��p�^{�xr� �� ��w????yHw6-Vx�eXԩ�=��v|]����ى�z�6ݏ+t���c����ΎM�Ի�G�>�NUw`�:�n0�٭UA�Y:G`��U;q��ћ#\г$��[����x:5#j�:��֬��ֱ���םk��=Kсs��Π8n�A������NbP�<h�[��{2v�H����f�y��D��[mۮ�����G2�=.���0�t�ݹ�g 몛�MѠ�:�U,<�lr�4���"�F2IN�q`��vnM,fmՁ��U��wI!�:�SY�^n 9ȩ��<����/�H�z/!�����29Vw}u`s�-�nb�����o376�kol���@s�-�nb������3p�_���ȥ:�m) ����(|��=}� �Z� 䒎NԾ�r�]"ɮ
:	���V��!F/]��)ە\[[gq��=qXgL����}�� 9䖀��1 �a*�]�wWuV����o���IrQb��^Ȉȴ�d�]�p>ެ��,g��DqD�#m�*��=�`qnk�;��Vw6��9�E��6SrJm�=q�@s�R��K@K�I$M�G)��vsv�����XǺ�-�v��ؕJ�R��s%�CE�[�G96�#���{U�5��j��iM'����29Vw6���=�`qnk�;��VwI�6��Q��Hy%�=q�@s�R��V��r��R�9M�"�^�;��g-�AЁ��_�M}߹Õ{�}�`o^#hN�)��"n;76��|��� =q�@G�旵�^����y��|�<���K@s�w�o�󿟏����fV�=!y�3AC�U+015�G7R�C�ڭ�Q� �7s3/6�㘀}�Z� :8���^�&H�a%G"i�`g^꽤��ց��H�������d���ݎ�9N8&�7���ͺ�1nk�3�5X�b584�M�4��Xz����~X��}Z��	$�J��ꐈ`��T֟D9�<�Õ~��lm���B!G%XǺ���Vsv�����X�����$���	sZ�9�~���m�9vr�v�v�D5�s;�$؝a�W��5�%|��9Q6��@�����`s�R��Hy%�'=��^V����{�����"�����K@>Ǫ�}�F����!r%*Q�`w��<����@s�R���76��H��NU��{��μ�`w7n�=�.�}ʰ1g��	l�AH�qX��`��`z�`/]`(MR��A�ᑄ��ƹ�mp�rJ糣t��Vں܍�nk�e�7O"�:iv���ņs�I�)��-Tw-����Mp�q�qA3Aۊ�1j�<�������>z��ҴS�m+��1��u�k��z`��g��_3�K(U9�ˣ�	u�I�]���+8�yE�d�I8%�Y�����h���[���FA<23���r���w���N�Fu,M]T��t�a�mU��M�j3�rیձ�rY �P�D�ԧ)�#n>��]X�۫������~v��_�I�%"t�n���@tqR�s�L@8�����r���(M�V-�vϛ�>I(�Uw��,��b��S��T�s7C4���-�� qR����5�܃��JD�B&���׋ �J?�����}_}8ϛ��[3a.�P�]�Vȗ��,kXV��k�2�Λ)m��h�l;�sK�Au����Hy%�����"�[�Q(FH��r���W>�������@0�EpS^*q<й^���r���Չ%���s�����ic��#��9JF㈴�Z��|�Iw6]���y��+�I,��E��Y�l�9$u)ʑ���I{��}����Io�~�s�%ܛh��X���Ē�m�m���:n&��ZI.no+�I.��E������$�se�i�7��뗚�,.%��e�Ne-��PV4u]�dqh�+�9aQ�����ʭl�8�	�+�I,��E������$�se�i$����q$��U��+����I%�7ϜI.�ˢ�Issy\�Iw&�/�m,���I:��J�J�G8�Y��\���;�|<�4^�RO�c�c�2?~e(	��$���lN��5�,�&׈H`c�U���� a
PBɋ&)&$����l2�#�e0��k���0����r���Z٥��,SI�+��
�<&(J��f��h�i�!�a�ʌ$X�q,CL�#$�t��C�N$2B@���Y���:s�'� �g�B��;�
y�<�GB!��*�D�}]=U}z�+!D%���-��h�e�I�33�����)n��D��Qȓ�D��K����K�6�i$��5�/<�_(��]z�Ȏ(�#$ci9\�Ic٭ZI,}�|�If�-$�77��$���K
��(�blmV&���%1e'\��-i�tZqj��\�6L��"�� ?��8�Y�.�I%���{��U�^�[-$���~�'$��9R9#��%��贒\��W8�X�m��Ks_8�Y�i[iIQ)c����K����K���ͽy�|�Io�.��M���%~m� 8��(M�\�K��|�{�e��כ��$�nˢ�OҾ}�;��+�I!{�z%wW#d�Q�#8�Kro�8�_�������I%�����$�=�e���5o tJ��j�AZ��)p��R���諔��<����d�4��z惛k�c�� �~~_v�\��W8�X�m��K;3W8�Z�l�
B(�NT#r�I%���s�����y��l��^��˜I,ݗE����K���#�(�$ci9\�Ik����K;3W8�T��z]�K��r�Ē�Ѹ���9JE���Yٚ�Ē��tZI.no+�I,{��If!!	RT�BH�nـr��ߗ��b�7ծp
Ja��*�����[�y�Y�o5���CBD�gm�գ���!�p���Vm�0UDn��y�V��MV�\`�f�]m��P�mSRZX��R��le煓t����z��mە���j�i��YN�l5�`4k��N�l1��i���*U�%�9H���.ݝ=p"ix�X����14�uˍĪ����J�;��+�\psK;6���9UnGWlLӋ�����}��g��֊-i�C��)�b�n���i]�(�g�.Ru��k�7`��1&���68�!�{=�Vwv��μ�`wri`su)�m�u#���% H� ��G�@z8��
����n"@Q�pǾVw&�76������޳6�u)ȕ8�N<�%��0�ذ�x���� r�b�)��HB7�ͺ�3��Vw]��ɥ���6G�q�e����Q��nAn&��j��m�Z�bt����(�R�m��X�۫:�U��ɥ��ͺ�8������H���Uy���4�t���g.����w޺�3��V���FHBT�)���<�ـ~z�a�D(�{݋ s����Z�iIQ)jD������o�V|� ��G�@zK��ff�V�V�m��H�*@;�1���۫ �kj�⒔P$m��8�c���N*��٣��jN:��(��w۾���w�l��nI]�}��ܚX�ۯ� �����6�u�r%N�ܑ�ݶgBJ)��� ����u��D����
B(�REQ�X��������SJIB�P��_��<�ـ���QAʎ!�V����n{ܫVo���ɥ��ͺ�9���$l����n���u�|�F��?�}� �7� �Q	�S�+�n.j�ԫ���\�б����`�l�6��䭞��wmͲ�@Kf�i�BT��6�|=�Ł�ͺ�3��V.���ji��$�mH���9��g�D)��v,ξ��m���oX۔�GRH�*����X����J"gy���,�by�3���iZ�EUݯ��DD(����������c>$�� C�߾uU_D�yVQ�I:�r$ȉI�#@t{��}>�x��R�9�W����֕U������];tD:��L^6HN�m�K�<&ғʅ?�ww�>���h��ܺ��<}>T�}"��s��9Ս�#�(9Q�Cr���Հ��G�@z8��%�����X]����6}��=�a��Q[��]X�߮�3�����$mH����� 󘀏D��I�ڑ)!`ssn�UUUV�w��:��=�`D8!ZQ|�!D���$X�T���y��YF�	<�Fm� ;uR+���Ӧ='68^��v�U�7����ǯBp�D9�jN��fi��s=��$=���P���������<��|��J��\�p��jmn���vm%����	�����zp�۱3���;`�vXP,V�v7��Z#�Yb���}F`IY�A�Uc���;��2ʫ��іGs����us���h���qt����ա�+v�Kղ���9�ku��b�㋷������nu#�HH��������^o� �l�`ssn�n���+��u*1�%p�}Y�BIL����=ϱ`��g��76�u)ȓ�Q��;��K��u`gwn�]�v�͐t����$UV`��X��Xϛ�����ŀt�~DqER�	ʰ3��V�����H�-i��ei���v�uĒ�a�ͷF�`ƥ�u�9-���	g�Y]T�k�a�����~?`��f�DB� ���n��.�J7N;��K�}��:fn������X���ǏSLN'jD���<���7��âe�wN�� ��OXێ�r)	�a�_}UT�=�U�}��:=������_˴�n�Vmm���^<��@t{G n�X��i�~�$��MƛQ)II��P:��J�M�B�.뢀�;����)�%�}��̉:�G"����`wsn��m�+�1n����Iʊ:rA$Ӆ��ͭ��R�Ih9�_~]�g�nl��]\ڔMZ�5�ŀo���ʂ(W�*�Y;N�`��X�[C�.��䨠�`g^�9�4�;��V����=��v���?8FHBP���<����Hn*@>�-�6ik׊��%IvD�>���Vr;9)�;[��rF�ggv�5��p�T�� :8���H�%�<�� t�oX۔�IQȤ���u~�H�{�`w}<X�۫��G�ʽ�]�ȝHD���>���h9�@tqR����f�N�9u*0�Ea��.�Ł�}� ��Ł_��DJ^�W
1��N�~h�'*(�$iAH��mՁ��u`g^�3^�3+6�(�H���y�'v�f��E��聺6��ve�j�/4q�QJT'*��ݺ�3�uX�u~��� �o��Z�y����R��:�U�H��x�3�<X�۫���!	C�����{����هД)��ذ��8��74MYq��*G��ɥ���u`g^j�3^�n�����B9RH�,m��7�����<�ـ~_�
"�$�)�4��XH���nԒi_ϋ�ѭ�����͇/ݼ�)�f�19�XkY��㼶3f�ݑ^��z�+ܔ=���D1���0����	JBK�!�$�i4�4B@�(�8@?�%�¹������D�PN�߶����wsۭ�ߵ�U� ��u��:A���:P-�ƕ�ᕩ���d� �5�n^�[ɣ�������Y���D���3�h���c��y���ҍյ=��Ɗ�5Ҵ�[�@��S�����7X�F�r:,�9nCeq��йYÊ^�K��Mk�Sk9i.t�FQa�	V��eZL���
j0��t�t��T݋v�9mҐa+9�$d�	�� �6h��V�ð큮�m�[�v��v�TYM���Y��z���)tA�ص��Qk UWD�<�.��!pI*���
�݁��7��!qqD/m�Dee^m��mBʭ�j�W�%y�iV��ڶ:�b@ZUNͰ2�	�������6A���SR���2���y6x�C��}��U��b�c�ԭ8�&�V��4˖���r��7n�k�m�U�b�m��y)����׀z@ō���md�4M�~��&��%m������s�\ؗme͹c�3�E�M�g����S��Gk:��n�-�>��0������*��m�͡��7Dm��u������k��d�먥�y����qk&��,������Ț:�3e�㬼F]�V1�: -�;F�-'�`�D�i�S��^��՚}A�{Eȁ�V���]<�w���5��Rv���f�+8�R�:UB�5j��Y�7Ȣ��j�Nfp�*y�h˞���C�A.#͡�F�8hڠZ���4q�Zj��u�%Be@@�U'N�ilm�v�,��K6���Ԙ��3Nr��H\+ �7;<%T;�ۗc���Ѓ2��Īv�8�Uw�ٙf�O.j~~����nq�W#V��p��prt�GT�A��V���nImt���}����N�[��"�s8��]�fv%�8v�U�
�2��4�q"Yx�P�Qܢcl�<Q��&JѪEt7���m�m��d�V�R�T�h�<`u��"������^���8����X=M `N&|�� ?<GH����CJ�����6�ß������{��ֶ�uV�S��'W7&���ynR�%΀���J�Cm[v�t�͌i!ݎ$�|b�;�B�v0;�Z���лx�����@GI#S[�{pv��n�������p�����=z�-�M���n#5�nyc�c����%=i:����YǦݩK;=^�RQwR�=�C,F{����6N��ɱ��c��[�2e���{���w��}����Q�I]r���O=+]yț,o�N��Ț��b�h��M'뻻�o^^�wW"u!7%����3^�;�4�3wn��3i'R��:�G"�5�s��Jɼ��v,}M�u}_���}T���6~��Gd�()��u�`�Ň�L����Wt��v����%97v��ν�`f���DDN��0�'uwu%�Ysj�j��|�`Do<�����7��;[�EDR�H�'���!�:\4�ͺ�W�h,I��U�K9��[d-�2Wef�{���`��{� c�`�j���$�mH"HXܚ_��`>�z� �;ս��Õ}�}�Xܚ_���?1�HG*I�?�T�}�Z�� =�:]L?�1f\һ.J��_���$�+�Ͽ� ��o��qR��*�+k7n�+s6����� fj�;���>�J�jFʕ!I8)�e��*��j�f�T�qk)lr���e�1��[�.�eM՘��kŀo�\�(�U_qs�ŀa����R���`{��g�	L�i��޾0�^,��f�I(�	)�%Xך�wf�`�w�߼�8r�߽�Q�}#�M���E*��5w8DDB������O� ;�T�}�Z �r�0���jꊻ.���?=x��D-�ظ��+��K��:i�:N��$WS,两��=AXgv�]	b�B�er���}U��򖔶6�	�HH���] c����G 'K���I\ҵV���_�{O�?�!)�y���Ձ�ɥ��fm$�S�'R��V�m���B��;� {O� s�5�ܨ�l���p���|���*����7ծp%BP�������v���R���`sri`~���&�p͞,nmՁ�ԫ^ҥ�D�4�,V��:6�)��)8m��m3u�$l]V�T%��I(�J���μ�`gri`ssn���Ձ�կD�B�NGI˜�m��B����w� ����s��#3|��8D�t䂄p�;�0�x��")���p�|`��yRی$#�!#p�3��Vu���K��K{����wWq:��nI\�>��-�~��|�,RQ��U}�����!ƐSQ�IB�=�>nmE=&�Pe��D��t�[���VɎ��'g�$+d7/b%,ȷ#A�v(6	Z��/V��vq��J���ԆnZU}&\l�wѶ�/,�r�g�@7=��Q�`�V�4��]���] ZE�ͭ'��M�4�kj��@�����~��a|�e�K��u�U���G#3���ֵ�J LM����,�?���(�O.�\�.���%��I&v�o#\�^���;=u�vd��h�v�<�G�@>�R�9hr�ܨ�l���p�9�4�ԑ��]X��Vw&��3bQ�jQ%9���K@t{G�@z�5��H�F�S�7:�U��ɥ��ɥ��˾��`ub��HBP���fm�=��� =� �$������s=f"�ML���LU��u�j�T�s�NL٥٨�2<�NAO3q� :=����K@>{n���5HG*I���ݺ�W�}_R��P�G:��y���0���^�����B��������ɥ���l�`n{�V5��Iԧ"l�G"�:=��� H� �$���z�nTq'D��p�;�4�=[��+�n=�;�4�:�sd��r�qGz�{Ҝ�D�9���SmP����bEᐼl2%QF�QC��3��Vu���K��K�W���z2I(S������������ <����!	C�#��Vw&�76�l�u���������,ǞVf�V���ӎR��G =� ���@zlmm4�A!�$RU��ݺ�3�5 :=���H��^C��ݽ�^W��b�3{O\�j��>�W��ය�<��ɵ�C򻫸�Q�*�Àn=�3�4�9��Vwv���՛IJ��Iȓdom���*@>�R�9h�u6�r��:$n76�����Xך��M,qnȔqE�HP�DB�{��`i��{l��	%�N)��D�o��}�|�W~z͌�GJ�9#����Vw&���|�,�DC�WeЮ�����6�X�YJKpN뚚��̡�Ӻ۶���<�dԊ(��!	C�#��\=�Ł���*@>�-�˻X^i�{�Y��������T�}�Z��X͍-���$#�$������X��@t{�� %˩����-���ۼ76�y>�G�@z=���V��JT�"ND�#qXܚX��0�m�����c�Ș�
^��,=�]b���2�-<�q���gQ�+�9k�}�&��¶IH�nɵ�t�5���˫L@\T9� �6��Z]���1̚vK	�sr�c �g^s���D>qH55�p�Hu��<�Gp\F�>:L�O��%�"��R㮯Hp���NU�:�����c�R31-R�2[�sة���F���ɺ@b�Yo6�7��r�јkqf�kz���"qE�7̿f����TZ*z�x��:��7U�^��/f�	�T�M�':����r��n%��m���� ��ـo�\��A�0��]ʎ(�R�
���ɥ��y�������������mG�	Dq�%X��@t{�� H��˗�t�h��ܬ��@t{G�@>�U����[��V{|��'���r������T�}�Z�� ~?���%����k���"�.sz� kzNy*�&�Pn���[�'��Hڴ�R'����x���x@9��X��yz��G �$��7���U�Q�T$��0B^����� ��0�x�-Y�R�IQD2I��ɥ��ɥ��ݺ�8�5�͚�r���ͫ���� �EH�%�:=� �n�iGQ��!B��3��Vw$�G�@t{ �2�nm]i�W�����%:��m�Ar�Ժ��v^֎�Bz9&1*I8�m��BP�i�Vu����`�}"��.\3�M�+7r�3m��� �EH�%�;��+bp�H��*8�`wri`s��/s��U���0��M�5� L$%~�L�kA��@�� ��f�!��хkh"6fXQ�YZ���kZ�;������ I����mb�3)8!��`�{�&C �OD/OpaLT���!@�l���	"�`IfJ &`OɈ��$D��������I@�'Sc�U�W�s<%$z�s�|������B����?~������S<�iDD�G"p���_}T����+;�K��Kt���뫹��Ui�#���=����`���/�B�:X�v*L5ʘק�$�,�A�n�ܚ�'gpSa9h��Tf��6f��� =������}hc��r���r����ͺ�9�4�3�5X�&��꤂���iGQ�mn�^m ;�� ���l��V5����%
F��`g^j�<��`��XQ�(���\�j�*�U\����?s�Vu�/��:�:�ݴ�� ?��O�^�>T�}�Z��᝿���3v+7V�g�:H�w �ݰ�I�p�[l��IxgF�Of��晢��H�*@>�/��a��<X��/SMDD�G"���m����<�Z�տG�@y��?��]ȥG!$����+7	���ͺ�;��V��B�*I���`c�ـ~z�`z�`(�脫�wӀ?����ܦ�l%JQ76������7ծpz[0�(���w�)W�	rZ.�'�:��uei;"$v6Ӯ�L(�*����,qu���za�IOd6B�9ރ�n˕���;z�Vj��"���Y��k&�m��'�STX6s�XΨ7$k����\�|*�����aL]�=V5$mIL�mؘ�P�unN�n�I���A�moם'�tP��Gad���ma��/�l��Ϋ$�I���i�Vom:��|�o�y~��ݼѪM�u[<���0f����u�D��n��Zse�j�;$cZʭ{9z\�ē���?�w�>�- �6G 'd�{f��U�jf�j����s�#�_��,��u`s�jѲB��'"�3t�`��XBJ���X�}8��R�z�$tԕ)A�����X�۫:�U���������Q�9Q��� :8� ���� =T��z��d�R
F�)8�p�]2�JH�A7��Ƶpׯ&�^�'T쟽���L��wwk��g߶�q����T�7��)R���NQ�VnK߾�}�  �Av����<D����ܩ�O� =}& :d���mfm���홢��H�*@>�-����4��Ҏ(�T�EBr�� c��q����ҿ>{��q��BRR58��+{����׋ ~v��$��\����%]�@\f�I-:]�)�n���j����:�S`v�c�DQPl���:�Rr.��x�9��V�f�u�s4J�U#���zf�G 'M��9h	��_>��ٳ�G���	"r��IV���*����r�<O<����O��\E(�����;�b�?=��s\jF�#nq��i`ssn���,��z��*9MO��X�-��^�ߗ�;z��7ծp�-��v÷�ޗ$fخT��5�)b����2�-n�p4��z������*@N��r���@rkJ8��jT�'*�����μ�`op�X�۫{�[��GJ��') ���� =T����.-$!(l�Rr+7	���ͺ��w���i���M ����+����g �=^E�Q�tӄPp�9��V��}�~�>�^����g���<�(�$WS-D#:���a���v�b�ZA�vE`Jn"ɮL�j��Cw�m���v,}Z� ץ�������������		$��:��vnK�ɥ��ͺ�ꪪH3ڏ"T��q5*T�u�>e�{�l��%3������:�5*�M����p�;ܚX� c��q�\�˽ͽ�//U�Dݘ��X�����_�K+��������LBt���wB�x��:�lq�p�N�狨:��\�޸�`��=�y�y�7e�۶	�5�3Xƙ��y#/-��E>�Z/;v�i�=�ܽqۤk�6)�i�nl�+��n��W]p�g��OCӓu�ҽ�&��R��،d.���WR&D��lޫ�a���.N	��kӨ�6��$v��0c{X��nUHlß�u��w��E:&���O�f��f��kz��z�r'F驔�Uj�K�X�mQ0tE��b�뫊�cM<]��߽�����`ץ� �������ذmOOJ��h��۫��@8͂��U`g^j���Gk}^e�Q�t܊88`�|`z�a�J""&^���2��3�Dm48��r�Nw6��}�Z�l�`��.����RZeHH�NW �{�`W�[�/� �x�7�4�3Z�V�)�D$��)$t�f�c]I0�Y����S�΄D�bJv�uۛ�E���h	�� =�:lך�]�J��Sq7D��,w���\%\T`�@���	E�I,޾0uwN ��� ��Ҏ(���%	ʰ7�4�3�uY�K٤�`g��V�f����Dm����9h�@z8���Hu�Z�R�'R*NE`f�4�8����� �V��?�%�mUL�*.�.��.�TX��汜̃�n��g���:�G o�Ν����%H�pp��ߪ��� ���l��J2�H�9R)*�����μ�`op�X�۫q��/]]�Ԅ��Àw�w��]��ܺ.�?�؈��>EaOP����������\���F�T��G)qX�&�76������������|�	Ԧ�n�Q홢����bs67�������fp�<�����Js1쥑���m��؃���t��^���\�|��XM����k����� =q�@Nf� �˫{�[��GJQ���Ź��R��(i
!%Ts���ذ=x�u�Z�R�'R$܎���i`s3n��%��]X[�v4�m]5*EJjʛ*��BU��y`���w^�X�� �(P�q?�W�����,���=C� �INT�J�:8��nb�ln*@�夸k�v��p8X,��foClj��>9��6�ݺN�{Yn�o,�_{���B�;����^�������J�(Iz���� �y�R��TNS�$vnL�DL�o�`ϱ`�u��z�QTJn&�AF8X�۫{�K�3]���i`;�Q�R��X~���;Ͽ,��V�Kf��7ߕ��z��()I@��!`qfk�������]��7W����*�Q_��Q_�DTW�dTWQ_�@E��*���*��ʢ ��"("�1"(B��(#(�"B( �� ��� U�� U�� �+� �+���� �+�pTW�@Q_��
��� E� U�h���TW���e5���d1}� �s2}p��@P   m@P �            �|�
 �H� !H 
  
RHT� (� R�@

 @ B(
� �
*�   ��$ ��b)����>�//��דq���o�n_k� ���,[��}���&�}������ �Ll��-�� �^���}}��.��m���|������ (�K��]�]���r��� � >�    *�% 1Px��;m�7X�e����} �}��ܰ�n[���ozM�[�6� >�;ҫ��}���zxz�=�k�g^�x u�;���^M�����[��zWp} w����{s�ov���7>m� �    IJ��4
����{Ͼ�y��Ÿ{w�o�k�E��>�x�� }�B����Ͼ<
P ����t ��r� ��ҝM� 7k��s: �v�)c4�4�Қi��:Pu�:(3�� 8�:I���.  )@P��� ΁A�Ί
q�@��)�"iJQ��BΝ4���JN� 6�t���;� w+�>vz}�u� ���en��<>x�\������c:}��|��o� =}�ӽ����շ{=/�Ͻr��(  � 

�����\w}k�u���vu{g���✚�s���}��5�y�W ���_n;��}�}� ��s�ۼ����x }}��}���}��ow�����_|�W�}�>���N�:��|�Bf{�� z�)�*ECF �������)P  "x�T�U?ґ�����UI�R�	� "�����R�� M))" ��:���_�����_��m�,�����4{��eTTW��_�QQ\EAAS��QQ_�*���� *��T?�"?_���?s�Ц����Q-�No�v c7:�CV���$��5���2�SI�c��`A� @�� ����4��$Z��$X�I����ŁBB:H	 `�@���M��J�2�L5CP�
Mҿws;�[�6�����Z)LЪ�N%p�p����0#)��x��Llܲ���9����d!u��8R%e��B�#��*I;~c�7��w�Jk��T�p��ߐ�$IҰ���I5c7>�W���~�`I�`@��r],c���#'0�S!�k�%ӆ�SX��%5��у�W[4��+�:VFю���᱃D
�M8�bT�4lH�`��pa(PMe�E �N	��&�U �Z�F��F�1:�i\B�J��%
�+CC�F��i�X�Dj���C�v$k�
|���$bFF h�X�t�)���{=>ٰHW��1�Bb:H-5�6ƚp]� �{��0(@��M|M�O��޹�����}Lc		:B��$
��!#E� ��$k
�]$i���i!��c��$��H@���T�B���Ժ��44� l�9n�%p"��i��kcn�Xp�&!&�v�����������F��a.;ݐ�f�SZ�\��BP�CEH.�RQ�H���j3S���,���C唆�c%2�������F$aL��ṉ�,�	.�X�5������A.�l�߉vP���R�*�~��ۙ�rҟl��Q�dR	��T�jդ��R%UWe\��˺Wl���A9wͿv�[�p��t�gH�w�bq��H��t�Iwv��k��hS
?�8�J
�8Jj7����m�@����7$!v|��*F�9���s|
}�	ɣ%H57�٤�Vݛ0v��g3�Ҝ]��#]8�w���6G�8��]Cb����_h5��K�%IM2��B��K�P�4�k[�����a͐���E+C���۟�":����4:��-)C�A��RA�`�hF�.:�+�cH$|s��7X�e�ܦ��T$��c]�?4��%4cV!��ݲh�bA�WBF�(U�F�j`�3���!�A���` �:��5�B�6��E"h�!M�)��D��B�6�C�R��s{��X�7��C��x.�m�@�!��m!BHQ�>�ii���ݙ��fS��.��9�k\3\$%<HSU����i!�\�&��KN��S,���j���>���9�W6���2��V�E}e�B��p��Q{�:o�P���˭ND�SZ��s��h��o�(F	�Ʀ�w����gu��7�1b�/f����%4�˳����F�%,>ֈ蕉��o�7�WA��(�*}��t`�����P`V��h1��~՛98CD�HÇ^D��	��Z;�݀E�_�d4����ɕ��~xF*h�R,�����a,�]��.��l�!�Ѳka�D!�*h�!CF���q0�ј|�(:P�fFB�q���e�%FA8���q�P�CS%!��Kh8Z:H�р(D�r�n�� Ӂ�Db����SXCrB���8��6p9R61�#Ma�aO4�P����|��l١�Ra.�d�RJl�����PÇ/�����ܐ��B$B�
�b�Ø�:1٦ѵ�])�pW[ќ��!
�$j]w� "��o���4a�F0��0�����IMN�;�3�p�ad*�10۴Ǆd.�6g˒$I�����!CFCRf�}�M''���jtӶ4l�3Zn��HׂoF;~!F!�M�fl����1 a��u���O��bm#M'ې�M��J�5iVcPѨ�4i��D�E�6�5�)�3]0%��vF� Qt�+�"Ѝ��h!tjV�vkp.�k½�a �Xߙ!SJl�R-b�G@�c��`L@#�@!�.�H��	���7�{���#",)��ҰH�1�Hˣ�4�
hL~cM�F�)����f̧��.�����+� D�i�3 ��,a ���|���k���>�gX�H�`,�@H� Ү�B�����
:qčR+ `t�8�J&��RK�i�4� ���SK!��FAБ DH@��P�0�@"�B),��!U�! SA�#�W@D5��]�(�
�H٫!WA��a�MS�.g�I5q]($��m,��A#��u	SLCF���B�au8CY�F�� sT��<Xm���K��0Ѭ�aF,�	��8l�5�R�
P#WL�֝�$�9�M `�	>2F�B���,*J�]X腁%0v�B�2]r|JDӉ�HG7'!���Üq�P�a�͜&�5]ID5!56ܷt��D���>��@, ��� ];1d���c�T��CZ���ą5l�dԐʤ�P2��/�J�M}���^BBHH�)�	&�6ZI*JB��D��jFJh7I$�ŉ�јK��1a3��p7��q�r�C�T��l�At�bB�7FbT��&�1�T%Il�J�$(p1�GHAhv�!�ܮ��X�F��8RNd���
´�HىM�#Q8�` �#MnoX;bN���Xj��B���Ya*RR�V�5
[ICPa;�4t�aSf�9��̈́#�j�f��!�lւ_��>��Q�8|�Z�99i"�͇	��J�]4#n�@,c�|�IZh�K�$00`��4�OF$�I�� �CF7f����@(F� `��۔��9CA�vׁ�aMaVB�@�dhː՘1���SV����yB���M:�&�턄L;���Jfo,8RF$X��:&�I��BSR�3lt�ѲB�~jaN�0���lʹ V��LvL6}
��G��Xr&���m9�.;���*b�4�#i�[aGI��+łWL�$�V��0�
h�D��IM:*�4�A�3�e��3XiH'Q4����'~�����v^�M#"&,�A
�"XP%4|K4L�B<>�ua#n�m��Yß}$}GZ��#;��]��$HT��
iI͆Е*�j�!;���.��.qM�]D#g��K���m"A"�F(C��@(�(X��5-@$�e�ըF��N� Q�D��:LB4t`�j$�UtF��H�D��9���jǊE)59]jЃ!�i��4a4�	d$�0 GRlaCA�4o�?,J�vC��I]H������t��pY��@��&n��K!�Wb�B�ԃ��-M���CD4�F�tF;�%$��+�FD16NHBD�����f�@�f��u���7-o-d��aD�t9
��V��	l4�dV�`��0�R�;%N @��kIӇ;�٩����)ROe'��W��m��ٳ��-� �  $  @   �h     %�h퍕#cm� $Ĳ����띱w\�S-nTh�� �W6�GI������UA�lZ��M�Gz�[� 0�'i�ҭF��Ev�J��� 96H���f�Nv��4P8��������&n�'��6^��VA���^�A���b����� 6�4Vݵ� ��   �-m6���n�[v�U�X *�`�1��$    8 ��   �u  h�vm�l�-m&�!����mD�l[�M���-� $  �   �4�l�]�� -�۶�!��$86�N��8�ºNB��ۂ���iz�l�      l��	 @6��\��m*�;X�-T�K�!�V�8 ڭ�,koZ^�9e��i1 �ڗG�������U<��bkM�DP����gK��m�N��@��V�lGL�X�)#v�L�Laj�b�*�àA*�Є��R�\��Ѩn(�@1���2M�J�K��n   �`-��[@l b �6ޖI���	Yj�q��v�[��8�-sb��{T�	�gkk�8xV���W����*��Gr���f�ID��t�5v9l6��c��[Wx�̹��v[Ki� ć��kh@  -�Zkm�[:���8[@6�kj@ m� �[���mi���[R �� m���m����m�  H -�v�-����mp�-���c�9  ��[��[��l�  ï�f���8K# ����i����B���᪋�B��,] �s���uT-[*��7�V�׶t���ړ�U��.N�����HI$�lm�ͶV vYm�X��UuUn�;(*�EqU*��{I�6v�� 6�Ãm���'nq"�m��v1�H�6�� ls���6�ڐ �� +iҭ]usa�l��� �e�N��u���
T���e3/~?:��U����۶�m[���L�$ �UJL�Px4ҭl�hl]����Ӧ۪7.�$��|gt �D�m�۵��M��m�h-� l�m� �gm� H � �  ���� ��l$�����K��� �`  m� �� mim �`-�����UԫpR���[gf��  �lA��O��;���h	�m��v l �E�u �n��;H[@۴�! �mċh  � -��Ӏ2l k�H�@  6� rA�� R�@�  �m��  �Y( ���>�mw�շ^ i����8  8m��s�l� �[@m�8  �`$8 ��[@D��  $ m� n� � l�`  $·m,�9��"�N�j¤���`� v�&�-�  �������Uj^��W,� �@-�I�۶�٣Wf�ja�l���ņ ���[KM�r��V��:C�,�e4�Q�r���TURD�vũ�[J  m�Li�7m!��an�̤t���ڌ��y��ݴn�օsd��ݶ�;$�֤�$8��  nK�%�h86��	  $�m-0  H  q�Tـ9��ho�m�6ؚ���  $m�m�[��6��-��m8� 	6�h -�    �6�-e�T���HUV�-We��.�kk)��`�h��nˀm3���.�EϐV��i֥A�!5T�J6,8��ꨶ�-al�mI��	8$�^ä   ��lԫVʸ���f��5@�y��kj�ڢݝ��*����M@$Xii���lm�]"P�f�Cm�6  �a�Ͷ��ie,�(��X�T�e��F���ks�hH �M�����:x�)��mUTr����UR m��l���{2�N)D��6�`J�jl���ʵJ��V�z�sUU -UuWJ� �����|�jG�r]-C���d�v�E��:�pm˴�+m�rΗ&��N�D�!�$8j��6�md����&� -�m)��ְ�`,�nm�m�.�&���|$�m���  ���Hn�	�� [`�5�H㵷-!:��  pi6�H.���g�Uk��U'+. [�������m��&�  ~��- ݮ �g���R �[��ɢ����&l�i��H[E���oi��I��  [[i(h�*T��@*Ը��mSG	D&�q��&�m�Mop8 R��m�m� �   q�m&ͳmi��Ͳ�i�����n�%Z���T-C��
�8�;vU@�����Ii�(K(j�t��7���L5��'Am�t��<�٢������|�D�V�mU��Nx��Mh�ȩ�608�ؘٕ���i��}�ַ��K.�[�i����a ������6�]UD�i(Ȩn����@$   �Se������2�*��TJ*յ ��utu��$b��X
WP�T�ְ�`� �m��d� �l6�.����	: ���q�lsMq0�qi�8���\�L���U�J�UV�UʻR�U*�l�Ŋfcl�m��  8�@հ�(|��|Zl9m8   �[\�k��h9 p  Im��-��,۶$M��ͤ�m  � �  �����n�� �< [D��kX[@mu�&ٰ��6�m��yj�ThSm�U�
U�٤�ְ<  �&�ۀ ��6�T��_�>|��6��[\� m��ŲPsj�[p9mi�k��   � �h    �@8 k�� ���� ���������p���m��ām  m    H�[@6�  �8    �m  [@@ t  [@ �m[[%����hm m   ��&������i6m)n �f����k�' �����sb�;f�fؐ5�l ��l�A����m� PEm�m���۳l��� m�$6��IŴ� �yj��%X
�v�遶��� H-�� �  �H [dp [KoH� $z��Zl  �l[R�;m����mm��hAa��l  �`  �  m���۬� �  �   �   H   l�� ��� 9m�5����	�( 6��p/[ml�5�[�� 	
��5�Ԧٶ*�BB�k�;1d���;bImsIk� -�-�m6�BC�H ��e��]��i$�� 6�bK��hrô� �r�m��  I�`8 $9$�� Ml�S�sZ l� �$l��߄ �pm�`l$ 6��n  	 m� 6� �  [D$`m^�@�Ś���h �d�A��4Ʀ��3wŮW�X(��K9h�0V�l�<�xM;*�u�.Ҡ4���UU*˲��   8��z� 8��l-�,�U� �� ��&we�
������'X`X`      �-���  m�m�6ؒ� �  m� [@ �`     �' ��� >���U l9`�KM�h ��`[Kh�	�&�U���!7T��-[@�"N[v��l� (i.d�~�v_� ��  ��   @  ���� ��m���m��    $sm�  -��ׯSm�ݤ��a�8k[�m��d4QMI��N�Y�ˀ  h���m�� p *�
�J%U��Ta!���PT�T�UH=A�x��΀*�e���YY������̤�͑��N3ϥ�9�sA̽�R@�i�J�On3J��lm� �ټ9�eEy
[�e�T
^ej�6B�.ܢ�Q�� [@�l�L��8�vl�mt� [W���U�b���( ���eW�yj��@]�Ωj�动�^�O-瀪m����� �&�����,�&�JOϾ���Lݷ ��  �[mc�d�i#m�  [B�eg����Cm(R�mP;m����G��J��lp���)'ط���[��͚N����5�PlU�`�XV\�gd�K�E��`$\����� �kj������j�������(?��)El6�P�G�"b�* CH�C�KAԨ�$(�W���Ѡx�y�'�%��B0M�b�u�V����Pxpj���VG�<�>W�X$�9�HG���ث�D@<�|�+�^ ���Ӡ�*�"8 q@��<��8U07�@��Юt��k��k������|	A��P�2H�!Ȇ�,U�U���Z�C���v���Y	��@8���DF@�RD�� �B*��j<�QQ�T�T�X�>S�Z�@4�U!Zh~�"%N���A���(����^�	�XlppT
=S}��F��J��t�T�(t~�A #����U,x��E_�xO]��D�1~�� ����@�/��D3g:{�P����h� _7�G��O:~�:t �h�b�� >zf �X��U��B���Nl��E���+��b�A<'��Cb�"���>T�(<8��uTTW���� ��0 ���!�oZֳ33Z�@UW)7<$A&y��뉘����㰀��Γ7O+eZ��52p����#m��K'�^Y5\��m���3gd#c������;2�@Ol�^[�΂W���[JE̲�&�V��[2fm���#[n�ch5AY�2����a0S*K�P%� Z�b�lT�J�ka�t���Y1{��X�8{b5���q� R]Ν��\���go@l����ؽ�Bs�#3�DC�e�����g�V�lW���6�����iθ�
��Ua]��6+��kvӂ����m�6Z�#![�tuR�&E��퍅3��X)��r��N�x��g[��V��%�ܴ�_\iQ��VM��T��khp���ڝ���bn�궂 I��J�$��=�5qE�d@읪+�;b�6!PW�*�c���w7һn�\�l�۷P]8M2k�\�(�'����f����hx˰!��9���qi�G5	�3�:`�ѝ�������k=[��N}����s�q���hs��Tۓh8ɍ��rz7AdO'&�s+����\q�m�婞�]�����I���qV}*v�(����l����B���dR�]!2��H�m���R�\j8 ��&�\�;��vi��,�8�O#��n�jҍ��훣t�z�$`�J��U�V�ݘ�)!�uH`��cm�d�nY,m0rm\�pʬ2gf��<e�Ѓ4��j�Z�y�]WUPR��D��+�L��T�l�j{,]+(8�'�9���]6W�.Z5sz�6q����:�muBi
��ys�c�c���ggX闩V�6����[h��s`��6��s��c���Us�h�ym��2�m�V��v�7P+���i�*�n{x��vh,vHt��Y!�֌����ڇ�:4�ڄ����Xj��㧧-��mĳ�-�wk��l7E ��<¦��vA�1[�m������w���ES�
|�;���U�E;������i��P�0���KoXK��E��e{c��ֹ-��\0K�Tg���.Hֹ�ꂲ��2��n$�XŘ{=�s=ըb�LEV`�n��IӦyz�N�җ�$ˣ$ZsFt��l�β��JӶ�����ܗd��ǹxd[azwZr6�մع���E��m��e�:�C�F� �ƻ5�\��%�X��;�o>�:E�/&Z�]fZ]2"�^(�(�x�N�\��2�g�`ɍʞ\raw����\yELgN�b�عG
�v�Հ}����_�J��C��ٰ37U��eM0R�*��`�c�JB�B�TnSٰ;�ݛ�g�t�%8�%'�rX�zP�ܠ�� n�h;�����#q�(�+1�+�g��,3�UR퓕���t�Du#�$�V޶ �� ���v��k�LU�.9�5㫜��!F��n�؞g����2,שt��A�f蝸l�>�Oַh��P�ܠ���NB���3-̙���f��]��DG�0*�D6yD�%:�A#�CU�(}l@��:�9�wr�tԃ��,�ܬ͜Xgt�;6q`v4������2)�ٶ���~��߄m7(��IqvTӂ[C��X9��$�;�V�q�+{z���:U�:��F���q3Of�����7=�SWn�a�@um��E��WiN6IR	�����Ł������u`���>��)7M��R!HX�ܠ9�P�7[�}lS�}2v�)�	�8�JE`wo]Xgt�������T��b�*DЏ](ל�{77$�������t���IR'��fwK{gc�V��,��P�eH��r����؀ݦ�ϭ�u�@{�������������b�d)6c�u]s�����/vݓgӺ:��w��NmqQ4ӥ!�|������u`�����Ł���Sr48ERH�|�/DL�=�R�߄�7(�p�u ӁJJRU��;�����=������kvl����S�M��WH}l@n�r���B����E|�ڡ���S��'*s����������&�r)�,�ܬ|� 6w� ;]�菽ޕ�"f�*�x+�pk4�^���-�����u8ݣHN�:�����zK��{�/�#a��ͷ���Bg[�޶{ﾏ�C���@w/҆�%H��U��;��ٳ�1�+�z���|���T�HF�r�z؀ݦ� ���ηHu1�5-����)�9l��P�!*�ovlgz��ŝ����Ł�Үꔜ�4���s`g;���������=,���]�7���5�:�S^T�ŋ	�n���r�ߒtз16��v'y�Oa�GN0�]��yu�rV�]3N�Z��k�'^fGlK�]!Ȧ���vJ9�Mt�Mh�Ol��u��Q������:�n-��<LC;��/)]��#�䣳�c<���),n�rn�&�if$��Rd��؏B-V{g6�������k��P�Filt��,���Er����@7��8����Ѻ;4��I��y�wqt;�1zyjf�=
�ܘ��ؠw�'�wOe�!���.���sڔ$�S��
RP�%h^�� 7i���2A�j÷Í�����ݜ_�$n�yX�z��ŝ��>��)7��ȤB��7i�@=mBg[�� ;zm�6�	5#�$�VguՁ�;��۳���̝���8�R��"�*E�:� u��M��j�";�����ߖ��Z[Jk����v;�q�k\����IӐ��ak����D�7e��YE�]`n� 7i�@=mBg[��ʻ�JH�m��,�ܯ�D���BN��TM�^�/΁Njk����>���nI��=7Qm;U�R����jB��X��V,�vn�,�ܬ�z��R8���mXlB��wj��ǥ��Vd��˫�:uD8�$Q:�i�`v���؊J";�͞�ݵ`s1�;���]\��d2C-$5������g�WK��_Jm�1���gVX�a�R}$ݮr�zڄ�ݠu���wN �N8�JE`vw]_�~H3}�`{�x�3�>�'T��	�QI*䓟{ٹ'���ܿ��A�1? A?
)�U3��˹'�~ٹ'oz��7R%!�3�3�>�� �;����]å$M��ەuw(��(�� ���\�������9@Z��l�gkڹ��n��G��<!�y#�ͮ ��L���{��|,o�:�I�!MȾ3���>��`f=�`f=�`f�Qt�@c�RQ%X��,��(��(�j���"d�z�%[c����k�+1�+�޺���X�>�Dr8�R�X{��
!&�(����f��3mX��v��RD�#�����R<���vݤ�I�m6�D����7��U~�Y�����Vc�V-����'�h�\��a���k��z�>|O��秶͇��8��a���^�*���O�����6��6��7��O8)�U�̶2�-��Wro�'
!(�9�͛s�u`f��>\��t����#$*�P��P�� �v�ͮr��iWuJNF���
��`}��V����PW�Gӛ|���T]�U�U�U� �v�����8�?J7�j��	*B�Ing�jI�0���e�ˈݶ��v^M�O7OS]
��I�Օ��8'i��tNiš0i�ݫ�K	�7jfz�[��]���s�kSl��zҗ5b�m�/\�V�atj%���4���D��vq�B�]T����b�um]�&L�z�?ϟ��5mj�P��c[��:�w�&7ccv�a��c��ɶ���[��ó�3zR�.�=�~w��ߞ���e�u��K���#�}�Gd9�u������*�㈽�ڌK;nN[�p2�H:p�p������>�� �7��n��Q�G#�H�$����@f�P�3y�6�ʯ��#�_�p�6�D����޺��zY����K5���������uJn@��*Eswp�3y�6��6��7���A>�BD� ��������ݝ���<X��,\���2R���[>m��Ņ�N�N#��s�-�����L�o>����sg���B�h�����@f�� f�~��$7��P�f=�NF�I��nE`}�8���R��~�T�7�X��X�yX��]:��N\UX�3[�ms�T}�DL��9@fl���N��'$�4�>ǽ(��(޶ �� w:q7W36��:tʖ�����	or����K�g�{�<�<��T�j6�*z��0\e�i����B.B�'aes���r(�R9�M���j$�_����>��`vu�(P�C����s����ܡ���Ո5�^��&Os��~�޶X������;6q`}���Ļ&��!V$��a1�Hv`�XA(�B�#,��#
Z޻��T�V��#:FA�Ю�̨�bf�4�`�B&("h�`�H]H�����H{�C7!&k06�ărX"������۰��U�cFA�%%��B�,�iR!e0�KA�b2 H��I%YQ�J��D�+$�*�!�{��0X@O���@%�# B�J�$(J�$F)�(@���H����0b�hKb+�^�&�E`)�����F)�X���}v+��tQC����H�Q�B���}�98�} s7]�	%2sjV�Զ�uN�ʖ��B��^l��zjJ#���v|�(�LlD"����7*e{ɩ��i��9?"�3{��~�����B��߳����q�`w��;�����e�ӖIUR֣�6�Y\kU6�Δ�'ukj3uڴbBXr��塪M�SM�J�}�
d;��>������fϒ�}
"gٯŇ�DD�O]yLӥT��EM7`oq�~P�Т"Q�[��
"gٯŀs��R�yB��w��.�̶���-���Nc�M��%
7�z|��6"���=,nZ��QRSU��S���=/TBJd9��`|�B����L.ǒ��H"?�LqU:����s��~��2{pz��m�e7L�>Q<�x�<���d�u?J�}l�1�,���n�v���v'9֑Pf6�Ѷ�]rth2H(�r<V6�*6��i֬5��<��u?J�[kv��Sĥ$n�nBA�1�+{z��>��`ol���iWuD9#�7U%\�9�P�3[�lL�v��s�n�N�)�PN��J���X�8�3�7�������q�c������؀ݮr���BD���h��{��v�6�����_����ƜK2ц����v��<C=(�j9�y�5���w3x��n���7�\�b�����\N�#��	�09'N�n�l�9L7X�ٽ����b�r�9�M�1'����k��g��^,���-��Uc���V޶0PqŬJ�g.8Eح��ѱ�m 	(�e嫢-�	f�n�:I���:7[Ck�-k-�&L�����M6� �Sʻ�;�5��3b��Rޫp^�������$9�M��Ȝ�fٻ"�
M���՝���%>��ɰ3smjJ>�9��ߤ�DD���,�қpƇ)��W�ߪ�;����~��~d�[��7�_�✔H�T�7%_� �������� �}�`w��V�D�qER��H'"�[��P��A���� {ҫ�%)#r7 ԅ������=�~?����,oOi�>�NS�$�R�H2�F͖�te:1��vܜ������e#J��S�:����Vf�,��;9ׇ�">��k6lfj-Rl�l�5�ɚɹ$���o��+�{�K���O�oq�z�Na��I��p��jI`{zx�$f�������ֽ���;�Ǫ]B�m:ں�>z�� ���7������wM�CN0i8�͜Xٽ,μ,�]ɰ=7oJm��5)�M��ŮqAoQ�JWA��`�{t-�d�Ȗ�$y��QL�J�ܔBQ*D��� ��K{g������u`z���~��Ll�����@n�9@s� f�h�Wq)I�)9��3�7����@b�Y�1]q9��2X��X�*�S�:��ک%��[kv�����7(��E�M�.�T�K�X9��Q�y���ń����؈K����ST����^��鉥ۭ�vs�5=W�f0��N�"-�:��'���#_�o������1�+�g�wK3gR���G�Rc�V��,3�X�yXv��6�q�!�X�8���ϭ���(�[������%H�n�wK{gc�VTA�	��."��,�2�[
� 塪&����؀ݮr�����ݣo��߿B�y%�s��B�d�3�;,��W]��NԒ�&�nӺ�V��<T�l�M�݈��(}l@���[�*�S�:�!O�H��X��,�X�yXV�Qt�A�8��ub �n�k��7k���������ԑRi�`ol���{����Ň�RY���7zz��
$ �Q�8�Ǽ�͜X��,Ǽ���pۤ�eJP#��I�)'N�óY+���P�h	�`Rjt)uQE�-�6]�T��u�H�;rO5�Cn�nQ ���Dm�=��Ḳ�n���.T����Y�K�=�9��5�?�G��!���@����Yu��/N�-�ki�)�컝Ҫ�f8��9�ۈ�egu����lE^��,�!2����>�G�NTN�d�5#lH�����ى�n
B�梫����"V���nͻu8ݮڝ�ˏ8y�mўk���tӐc����� �n�k������~�6_�7%E��&�,��ꪤ�k�+u���ٳ�s�Ґ���D�IWv�{\��M��[�v��ʻ�JH�"NAF�,=���=�`w�x���`ol���iWu��ԛ�o뻹@s�b �n���@n��|�o�߮�fN�Z��{B�7�4�qAo6NꎇN�ڐ 9����9K�Wk���
	�� n�h�l@n�r����s	u�K��)Sb����̵jQ�$B�W�U�����[�ܓ3g��,͝JT��"���@n�r����z&N�z���މқp�ۑD�Vv�,3�X�e�P�{׻63G�*�NX�e����@��ϼ�`��J_5�����^>ss�Z�eB�!8�����k\;�t�͒�=��:s�r�1�e�b�(��@v�bv���j�r��ʻ�JH�"nA��X��_�B�;�����vy���Y��luI˒\6���� �3�
PD|�+��D(/������.wj�c%@�))%Xgt�7:q`f>�`go]X�(�
:��Ӑ�7%��ш�nP㭈u�@����*�����0W=V��V���d�ӭ�Nx�n��,�����\z���O����nP㭈u�@v�b7���UXq��H���ŀfwKs�c�V���Cq�P�)t�,u�@v�b=3�^��;���8v��"�FR����Ł�����w=7&Р���t�3���ٹ'o�^�J[uLm��e6X�fM����-�� 3=�`w��>μST�tIRS5K͹3�^�痩�7��Gܖ8�{6�.��ю\sI�MʻCM��Un~���`�c�;�xyDG�A�^��Y�E�M���U)�,��w��"����`fW�61u�{
d��.�Itʒ�4�*��3���9�̛<��GSy�ߋ �����u▛���Sn�m��)�^��ՏK �3��!G���}���j~j��S�t�Է61u�`lD)�w_�gu�`s��6Y4��!BU Ht�!T]) XEL��z���� ���*D��,J�`�*;ьbFP6i���2�" �a�JiRb� �2 2
��M}��֐&�֍�H''�A���	�$$HH�F,�`�}�`�ف,�ѥ�#�)bh�B0FƄ���&�A2
�!¢V��D F�1R`�R�	��Y`�d!H�|� �!����A�N@�����XH"A��bD�@�B,H�"H�!�H���;��ͫ�� m�m ���[7'�c=rO3�n���;j7K�5��Sl���ٵgs�c2p5Y�5��Ź��Grm Up�AC���j�N��X�1Ԡ��(���n�^� �d�0��2��{hYa��0fCS-U�s������ZS�m��H�ĸp���F��[Y�gh�@u��s���*���!@:��Ʈ��nn��YA#�[u���ͷ��K�ݸlu�Ԝ�����s�'o�������xpt�;1��<rpҩ��fG�cR+ :
����5��m�vP-9�\[l�ae����h�ݧEmUv��w��	Tr]n��U *�,`q��X)�D��yѹ�<���s��̴�i��c{�;V��B�]�tp��nEY]��\��8�UŜ��XpP��n�<d,=]'X��F2��
�Q�F�h�Ly7��f��0�l\yt4�����3�4��`�)w&x�&9���|�|��4p��� H�ݡ��؝j@u��.����գF��*����Up�˞�nؖ�;b�E�G2v-C��,σ�q/�9lF��õv�oo]�u*�m-�#�>y�-�� v+ګm�x�50��y`�V�h&'���ڛ9JL��Fr�=����z��� n8�q�_b�:ᩂٛ�&4�vU�H�+��-�y�M��v0Y���j�;v�a�9�v��Y��6��wC��2�3��9Z���ȪY�.�96����us�[`�EJ�����bM��j��J	�+n��]l��М�Q��!��rʙ㛶�8*z:�9:֣-�]	��`��.ݑ�ݱc����s˺Q]�*L���J[F˭�Ӳ`��^M�m�H�8��Vč���^�k��lq��!��ݲ�J��
�/��M�n�r�0;`���;�h���u"n̹����6������ɵ�&Pg���s�:�uS�;v�����:X"񆭭u����CaaۘA�l�3V�f�]��"ʍ�iSn�`D(�j�G��Px�T8 ��CT��k4I�(Zѧ��ڿw�7|U7r|��&��&�������Oi�c��v��2�0e��2g6��U��7[v��E��ק+���J���t�9�v����sԘq��y�g$��.�96��(W��!�3��}�ֺ��+��s4Y�:��&�e���[Uӝ�z-��r��f	� � j`�aۇA.-�3i\p��z�W�9��{�����KЭ���v���Ƈ��;]�mI����_;e�b����a�=��Yw(n:�D�"N�� {���X�8�s1�%��ǥ��ײ4�S���Ze۰;�x_�BQP��6��3�� �3�D)�gen���Tܹn�P������З�EQ��;s�Ł���4��P�jF۰؈�����;��`w���S=��8���T�nA�U)�,��v�����b0�޴��b;��Yp]��kP��S�`9����0[�ң1��9�;�7+߉b�У�QElnO����`�c�9��G�@f{�����-7iʪn�tՀs����J"SV�
!	D(���۳���`��`w��(��Nw֪��6�m�t۰;���ݣ~��{�� n�h�[�*��*�JD�7�}�`w�x���a�	D欽,�����#L���ϭ�u�@s�� �����~���tl�R��ݱ�O���6�kup�hێ%�kk�`sw��G|��*Z"R5�����7�g��3�ꯐot���r��%HH�Q�Kz�ؽ2�����@��#����؛rR�N�`�c�;�xY�
"��"l�ݠ5ö 3�t䪻�&�!�7%���u���zXճ���y�36u)R~$��9#$��}���ҚXf��7:q`o��̍ÒIJ�]'B`�����f��4qԜ `�xc �E+�r��Q:���m��{�}�u�@v�g�;��@k�~�*���9IH���`�����q`���ܭ�X�9Sq&FA�I`}�l@��6g�.؀7[��0�Q-��M4Si��$�)�^��ՏK �3�����D!'�_7�'��(�!#tF�r+r�q`�����q`f>�`u,މ�*GHiƤ$[���t��5V�ΖxDޝ�I�B�lHcS���TJu!RD�5Q��3;���l���}�+��'�t|��lQ�������ި���Fe{�`n-~,3�X�:��?�(�F�3r�7+gy#wޖy����mN�ۀ(����`nV�,3�Xs�V��=�`o���7ENRR$�X�v��7�F�^��5�5�b"�� !1����j~5rdћ���u��~?��-Rg&�i�����Uq�%�Ck2d��L��iu;��Ƴ��enn�X�u�T�;G���=X�y2��-�'��@փ�խ�&�H�]�թ3���7^�k��*�7t��>L����;���<v�z��e�v\�+>�2��|'�\���*���v�(���kjk��=dr&��,�9��Ͱ;\Ա�W
!B�i�_�-
m�m��eٹ��	��gF��\���aG���!��%��%�D�M�H�)Pc�������}�`sr��>�;��`l�Ҕ��4�M��X�fMꈈS'ufڰ�u��8��H��^�J�q�%8܊��C��ݣ�/�~��J#y�j�bt�5*�6Ն�D�{���,r�&�RJ�Vo����f��m�MKN��n��1�`j�
;׻?�Y�V��,�TsG)#�rR�!zm�{[�m���iY��ͳv0Em���wϗJT��R ��7��~�3�z��9�Ǳ��C;�K�����`��U4���.�J�FyD(�����~,r�&��QGw��ES��SS-�ҦՀf{���1�f�Q3����՞��7:r%Jn"D�*rK~]������9�@�� ��6TM��2Zj�L�>�fM�仫7��{���N,�6.qE �*I��D�U�˺L��[\F��F5rZC���+k���\�::���H�D�?7"�3�z��37�����Vd�.wj�bt�5*�6� ��k�D}#�_��{Ҁ�� >ӣ�ӑ�M5*69%���u`}��l��	�b\_}�N�X��;���R��:�r���1�+:�����v���X�n��`ӡ�vMܠ5�55�@v���\��}���i`�zkKn-s�z�JD�m��m��#�v��n��N�ۊ�h:lܽ�1Uw5�@v���\��9�@nt�J��QT��S�I`nw]X�ܛ�����f;؈�6vV�J[uHpr�	!`n��3�z�������;}<X-U����mSR+�����qXs�vy�	�(Q�DF�3�l���Z�9R��Jn���5�@osV 7k��5�[��������{���f����=��ҋ�73�E�e�N���UJ�9��o���ᖦ�K��j�@���Bv��\u��d���Zw��J���J)IHrU�����#|��`��;��W脼�����*�`9d�í�Z�X��vy/%[���2��`}�4U:NU0t�R����w��@>�� 7k��5�[�9qEQ�!M�%���u`{���^l�uc��>�c�.�%�Y��������%r�Hy�pv) ����[�5��?��q�HuF�ct�RC�Æ���9z,v9��g�6,�)q�cAbݣ������4ָR��D�vR��v�Y�����>u�=�'�Ҝ97C�"���b:���Ͱ�i5n4[΍���\�)e����ݜ��L�m�Z6���X��ѭ�;����e4Mf��4ɟ�A��@�ߎ^�ٕ]|����ոwM&�9�nm��u��#d�)ny������:��*^ٵŲ��n�l��ׅ�}�Ǫ">���ڰ1r�x%9N6�nB��Xճ��UR�wu�G������ٰ>�q��T�cR��4� �����3-Y�)��������,�����ӐM'%��$�;��;�͛���ԡ)�wޖ�OR�'�$E)�J�3�5(K������vy�j��,͛�(:ӷaC�o5v���I�svݛnD5��mN�@�n8�mӱ\��΍u�~m���� ��h��~�>��ާ�@k��������UL���wJ1D&��ʱ�	̞��nI�u��rO�vq~������d���Ӓ����Xr��g��䢫<������9+�t���))(ʰ>Ǽ���ŀ}��Ԣs��+���P�4�T��lU-́�]xX�"y�����V�{��3���>�7$rF:Q:Cw�2�v��y�޵Vä���@�T�M:qRQET��Jwh�Lr��m	�SL���vy�j��+�>���B��Pg��t�ITۤ�*tML������(q���ݯ��QFf�)i�*�29j�mX���������P�8�!$��! ,BV{E!$�����"7[6EMH�w��4�p iWl��8����9ͧ��f���1�a�����{���:�D+d�4��h볂	�U��n����T��^*�W6�j0�:�#��zWO��f_5���:Vb��C�#%�Nl6J{�/K �w]��fZ�9��V���Cq�T�7 ��X��,�����/��k6lb����o����e���أp��ح�Dtl��1h��&�S��ۗ���?#|�,��j��o�n{֬r��`s^�IW��\`w=�`z}+<R��T���M5`n�9@wG[kv��څ菢d�ʽ�%HHډ�
jE`wWO�v;<�]��j�̭���b-67T��uV ������(}�~���Ӿ,�c:��ICq��NKj����~kv�3z�~���Y���)��g �Hl����h'�|��g�7YN�N�=6Iy^�蘭��r� �����7U`Qqqd�5r� �����1�+��t䨩�nASp������L��s�tu���Lh�uC�*�7-�D)�ٰ;�͛r�q`gt�9r��Ғ6��*��P��P�!�5� 7��@c�s`J���DA�A�\�RMk�d�4�4�A0OZ��'aL�lܛ�yF�䋍�˒5�c�und.ܯ���o�5�ޝ˓&�q�҉��W:�kp	���ծ2�q�ۥ�5I��9����d��`6��=Q�q��Fҝ��C�Zh��-{a����)�@泰���6�9*�*��[9Ͳ�6��i� ���N�瀧�[�m�$���tv��u�����rn�+<Oi:~�ǻ�{��~7T�g�j��rg��痪�o=8�794[	�6�..���#�k��MD܅5"�=���,�����������wQu!#`�J)���ݭ�5չ@n�9@v�[��qNBI��$�����������Z���v9׊Zn
m��)�`f�9@wG[o;@cmB�M�S��J��qX��� �7���w]Xc�V�*�҄�i�
Q"����� t��޳F2��?~tӫ����fi�6�[����M�����>���{��ݭ��z��7(r"s7$��?���Q�<S�r{Z�+r��V�oK ޮ�Ғ7BR\MU�6���9�@����-U��G)��"��Xm-������q`,��@=l]�uA6\M�QWp�3y�j��Pѽu`}���	�Q�$N!4�
J���c�s�<��_,��6�sqn�[�]r�iD䉤����u`}�yX��u`f��>�g)R~�*�P��{���jo;@cmB�M�U\C�#�L�s`w��j�>�q�0�T�"�� �DH��P�d���u`v=�>�'@nJ��4�Ip�3y�j��P��Bj:P�lP!N'%��w]Xc�V�o]Xٽ,	Z�[t����R�p�μjÅ�F�;N�:�cN��v�6�`suF�AҒ7@�)Jm��׼��ܵ`s��/�9����J��t�*������tsP�3y�j=�ϼ��x.�lJ)JӒ��ވm�@f�9@wG5�t8��*۪�N\̶�6"S���X�f́ޮ�f�(ƃ�Z���nIϧsŕ%IC��J�>Ǽ��޺���XwuՁ�F��T�j6��QȘ/�����2�t�:fK�a��1L�VQEGN���ݭ� �;���w]{��7_yX�'�7%D��$I) f�h��@n�9@>�j��t���QP�*E$�>��1�+v�q`gt�9r��I	:��:���s�tu� f�6� 5j���*9N�e5"�7kg�o�rN{�ٹ'>�}w$�Eh|�������c�2�]��2�m��H�����y�-˷�D=r2��g@���јg�1<�W�	k"t-Z��3��p��s��/F>j�4T���g��魯WN	Jv2��i��1<[lX�Q�u�1�m�H@q�[�]�j�1�j1�չX�^�r���Z�����C���=\f��=ɱ�l53M&9�G'���Cɹ���藯fg����wn��n��r~t�<dd�F9��+
���Jt+��۞�c����N����RD�J�q�(�&�8h�}hm�@f�9@wG[��qUwRۖ��ɚn��3-_�L��f́���`f��>�gR�%4��SR�%X��P��������@=)���(��ӂ�X��� �7���nZ��μٰ;�=aT�sL�n]J�� f�>j��P����wJ��V��Shm�m��TM2Dܢ5���mj�:�8w[��7>,��Q�*�eAW]�]��ߔ 3k��;c��7��9r��ITd�)'*�����W�TB�U��ֺ���vs2Ձ��]�*Tr�88�jE`v��,��vy%���vՁ��l�NN`4�N�fn�&�.�@�� ����(����莦�q��F$�>���#zߧ n�@���s�����56Vŝ�����5�g�pl�61b6LB��vl��T���;Ztv��蘭�\��l@�����7W��(�8)��[8��zXwuՁ�=�`}�N�ܕ�H�G ���`}����	%���J�E�S�;+���ؗJ��H���NKħ���9�͛�]xXyBS<�k�<���$��$�ە`}�yX��5� 7�����u˫�����+0aj��Yɵr��5#�Z��^.Z9��7�z>���]7<ٝ�G����w��������(�����TL�jjS�XO;�~K�*����X����ݭ�XoDu7#mʕ%H���6� 3k���DL�� 6y��a��J���TcR�%Xz�,��V�{?M�9~ﵹ6�� ���Q�{]�X��JN@���'R)��[8�=}��Հo����(�n�b��;b6NnI�]<Ymr�[��7ic��;�;�O�/�9���l��͆��ͷ�����6� 3k����$�~�s>����JIN'��t��������Vut�`|�y��G��{�D�:J8���5`s��6z��ВQ3��mX��V'����jSj��Ksa��Mx@l�� 1�����"w��P.}�� 㦈�&�8X,�v��ud��]�ܓ�;���|�)�ԁ	#F� BH� �EP8���F
�m]#��g��	.����A=~�}�uv���1�H���k�d��	c!VaX(����A��Y�䄨q^� �t��"�L�`D�a 4�(D	�*��	�6�j�0!�����	Q��D�@b	  BHA�"��$HT-t��H���HMQ)f���D�:4�!*B��JV��!Q4Zb,`�} ���BA�&� �#c �D�!"|�1
KC����a���E��!0sZCB��$��u�����w�?_�߉���;m�3��SF8��N�t�,0��q�ˡ�$����VLJ�;;N�[W.��D.q��<�`��Ӷ�8� *�G8�AcZ��;!���1�9�v��F9e�<c����fE��۵8ٸL6d��U�U�Dw��^��m:.[X�a{Z�ۍ����l`�y��pAgtf+����뭣���z���j��ҾMt8;g�.u���Q��l����V4�K�䭲)��M�k+ZX���̒�g�^��J� ��q.�#�ǈsv�8�f
�v�z�\�&F��5��mTi���U�j�*{*�[+j��U�X�'4YZ�۱OZ�=,m����;8��Z!�6����Y+n�I!��1�+r��^���b�z���Xt�U�+�1����7���I>����;1�"���N��q��1i���}>��-lv䨩y���%�{�#��W��*`����)�l��Ǉ�:Ԁ�ب�)I�+r��P�N�Һ��ӹ��6y��Z�(;�ձ-[�B��`�u)���滶��Y3�.�`; ]9�yW+�����K�![�Kns�[SW]<mI-s֕^�V�WT��\��n��v��ݠ*U�TJ� ȏ��ce�&�h�[]������Z�K�t�����;e�V�<4�5F��`.T6�s��y�v�m=)�j���i�&��i��g�f��e�S�vzm�lٷ��6�-�4YSv�m�M�oMT6���m@�d8�k'dN�C��8�g�ɑ�����\�N��W����W6�Y��p,:f�9���M�S��On͓nlN�$�u�ͭ�6���Z L��g$ꎶ�$p)L�ͮng�@�ч�dK��"tA��S�58sm�t�r�<�$l�˲�b+����6�	�J �����l!�B�W@�\�NCg]Z�rK�Z�1;�FYM��R�n��(km�Ϥ�u��٠�GVx�����=��`�]���4UF��:�� �G�G�Q;NtT]�P�"�Dԓ���4k�2�j��bt��Q9k��#p���`*�ޒ��[�q����.�{q�.�}�2�;i�b����5g��(�m�Ѷ���q��9.�uւ^eK�4��1#4T���ì6p�:Ct.:�e�����.8\]��s���jSY�����.���@q�gV��N1a{5zP��q)��,���v��sF�6΍�%{Z(�3���zw���Őf:��cte�m҃�d�ۭ��ܧ8�uHmJ�EӶ��;���O����a�qfiց�ݵ`}��M�ޮ�6!BI}!Ž�`f�=JT�Ғd��V����ޮ�,��ʰ>��W����G�e���hBm˚M�s`n�~,���`}��V�����>�nJ#�H�&��j��P���ڰ;��Vܮ��j�Q
z��f���֊n����mS�t��mB6��ci�@d�:@~���{�����\z%�u������k���5�9gv�H*(�kn��_N%������y����*SnV�����}���f�3;��Z��%H9J����VV>뽟!�ʃ�;jxO�GY5/�U����`}��M�B�99;��e6�JT��qX��vgu՟߿R[����~�>ވ]NH�q)*D����(��w�`w��6+2l<�O+��`fk�-6�e�ERpSj��+�6�ul���b�y���V�)�SR�9*SQU̻���<kq��vm�V�� .�x7��I�I�E$Q�E"�2��+�������� �}�`g���ܔG$�SN+ �;��U~���z���}�`ec�W�T��藠9# ��"r\���훒s�w�rb*GD������kvlsq�NJ�*Fۤ�Z�����5(�^J�����+ޛ ���`fw]X�WpJ�r��n~jE`dm7(N�����ms����)�oO-MNx����y{Uü�w3��㳛��:.���G��V�Ve ��>m��v��mB6��ci�@g;��9�Ƥ���gu���3_yX]�ٰ��w�P�&L�z���L�©8)�`s��6+2l�P��Q��;3޵`g{/���&ܺ��nl==]{�`�k�9��V������# D�#����z��_�����X���SrQhrG(N+ �5�u���(������c���av���!3Fy�68+�g���]���nq5�q�W9gZݴ���so��&n-����ߔ 3k��66�����eJ���C�ӡ��j���ܛ��%Tb����)���v;�j���V`5 �'n~jE`ec�V�oK?�U%��]X����.�� �j5*EI9(7��3[P�ͮr��D�u�J;���M�:��rXguՁ�=�ܓ��w�rIϽ�ܓ ���^�����ĿO�"���ǧ�:��.�����،N��f�IHݩ��i1���Q�.r9�ص�[hE�Ԍ��D�R���!k��7nx�km��s�tE=I��F�8�X��-�,��{&���d���ծ���wj�r�5�J�;s�մ�m94sw(طk��6O�z�^kq؜܄��e�e�ks)�-�^�w\���4Yu���fasV]B�zT���??��R���Z[�ܳ��S�Z� ��V��W���,��+���+�붛_����.Wrl�f?B^�\���Z�=�/�US@��3C�nl�+2o�DL�;���6Ձ�Wroc�T{
���(�49#�'�oK3z�ͪ��_�r�>�m:M�2�m6�z#��o!�^��66���ݠ1Ԭ���tK�覦i��������~�y8(X � ߻��lA�lll{�o�؃� � � �������~�����KS�Y���xj����<�.�8�ݛpM�qQ�l>#�k��n�f]�<�����s���A�A�A�A�w��؃� � � � �����B
��A�ll}���v �66
Q"��+g�CM��L��ʙ�6�(�lllo���6 �#�b�H���� � �����A�A�A�A��߮�A������؃�
*CPR�%(J;��<����i�ʚn� �`�`�`��~��؃� � � � ����b �`�`�`������A�lllo���6 �666>���.����֌fk&�A��D,{����A�A�A�A��~�v �6667����y���6 �666?���kZ������\˱�A�A�A�A��~�v �666����f�A������M�<����{��v �6667߱����f�P�)��y�oY�3p��ߗg|M��vY��(���&�Fk0v]e���lllo}���y���6 �666=�{�ڨ������߮�7APA�A�BQ�˙��6�m��iԶ�BQ��������D�b!� �6>�~��y�?���A�����߳b )���PA�l��r����t�-�4�l�	G�A������b �`�`�`��s���A�� � �ʁ�C������u�ϳb �`�`�`�����M�<������?~�ɬ.d�X�̻yB�����b �`�`�`�~��ٱ�A�A�A�A�}��b �`�`�`���]�<����u����fMf�5&��e؃� � � � ߻��lA�lllQ���6 �666=�{�؃� � � � �����A�lP�H�(�BQ��ߛl�ے]9����ҡ�1C�S�,ע�m����L��ge�a�f]fe�d��WY�y���6 �666=�{�؃� � � � �����U�lllo���6 �666>���.����֌fk&�A�����~�y�C�D29~��]�<����￿�b �`�`�`�����@S�@ ���P�(�BQ�ٿ5ULM7UR�[�H<����}��גI�~��>�gc�V`��n:#�H��V
g��v{�K����(���BF��
>�IWs�l��s8��mS�*���n����菻��p��� f�|׍�7�����?Mq��MSO����)�U;m�N�I��zм�`�s�7qZ6ff�SY5p�̛ND�,K��z��Kı9�{�iȖ%�b_����9Q,K���M�"X�%�٪~�&�ɬ.e�X�fZ��bX�'>�z�9ı,K���I��%�b}�w��Kı;�׭M��TT�@�%���}O����̤P|�~oq��%�}��I��%�b}�w��K�T��j'���jn%�bX�w?~�O��7���{��߿rУ6��}ۉbY�D�}��iȖ%�b{ٯ֦�X�%�ϳ޻ND�,������4��bX�'����a�nau��ɴ�Kı;�׭Mı,K�?�W�����v%�bX����4��bX�'�w~�ND�,K����ʃP"�?g즬�Zh�d�5m�汑�B[�ϗ^l�^�0.��/gV�u4ݚ�zʶ�Z�wf������z��S�����p�d̽�c��� �PaJ��ծKe���u�3����g�U��D�6�:��i�$���q �UMp<�h�:�xi'�6�=[�n���ɱb:b�ֱ��x�i	��(�v���nv��=���k�l�nAa���w���[��o�Ur̫v�CnD�M=e�wM�׍`ڤ���ڶ���lU��v�����Kı>�~�v��bX�%��٤�Kı>����O�j%�b{ٯ�������ow�����vY�2%L5�r%�bX���f�p�@��j%����ӑ,Kľ��eMı,K�g�v�������bw��kY�:eL���B����$.�/K��
bX�%�u쩸�%�bs���ӑ,KĿ_{4��bX�'=���Y�����I�.�&ӑ,KĽ7ı,N}���r%�bX���f�q,K��5��?M�"X�%�٪~Ф�MKd�4�m�+!I
HRB��2�9ı,K���I��%�b}�w��Kı/{�eMı,Kƻ�>�jx��Z����)����;�=,>��gGNz����zmr/��������7+�۬�O�X�%�{~�&�X�%���ߦӑ,KĽ?�����*H\�ݛ��
HRB�snGE7.��95�j�3I��%�b}�w��4ڠ|�4�b/� i�MD�/���Sq,K������r%�bX���f�q?��MD�=���\3[�a���M�"X�%�}�~ʛ�bX�'>�z�9��T��j%���4��bX�'{���ND�,K���a�f�Z��Je�ʛ�bX�'>�z�9ı,K���I��%�b}�w��K��EO�F�L��_�Sq,K���_�*�!ө����sp�!I
HS�}��n%�bX���6�D�,K����7ı,N}���r%�$)!lD-�Ҫ�7i�@�m���TK��qu֌E���$��۵�ړ��Ր�J3���q1�&��T銪��[u�)!I
H[���iȖ%�b^�^ʛ�bX�'>�z�9ı,K���I��%�bs�O`�m�eT�SM�����$)�k2���Pc���b}����9ı,K���h?�Ț�bX���m9ı�{��;��g�����G����d�9�{�iȖ%�b_���Mı��tF	H�4C�Q��C�|�Ѐ�"@����M#$�i�,�AXhq�.��nT�SuZ ����A��[�}�A�@�(&�B`e�c�b;h X�:q"B$�q�t� ��W��c�5eID�!��g~��T�>�?�Ъ'� |�xT��E�>�?��+����x�iW��:(�(��O�s�o�iȖ%�b^�^ʛ�bX�'�����2k54e�5m�]�"X��D�o�f�q,K��}��iȖ%�b_��eMı,K�g�v���oq���?�~sR���d��n%�bX�}��m9ı,?��T�{�����,K�����9ı,K��I��%�bt�v6���as.]9�[�Z^��Q�=X�q��`(-���3mfkuW�7=>�~Ou��=�{���T�Kı9����Kı/׾��E����%����ӑ,K!It�m:m)R��9�����"X��=��Kı/׾�&�X�%�����"X�%�~7���aQ
H]�/Z*�!�u4�9nn�+ı/o�f�q,K�����ӑ,KĿw^ʛ�bX�'>�z�9��{���}�}떺�p�����x�,��@�N�߾6��bX�%��*n%�bX�����r%�b�wo��3��.�@�,�Nn�y��Kı;ܧ�2���L�&���r%�bX��ײ��X�%�ϳ޻ND�,K�}��n%�bX�}�p�r<oq������{~��Cs��0����2m\���H�i�N�w�����f�=���wϛ=t��-�*=���7���{�����ND�,K���bX�'�w�6��bX�'������%�br�9�i��&�T��ӛ��
HRB���٤�?+D�K���ND�,K��~�7ı,N}���r'���{��~s2�͵�}�7���%�����"X�%���jn%���MD�����r%�bX�����n%�bX�v{~.���0�L�6��bY�"��O{z�jn%�bX�w?~�ND�,K�}��n%�`�N�7��|B�����m��ST���su���X�%�ϳ޻ND�,K�X����r%�bX��p�r%�bX��k֦�X�%��bIOʨ����v���ͫp���[l��*�n�u t��٭8�F�1�֎�gf��]#d���Ɓ��S���\�6�#�s�+UnyD]�e���9���=[Tˋ�q�g<�i&)3����#v���x�q�����
]��k����6�Jm��7b����K>�4���c��>���Y���mC���BjP�v2�;\5��T2���)gb�J%D%E��Ժ�CW�#d��x��dl�k�7l���.؃�;[[�������6n�j2��{�s�g�ı/����Mı,K��ND�,K��z��'"j%�b}����9�u��=߿�Y��lvd�(�狀ı,O��m9ı,N�5�Sq,K����]�"X�%�~��i7�:��RBxr6�2iKM�t���Kı?~�Z��bX�'>�z�9��!���{~�&�X�%�����"X�%���=��f[�c5�jn%�g���O��߮ӑ,KĽ��f�q,K�����ӑ,K��s^�7ı,O���ə�ur�5m̻ND�,K�}��n%�bX-}���6��bX�'��?�Mı,K�g�v��bX�'MzWG�.�,�1ל�6�˦��5��ǝ��ܧZ�c�n��m��n�Ւ�e����}�7���{��}�p�r%�bX���J��bX�'>�z�?�Y�MD�,K���i7�RB�p��-6��6L��髅�
D�,N��M���x�D�����؛�b{�~��r%�bX�����n%�bX�}�p�r%�bX����ְ�j���ֲT�Kı9�{�iȖ%�b_�}�Mı���MD�}��ӑ,K��~�7ı,O�ٿa5��̷Y�.e�r%�g�Q5��٤�Kı;�~��Kı>��J��bX�5�����K�q����7�\��ۆ���w��7��b}�}�iȖ%�a�(Ǿ��*r%�bX�w?~�ND�,K�{��n%�bX����Nd˅r浙u��d��m��k���5���`�r&Mȶ�=k�7d�/dY��������fm9ı,O�sҦ�X�%�ϳ޻ND�,K�{��$�MD�,K���m9ı,OMS���f[�c32T�Kı9�{�iȖ%�b_�}�Mı,K��}�ND�,K�������U5��~��ufa�P|�~oq����O~�&�X�%�~��ͧ"X�%��nzT�Kı9�{�iȖ%�bw����Ni7I��T�����&���Mw���ND�,K���T�Kı9�{�iȖ%���Q5��٤�K�RB�z���:���S�[w���K������%�a������i�Kı/o�f�q,KĿ}�fӑRB���B�v�T�j��I�m�t�.�*5������WnU�ȥ�k��q����=�o�K8��[����oq��߷���r%�bX���f�q,KĿ}�fӑ,K���=*n%�bX�{��ES�&�U6ܷ7����$)��٤�Kı/�wٴ�Kı>��J��bX�'>�z�9�uSQ.�d߽r�3n�4��oq���X�����r%�bX�v�Mı���j'��߮ӑ,KĽ��f�q,K�粞��335r�Xeɬ��r%�bX���J��bX�'>�z�9ı,K���I��%��c����q�x%�K���m9ı,�У�R����*��
�RB�����6��bX��u���i9ı,K���m9ı,N��Mı,x�������Nf�s��T��2��9��P�<^7#���k[�vL�l*���k�35آ�g�%�b^�߳I��%�b_��iȖ%�bw�=(~��2%�d.�����$)!Iw֜�sI�jf����&�X�%�~��ͧ"X�%�������%�bs�{�ND�,Ky9��YQ�U(A�n��MMUL�Z��A=�҉ �&���n	"~�~��i7ı,K���m9ĳ�ow��ߕ��`�7c��{��2X����ӑ,KĿ_{4��bX�%���6��bX������Sq,I!Iz=�U:Bm�6�����$)Ŀ_{4��bX�%���6��bX�'{sҦ�X�%�Ͻ�m9ı�{�;�����|�Dqr���`e�4��z�\�n6�̽�����]p���Tբ���mr�:������x5c�f��d�#s�I餓6��Wh�96Ŏݒ�%���td��9�b��N���&-�m�hb�T&6"���qj�|�%��n7�O9紼�M����N'=�����=�m�팍���]�wObَ{3�m��/�o�ܛuas��9�6;ٳ�F�P�fϊX�g����'])�����s�;2u�
7��X�%�}�߳iȖ%�bw�=*n%�bX��=��Kı/���*�RB����+0m��*����v��bX�'{sҦ�X�%�ϳ޻ND�,K�}��n%�bX����/�[0��$.�+t�t�l�lC��7ı,O���]�"X�%�~��i7���������r%�bX���Ҧ�X�%���}�,���L�-�Yv��bY�_�(dL����&�X�%�}��ٴ�Kı;۞�7ı,N}���r%�bX��e�32��f蚺��n%�bX����r%�bX���J��bX�'>�z�9Ĥ)!O'1�+!I
HRB�,���6RK�d�#\�E���sևc���7U���J�zK���>�ﺸ�ص�(�{�s�bX�'��?�Mı,K�g�v��bX�%��٤�Kı/>�iȗ{��7������d��uSc��{��%�ϳ��NCȤEO�r&D�/��f�q,KĿw߳iȖ%�d.�^
�RB���ޗ�N��t����]�"X�%�~��i7ı,Kϻ��r%��D�Oz��Sq,K�����iȖ%�b}�񆵘k5��Ln[u
�RB�lB�	�7��|B�,K��Ҧ�X�%�ϳ��ND�,MD�n{4��bX�'=����3,�ѭa�5s3iȖ%�bw�=*n%�bX/�׾����Kı/���i7ı,Kϻ��r%�bX�MC�&+g��U3�Z�g���<����j�+�&�ܓ#j*%���hMc��m�����X�%�ϳ��ND�,K�}��n%�bX����r%�bX���&���$)!r�9��M6�ԍS��ɴ�Kı/���&���&�X�����r%�bX���Ҧ�X�%���x\/�RB���ܴ�m�*m������n%�bX����r%�bX���J��c��:��o��K#m0@��&�~����ND�,K����I��%�b}����f��Ku��s3iȖ%�b}۞�7ı,N}��m9ı,K��I��%�b_��iȖ%�bw��asYin\.�Xf����X�%�Ͻ�M�"X�%���5�_�٤�%�bX�����ND�,K������%�bw�;.�hsb�Q@1N��+z��3�{)F�:��n�7n�IK��ۚf�-�{�2X�%�~��i7ı,Kϻ��r%�bX�v��9Q,K����ߓ�g��u����7��Nԥ7ı,Kϻ��r�D�K���T�Kı>��m9ı,K��:�d-Q���D)!s\��i�#t�2��\��r%�bX���Ҧ�X�%�ϻ�M�"X�)D�K��٤�Kı/����r%�bX��Sޚ���5��L�J��bX�'>��6��bX�%��٤�Kı/>�iȖ%��T��·q;���Sq�7��������S&��m�����%�b_�}�Mı,K���6��bX�'ݹ�Sq,K���ߦӑ�7���q��Ea���Z�U��J�t�|Ɏ1{��M
ic��7�l��X�Z�ѫ���f�q,Kļ��ͧ"X�%��nzT�Kı9�w���Ϣj%�b^�~�&�X�%��O��\3Ys,����fӑ,K���=*n%�bX�����r%�bX���f�q,Kļ��ͧ"~U�MD�=�����Iras5�f�T�Kı>��m9ı,K��I��%�b^}�fӑ,K���=*n%�bX��<�U:B���U2�|B��Q
�&�}�4��bX�%����ND�,K������%��,�O��~�ND�,�Y���9���JQ��Ou��ļ��ͧ"X�%��nzT�Kı9�w�iȖ%�b_�}�Mı,K�7�(B�WAZ��))��� ��p�!��h
���g]&���`�*��(�2�Ie&M�/�v����"�cAAh�:�H�@�@0 M)��	 V�A�Go� 8-�m�f��L�TQ�ڬ��,3l�=l�����g����++�ٹu�BU�,�ϑ�`�T:��nr��]�'���<�檪��rr�B�Fԝ��ۓv�v�W[���e�״��C��=�67 a��D��T�O=\e벾����u��Tv�h�b��;n�!�93r�HkJ�(�	����YwXw-s�2q�/E ��v�^��T!J��3�Q��t���Q�m�8�X�h�i�r�kfV�g�'Ғ̺Ȼ��m����c��xƭ`�JV��QX�\Q2�N� tkf����+v-T�s���T<��l�<I��[�n��l.�6�g�����j�w.{p��7o$�7�P��,Dݶ:��[c�/���I���̒ʲ�Rj�l��iZ��vk�c[�T�a�u���NG0YFR������3:V�0B
�@�.�U��MD��/.4�-y,4�l5r�&�����$�٬L��3��Hv�é����"f���NJ���X�W��mt�.�P'�����bƑ䝗�J�����cU�A��G�Sӽa�g��z��w�����s�6�9;.-�m]�1�� ;��X*nQ�H��]��R�S����6��vy���u�� ����ZλIme j�U�
f��Wv�n�N�U�JGQ�lI*��6�Uڨt�1>#��]ʪ�v����x.j�`G�۲��g�[�����,�C�UJ���v���UYF�P�����mc�mXW�r�U�W`p�m�r��9j���S�Q�9���V������"��������T�8N*Y%n��zK� L��^�p�U]Q�UC;�z�,�a���Ⱦ-���ݨ2�6�t�l�mrĽ}�^<�[K��wkZ�Q�t�&�
������Tl�z�6X$!�ᛋ[��<��yc�T�#��J����]"۷Oo=�!���������fe�ɩ�� ��6+C�>�q�U@�DC��@0.����À�_�4�uUQ�9��-���Lԓ2��$��;���!�3�n�S��nAɛk��T�� �&�݋Xf
^�U��gJ&l�W:�V����5ѹ�6��l��[&�M^����!,��M�7Tmr��m	Ƅ��l�e��ݻ,91�*��:۪�������W��-��B�y*R��[r�۳[ڣ<�4;kq#b����tRw5cn@:9�׋�tgu�[(o�w��w�;��ߟ���c�ښ���\gP�#Q���8�R7�b9Kvu�����	W�,ׅ�sW3>Nı,Kݹ�Sq,K����]�"X�%�~��h?,�MD�����w����$,
7J��M7�Z�35���X�%�ϳ��ND�,K�{��n%�bX��{ٴ�Kı>��J���uSQ,O������a���fm�˴�Kı/o�f�q,Kļ��ͧ"X�%��nzT�Kı>�;��Kı;�o%�ff���hj��s
�RB��J�U��%�bw�?J��bX�'�g}v��bX�5]��eMı,K�����f��%���u���Kı>��J��bX�'�g�v��bX�%���T�Kı/�{ٴ�Kı=��ܽ���fU�롷"v/a�4��щ�.�1L���l��$:��΢ε\3�%ND�,K����iȖ%�b_��eMı,K��{6��&�X�'}sI�d)!I
HY��ES�)�4�c*�m9ı,K�u쩸|�t������ ج�Ȗ%�߻�ND�,K�\�*n%�bX�}��m9�����ժ��sBt��M�+!LKĽ��ٴ�Kı>��J��bX�'�{~�ND�,K��{*n%�bX��Sޓ̳T��r�ֳ6��bX�'ݹ�Sq,K���o�iȖ%�b_��eMı,K����ND����У0�t�l���L+!X�%���ߦӑ,KĿw^ʛ�bX�%��{6��bX�'ݹ�Sq�7�����������S�FJ�`��]a7F(�ӥ=]��u��MnƧ`�$c_�|/��өn�t2j��]!I
HRB���V%�bX��{ٴ�Kı>��J�3�5ı;�o��r%�bX�����y���,�������oq����6��bX�'ݹ�Sq,K�����iȖ%�b_��eMı,K���\5�V]f��Y�ND�,K������%�b}�w��Ka�c	��CD�Kߵ쩸�%�b^��ͧ"X�%��{y���r��a��J��bY�E�����m9ı,K�k�T�Kı/>��iȖ%��E&�w��Mı,Kޙ��5�����̙5��ND�,K��{*n%�bX��{ٴ�Kı>��J��bX�'�w~�ND�,K���֍�39�0�7bU�WK�E��m��ФGV�x��c2(�y��piQ���{��X�%���m9ı,O�sҦ�X�%���ߦ���&�X�%��*n*HRB�5���rT���˩���X�%��nzT�Kı>�;��Kı/׾�&�X�%�y���NHRB���f#N�m�M�tɅq,K����ӑ,KĿ^�4��c�!���~��ٴ�Kı;럡������ow�����n�Rΰ1��Kı/׾�&�X�%�y���ND�,K������%�#b}�w�iȖ%�b}�o-�3Y�e�0�kW34��bX�%���m9ı,O�sҦ�X�%����]�"X�%�~��i7ı,N����7ښ�.e�����b2�Tz�V�ʼ�Od�I-�khv���U����:A�����7���{��۞�7ı,O����9ı,K��I��%�b^}�fӑ,K���N��L��.��L�VB�����g}v���Q�&�X��߳I��%�b^����r%�bX�v�M��%S
�RB��*�!M9�m����}ı,K��٤�Kı/�{ٴ�K�D�N���Sq,K��s��p�!I
HRB�b�Um9�6��m�n%�g� j&��߳iȖ%�bw�?J��bX�'�g�v��bX��Uvs]B����$.k��6䩢���5�ͧ"X�%��nzT�Kı>�=��Kı/׾�&�X�%�y���ND�,KlU�b����ݎy�[c�=��ݶ��)��`�W�Sι�˸�٠�V[c���'�2�E��F�-�]*FKu�2	�2s������G���t]=�{V�ҥ ��ܮ�v2��&)��M��v�І�W	��$�X���:��(��눉9\cŶ�%��I��q�Ck��e[���i"�gI(f4/M�G;�q@<�GĘ�=�ux&\����w�{��r8�-�#T����Ռ�WU�1��[�mnk�0�$MnA�,&���6�FK���u�bX��g��ӑ,KĿ^�4��bX�%���l?��MD�,N���aY
HRB�+gu��N��T�ɚsiȖ%�b_�}�Mı,K��{6��bX�'ݹ�Sq,K�����ߛ�oq���?�~h�I3Z��*Sq,Kļ��ͧ"X�%��nzT�Kʌ5Q;����Kı'������$)!s�^��4����fӑ,K���=*n%�bX�}���r%�bX���f�q,K�s���|B�������t�
dl˚�Y��7ı,O����9ı,?�:����r%�bX�����ND�,K������%�b~A?{�?u�4u��;�qzZG.�'\m��L{197cG�m��/IT�,��������bX�%����n%�bX��{ٴ�Kı>��Jȳ�5ı;���p�!I
HRB�j�Um9���K%�I��%�b^}�fӐ��Y��$dL�bw�?J��bX�'{��v��bX�%��٤�Kı9짽&�f����\��fӑ,K����*n%�bX�}���r%��5Q/o�f�q,KĿw���r%�bX���~��M���q������ow���ӑ,KĿ^�4��bX�%��{6��bX�'ݾ�Sq,K���>�v�̵�|�~oq����}{��n%�bX~F:�~ͧ�,K���7ı,O��z�9ı������CF�5\u�e�e��]m�Վ�}�ΓNr:K�u�:D"�5.-�[��Mı,K����ND�,K��l���%�b}�{�iȖ%�b_�}�Mı,K��l�p�ԷF���K�ͧ"X�%��o�T�?���"X��]�"X�%�}f�q,KĿ}�fӑ,K�ｼ�5��[5�.kfaSq,K�����ӑ,KĿ^�4��c �C�$? �&�ı/��ٴ�Kı;��eMı,K��߰��RR��˙v��bY�Q;?~�q,KĽ��ٴ�Kı;��7ı,O��z�9ı,OǍkxe�S32R]f�q,KĿ}�fӑ,K��nzT�Kı>�=��Kı>�����bX�'zv�S�j�[�d�����d�y��sWƵØݩZ:�"��:z��vJ;������TemYk�����{��7��۟�Mı,K�޻ND�,K��oI��%�b_���iȖ%�bvj���p˙35n��̕7ı,O��z�9�+�$����L�H$�~͡"�'�^�ȟ��SQ,O����Ii�J[�t2f��/�RB���n�B�,KĿ}�fӑ,K��nzT�Kı>�=��Kı;�o-�f�e�e�	.f�q,K?*�������m9ı,O߮J��bX�'�g�v��bX"uZ٥@�7Y}��n%�bX����K�kR�d����Y�ND�,K���Sq,K�����ӑ,KĿ_{4��bX�%��{6��bX�'�=�z�S2k9�����������8�gk�We:4"����S�[��d�L�73c�����X�'{��]�"X�%�~��i7ı,K���l?O�j%�b{�?J��d)!I���U4�
�����_�KĿ_{4��bX�%��{6��d)!I������+2l�b�Um9�Jq8'%�fwK3gc�V�wK�j��T�	��1�,͜X�fM�}��a�3�����F��2&��'1�+ �;��fwK3g��P#D4�� �)E**j�e25r�+J	�K=kzh��ԑ-N��#�/I��"bGg�
Ri�����d�V�����&֔y^r��t�d���q���B�c�ͮ-�Vc�s���H��v��v�:�c��NְK��ֶ&�@;v��6듭Ͷ��+c#��Bp�l�y�λg[��g�lg����B�l���t�ܽ��uF�c;������{����1B�N���s�״�yz+�y��;����p�]u �u�p���S�n^(gX����s1��^���G(3+ޛs��JT�&ۑ��NK ��f�Ձ����}����:p)R16J�F*n���xX�fM����(�;��`���`gl�Q��$�ܧ)G1�+ ��h5�@f���Ż����$�)̷6�;����	Ws�|����3�>��9C*D�c�'T�h�ɻٳ֭�W,�y�X�����1��O��-TL����>��`}�8�3��zXsU���MȔ���>����tMg �U �� ���:�PE~M8�gg2��`���>�c�BID���[�R����?	���}�`f��ԑ��K7���k�М��H�dqX{���}U�߭ s����l@n�9@v�bR��NF*i9,��f�,Ǽ����w[N	��N9	.�N�FtK�Mۑu����9H1%��C�����ެw`�H��Dj4����Ł����}���>��`gl�Q��)#��T�X�ݮr�3y� �n��l^�!#;��M8��qGqXozX�{ٹ�IÌE�E�$?t�B#��\X`R�F%P5~��Ѡ�Fb�5"TP�P�e�B�T%%H�A�h�_ }��(JjVOf��
Hb�i���4��H�6H@!"��f�s�pe�n�8Uw� *)���� (E_�|�"4<�C�P�*t<
��D��p�@��6�yqBȊ�ؿx[������^�9�]M�Dj�pPRK ��h޶ 7i�A�w������
���)i�`}�8�3��zX��,���m���J�MG$���"k�j��ɫ�H[֞E��ېq[v54c7qZ�"�$�j~��n���zX���G���~,��ޤM5T���C&i� �n�kv����\���J��i9�����X�8��n���zX�N�J���N7N���k���� f�hD}�؏�}���Xw�J�ƩI)�I�X�ܛb<���> w=�`s�xXfM}R�qb�Q���3��1<�֫ғ��q��X�1,�^��b��r1ۆZ���o{ր3[��[�ܠ���m�US%�M�9���!$�*��~,����>�c�B�;�2n�Sa3Mґ6���Oc�V�wK ���Ӹ��Q�R�?5!a��g��7ޖ��,͜X�NRt�N2
8}�I,}��I%��>�$�\�n�o�{~���
T򦚊7�*����s��S2\��I�30�[����������<0O23m�+���
b���t�8מË��ϛ��!�{:�Լ��v�T\!�5qͷkG3���`��F4�M����(,q���kt�qcy�ɠ�m������Гr0�s�	��ږ�"2�N����HGm���gf��57L�Ĺ�;�3�Ć�4��nz��:v2�eh����ww���f>~^����Z�UnUt�|ɎҔxl����X^��6qrZ�mdB����$�����|�[�p�$�g_|�Ktv�K�:�J���R7"NO�I-�8V�K3���I%��;I$�;��$�w]ʍƩ&&��pV�K3���I%��;K�Smn���K��
�I}�_JMm' �R/�I%��;I$�;��$��+I%�;��$�SWSrQ����I%�wO�I/UwK�I%�;��Ic��Is���
7Ni�O�#s�r�j6ۧ�a��4I��$N+��Ո5l��1�m5������| 3&���X����K��|�X�wk5��5�r�%ݶ߾����J��������\��v�Iow��$��+I��>�{��	u������� ����2���USu~%L��u�Nd��sP�u�N9����+����ߟ�~��ZI,ɼ��$�t�$��u�
Tlmʑ�����s�i$�&���YӢ��K��|�\��rn�J�8�v�tVܻ�x
�Y{J��1In1]a�`�Z������d�p�g��� ��������i$�ٽ?��K��
�Io��J�n\�`��� �}����ww��Q,�z}�Iw9�ZI,ɼ�������^e?x��1��v�If���Ku�����{���^r�ou�f�jK:$wrn��9>�%����>�~��ݝ���$��Gi$���>�$���"$q�J��pV�K2o/�I/�߁�s���-�߻��s����=.��'��Ϯz������轉,k�:Q�=Y�s���Z��jwb�J[L���N��"�I%�ގ�I/��}�In�´�Y�y}�In�ؔ�&��D��đ�s����"dn���OҀݦ��;p)Q�I��'%���������Ԗ����f����w�Tn5I17(t���R^��U�{�3+ޛ �����Q�" ��c���TH�j޵�Vw�$��7*D�Vc�V菾��z�����\���U�/��p��7bU�[u�����n����5�˭��98qDW���w�u|�k����m��Zv���s��7(u26�	�G�3r�3�3r���XW5�DHゔ'?F�9��M��Vd���yDEQ�����[�>ֻ�	�n���A'��>�`gt�3�3�7{�JT�(�7Q��U�5�@{������;��P�=7$�TP�+�������%֬75��b�lM ����Ds��(@����V��KN�!�s����������N�)��,O�|w|��Ի�q���g����-��U���V5����9�Vd���B�g�ckn��d��ݜoK���3Pvk#\�v��ܵYŰO$rDN��^��*[�v(��� a9�r땎�v����7V�3Ha�
1.�&�"j'�0n\Ӧ8�cY��x*=g�7E�ܰq�p��Sk�I��]��$�4�Gr	��f?+1�+��ŀ}����w�R�%I17(t����{�~�Q�Q���`�y��w&��:<t���r�I�`}�8���X�yX�yXX>�nJ?F��qXkv�ݮr�ݮr���ӽ~��;�#���#�rX�yX�yXc�V�wKv��H:I�!S-�Y�fu�t8s�r6��2�k��4�v����!#���$���{���:a`s1�(��{Y�`rrwZ&��R�ӑ�4�����^T�j a��������}�����X��m��4�,��v9]ɳ�DL���6;�K��cN����L�vQ���6l��+�{��3;����r�q*I���X��Xc�V��,ǿO�o�߷���:㖴�滊'�8�U��:�v�8\�b9-���chv^����{��|�p��'I9Q�����+ ��c�Y_ �ܠX>����8�A8�3]��[Ҁz��nW���d�T��97�ڒX���ΜY?~�_�%%�B�%
*��2l��v�R�#�8F	��ȬΜXc�V��,=
!z�Y�������&��RS�EUb6��菧�޼����Ḿ��0��H���H�&��v^
Nw&��^�X�}���K	:tv�m]"	k�a�$����3;�����������>�`}�N*HJ���9,Ǽ���(S'{[�`s��6�f;�P���Ͷ�8�	��IȬ��+�}��3;��������:SN!���qXy$�y׻6�������y(pB
�^��3����I��5��ֳDnjؔ��3;�����������>�`}�����p����R5G��n+��W�ܖf���::�|�χh3l����U���v��u�����}�m��;��^��n�1ҙ�Ḿ�c��M� �n���P.[�����ME ��,��+ ��z�W�����+w�Ł��bR��9IJi8�u�@n�9@n�b6��p�L��J�r��3�3r�>�޻�O���rO�#�	!AC����n�f��Wb��+~�΋F��M:r�#�4ک�#��0�B<�B	E����Ga�L�j��"Մ�Dv1��E� 4b0�~a�s����6����ə�ֵ��ml,X�u�{iC��sm8I-��]��x��=(jĮ���U�u[c'	U���(�n�:Dםm��d�vj����ѽ�p檩b��(dݳ���y�m����(��_�o����v�;[� g�lQ,�E�V-��}���Δy�.��8�ض�;Y+�nz��|~z��*�h�i�$��vFc�b��+ڧ��F��Bk<g�������,l���g6����h�ZD�5�F�.�#�� d�؉c�΁� ��6�H�\᭻h<Q�u��h7!�2M��LlV���q0
�B�hFE�@ƫR��P��X=Pqn�HD�YF�.y+8�:�Ͳ�&r;��0����m�:�g�`��!��\�ћ�oJ7�c����Ru�=*ʵ]�nv�t�����R"����<1�lGv��qU�s�D5,�����Y^�������A���kMv�<�r�����ձk�ll�k��5�1Ѳ���n�;U������]�V�G�
�3����= ��a��ӻp�G�C�q��=D�.6�\�on���c��dŻt��1�h�;H<�!$���6�+���s���Ѿ"��������cs:by[����4�2����Ο@TS��g8 �.z @��ـs�ݘ+F�����Z���ս���ڥ�� ��U�j���U�U۪���E�(v�Hn��!�Ju&ݰ�t�WZP�s�uHA�t2g5����XA	��J����ae���R�7m&Y�i2��e�6L� x��vW;��C��1.�9k���uD��(Uڸ;jD	UWj�&\�f�f|^�w]nwי�2x���mns .�x�&��L[\V��AX�<[l0��m��"��U~|>7l���mq]7�����[H�xŴ�$�7/$B��ɳ՝�EWl�N�3��:A�N���f�öֶu��)����ΊyW�`��ۭ����tX]���E�����K�?{Sd@v*�?B:��ҁ�3Jy�G���v|(4�G���5u&��jj�X+��-g��B�np��=�si�鞭���ڝ��Ж�v�,u��s(vd6���쫹�{�i���$��������-�Zyxd�3�J�dz��c������DRa�L�iյ�%�v�)��4������$'�s�ل���V6E���^@���t��q��p�b��pm��T��Y��Cgn�ks�Żs`�=A{S�{���{���~~~%�l��\3!�ɪ���n����tk
���<�-��_�w����|���P�RD:NE�{�x�>�ܬ3�X�yXn��4��QD�NJ6����ﾉ�����OҀݦ�~�I(S&���M�%�˙dӛ �w]������_���~�3_�����	2T�Ɯ�c�Vc�V��&�Д%�{��`sjV�Է.�:��~�E`f>�`Uf�y|��K1�/�oϯ��-Mgg����7={V痢�w��n��ێD}�F:��1)��U��<fը���m7(u�@n�9@n�r��s,�i���i��f��9��#TBO���W?� C�~�r�I����l�]ɿ(�9���Zt�M:l�����~��7(��(u�@osW�̢UKu#SM͇���$��{�`s���3�X,��VwҚr�M5LI�`}�yXf��>Ǽ���/�o����k��ڜ��6+�g�uҩ�/�gWh.s�g�u���u[-v�$��Ks`�q�r��`}�̟%�|�5�����=�n@R��4�3k���L�޿�~�����a���M�%&���V�Ӌ�{�ͪR*����D",6��������`f=�`|�wD')JC��T�2�c�
BUܽ��f��r��`ft����D��J%	H�5�@~��︷��;�~��P���Z�X�B6�1Y�C���g�Jv���x��h�rt��w���w�Ϧw�\#��SI9>5����Ӌ�{��3;��f�IJ8�c�%)C�X�8�����#5���n�����>�'Ji�M68�7�{��3;�������f��7}<XX>�nJ?F���Xz"&{��`s��69�J%F������BQ��DEc���>�L��T�T�ӧN���>�w&��P�׻?��l�gt��M�����MG$�"h�v��<��x��wS��!ۚ�וӶ᥇u^)��JM��Ȭ�ܬ��+ ��������]҄�6�u�4�>Ǽ�ВS!����ٰ9�̛�$�d�ݱ)RJ)ԩBR+ �����=�g�%3�����f́�Lk���8����ms��7(��(u�@��R�$�%INP�Vc�V��I.u�����>�w&�ꈨI8�Iz!-͙��ә�4�	i�A�$æ��� �v��C2���s�[7a��<ٍ����[�]X�]A����:�F3��C���1��S�a�t�V�b��]�M�2�l��1��W8�۳uٽsa�V	���f#�8��e���p�r��-i�c3;a�i�n��l��٫���'
��:d,ȭ�ې��u�[���,3R�5&��&���!�$�|���%�E.J�3����Ф	I��ĸ�^Ӭ]xn݆�@��\�@7?������7[�ms��7(V`U6�uD��Ks`�c�҈��9��+u������UUI��rQM�Q�rX����ܬ��+ ��sU�(R6�	��Ȭ�ܬ�]ɰs1�z"Sμٰ7�2�Z��j')�8���+ �����������>�d�#Dn7!%$X�M���y҆Җ�!K#X��ѭ�k�[�l�m��R��V��,��+1�+�{���N�ԥISI9,�]ɻ�脕(�P�L�����Vzl3�Xn����&INP�Vms�ms�~��{޴�?J;�w���dR8�qXW��K6w��f�����3�:�}�ܔ~��%.Pkv�����N�OҀ�� ���]����]�j�\gP���m��$�lK�TgI�Ru�NҦu[	�:r8����ms��s�o5��}F���|�3�+�je��d�M8t���f́��B �n���Pjf�&��J�TT�6��Z���숴����D �D���ȩ��`t��k^�w$����'{�d�M��JSM�VJ"g��v:����{���7��ӥu)RH�"�T���6��v��7���ݭ�����}��$ʶ�tW����5�e��^!biK	��Cph���5�j&ʸ*�p�~�o55�@f�r�>�'Ji�M7�D����7��5�@f�9@n�9@8қ
��>��D�$��o;�{��~�I{_yX��V�S&aSM�7#c��:��(Jyכ6��f����V�$D(I_Д�;*�q(K��sj���+q�[��KDݑuw(��P�� �:@f�9�6"#�e�V�Lt�f�Kcr3R27:x�db�.��W\s�	Rt��z�I+��X���ﵼ��q�8���X����Y����+��+w�ĥH䂥*RD��;ΐ��Pk��3y�_�d�z�ԥI"�$�Fێ��}�`v=�g�RY���{��3w��ISqF��K���(�jw� 3k��3Y:SNRq(�m8��z�����ͮr�{\� �?�>����S��	��t[L&�kt�7�6a����ͱv ��L&��l�P�6�,��[���k��h�$�G���6���p��]���6�7��\�+q�q{5�e	a	nzb �g�,`�n0����e^�e;%$���;N<q7nv���|��F�z�v�<��tK��B�y�떕
����a%8;[�	��<7B^uh;���r�ܳ��ֵ��B*����}�rf�ٽf�Dm�:��۶E���8�U�qAA���p�I)�nJ?F�������v���������o]XsH�rQR"B身�ms���艓�OҀ�~P�s������U�G�M�R�!QȬk����B�s�ms�ms�&��iʃ��7��X]�v������oK3vɖ�m������VOs��޷��=޿�j5��T(�#\��L��p��fv������t����p�"�֫b� n�g�m�[��n�Xfʀj��`gt����k.j�	��rO}�l���B��F&>����#�Gn���H��+�}&o��M9HmĜ�)%X����ms��� iM�U�]Q73e���s�ms���(�jsH�rQRR����`}�yX����w��f���Y���7����*K���kMz�I�9�gi�c�7jܦ�T�&�z�����rV�������>`�7��Y����+q�[҄�hq�*8��z�������;+�7�"&L��&Zm��R�S#mX=��nIϵ�]϶$�)B1��AH� � E@�M��,�D��"��E���y]� �D��8I�,��2f�;���j9��]}����M�H1HSNF�"���T ��It�u�%ED�d# �Uv�d � 0v�%]!,5�6��� E�A���H�`�F,�A� H0� FD��E�ȑcX�:D�b�Д4;@�i�� �i��P��| ��"��M"�&�b��U���}7$�{훒|wف4�n\�i���ua��O:�f��箬�z�����3w��ISqF�໹@=�b�}o?d`�~�mo+{��*6��*Sr�S��H��8�h��q�gհ��l%�9�=ɴx^�S5�ݲ�U���� 3y�@9�t�ͮs��C��Ձ��n�Sh�J�Ա���f;�Wrls�j����W�B�D%Tw�2{�NJ*DHGrX�����޺�>�� �;����wJJF�%)R$���B7���ݠ����~��b ���a	X!`��Sg��جƕ{���Ɯ�7%Xf���y����f́�w-X��̧?���%\u.��C��Ps���t���ɸ�����v�vΑ��M�l���Z6��v��7���;���m���5S2۰>�w&�
!)��ץ��޺�����������*r)3W��{����B ��h��6�ғr�8�$i7�޺�s���]ɰ�	yD(���`ya^�S����#!$� �ޖ�����=�>�rՁIB��	>weT��EJl�Z69݄#�;Mgv��g�8���\j۷�h9Z���<e[n�B��PE�����e1&Mj���`6��N���n���izY�7N�E@�e��:��r⣦)��7[ccŠ���N��:��z ��WH�GTW-gG*yw�����t�D�J���.͝��u���ڪf�؍��ǍF��R>m[<���\)&"��U?������NwVk��V�nk&�D�]�o;=�
���#�,,Y#'4�V��J!!��%%)	#RM�k����+�޺��zX�Wq)I$��GWwr�ͮr�DDɼ�� o?Z6����]�)9iʃN+�޺�����艝�~�u?J��L�]�q�!)"8X��,��+1�+D$�������kT�m�U.����n�ͮr�ݮr���b �n�sv��s����-$5��ոCnz�ȼ��Wh�.���$�*Up��qQ���(޶ ���\���n��4T�i�34����x^v(��C��ګ�]��P�$�}�nI�?yX�yXX>�nJ*���p����\��\����K�|4�DF����������ٽu`gt�>֫x����$�ENI(��(D}�~���z�k��?{��?o���S��j��cs׳s��ܛ�N5����j}��A(r:��T��q��L��YSW8��B �n�k��7k��7{�JT���(n�ԕ`gt�;+�69]ɰ3��W舙:�Z�4�t�K�j�f��7��69]ɰ�	�^�,J)D(�J"�)��� �n; �;��n$�QĤ�H�Ǽ��g�wK�{����:Rn '�4�����b�}��{׀oS��7k��6_�}�w@��-ѵHnxٝrnG9�i�u�â֗ui��0�%�M��۱����ݠ3k��7k��3z؀���ܔ8�BHӒ���3�>͜X��/�I��%)"c#�����@wS��3z؀3[�ms�c�R���Ɯ�4�>͜X>��rN}���OP0P���U�u��mWrlgvɖ�%4�uJht� ����򄗻����[�3��V�3o���k����j��#�^�艹K�<�vV�<�V0����Tܒ܀���~��7(��z#$�z�{�%&�I�8��I�����ٽu`����{����:Rn *p��3W(�� �� ���v���I҆����rU�fwK��+��ɰ؄��s~Vgd7B��1ʐ�4�;�?�v{��=�� �f;�1�,�2̙�*�jZ�5R�\��I1��r�rٌ	�Mێ
������6'��)v\ʆLʃѳ[�۵:h�ZKs�r�8�u�\�ݭ��n�cr�]�Uj*Nh��K��{*�*��;���.�Z�����;s�ǰ���>m��§�7k`=���v0��=�!aq�l�+�v�������k��n-N��-��豴-�CnhŻlZw��Dcs�\C��#� z. �JNs�jj����3T����ٴ���H[�� 1�lnQ�����#����qP�����o�����s�j�9����}!��ٰ7�I��'#C���R+��ŀfwK��Ł������bR�H��7I5%X9���^l%	D)���f���ڰ>��]M�'J5$��rX�8�3r�;7��3�Xݽ%&�I�J\v 7i�@#�����ր{�Ŷ��a7�K�C1��=��^J�ZhR���|�\�qlj���쳪�5���m7w37s�{�� �� �����2C���`{�'��D9�J���wEx EJ��+�l:�\c��=Y~u�J�5� �V�JBHӒ���Ł����K�޺��zXkU�JRD�tԃ��,�nPy�@���[h���9"�"�X��V��,͜X��X��iGN m��$���(��Z���2w:H��F�G���[u��r�H&HJI�*�3;��ٳ�1�+�z������%7QG%4���{���7(�� �� c�wN$��Ƥ��X��X��V:���I�G������(4m���f�?���X��Ji�a$Q$�;7�X9���^����{�`n=t7�NF���3�X�8�3d���TF�-�.�mȩ��M��ӌ����4d.�7T̅Fv�nֹ]��������r����&�ޟŁ����ٽu`����Z��R�&���T�`s��7�P�DBJɽ͵`���;6q`v1��u$��[�9ܵ`�c�aD%3�ǥ������b�l�-LԶ�6G�*��y��~,r�&�z�B�"#������DG�Dl%P�U��`gO?!�t����&�����Ł����ٽu`������"N&��7�#��e�<oYn
��U+�=d�`�� ���4���Se��Vd��� �3�B�^���k�`nl�4K��r6���9��P�7[�޶ 7i�_���<�OJ��S�#q�V�ޖf�,��+�z����;�n:*TRF��DD)���`w��6s�j��g�ݖsU�%)"i�jA�rc�V�DF�7��ݦ~��`~DDB�������������ʨ��UEE�U��TW��TTW��E?�H
E `�E b ��,Q@��E `�P(��1E `0E `AAH ��U�� U��TW�*+UQQ^*���� 
��� *����
�����
��� *����*+�TTW���e5�� 8�� �s2}p{�            �    
 @  ơA@T 	P��J�B
�B   ��*�( HT      �� � H(@D&   � A*P@�4��M>����f����zo=� �ngݞ���v�{�r���}nW�x Qǥ��W�ܻ��ۥ%�1�g F�+�z���y|�v�t�sd���9�d���o�Sqwm�w��<   � R�@ɥ {ʟq|��y���Mڷ3�[�>�ky��{���rj��7/}�ǹ�\ z;���X��/>��V�t�������m�K�8��}�rt� W{��M\�un�y_[��z/� ��� P��J
@ w��w�{�R�����rt,��̀ɯO�[� �     �w��|s� �-Q����z �>��-�ی�nm^�{�>�wϛnf��Y�n�M*�4���� P ,��A������쫟n����us�;��� O>�w>���y�U2����<� 9�LJD 6   E�� � �N���  i���J'@��� w0 ���( lP  

 
� �` 1(@ 	 "  ��  P+@ �b�޳� c���Y��y� ;u�k���6�� ��MqgC����s�{�CO����y�y�z��jvr�f� 4�6ҥ* �S�CSeR�4� <z�RMB�  Ob�Q���L�O�BT��*T�� �"$�JR$@�jz	�����g��c������{��|��EEz?�EEpO�EE�
������(*�����ЂD� R2 P���JdJvS:$�2(��QdI�20���"L$0��`P�M�+��\% e*0�3"nT����F����4�4�jd�7�4d��a�K���7y��Q���S�?K�Ӌbˑa����?x~�"el$��i��$\v��������d$c8x����J�fL��I�я��$Ho�l�6�(L���I�I�f$�c9�䐙��*y�L���\<$�"X$u�k)���셗-��MHH��42\��7]ٰ�e�Mvѥ���L
^B�<�<
f�L1i�S	Np�	�n�@�9�Js	I�
��>��<l�d82���M����J�=����=�� !�MOõcD�z~G��a��cE�;'<f���fs���5���{!��s�}�y�%�S��O?$(���n����C=@���E��EZ�J�kB�)ɭ�d����,�ݑhd�8)��lx1�4x���
A��<4�`1�&�$IO_�@��'�?7&��1-�rBr�HHGB,Z_�#���,
��H,F��b�L��D�XF2Ж�F�r%�$�`\���������|��$3y&���5<�Á	#�$����k͓��m]g�I
��&Bف��mw&r��<4��JrFHW���6��t�1�6)7��C^B'�e��D��k蟒RS4�������ŅSՉ\�"LBq�� �P��Oj�|c#���VD��^�&�Ѕ08�hA!�����
a�@�XC5���p��B{|x�=5=��$�R&�O=�dH�o��@�� ���#�b�1X� 
f�\�"b�k.s��y�9燆y���k��dhF>�$�h:�*�1"�bňDl��
�k�*�K4��G$���e��$?r�Q���e1H��LH��X�AHP�$
�$���0���*��8�#)���$:!��@EB�#�F�X�"ŠF��B�h@hb�j�A�A(1�.����� �&�$�k�ً ��ō0ӛ�Hi�BH�hxB�H<<!G5�B䜜�L��eЋu������ѕ�И�2V�!f����a���(B�B���,vbB�ad2D&L)��Hp��$фͨ�3[�� H���p7�jbhq�t�B���H;�H�SN@����,<`A�Ƹ�MR BQ��@�C  S)@`� �����!�zAl����C��fo<��!����XԈ�?~9.�t8 ���״p�6F(\r�H��OX�򑠱#� � Ah����B�@�T���\�ȖЍ	H�6B�bD�0&2!]F0%�SYr]ЍH��c�"B�H��g�:G�<a����2���B����g�!�����%f
��FF��!b��\�o4��ah��bJְ ��Zp����_��VR���i,�w���N[��RQo'�3h@��dj�'��(��cLj���5�C�I�wІ�����2��0�n�9�䵥H�5�t��>f�||wrܗ���B0`D��P� a�$cR0�NQ#FƔ!J�Ƙ���y��rH`�1e°+
<1�X���i�@�\�q���.'����)����
� E�����bS�K�@�@�(B��d.���0X%�&hшB5X�������
Y�x�4�1%2D���4-�j�\@�rÆ���1���m		�k`R4:@�
�

~�	�Hq��	��>y�p��r�p�H�Ӈ4�d��B5%�� �B4ᆜ��T��$Y��.��(I H&�!GȔ��i��P�"��B���Fa�XE$	@�
BD��2�^&Q�F(&*=1Wa����R�!`p'��8k�@������)���d0�&�)-w������U��,�[KbH!%daYI�^,�+���Z0Hi�d��ܟ�?l�4mġ|֛���~�0B#K��I.a�$H��H��#IM�X���_$�1�Bia`�B
Q�S0�RBYT��A��㧌h8:D��.<aVSSș�Q�L$W�d�"1�`9�xP��I�I���\e��]r��Ƽ|��3dO%'��7�L\�_Fs5�� S4��-���3��e��M����zK�����;T��瑅�� ��O�����6�64��B�����O/�1�x��L���A�	�h�-�M`daY�H�H�&X[��jc���Zb�쌄J-��V\��+����B���@�5Ē50 @�Ywv�
��I%1 �����%g	&o.q�:����
f��5�2�4<cu���ġL4cLC`Q�-\	d�%�W@���łT#R5 �#@�C]aL ��7X����7���;����s���XnY){
~)�m�p�4!L|�~�&�6y��.��ny�6y��B>�{!�N����"H��$L˄1ӝ$B3�FH�L� �
᰼�	$%vM�M��t8BJn˞�����H�p��$�ÍQ�p�,��2�Z�"@��L�kLs���.i��$/�4�(rG���IH@$��Dbb��$��ږ���&`y�M�rA�vM9��a��7���׍�a"X��r����ON��$�*�������k�}z.){�
j�i�i�8�r�:�箾��t�\`�4���X%H�F5�I%L��rIqі�d�̙mb�����o���y�V<�c����3x�a�S2FB�XG��d=g7��O0�W�P��������aV<R�N�/!�X��<����?��Jă�&x��Y����22�2�	+9!,+��c�ǰ���^r��p#
�! �á���1��LwL(D���	�M���/���&}����>�r�����I�'�xP�����&�w�o��xbB���7
F��Yr�K�(d)P˙and�i���Iy��9̼%ˤ��e�BA����E�*�S�)���c�x���
s�d��"K�����!WW��K<f���P�	H�VXa,0 �����y�Yc	FY���6�%³���G��ar���4��%��P��@ 4HҸF���W �"Q�p�B"@�!\��Bo<&x���E�SO��9w�2Ja��$�`�@�+37M���,H���@���,'�8@
�a
���]�N@�0#K��I!C�XE ��n��1t�*Xf��I89�e�BP��zp���H�^ D���R;��~�T -)�a�F��66aaxB��	6y��y���I)@�D�!��Ӟ�F�<�9
p�H�e�ד��NC9���aOd%���:C�^���4�n=�O<$WA �?E��@�&�{bI��=:�F0<)H�1!-I4�wN�� �         -� I��Y�tE�ʩr�"���eV�b�]����M�  �*����_���U[!;q�����9�ͮi`51��)V�'`�꧕�����$�-Tk��.�]6�H  �iŴ ��^^����ҭ���m5�
��l�p��"2Uj��dw((�
��0e��ʍ�TqsS\�n�t����h�5��fG@�F�[/*6:�V����7ɨW�m(
�y��d��v㕪�8nU��+)��+�LKu)���q�1�����X֥�k�ev�嗖���U��'e's�(�mq��m�Ru�5�����m��RW��e�j�W�� � r��&պ�jԍ� ���,6�-����HN�[��0m�v݉��l���-|p IKi�ć	 ��j0���-VQ�j�ݥf�m[�l6�  6�`���M�f�$�,�ۭ���e��@ m��m��8��d���  i �$�[)���"� �+v�iz\k�KM�C�l�g���m� 	�E���\	 �a�� 6�5Phڶ ӆ��n&� �t���t�lzl�jp  �l  �i		�ɶknN�VԜ�`"�u�q���
���5J�����+�K��[���u�Ė� H�j	�++U�LkҒ�\ͶY���[D�    -��  ���  ��  ����n�� �6�( �6��t�[%` ���C���EZ� �E���l �����W�i�=��pմ��PO�c�#[l����zv-�e�r�K��WV���� ����m�  րڰ��85���l[xӋd��J
��n�¬��[Z�w�u�۶�|�[�� /�H�bmp�v����[kI�-�^�� 7m���u�c���6ͻu�kRv&r��u���V���v�۲,�P�ЭmUWʥ���e]��@m���F�-����l�X[��K�  	)C�KZ��յ�v��	 H	6����[�ү-����L�/#�m�TU����XK�U�*���tU�UW.���D�.�1)-�]K�� *��1<ݺ� �'[Y0��&� k[m�$�� ӃUTm[�����&�F�XHl�ڪ��n35*�-�� J��nV���{h&]�	�V�h�6K.����U��򪪮�e��m�8�/JM�e�%p2H�IĀF��9��&�+{L�
�j��aʪ��+�Y�:Fy���Wf�Uc��ݧg0�-�� +j���;^�;��u����U�U��uv��Tj55�)-+����r�S�&Ba� �IΨ9W֩��� �]�u�Rβ �Rm̋�tA��q�i1 �KҀ�۳l�ݯJ:�($��hm[-��sk̀8�*�Q�H�pj7E*pm���6�"ؒ�A!��-U*�UU,pdZ�
����Tv�¸؛�� �i0$�� �I�m�Y{f�uȳ�/V��hp �/N׳[v�Y.Cb����: �t!+G�s�HOclx؝�v�B�a�u3��r�V����2��
Z�a	�@ �@8 �t��i�N@p���H �	�_��| I��Ӭ[�	А:�[@ 6ض�  m�����-��` �i?/��m�6 ��  ��W�����  	 H�kh	  8ٶm� �`mH�@�pޠ��׭A�*�u��s�> N�l����'i1h 	[~�`��6�ٗ������$ ��   M�o`	j�RK֕�(�צ��ht���f�t�Am�@   m� 	�� #�ض���;Ͷ-�����kh Hp    K)�:v�,�8m�HI$��Ͷ6�m� �V��@٪�`jm�Wm���`ݶ��6�-�һH  �m�`H6ؑ $�� l�U�m���v#�Q�#��E�F�l9k	oI�S�-�I!�� -�a�;m��$�N����L�Uҽ/2�ڰ�6SkkS,c�v[t[��[d �&f�u��M�m�A7nU�έ����Z�{.�HL�@  8 �c��e�`( ]�R�A�G'mU��`�UT�E� �
�▩^j�0�C-tq��$�$6ͳm&Kz�m��'-Yˀ�>� -��m&4V���p  �l  p  [m� DW%l�\=���v����d+~/]z�۶� ����^8�Β���-m#&l$	�4�v�vJ]�m��jV�Ӏ&�7`m�s�͚n��ڶ��7h��	Z��5@r��	��>�`8��� ��@vź��	 	m @$H��m  m��x� X  $� �V���&�ۜ�h   �>�   ��Hm� $��� � l� J�  ��A�Uє-A�u/*���%Cb�����6'�R��C��  m�m�   $ �� ���,kY8	�  m�@�.[�ݵn��^�m� �-��V� ���n 6�e�p-�6�I�N�v��8	� �b@ [V�h C� n�H  ��)t�J��(ꨤ9��6�64n� $���e^�V��X�n,���� dul6�m8 ���  ��  $F�H�  �m��	 6�5�   � �6�[C�E 	 ����V�    ��  Hm� 8�	  ��      �>		   �	 -��  ejڪ�*��ܛ[h�VBR{*�u:)� +�q&�l�I���      m�� H� m� `�I�����k�5݃m�m ��hH����}'ͷ�j�K�&�`	�Ŝ�	 �	��N�a�m���q�z� [C�l $=m�� M�`�I7J�"�sm��Hm�m�m����g ���-�� �a%�� 	,��>[u��l��(�vl���q�WK)d5$����Wk5H  ���qm [@'B@%�o  h[@   �c�� h p�   	� #mm�l[@ h�` 6�m�t݅�H[Z�p8H��;sSl m�[vض�  �` �I� 	�ml p �Qmmm׭�d��-+`         ��6�IU�m�� l��m[`�J��$6�t $� ��damH�n����`�m� kY [F�"��'B��
��\"�E�埩�϶�U�u��d�  8ݳl zK���( ��  @ �  kn l -�ۛU\8����%��F�6� -� -� �6�ɧd���Ĕ�Xm�M����    ۶BF �e��c Y��盁�n� ����\�\�K5�n��8���p,kx�j� ���YԤ�tZU���p
�̸ö�P -�d�Hf�\��5U�)*�fF۱VtpfK�k�!��   	��e�I��[vD��֒��V�H$��m{v�0�6÷N��6�t��	-�k �m�m��h�-��ڰS[U@Tٳ�@毁����Zڃ=��>|���^@|s����9�Kչ�RZ�[[��Poc2��x᪜�������m���s%��ԑ�l�P �a��mv'[I�����)��q�slV��q�`����	±� KN�2>���E�hZ,. �a������.z���mF�d��Q��[ebM*D��-6�E���zΒm�$�T�p�U����ۣV�@$K.�[��#]����I��$�3B���k��ݶ�m�h7m٦Ś���t�e$��ݣq���&ڹV��҄�U!@�@mS��R�q�@� � p���+H���I�Khڶ� ����:�Sv��q�  �N��t��Cm���Ի�ª�V:�4�
� ו��moV�Mњ�h-�մ   ��t�6�0u�.�'\����j�m��z�����5T:�]�Z��'K������ VN��U��U�rǳ�+HI:�66�s�(UT��ᚪ�ch1A��ێ�24/UUL��.����	%T�ڧn���0@T�k@ �#Zm&H��Yf�  ��[@ ��fH�`�F�ĥ��児��:���Uv��m��஦��W���	�;u J� �:F���Xs2���,�;K�ڐ9vv[:�-ěu��͖� �o�������PO�(� ,`�B
?����~��N��D��"1
O�P^����+����apbE`Ē�C��b�T�TP���?1@�  x��Aނ'ފ��=�:�0�!���' � @��|�U���%�N�� ������}X$�H�c ��!�H��I�1�$�AH�@�B ��O�P'Qz�q1R�t=�@���OQOQ0D�P�:(=A`�Tb� <}�T5@7�1c$#,��$H�bD� B���~�1�@މ� ��z� �(&�`~ �]T y",��R�"? ��E��F�	�'P���1���^x��x��*`a��N��)��Q�'E*u��>(>��(�T� �  �:���*h~�� j�E<���-z��"�?�
���#��F
5
{���=�N�O��� 	�I�m+$t�@�y�cvڱ7$ruQ;�9�UWnUw8��ӽ�V8c�le��3��0B@p�۠���f�2�b$)V"u��:/Z賮��ɕ��V=�[]����iԍɆ{.�N7ZK�{$$���ɸ�8���8�.�Y
�u��i�pq �jL�u�ʲHD���n�ܹ9��q��6���zu�b�a���E�
X��	��5��F㋣<�)�.�T��t֤�:�Ai�x�W<�tS�n���v�l�������]���k�\Sq(6Q���ƹ��ݧ��a�>Q :�u�3���7�:��.3��C�.{nKd+�2�5�v���%̽ͺ���_7��]kl=���+s��lDӢ�����ȉ�V��k/'$�$��s���q�JZ�e��;i�sڻ��fͩ^-�v�"�M���J��5:fM˩��w�9�W��l��N��������a���D,�sqr���Y���c�Tu�US��[6��pq�k�Z�X��l�a䰕�Oj�xml�,�e@��Ӗ�[[���`<[N�ݧ(�=TglX8Wj��ܒj�L�h����A��6���`]<���:�����[Gc���o$�hMD�h��H�mOԭV���u�%Sa^��:�8�RZ����`��R��a��ԙ6Uݓ�BĎu/h88e�k�q]!p��d�go	Yu�� Es��^����Y��$�ԀW�8��$  !�Jv�&�9��ә��%[�,���m��!��r,��Cb��l�T�*� �ýW� ��-�k�'V���Nun��9�t6S�e��T�q�ǭ͔���n����\��Z��������R6�$n�����XT��k���rf݌��GFҬ�84��]�����,[�k�Y�Og(��s;gg�%u��˂8Cu�c��+�]
dʨ��7K�6�,g���^:v��+ne��Q: x����(?,���X ��D*�����4X#�;��33��mʹܶ�=j�Į59��H��<L�\ĳ���Y.C`�T�&�lqN��5�7kxN�t�e#^�\1{�����L&:����ǙL�^��\e�s���ii�m�ƞ�׋m�Ii\�
��^�����ՠNw]�kcq��KUk�'l�r��m�
�<r���;{�V���m���0�F�X�Kse�鹤� <���9+��
�A�.w9N8���=�q�P9�)�۷'gvL�a��.�fnV�|� �z�o?�諭��m�h�}�D�I�F8�շ9�	(I�QTl�u`o� ���9yqqH�E?��,�C@��נ�f���^���M �⑷2$��f�� m�@u�1�6W�}�+�?s�)2dd��iɠywW�~�S@���@;��︊�� y!:"̐�ѹf�]�I{I��)�9 q3���n�	��L 7��$���}>4\�nj�sì�s���+2iw3NI<��s�Pp�~�C�u���a�OP�L@zM�v���1L������@��^�ff%ﾟ��|�����m9���F$��gu�t���� ��u`��7�7P��P20�G�~�S@����;�nj�s�,�}�eny��H��yM�Z�(qr�N�w4>�<�b��	���N�f�Bb��)�Y���[^�wu�.����� �)qH���8�sq 6��1�"��I�>�ď���2L0����I4^��w����H��QT�J�aH}�(��{��I'w����7��X7��$������mz��h���*"��$�Vnf��$� ۚ�v�����o��{��~���4�^f���Z���'J��m�4tbH͞6��{��?5[;�Cw����&'��#�_�ۚ.��׮��[^��r�q����j&�9�.�Y�d�>ŀz{���x����$����h.����x���XTBP�w�w4^��^\\R<�O���}-��7u��6w]`J�H��DD���4@��"���߼9$?q�qH���)�N8�.�XͼX�۬�(Ms1QRq*�mڨ�P��y�v��/OQ��RvNvYq�9����;�;����W�V�Ґ�+]��9���>m��>��rQ�o�`���/�,QxH��������˺���;�O&A<��s�& qR�s�*@N�x�ȅ0N'�A�g�f.�_٠r�W�~�w4���{�[���F�Uլgu�В�w|���Հn�xrI�c���6 �$`� �) ��ٝ3p�f�n�"�lf�l<ն�����{.�J�͖Bb����z���F�V}p<b�b��wB�WVۻDػr��W>mNأl�mz���g4���G�:��mkjk��	�E�H[\�%�A�l-�qD����E�ƪ�m4U˗�'a�g�~=v��8Mm����S���k��F�o\n��%��^Ɩ���\��ݷ-�[];��K�x#v,����[z�'���ʺ��d��;Xm��e��%�"��v�����}� ����7u��""#�M:�^\\N<���1E�9���Zn*@u�����R l��ݼ��B����ݴ� :㘀�qR�J����$0J&���nL�<�W�z8� �$��UW���R �32�TX(��$���]��v���V��u�~�	D��t��$�B�������4��@d���Y�^���ڦg��j_A1O��A8
73���빠yzנ~�w4��Ɋ	8��-�{������$E�h?�O~A�D��I�^���ŀ{����DB�>��[���F�6�&h^���w4yڴ����+�D���cȜ�G ;�K@>�R��������q�M��ӒO߳���|"8��w����u`m��j�C��V�j�����_/cR;��/5pKp�vz�
�t{j��9��c&)�c2!��h�S@���@�����Z���$0�;.�U7V`�7YВ�7��pOwV�e4��oȰQD$�H�\�o$�^�����AS�O"��Q1�'��� s�Հ9��B�1A8
I��[^���h���:�V�|ñc��܍�7��� �1 �Ih\�Q�Y�ǧvi�s��#E�D�����d����i�2<�	&�w-����w�?7�Un������s2K@z䘀nl��bH� Ly�@�v����h��߳*-_bq�#����_�߱ �� �1�$� �'K��f�f�ớ����UQξ��ϟV�M� �����$�?���_���ϙY�%�G�s2K@z䘀nl���K���&���ګ�.#�t�Iq�ͤ�XN�q6�Dsl�ʯGb5�񪟘:d����1 �� �1,�+1I��Q�h�������Ď�)�r�W�z�M��b��S#�$n�n ��� :H��b����m��9���r�@��V�Ss�*BS�����$����E�W5u�y�f�v����� �w��'�~@� ��]W@9�coٿ��\w��g@�ו�����Z� p��BYu*�b�377��uϵq]9. ���맱�;\/S�;&�l�$#��݅��c+ȶ��B���nЭ�x�[J61g`E�c-.�97J�'����@d�۱&��Lq�#��Z:4Bln��[����H	���wA�y/[sF�൳u�.�]x�q���@��=�a뱗�rܹ.�nz(&��K�M�6��jL�v������^�v��G4Hv��g	�X/[b.�3���m�������S@���@����R�NE1)��E�wYM�ֽ��h�j�����H��\c��A��G���I�@wd��o$�#̺�E�b����G�z�M�v��ڴ/Z�
��r�#���B�C@��- �Ɉ��&�;
uy�u�٫,�t1�]�vd�ٷ\�.ܧSb�[9��p;qE����k�S��Ձ��s`���1�l��=��ᙗ4ܹ�-̹�y$���s�ȣ���Q��*@wc��}6�^+*�4)Ly�@�빠{Ϫ��g�b]_U�yzנ�W����LMnf�ݎZǰ@z�L@8� �	JdMI��n-�e4�y��?�o>ŀ{ծpI%<�YvMR.����C�z�FY��ϕ۝�F���C����ck�4�1�(��pXۓ?��|��� ;�˺���`ۊ�陕0ۣp��������������ֽ �#��0��lNf��>�@�v�=	b�"@D!}�������JIa$	IB�B¤���
����J�$L�	�IT;ၠE�@ՋbB2�x��!$��P�)̱?0�����#OFR��B$�0����I���B##W��n�x$t�"�� TpbE�dxq ��<�ɶ�$)C5&��C��#�a�`�! F0(:��0�
��T�&
��  E�WN��� q������(��� �q����#���ξ���s�Y�P�N������v���wW8B��o��ӽ��(_Hn�b��II!!E7�Ӏy��32曷2f������'���g>PKd��{�_%
�ݧӀn�b�$������w�s�`����6�I᫧�Z��FOfj�M��<-�^@�C��.�ι�����W_}2n�b�>����}?���G֪����}�������7�1�����O�:���w��>��	L�w����]
%��J�+���6�j��l�fۻ��x(���9$�Es߾π��ŇB��3�]Ӏs���dܪ�%t(�����;�YС)�w��)����(ȅE�0� pQBw��ß����٘d�M�v\,۫�����4���}!����@;<�!�9	$X��d�#�tv�p��.�쩤���n�#ۣ$�5�o��|7αP]U�USV��&M�����/���ua�>��X��jx����j�J�ffO�n�ŇL�w��ov,ޭs���>>��s�cQ���}�ߒ;��sJ��|�z���jz�N<!0�"q�;�T���-�������)��w%E�����V��=�x�(_Hzw��>Q�����?(�P�G�Hx~�?�VNχ����n���7�<�-����N�:�j.����`ϓ���֢N��JP��9��"�[��¹2v��8��n��=N�g��)���X��Q�[�ۍvu�i�n�S*��݁z㝰��K�ZV_IZ��v�݅h��t��"�b˶Oi��N@�9�ֈ8|q�$�>�^���2;�Zt�4�����ͨo�7��nBi�B��Ef �z�n��ژ5pl�z�ngݱ�'mfɜg\]Y`�t�c�o����~��?� ��urI/�=�؜}'�B��:po�}��Qc�7&oٟ�]��@�wb脾�ݧӁ�(��}��}UJy\��vL�%��gB��=�ذ�}=
#��ذ>P��V�V�#���t7h�����&M�}8��]�N�V����}��;揱|HҐ��h�E��N������>�x�z��/�=�z]�<��x�[�:s��u�tl�l�]�R�J��L���O-�b�.�i�#R����t����;�T�}%�,.n��fI�79$��{ß⸑ DT(IBQF�>�|�����P�S����p�@G3@��V��uՇ%
�	EV��V��� 7F56��ĞG�8�.��z�����\c����dnL��1�"��I�� ?~fܫ��i7t:ӡk�%ۣ�U������VS�'�=q�Cq�V�dU��ڱ(��7{�`N�X��,Ӻ� �AȨ� ��@���+��@����<���=�w4գ�RF���RU]`�x�N�K�
�	E�`�@$bH�X,�z�" x������y[^���M���%�4�hys}1�6\�ȩ#��ʼ�S7rAsWX��`�Q����~�s@��^���f�O瑀��L�7i�:�\c=d]��hM�B���%��ZK�������4����w4]���S@;�\S$nF��=� �1�6\�c�V"�G��3@��^���M����~�m�b�M"I��7� �[u�{�����"�P������� �|��A�s4��������R��+%�n݁y�*��������l���]Jn�_s�8>C�v#���5282D��w�nhۘ��R�$���0�ڻ���7v�i �� =rL@wH�@��f�'I&!0�Ǡ{��h������_�4
�~z�ܮ&��6�,�si�b��Hm�@{�����"�1&��z��s@�:o��=�ذ��X�BP�X2��4y/,�^�}�z5�ܙ'8m�,�`���k��m��u�Y�*�ʺ6ιhv���t�Ӻ�����I�v$n)��z��;�η!��aq�!�ү5%��ɮz�|�q�x1���Ύ҉괰�J�f*U�,��8�3��8�d��,qm�ێpu��1�����w��>=�.m�Q�.��l���e�/{���=��}w4���&8�<�O;���fl���q�]K�����.�?υ�ch�#�g��;�Z���*�����~�m���a$Z��,�$�_��������� �79�'�9}��F������=޷s@��Z�n�գ�RF�&ER)��[��uv�޷sC�_�|�|_����D�$���:�V���M����w4g��Y&4�f	�E��Nz���;��zY�C��3��t��#ě�%I�bq� �Z�e4Vנwu�������}��cXH��G�9$����?)�^1\@A�BP�}�ذuwN�7� =�M�sV\UT�+���=��`t���!D$���s@����=Ϊ�Hb �2%]��۬�o���(Jw{�X��o���8�z������~� ��ذKn�K���$�<�6�*ۛJnn���k9y�AŖG\�s�ZHI���)���qnf�˭zt��rL@wH� �X�ớ��U�\��]`�x�����߫ o��X�����n6G"l$��9�����x���G]������Xz按�yH�`��@����9u�@�����w�wU�&��2ch�9�'& ;�T��Z�EH�n Lw\�5E������5e9��N7��Il�j�R&o;���|�W\�c��������H2K@wH� �Ɉy.Y��J�E��U��<ݳ:d��ŀ9���=�w4���+�a?��H!�{�T�w$�t��M�Xu�av75r���K��w���9&�&� I�� `A (T�OȐ�#��~@�7�7ӒO?L:_��nKY[�������R�}N^��"�.��-��qH���rB9��H�;�@�g���Nw\��΋�z��r��ٵ˦dO�$�L�=l���[��r�_ٙ�w�nh[�f�'m��4y�Y��Q�߿V ��ذ7l�{e��(@mG3@�ֽ޷sO�f%DB�}w��݋ >�cSv\ݫT���SWX�w��ou�{�����_���~��~��Qj�3TM\U�]���0���|��X��,��X�DIfh��#ŀă�1]�v���$V������,"#�#  �>(��(
20����x�O$���0 "�A!܄���J�J1��ct�I-�A�1�XIr�0	�1!	 �Ą���2����#	=���-fJB�.b���`B���8�J��C��TK�)�a�`0.1 @��Z�1%C!	HY$�p!DZh�k��(��F����xAͲK��8����b��O�G�1<�I!��_ ��CA�W�p�Z�1 X�B
��a?Q �$R1����"�]�| ��.��� H�a$�,i�Lbas,H����V��1L�`�r�s��?n�������-��č���Y�<gNx�lmwU�v�3�֬H�� i�rv�.l�y�v��,b���Cp:���.ζ����օ�"y8m�++v�*������Ql`*��F�ֵ�gE��Fv��8�j�	��8��j�L�[�uhӢ����pl��@�L��V���9:�<lL�M;gCH�V{f�L�s�PS���6秡鷋t�\�:�;d���T��j賮wc�F�eθhj+k���E�l2�뛎�]nc	��[�h������Y>+�=��8p�.�kYLs-��%����tm�\sʕJq�vcҩ�K��m�κ�9m�j(8�u&L�:��n�9%WR�'8��)��llA�Z�mu��� [^rC;f��l���ɋ.鈋����j�v��n����*gc�udP&�f���;gj�s����R�÷E�㋥�\��%C��v����;�k�m�G�K���M�z����ŗ����٣i6�R�l����KS��Xm/!���.9�wlѤҙl�keT)+Z��yl���6�6�E��@�D/d�p���R��^�Ѻ��{a�5`ۄ)&m2����9�p�v�fu�i[�Ͷ�P��Į�Y�ؑ��'��.I���H�ٹ�kmóV��jk�N+�.�7@u�W �T� m���;pb9��qN�Mr���dM�kk�^� z+�l;�d�ɗ�=M�iPMl�M�tR�UUR�J��8�N���Z��r�9�#��:_���䁶�t[T�n,Ut=��ۥj�]��c���N�fލv:�f=j�س��j��m����Nv��`�������񣇉��kF����c���g�ڕ����^�X�e��Hch#t��\q<��XC;�N�G/X�6��ei9��3R��r.V�c���L�66vECM�e���2|���>m��Z�b�4O-<���|N��u�Ms��;=>J�N*�TC��O����y�C��z��﹃)�ɛ�`������a���V��g:��RQ����M��k�l��e���=9C�v��A����V0.Q��3ڥM��y �S�9�q��I�DFɏ�v49�v�L�+�y��:��u�t���6�s��.^z3g�z�-����l��h����K�v�Ֆ���p����.֔a�fSF{v�p=vwNnگ�����;�3ژ{$M9I�M�]��me�ml�b�2�4GWe��)�a2�H���}���9uu�{�����_Hl��
n�ʹ��5V��n��
1$�+��߱`���@����:�;$q���7#�@��ŀy�f�w{�`_u`3Y���D�d�)3@����n�˭z�n�{�f�'o$I�JC@�H��UT���t��&� ۭ��^`b��F+r;��y76^��vDn^e{g�]&��<����N�ŭ��n��ۓ�*@t��� uBUݛwl�ˆ̹��'�����PI DQ�R!D��}WO���� :=�ۓc�f�I�PN93@����e4�b\��@�빠���\ L�`�,�>nـl�u�n�ŁД%��Ɓ�E���iŊ9�.���*@t��� %ϞsoC4�F&�5�GaӅW�N��m�u7n.�<��=����ō$q��#����;�w4Y�@z=�U}�y& ;�Y���^V��n� :M���ܘ�|�,�JS'7�FD���+.n�f��=���6[u�˚Q
3+b�u� ;�X����G3@�ֽ׮��e4;�܀����"�27������{Z������T�w-z޶	�&3��H�Q��m�=-���k����r�N�m�z�=X�]vyH�n'!!ԓ4�S@�[��r��׮�~���p�?��$�Hh�w4rL@tqR̒������ߍ�nT�Z�6[u�y�Ň�DL�s�w���:�v*8�I�G�Ǡz�Հy�s�|�ف�&D%jj���>���lRF�Q�$��ڴץ4nL@>qRѐ���]�����\�י���a�՟V2{4;p�-�����ֻ�C���8�J@QŠ~�)�r�^��������W*��ubj4F��E��0�n���S#�ذ���� ���!I�M����빠z�V�����˭zWȸ�26��m���� :d���{�& 8�@;է��cQ����;��h��-���M��%�� QB>O{>���K6m��\�r��,�����\WX�샱u��5���U1[wj�t=u�L'����ĕn8�Md���~T�>:���p�v� �q�:�d#r]==�,���Y�6�q���=
\5iĖ6����Wc���l�G�u�R���z�����.�m���A9� :v���۵�����n���f�ݡ�Qн�rZ2�^d��@�t7<��z*
�` m�fK�%3vBn�q]��j����JfkW��5μ�i���4��B0h����B5�s4/���z���=l��? ��ۚG����ƓDuj��� �׋9BJd��� �;� �ֽ�;&*)#I�$d�4[(��{u}UWn�L@>{n^�&E %!�~�)�r�^���^��e4��X��E$1H�)�Ɉ��:M����/Y��sة�����5�YDhNW$�M�d9�;�{�ۓV3nAu�h��[#?6ߝ�Z�� H���`�$�<�EWa2]�J��� �v�i(Ԓ�E�o�ۚ�ֽץ7����/��H�h��{�4]k�=zS@���A�Z���jE�s4]k�=�np7l���w��9:Z�)L�x�Sn=ץ4�ΪS@�[��r�^�޷��LB��I�F�0��u�vA�ٶ�.u��	�6孚�働��ols���$ǒ8�Z���=�w4]k�=�j�/uL�� ��ڐp�>nٝ
dr�� o����0��lMF�n,Y��˭z[w4���T�!?BP��Dǭ����0�qHE�d�7&D��:۹�z�M���9u�@���<IE��i�lr*@;rb����߹/�Y7t ��2�JK�A��=�i�9��&&$y��nx�c�m̫���p�k�r*@;rb�EH�%�%,�9\�2	AD��h�׳�#�빠u�M����9T���Bb���s��&��"��& <�V��VZ�v�]�wk��;ݜ`߾��'���9'�AȆ([�~�$	%!�w���:u��<���<ݳ �I{�*>��W�a��B���[�2��z�g&!9pnwi1�-��-�J�8I�6���w�m�����:8��l�T�;�J�ݽ�S���@�빠z�M�n�˭{�GW�>�2�,�bƤ��w�O�|�,:��\���7�b���RW�A��Hh<]�f��ֽ޷s@���ŞG+�!Pqbnbۓ� :M���H���G�n+�6�CM���� ͘D��ÝŎݰ=�`^&<u�UZF�ed�ɐ���\�=��A�{V kL󸗐����Bk\�}Q�p��xLg�t�烃�z;���;nmi��a��n%��=�r=��TN�Ur���jx��1+�
n�lR��E�<�d�>L����uڔ덎{X�/ovv�Y9�Dpftp����n�W���a��z��/�t��}˟�LcN婛�	�Lrm�����Ӹ�����C{��{�u/�\�+c<Z�Y������*@t�s��ܘ��m\7"S��I��z�M������*�|�w�nh��o��L$d`������& ;�T��6����IF���Z�z����h�������Bbi92'��7� �v��o����"��㝍�sӷf�ԀV���udW��S�i����K����<���)�iv�9�k�?߷���Rۓ�*@q���4%�)޷s~Ċ��=��4[)�\Y�r��%,ͤ�& ;���l�*@:T�tq�m��16��=�)�z�M޷s@�ֽ�;&*G�Ly#�� :M��EHnL@wd��u��ut��!e���v���Gc�h�\�6^y�J�c��N�݌R:�Xv�gd��"��& ;�K@t�- w8�ԑ�G���9�.�������h�������Bbi92'+ ��ŀy�f�.5B�!%Q"�b9�;�*j����<�`��Y�3c	0@+c�<��a`�+XA$g����\]8�OT?wD0�0@�*x-=�E*�E:: x�(Q�	-Q��}� ��u�{i��]ԣ$K$rf��e4{��˭z�[�����\�Q4�baZ�������ŀy�f�$�����4�,͉ҕl���a���a ��}2�&U�{�^8{v��8�je볿 K��b�"�I�@w8� �e:�H�&�P��q�������=�w4]k�?S�b�q)�������0y�XtD˗�X�v,�n���A2)�@jC@����9u�@��Ł�	L(��ـ��$�����E�nm �1�"�I ;�]�m���pSuϵT��s;��ؼH;vY�C�h�n[��$�jG��T)�m��Z.4������ :H��"��& =΢㑬B	��ɚ����"��& =�*@s3*Vh^٦��a{���qRۓ� :H�@�G\fHx��������9����EH� \d3sr�0�-M�]`y�XB�������`Oo{��<}@�B�� � F�n{m�.i.��4�Ɏ\�ۡ�[e-�j]5���V�6�ڙ�a� =6a��\;��)���+&[�NwgV�٦omh���7WR�0D:��s�E��0#�4A�c���^�k�V1$붶z�:Dq��p=�|�O?&0�� �(U�΁"�Iŀ @�=��dGX�w5��]�q�f��ݶ{Vݻp��:�ͮ�����l	��q(���������﻽��t�wѠ�E�a��+fi�E#C+F��S�=��qs��9������ǒH���_�4{�����޷s@�Zѿ�Ad��ә�{�w4Vנ~���[w4ު�R6���nm �1�R� ;���z����S#Cs�z�[��9"�s��䘀��Y��E�훷u����rEH� �1�n�~�F�x�?��8����4��=;p���si�rO]��.7�n�G�\����7��@wH� �I�� �s@��غ��B!ǉ��+k�?�:D8 |�<���$�����޷s@�Y�\X�M��b�ǠwH� 䊐�*@;�b�u�p�r' �9��ح��{��˹@7�v�}kF�IȦ9�3@�qRۓ�@t�R��*��с�j�=��ܨ�����)g�8w�J�:�/X-�r��v�1�f�M�n�m��߱�I ;�T��:\���pQ(��@��)�z۹�{�w4]k�=΢㑋�dD�d��@�{��~��xr|h��R
�$� �"F%D�����`��S�-��g$�~���O:���b��@HRf��u��9u�@��)�z۹�v,�..c�Xdj	��ۓ��$T��qR����~;��ڶ٩G�kuWc)�H��<��U�:��v���!��]�s2�*Eř��=�*@t�R����	s��@{���� �NA�rG3@��s@���w���X��"�˥V����@w8� �I�s��H� }�蒮B��	�wf(IB�]�X����X���KaV�[0�j��o�h���޷s@�n��t������l�$��	���7#l�q4�N��r�yY��ݳ/�ݛg� ��#�)8������Қ+k��s���+�0��%n�v��`�w$��$��*@:��..c�Xdj	�h��@��j�:۹�{�)�vW����$QLQ=��EH$T��{�& =�$$�$S�I�[w4{�4Vנ~����gB���7xA�;ѻ��_�o|2s�-�L@�姮���rڢ������73�u$Y�Ntk9�Mɮ�8�WK�5d�B��#gj݌���b���+�sn; ����	��1��[KK�-���ű����0vTѶ��L�d�a���9��Ƥ��L����ۇk�o#Л�"s��2�<�=�l�	�'��;V�V��.�G]?���{Ͼ�]�k�.�ݹ������Z���G&�m��Er���D�6��繚Ǆ�C�C/6�	?l䘀�=�� ��U�U�h��v`-����d�;��/�}��~�JhG���m��R(�z�;V��n����@�ֽ��\rc_�DH"D��=�w4��Z��z��Z��r���
`ܑ��h�ڴ/Z�s�z��ֹ4䁄�,R`�(�C:{u��U�9y4�v�m��c�vH�vM�-wM�^�m������<r�T���V��^\u��H26(�z��[��BItD$�%	,í�,�Wt�>m���1RH��'���Šz���?s�h�k�=Ϫ�=�7�H$����@y䖀w�b�9h�*@��C�$�4H�^���r�T���-���˼Uf�F�SW8Xpgb�e�t&��e�NQ�u�/�\D�c"���m�H�$q��s��*@y䖀w��앛�}�Y{����h�*@y䖀��1�� �R�XLSbnH�s4��Z���%	4�K�}8�v,T�)��'1�����^��}V��۫���;���ʺ����ʩ���<r��*@y䖀w�b9��Z����[�C��F-�x�ۛ���3Y6�1�8�۳{d���R��A����H<����@s�- ���$��&���;V���^��v��빠~G�b$Q�q���$Z�s�K@z8��$�Y�N6�$�2I�@�>�@�빠~���I����&�z�����y��ȸ���Ĕ�1E"�/��h�@K�1��-8ђ�:�L�Җ�ηIs����g@��LN�.j{Y۞M���k�����]�m���_r_9�v9h	�*@:�ul�W��*ɹ��0>�Y�(�*�]~�8�߱h�Jh����i1��z�Ss�?kŇ%;���:u�`3U�w7e+��T�]U�����`����]`~����o�p�yd�ss5D��Nf��t��W�����@��ÒN��HB1'e$�  �V@��Ȓ0�B���&����!aYpFЀD����np��`XG� ��u|1�(R �[E9��@�
����-HU�BX!B,`� *�P#�u���'k�ZKD�aX1"�5H! �T-J!H�&�	��-�P�YX3�C�tc�ZH,� $"�bBR�1�$ �J�(�����#cX�HF�H0c�X�R@�.D��1BP�@I4e!BU�� �_Jx(cFw�X_8B@�~A�T��� �	A���=��%fL��IIH@�W]'��h����""���$�$Ǔ@�)R�}����ݩV��vR���qrg86y������뭪3�oY	�eU#;�V��k���k�Դ]�B�H��@	����R�U�a��"U��M�������%���ul�UK�W�iLn'��$�F�����CkqĀ���Izh����i]v�)	Z��kj�svn��;j�	���д��9ݧWY2��r�V�n���]i�����	v�<����.^�6,�ml8�6�۶yr�u��.w����Ol��r\�ҕ�J6>qk��그�C��K������۰<�KrAkt4\r�ln����]�Q�g���H-�c�v�ZFge�%������.�ءE��i\�P	��z1;�@�{Z����-�kH�n�� []#��hӺ��K�/I��p�.�1i�:�'�m�YڥL�"6��2D�g��6N��ԀUuH�IA����ȥ��e�g��q�D-�cĹ���Ҝ=�kn����{V�+2�\�:e�<�0#s��M�K��/-�f�]��i睚����e����`�j�b�h�+��m��� '@�v9 ��@糵�]v	UڪU�v(�0���퍚t�&��Z�\���]��j�\�		�mq�ES��[I0���',E��� � ͷ#[w-����A�����UG�2i@��/NP
B�p�s�JV�d 8�z`���K��p��`e�,��+[p�5��������g���:�܇O�J� �m����In|��59QYQ6�3*�Kf���T����UuV��q'jb�r���Ӱ
^�.���zۗgPl��*�D�$���m��]��(b�i..�Ⲓ�-�smɵ�3K�����:%�ֺ��5֓"���\u�wP��ř7T�-�:�v��2�c�L���v�MR��ي�0l��q����P�V�ء6-�8�e�\8#��L�)�Ɲ3p��eĘ�Z.ά��3f]�������_F
��Q=OQM=�U�" z����*�� ��ٝ�po�W�p�9�.��E��ɹK�1�؉�	�7g�X�k]�j��Gg���D��N�9kr�.'<�<L�{�Ƥ�;u66{Qɍ�m�"ڷ:sѹ��ܝIq۲�N�{N�o`"���]'v����V�ڷl�1�;`8�e�s2[���gs��(n����u�k�m"�N�n���@[�Kѷ�Q�K�g�簠��Xܝd���%@��מ��e��z�<���q������K�[c�
��6��z�[m������6k"lR@����|��=��f ��%	}!��dnyM]U�c�$QǠ~�h�w4{�4
���ٙ��_���cȉ"ƣqh9�R����@{�K@�n���SeM��n�%�u�N���Ss��"'��� zR�,䦕�.U���_9�vIh	�*@w=�����{���W�sF4�Z��`^��/k'$�X���ɹ#l������֡�|9>s�C\]�����W��8�x�{m�Ϥ:v��|\���A�d܎-������P�>�	�����Ɓ���=���@�sY"�O�eTլ��f �u�>�����z�"Dؤ�	!��������7k�p�x�?(���0[�SWT��ڥWj�� ����:#����7z��*�W�u1�*y`�d�B�/K����2�U�nYMWU�a��Σe5�jꨫ��WUW8��X���k��?�����@=�W>a21(����{�ٝ2t���7k�p��9�d�)J��EU�%ʲ���:[��=�np�
F@�K$�T$�Y�]Ӏy�� g�:gwn\͙M�n�������h����{�S@�����LV)F8���@�v����~?��{Ϫ�;<��Y$Kf	ƔSȤy�lH'k�<X�E���n�����9!�X�t��6�7Z�YM���y�_ff~A�?�Z�1$�I�#fC@s��:��M�}8mwN���?BQ(:��'�&Lyȓ�@�|�����G�S��~��Հ{i�����o!��n-�v�޲�.��MS�1�	���$�߭��I�
8��@����˺��v��v�������H�B��N8�"�y4�i^z�����Y��+�mu�tsZ��w���,[��n	dy�<���@��U�_;V���S@��q7$��L�:��=�ns�I/СU�w��Ц[�����~���� Ҍ��8���h�����˯�@�|���5���� �qh���*�W�{�S@�}V�{�X�x�ɑ�	!�Y���=��`ծpy�0	��"���|��?��9��j��K�n�u�.w�m�c�=c����3v�l�%�թ��	lJ7ca����e��]�8�d�=�q��=:��d'F�;��S���ݎ��N����O'����	7M4��n�܉=�����(��S�aP�;u���n#�ƣ`�;���N�m��A��B'p�t=��g�{uԭ&ս�F�
�A�<y�+Susk���~ww~����o��&����j�����_,+��؆��wg\f�p��qխ��i.yms�u�U��oN �Z� ���С/�:u����}$N�#��Š_>�~�Ď�>4�_���;V�~�vVF8�6��=�)�U�O���z�@/�U�~�x�p�0��$�������h��z�e4g�\u�ܓ�28�z�e4�ֽ޲�����4�)�@9!`��j��C����Y8:�]�[b.{q��L�E$��77f y��v�g��DB�Cw����ƲH�L#Jd$�@����ĎNנ{��h�Y�$��"D�)2dl�Hhw�=�v� ��4z�h���&,�dMǠ~�Jh�Y�~�Jh�k�=΢�I��IɂmŠ�f��t���ֽ��U�mrx�?��8��̃Y	����]�<e���OR㦞�=0�X����h�b�ڃI94��M��z�>�@=z�ݏ.�ōFc��h�Z�Q&�>� O�^���9)������ܑ�$Ƣq��|hu�4��� z!����rI���H~����#Q���Hhu�4޲�+���h��5���������t� �1�6�s~m�??6-�כ�՞z�e�F��9��6�l;ڥ��&�<��w]�q�����Q���s�`�)�5�6׋�����4�z�e7���"����޾0����BI(S&��ύٻ��73p��ͼ� 4�������lll}��}8 ����8 �}��>A�����ߏ�5�ͻ3sw��A�A�A�A�߹����lll{�w����lll}�~��A�66
� @r8}����A�666>�R��ar]�˻s7g �`�`�`����g �`�`�`��}��� � � � ӿw����lll}��}8 �����Y>�!3wr�ܸd�t�c(	/��)�Ei��q�л
�;��pY:��3\��Ɇ�nnpA�666>���|����;�~�>A����~�ӂ�A�A�A�A�}߳��A�A�A�A��l�~ۻ�r\��7.i�� � � � ӿw����lll}��}8 ����8 �}��>@S�@9��{>�<ɳv\7s.i������lll{��N>A�����~�>A��H��A� ����|����>���x ���%��awt��wg �`�`�`���ﳂ�A�A�A�A�߾����llli���x ��R�A����|����������3v��34�ss��A�A�A�A�߾����llli���x �}��N>A������g �`�`�`���cD*��e�?�.�ws�@��ݲ����xnN��@@�3sY���-f��6WUZ�ō
)��d�cٸ�u�.j�{c��cUf�V�v���	��\�cF�c�k{\�όÑ\�t�W��\��u���C6O&7cG6�����E�������Jn���$���6�'vz�ۚz{sņ������e��F5�ܮ]�ܽqzՓ^k��{����Ϋ+��l4ԎjSr6ق5��a�NKV�μ��s����u�g �����ۗt�A�6664�߿���A�A�A�A�߹����lll{���pA�666>���|�������>0�]!���[��|������ϧ"?�$D29������ � � � ����|����=��o �`�`�`���J^ϋ��.n����� � � � �>���� � � � ���xpA�6664���x �}��N>A����=�3�ۙ��0��w3s��A�A�A�A�߾����llli߻��A�666>��>�|����s���|�����g��ܺfnn�ͻ���A�A�A�A�~���� � � � ����pA�666=ϻ�pA�666>��>�D<�~��s:�Y�/j�gg�3�5�r���qh�b�GW<�i�F��y�L�]c�v�q��w��e��v���>}x�_Q%\����u!wf���R�J>P$� H#�E������C�l�=�)�Uˋ���r5���q��`�)�5�6q�@s�e��6��(�4:���e4���?(S��� {�yr�qrT]ԩ����t� �1�6�sPo�}��O����57kW���c���x[Dv�8+���gi)6N'�{������úf5"��]��@����g�Y�{�S@�^;q8���N=޲���QT�w����e��Z�jF�"�	E!�׬�=�)�n�B��X4�D�����!��2D��d����dU�0�")�: R�?�X2�18��XO��E�@�@J�j���U�B0�	��!YȲo��>��@$H�"Ab�!�O��B|C�D���t�!T�?�H!�֩ �S@I�<�b*��? <0�x��(��f���5�f��̡]�ͩ��j�5w��)��� r�� ��ŀ�٠�ubC�$�4C@��^��%�$�����~�x�������i�3s��<&�+�.��ۛ����ƶ����؛�� 놵hN
��=��`��x��	G�_u`���$��1�1(�� �[f��YLg[��or���}3˕+���Q�Srh�O����������5JT���ʩ�n亻09DB�w�8�_ ������$��"!7��|ـ|�����]]���ʫ��t� 
�&�;���$���￟���nz����R�\�u�/3t�BrWk��e��]��[��we���1��<����h���=�ՠ{�S@�KMfG! �	���=�)�s�-�6�ɨ�����2�whܰ���$�t� 
�&�;���W..'��&�qŠ{�S@3�l�=�)�{��@�:��6Ȧf���MY�����Q�8�u�8�v���	BOK%wU���7���GmiwX�Gk+p���U����^�@{UR�K���/*yg-��9l�ɭ�jx�<{/Gct�󎖒�h۷q�l��Ku����ր�� �u��4�F�[�lU�"wnz88�b�%�	m��d�567UN�c�!c��{�*hѷ�j컂N�x��9ً����NuF��;)���+��) l���w{w/�<��շej���.
�`��\��z3]�8��k���mض�V�u�]�͹Uw���y%�=�`�+������b��pƘ�Dr�ڴ޲���f��t�����'$��$�-�����[4�.�>4���)�:�qBL��Hh��,���@77���Z�6BAa[�����Z�M]���0�~�I�~�>��� �u�@��L{�K	��ɑX��kG[r�t�le���;�M�8�[u������P�8�Hh�j�?z�h{���Қ\�����mbnG���O?w{9�+�
� ��6C���wY�{��@�:��$�FGJn����n�{m�rQ
g]wN��|h�\��`Ly��$��=�`�np���B�Z�� �T�K9MZ�UUv����=����{{8�;ﾚ�Қ�\���b#1�#�C�}1ɵ�!s9��#�&����7]�~:T�6�䉎29��NH7$_��}>4=m�����D$��n�� ��6��z�]]nV��{� ��j��䖀�G�:"L������5pZ�U]����7i�����3�f /6� <��SaJn�Rv`tBP�����ۚ�����M����nIyy������H� WI5���C��������rv���f��B���t[����rr�)�lY��:3�Ϩ���w��F�Ռ�(ԙ�����h�Jh�ՠ~���R�q�Ȓy��&��=�gD%
dn�� ���ͻ�?v<H�q9�ㄒC@�v����
)�s�u���j�V��'$�-����g��@��SC��C��?
���쿻���LI��Gp����m����"��>���;f��]���E7;�]��z��A6��wWFa��oS��8��.h�$����r5�c��4{�4�\�y�?D$��%�?߿^ ��Q-@�d�(�Hh�ՠ~����n�{m��QTt��UMLҔMUMN����sy�{ݬ@w���YrD�I�bOi�@3�٠{�)�n�s�Д�{8��\�Z��w3E�^f���䖀�M� �rj$�S����^͘f�RY.h�̈́�Z���ݍ�F۬�Ղ�':檭,�e�ɇ�0�tq�l��v!�+D�In�yܱg��f��7��{m[���
<�z���{x�n5e'��ZW�U�U8.��]��2�	�{vrR�M�rm�AC�F)�j��1Y�{v��N7gBd1\�zh�ɼ��&۝�F�6���(w<�؄��&��	�]��%�����M�A������~��2�3=�*���e�ŋ�
�w	����i�Y��u�tsY�}=po���u6���m��'�@{�� W95��g[��G#NH7$Z�YM �u�@��S@�;V���_FH� �܆�-}׀{�l��(Jκ}8����ֲ�uv]e�Wx���u�2~��lyɨ�����	2LI�$4s�޲���٠{�l�:!{�"�+U���ʹۑ�0�M�>�m�@������ڃ�;u� �^�du�72<I����ƀZ����M��h�QrA$�1'�4�ιȅ���f �k��;f :�eǓ&9#N-��M��p脔��_�/� ��S&�SV�U����ݘ	)�Ӏn��ε�{�S@�y\u�������6�@wM�Lr���2����V��`�sZG��ɹ;[e�7]�l�nsl�ms�s�t�@x.���&����;�� �9h�@t��I8�����=�)�u}V��YM 꺭 ��� �$Ęa$0u�py�0��#!J�KВ�	E/�3�`�O���|���ץ4.\\R7�%$qŠ{�`��-�61�@s�r�����BO��@:��@������Z�e4�s�Jb��N9"Q�G:��m;<F{Kt�G-]�Kk�6��i˶A��(�ra �Ӌ@������Z�e4:��E\ʦ&C"�P���;�� S�j�l��b���Ԑn8�z�hu�4�ڴ���=ܔ�ڮd�d��A W����<r�z�꾬;6E�z�sY	#�$X�L�@�]�@�Z�r�yɨ��T`V�]��H�v.�|���:�\�m���R��f�un�Z������`I"�=Ϫ�;���g�h�e4
�qqI$d��)#�-�u��~ �~���j�=Ϫ�:�U,J&G�������@s�-��r*@]��m^�R$Bq�}�ؽ�oƁ�ߖ���w4?ىx�|�
����Lnȣh�D<r�� L@{������5pF�"��)��6 $���A��XB���!�R0J=!!��V"�o0 B+�'qM4���4# ��@����o�<��$=�i�����0Ԅb&��¦	����	�a�\����~�~ lYd�mn����D�$�N��#�V�i���Rl�v�`ѝ��qYӂ���H�0��� �.�
E��&)6̈́8"�&��2�<'m�����;*mT��];tA٧v��[u��H�$���]�Z�sSs�Æ�
�t�W�Z�m�a�ñ��J��ss�u;nɊ�����d'mqSқػsWm�1q�j��eF���]e��\��rR��̓��U���Z�
lwVb*㥶r�lnY��i��v�l���S'Cs,v����vbB8S/V6{a�Y3ٷ��=<�]����^ٱ1H��e˪�7mt��N��an�`�#rf,j��N�<���138öl�k��qӤ�sE��`�t�vRV\�$��q����;k]� Cɫ�6h8�nx�,��a�c`��<F��@De5�t�1�9Kfy;vw���A�]m���N�`��FyH��r���uyZ�n���gq�Ӯ����mV��>1�����݃S�ON�3��M����ko6�`��/Cm�E
�v� �m�<-�M��g;u9&Uv����g�by�vm�c��L���46�C�vZ�� v�b�U�q��]�ְ�b������S�� �D�n� ���H=
	;<h��jk���x ��,qp�n����2��vDT�OpM��.�Z"1䋙b񓱷��"-�c�욚�ym6�v�$ڶ:Ҕ�6�:h:��q� �[v����\[3�l����Iq6�����ݤ�[4@���RV,�a��<�T��|���ٟc��c.;���m��h�\��ZMy���:9B=	cc�v������7c�m����Vm5n=�ڃ�.����t�+�i:v2��e'y�-�3U�e.�Ӏ7TYݸ��;泲-�B9�6vX��j.J���	�$�8F���<���㫗n,�Ɯ�r�^�0k��c��-��tuK-�ZK���v���?=�z*a�ExE�;�L@����_B��+��+���=��!y��b�Db�%%פ�tt�o�քl���nK%�T67���x2��.�^�D"VT��k��@���F�0	�kpY5���Ι`c1�����ݫӴ:k���V��ac��]WPpդe��ur�O+�-���I��=���3n׳Z;7g�tA�H��^6�����8��M���@����p�737K�犋��yK/�Ɵ-�f�anb�pt��O�s�Շ���a���e�Iڝѹ ��+t-Yf>�>����[��m��%�}8��jh9�15�'3@?k�?{�4s�8�׋:B�=�O,����UUXU�������9hs���& ޵�q`�G�0�Hh�31u��{_b��n��DB=�8��r��h�d����-���h���~�gƁ�v��{���4�2 ��H�eRnFC��grs��s�gv��9���;���wK-D�l�LLQ�3�����t���v����h�\���'����'�s���@VD�@| 	e:��� {v���������\LMǄțy#�@�|�u����M��S@�r�u���H��@���`�i���fBP��;��TLL9�15�'3@=��~�[0����m� ������]R���U9딭嫋�t@�c������sJs̘�'*nw>��������&�$-d����|��>��?/���`��b��H�I�}V���)���8��f~����ge�����T���n�pk�X��s�B���"�	M{m���8���.�Aw�q���h�Қ��?���DD*�߼���������-IV�����1�@{�T�)��������.��U7GR�On��i�<��ը�&��d3�:wnӈ߽��ۗ|��c�W7T��πާӀ}��`�u��}!��@��/��!�nH���:d���=���>��9�%2{��k�	0�$Nf�g��h�Jh��Z�YMޢ��RH�7LS7P�`���-���U}�Y�@�;�'�<i�I�v��6������2�U�Z�a�nrس�2��A�����g��B���s콺�bn��Z��ɚ^1._�������H��x��g(K�:}8���.�.�T�ڛ��0}��?%	(S'���>��m�?B��tu��R���6��u�o��Z�����I=���p���n�w2�ݜ��P���pk�0}���J}�8����̍I�F7Z�t������Y�~����� �k\��$�d(]$"�@����O�'�m�.�lm̮����=���?00a�z.����v�Vb���3$㧨�\��g�
�bHc=vq�>bpli�z
KN#�`�v��;6#�7�k�ų�y9��' %���rm�1�[�3\�\�\�6�ؓkn{a���Yn���F�ݠ�y�̉�h'�;�곮5� b�c���q��H��O�Z�K×9�!�]u�����{������O7[w�R��PR���ͳ����Z�O-�΋����*I�G�!�)
�_��@���?s��3? �Y�}oط�&6�ɑ�MȀ�=�����y�����:��<i�$4W~Z�t����Č��M�gƁW����,�wr�m�{^nj��?W�W�_�����D�L��n1�$4?w]@{���Z��{Yr��N�����]+�,gN1�lq�s���:�'���d��F���5�m��� �ծp���IG�����L��f�Lܹ�n�����o?���`�"���� ���>��0N�ꖪ� ��7Z�t��g��4�fg�^�>4W~Z콓j��
aH�y��s� <��@{���8��]�&h�5jj������DG������� ۮ�N�;�\LҐ��z�)=��n������,�E��[��1׭�n�I̎18�H���?s���M ���h�JhyqqIb�.�f�p���G�
��߯ o��~��h���Lk#c�Hh��� ��م*��#��J">�]w� �})�UNed��cq%�cRM�I%;�8�5�t�y�0{[�f�r�92(��x����v�����g�٠{�)�w�@�EFcrF�nj��$6�έJ��2�4�������n��ٟ�F���s��I��"���� �95��y%�<ݛW�s6�
�T���X ���j�"�n��5���'����������p���Kn].�3wP�� 9㖀�H� W���=�s5wB���UB.���
�J>��9$����9$�����:���B(��i�WN� �����YV�U�]^fm�=�*@�&�;����������go�z�ڪ��B��]�Y�[8m�=13�����
|tF@���=������S�q�3����@��S@�;V����hS�qțF7L�ܓ@��ـ{i��>�x�0�$)!I
W���<���2%��[~>͓7I�����wdND�,K���^'�,K������Kı)���x�D�,K�{͑9ı,Os���3L˺Ct��ͼO"X�%���٩Ȗ%�bS����<�bX�'���"r%�`|�"{�}��yı,��/۹v噦Zn�٩Ȗ%�bS����<�bX�'���"r%�bX�����<�bX�����"X�%�ꟻ;,��6
vJ�v��lDF�]7^u�֬���;u̵���.v6�i��(Yk�rZ�h5�����^in�z�k;��i�z1�mHɵe�a�I�p:��]���ѵZ���z�a\�1<l�9T���-�9�8 9e$��Mɒ�VGsUa�&��W��I�ݣi�����g=pD�s�)Mۭ�ËWo2s���e�w����u��n?^��������N�5�n]4O$�mp��h�D���ƧӞ���s�s���t��34�ݤ����D�,K���"r%�bX�����<�bX���f��<��,K���oȖ%�b{���K��Kspˌ���,K����oȖ%�`���jr%�bX����x�D�,K�{͑9ı,K������ٚe6���n�'�,K������Kı)���<�c�)��;߹�'"X�%����׉�K�q��߷�5Xr[�5k��{��,J{�{�O"X�%���Ȝ�bX�'��{x�D�,K�w�S�,C{����ߎ��GtC��{���d�,O}�6D�Kİ�R>�Ͼ�O�,K����jr%�bX����x���7���{��>�������K牎�+հЬ�g�FƉ�k,f���sZ���ݷmܲ�wdND�,K�w��O"X�%���٩Ȗ%�bS�{��yı,O}�6D�Kı;���饷f鹛�x�D�,K�w�S��@�A E('X @�B����T��'��D�%�O����%�bX���l�Ȗ%�b~�����O� r�D�{�4�n�ۛ&Sv��ND�,K��﷉�Kı=����,~DP�DȞ�~��<�bX��o�S�,K����vf䙚f��n��<�bY�,����Ȝ�bX�'�߾�O"X�%���٩Ȗ%�bS����<�bX�'��r\��[��f3wdND�,K����'�,K������Kı)���x�D�,K�{͑9ı,O��>�^�s�Tѹ���M�#v��a%�x�"�ͺ^�rȱ�k���������W2����Kİ{���S�,Kħ�{��yı,O}�p�Ȗ%�b~�}��yı,O��ݳwns4����ݚ��bX�%<���'�,K����dND�,K���oȖ%�`���jr'��L�b_��d�$˲Xe�6i���O"X�%���͑9ı,O�ｼO"X�"���,h.T3F*EF@DD@�!#pT"D @�X"�i���EA�<?C� 0bRG���S��		Uѐ��P<�zP #�� ��  `)�]E��b�P���=��MND�,K����'�,K��[zw6L��ws0��"r%�bX���{x�D�,K�w�S�,Kħ�����%�`|2'{��"r%�bX�ϭ��\�ܓt��ݼO"X�%���٩Ȗ%�bS�{��yı,O}�p�Ȗ%�b~�}��yı��=��w�:����Ͷ�X�i�-�Y0:���6����t�N�[Ӱ�m�
c�(�fl��ۻ5<�bX�%?w﷉�Kı=���'"X�%���������L�bX>��MND�,K�����76ə�n�&��Ȗ%�b{�s�ND�,K���oȖ%�`���jr%�bX���{�O"X�%��'�ܗ7̻�fk74�Ȗ%�b~�����%�bX?�����c�ș��﷉�Kı;߳�ND�,K��}�.�ɹ������'�,K?�H߹���Kı)�~�x�D�,K�{�"r%�`|
L����׏7���{�����K��0ݘ�IȖ%�bS����<�bX�Ȋ�~�dO"X�%���߯Ȗ%�`���jr%�bX�����ۗ�B�,�X��sOJ�*��]�b�=1YRuu��O&dl�9t��F��_=���7��,O}�6D�Kı?w}��yı,���ND�,K���w��KǍ�������[R��m�����,O��{x�C�DO�@
�M�`����"X�%�O����O"X�%���Ȝ�bX�'s���6�˹&鹛�x�D�,K�w�S�,Kħ����yı,O}�6D�Kı?w}��yı,_}4��٦f̺Cv暜�bY� ���}���yı,N����,K�������Kİw�59ı,N��Op��!��s)�wx�D�,K�{�"r%�bX(}����?D�,K߾�Ȗ%�bS����<�bX�'� |�ZN�T
��o�I���L�m��b�b�O���Y�S�	�n��B\��P��&i4ܳ���m�����'X��{W�n{v��h�ն��b��Ġ��Px�s�2�خݞ4��`8GYp���u���W5P�-��b��죓/L�N��A����m�b	2��u� 7��96�[@F�܇���W�U�v�{r��[G^Yw���k���]43��{���{�����&�ཚ�5�Z��Z9Jf�862s=/k��auڝ�V�6���d���swiwY��'bX�%��w����%�bX?����bX�%=���� ��"X�'{�6D�Kı?g���nLݙ�\���%�bX?����bX�%=���'�,K����dND�,K�w��O"X�%������.��I��|��{��"S�����%�bX���l�Ȗ?
���;����yı,~���"I
HRBt͡�U�$���-M��B�Kı=����,K����oȖ%�`��xjr%�bX����x�D�,K�m��4��f�a�wdND�,K�ｼO"X�%��!߹���%�bX��w��yı,O}�6D�Kı?u��\aݒ3v�j�Vb���sW�s����c8[�m����Gl.�K4�f�ssoȖ%�`���jr%�bX������%�bX���l�Ȗ%�b{�����Kİ}��S��n��iۻ59ı,K�}��<��P>Ar&ı;߳�ND�,K�w�^'�,K������Kı;�<-�si2��ܹww��Kı=���'"X�%����oȖ%�`��xjr%�bX�����<�bX���~?\D���{M���{��7� @Ȟ���x�D�,K߷�Ȗ%�b_w���%�bX�����,K��?_gK�f�ɓ7fɻ���Kİw{59ı,K���x�D�,K�{�"r%�bX�����<�c���}>�����l4�ʵI�h�XZ�'l��RS��ޛ�j��n���g~���c��\��]ݚ�D�,K�߾�'�,K������bX�'�ｼO"X�%���٩Ȗ%�bw;;��2���mۛ���%�bX�������L�b{�����%�bX>��ND�,K����'�?�2�D�>�o��i7t�Ɇ]�"r%�bX�����<�bX���f�"X�z!�r'"^����yı,O��8D�Kı;���:M,ݓf�swoȖ%�2�s�Ȗ%�b^�߷��Kı=���'"X�%��w��'�,K��ziN���ن���59ı,K�}��<�bX��ǽ�<"yı,N����<�bX�����"X�%�������fBl�[��X��1擬l��q<O1�GXvgh1���]jN�-wN���76�f��n]��?D�,K��8D�Kı?w}��yı,��ND�,K����'�,K�����K�v�K��f�9ı3*~�=��~�O��ݩ�s﹓S�3*dLʙ�~�x��Tș�2'{��92���������2��"A~�~�WݢfT�9��&�"fTș�3����?~���a�Sb}�3�T�Lʙ2��s���w��{��S��s��F�QnF�����Lʙ?��M�}�OߪdLʙ﹜��"fTș�?w���?~��3(������ o ���]ND��;ܧ���~;�l��s������ș�2'{��92�D̩�������L��S �w�u92�D̩����^�¢T¡D��M+�E���rF��Ӻ��3e�
�@n"�,>�<��o��q�䮋.��7�Os�2��s�^'��2&eL���2jr&eL��S=�����2�D�y���"fTș�;���vM$ݓv͹�����L��S �w�u92�D̩���w���L��S"w��YS�3*dLʟ��{x��Tș�2�M)�����.ݹ�592�D̩���w���L��S"w��YS�3+�؛�=����?~��3*d��d��Lʙ2�}�g���ԃ5������{��;�����*r&eL��S����'��2&eL���2jr&eL��S=��'��2&eL���}~8�'���ǻ��)�w�ʞ����?~��3*d>��}�MO"fTș�3�w��~�S"fTȝ�3�T�Lʙ2����c!@�
~����J;ء���0��sm�k��-ٌ�An��b�:;bhۂ&M��Icgf�$�ܮ�����]��S���a���Ge�:�]!�z�'(p����m��r�q��!28ćW�!��ۍ1Y�̎A+�������xjD#�ē�Ђ�kp�]rtV�!���tZ�O�����.usi���n�� ���
���I��o�������Ӷf�-���j��.����4���h�m�}A��וZ�������/��i��S ���ɩș�2&e?��~����ڙ2�D��g,�ș�2&eO{�{y���Os��{��~�H�
\�V���Lʙ2�{�{�Oߩ�Gbn�ȟ}��92�D̩߹߯��2�A��r�r&eL��S��ܝ�4ܖ�ɻ��ww���L��S"w��YS�3*dLʞ����?~��3*d��.�"fTș�3����~�S"fTș�>��\��B犀�|��=��)�����'��2&eL������Lʙ2�{�{�OߪdLʙ��6ڜ��S"fT��oL�5��nY�7v�?~��3*d�y�S�3*dLʙ�}��?~��3*dN���jr&eL��S��{��=��)�w�����3��樫/i�L�7(hm��kKrmmӸs'E���c�5�T�;.�C:�|��=��)�>���?~��3*dN���jr&eL��S����'��2&eL���2jr&eL���������x��TJ%_=����w�jdN���jr�^�92��}��'��2&eL��w�592�D̩Zۼ��L*!UL*!m�����-\p��mND̩�3*{�����2�A���592�D̩����'��2&eL���mND̩�2'��gK��ۦ��6K���%�g�2}�٩Ȗ%�b^�����%�bX���lND�,K�}�O"X�%�{�l�wne�i��ܻ����bX�%���x�D�,K���Ȗ%�b{�{�Ȗ%�`����Ȗ%�b{�yfL���jN�Q��2�V���{1��6��.Eqrvp�<��Z0.�ʾ�������,N�{�'"X�%�����'�,K���sC�A�I��� �	�s%��i�t�w3&]ݰI�<�����ؖ%�{��"X�%�}���Ȗ%�bw�ݱ9ı,O;�z^�[�6�r��<�bX��{���bX�%���x�D�Wb*�dM����Ȗ%�b{��É�Kİ}�zS�����fHn����Kı/��w��Kı;��؜�bX�'���O"X�Ȁ ��}���bX�'����nvn��˛��O"X�%���v��Kı=�{���%�bX�w��ND�,K����Ȗ%�bwݽ6i�at�.n]��r�g=u��d�������]f�D�g�<��:)�ۻn])3a7v��Kı<���yı,K;��"X�%�}��w��Kı;��ڜ�bX�'��}�.�m���6L�8�D�,K�����?�9"X��w��yı,O��m�Ȗ%�b{�{���%�bX����-�3��=�Ou��=�{����w��Kı;��ڜ�bX�'��|8�D�,K����Ȗ%�bw;;���7#��n����'�,K>�{�br%�bX���xq<�bX�%�����K���؛߻��<�bX�'s�s�M7sn]�ɷw19ı,O{�|8�D�,K�{���Kı/��w��Kı=�ޯ����oq���}���$�]�S@V�u։x��e�nՠ&�z�^����v�n�(v�v�I�ݓr͹��Ȗ%�bY�{���bX�%����<�bX�'�{���I�L�bX���8�D�,K�J}����K���7u9ı,K�{��y�9"X���ىȖ%�bw���yı,K=�wS�,K�����I����ssw��Kı=���'"X�%��}�Ȗ?���,��n�"X�%�{�~�'�,K�w����q��p�K/����oq���'�,Kĳ��u9ı,K�}��<�bX�'�{���Kı<�o���͗Mw2l��q<�bX�%����Ȗ%�b_{�w��Kı=���'"X�%��{�'�,K��~_B2`�!=!1��J��1���!&bL�A �'�!Ō@�P#@�`!�BF*����%��	��\��<qHU D�z��A(�%�`HC��x�0���!�`LX����������y�� m{H�3
b��oe�������-����� �W�bKc�8���fw�ط.�q����ؓ�sգ�s�hM]�:C�$��R��(7H�k�#��ζF�u�s� �����~|>I�4�e�M���8��(H�N-�ִD�1dց�H7M���Ck'`����[��p�1�/Mm�f��zu���mJ�;oFz�{��d�y֤��n�!,�x�3�y����*9�m�t��@�c22��%p��z۞,�Ob�gSU�h��O"�
�ѶP<�����ds�]D��+pm�-�ܯK�5� /d[�4���.kr�@Z��wnK������Gl�t�m!��k�M�P��O�W���mujN�%F�t���D�/����c����V�P�筓��HXI����)�N}5mum6D�tU�fю�����e��'�;�+�\���gm�҃t�;�X�n/O���;��6�5!T�0��)�l:��[U�m[]�N҃��	z��P���v�Gm�*�vW�b�[
�5RK@*R6 �i!2:۬K��d�ݝ�U��vŰ�mm[p�\�����ֶ4l
��Jn.��"F.j��ͅzڠ�9��e�$7^��HR2��HfCpv�[���)-�T�7%��2�q�. ru:Xڠ2���̎p-���V�K+J�qB��-���ol0�B[<�9@(�CjK��jc!pHo[.:�[M�BN;[v� �����y::g��rr�MO/AZ�;��*^8#���(	��lh�V1;z�5/.��5�ة�sы�oQ�v�fxv�M�+��79-��藨9�"���N�òl��A���s��=��֛��s��l>����\��iݞ��V�4�>�sZ:�[4��G-�F�� hԏe�ͥ��K��hv�%���K��*�u�O����k���c9�h�����6�`�C%��� ��P�TZA:�
	�P��<(�}DM���=Oy,�'�7s�n�P����{�Ѳ�	[��i2�g���] �U25h���6��q�s�X<�4���=��dz�qӆ���F:L�r�.��n�;ڝ�{A�t��n�	;�kW[4��B��^d-��;Rk���a������X�ݎ���m;cl�;���H}��������{|y��ʍP��_,���#t���bKa�?�����>�.�f�u���ܻ��n�p�,��3O/��d�.��]m�=�ޔ�X%�&a���u��Ŀ��}�O"X�%��^�19ı,O{��q<�bX�%����Ȗ%�bw;=�zd���̻���%�bX���s��J�ș�������%�bX�w�S�,Kľ��w��O� r�D�=ϲ��l�ݹ�e�n�br%�bX��߼8�D�,K�{���K�"^�߷��Kı;���,K���OK�kt�˒���8�D�,K�{���Kı/����yı,Or���Ȗ%���(L����q<�bX����w3sin]���Ȗ%�b_}�w��Kİ�cݿ}��D�,K߾�É�Kı,���ND�,K���7N��D�۩h�u���iܶ���ϡ�z�9�-���i���Ȗ%�b{���ND�,K�{�'�,Kĳ��u9ı,K���?��oq���~~o��@ܜ����Ȗ%�b~�y��� �� _�@ב2%�g�߷S�,KĿ}���O"X�%��^�19�ʙ��v�|]��t�n&n�'�,Kĳ�}���bX�%����<�bX�'�{���Kı=�y���%�bY������B��f狀�u�ϹD������%�bX���ىȖ%�b{���Kı,���ND�,K��ܗ���ݛ�2��Ȗ%�b{���ND�,K�{��'�,Kĳ��u9ı,K�{��y=���oq����W�36'JU��\�����ܣmg�D�X����e;(�]Y���nK&\���Kı=�y���%�bX�~�wS�,Kľ���� @��dK��w>ʜ�bX�'�/��ٗ4̷K��8�D�,K����r%�bX��{��yı,Os��T�Kı?w���yı,�:S����e�Iv��"X�%�}���'�,K��=��ND���|S�̷ı��P�H��\!Uu!�'�<�?xq<�bX�%����Ȗ%�bw��x[���f�s7w��K��C�UD��>����9ı,N�xq<�bX�%�����Kı/�����%�bX��;��v�ۦ�.l���S�,K����oȖ%�aԎOs��Ȗ%�b_}�w��Kı=�s�S�,K���N�0��Ƥ�ݺ�#�e�a�8��7`W�6焃������F'gª�������)7M�3O�Kı,��S�,Kľ��w��Kı=���'"X�%����É�C{��7����\T��z����7�ı/����y�R9"X���ىȖ%�b{�y��yı,K=�wS�,K��v{��4-�&�f]��yı,Or���Ȗ%�b~�����%��0ș����r%�bX�����yı,O�ܹ��f��ɗw19ı,O;���<�bX�%����Ȗ%�b_{��yİ?��S��r'�^s19ı,O�=/��ٗ7&K��ͼO"X�%�g���r%�bX�s����~�bX�'r��br%�bX�w}��y�7��ｽ�k�k�m��ˆܵ�C�9�Gɴ�Al�v)ͱ���c�:�3a%ۛ���bX�%����'�,K��/{���bX�'��{x�D�,K����Ȗ%�by��x[���sp��s3w��Kı;���ND�,K�ｼO"X�%�g{���Kı/����<��eL�b}��s%ۦ�m���73s�,K������yı,K;��"X�ș���x�D�,K�}���bX�'���:]�6魹vMͼO"X�%�g{���Kı/����yı,N��s�,K����'�,Kľ�ۥݻ�fm�ɷL����Kı/����yı,?�?m����%�bX��߾�O"X�%�g{���Kı?����~���	�tC���|�\���sӉ���c�f���Y�Wl;��6�
r���nI���Gh�G�����u�tX�d�V�㗰�'m�n���s��j�b܊���V�ۃ�I�В�2WVs��Ӄ��lUWE�������)r�ݮ���S�>�|B܀�]�SZj���6�znq���=W&w[�U1ѱUh�Mײt�ǻ��ۗ���k��JCWM�шp�.�cm�t#����k�9�٤�vr�����Dk����bX�'�_����Kı<�����Kİo{���Kı/����y7���{���/z0��de�|�bX�'����<���1ș��w���Kı/{����%�bX���s�,K�釥�:l˗L�K��x�D�,K���"X�%�}���'�,K��_{���bX�'��{x�D�,K����ͦn�I����Ȗ%�b_}�w��Kı;���'"X�%�����'�,K�&Aϻ�jr%�bX������.i����ۙ��O"X�%�ܾ�19ı,O����<�bX���ND�,K��{�O"X�%��d�!��Y���\�z��U�3�T�F�ݘ$�{].T�]=�#u�V�lS�]T����oq���������<�bX�%����Ȗ%�b_w���%�bX���s�,Kľ�=�.�m��3r웻x�D�,K������E��DǑ9Ŀ}���O"X�%�������Kı?w{���%�bX��{t��wL�ɦ�\���Kı/����yı,N����Ȗ%�by��oȖ%�bY�{���bX�'s��;��B�.i����yĳ� dO�����Kı?}�}x�D�,K�����Kı/����yı,Osܹ��\5�������Kı<�����Kı,��ND�,K���'�,K��_{���bX�'㾜)��X�PE�՘�F:6�ڹ��k��q�6x�yn4Y�T���k�̼�5G�w�{��ı,���"X�%�}���Ȗ%�b{���� #Dؖ%����^'�,K���|S�wv��K�����bX�%��{�O"X�%��_{���bX�'��;8�D�,K��sS�,K����x[�t�sp�f�n�Ȗ%�b{���'"X�%����gȖ>*���B
�A��'�r&A��Ȗ%�b^�����{��7���w��]T����D�,�P߾����%�bX7�����bX�%���x�D�,K�}�br%�bX��g���ɛ��˦ɛ���Kİo}�jr%�bX��{��yı,N����Ȗ%�b~�y���%�bX�����e�l���no"�����kl\��L�\&3!4�Gr	�%�ɗ�U/�J;WCK�����=�{��{߾�'�,K��_{���bX�'����O"X�%�g}��r%�bX�g{{��em�6�nn�<�bX�'r����Kı?w���yı,K;�wS�,Kľ���Ȗ%�b{���/I��[�Y-��ND�,K�{��'�,Kĳ��u9��@!�2%�~�x�D�,K��19ı,N�z^��e���.���8�D�,���2}�۩Ȗ%�b^�﷉�Kı;���ND�,��ME�߾���yı,��J}���Y.���r%�bX��}��<�bX�'�}�br%�bX�w���yı,J=wp��$)!I	���|R������K��[��>6y�sl�e�5��<&#t�����[�l�n�l�3m�nff��%�bX�e�ىȖ%�by���Kı,�{���bX�%��{�O"X�<ow�����WU�m,���oq�X�w���yı,K;�wS�,Kľ���Ȗ%�bw/��ND�,K���:]ܙ�5�ٲf��yı,K;��"X�%�}���'�,~ dL��_��ND�,K߾�Ӊ�C{��7����\QW4��j��7����$)�n��)˚n�6�`[f��Z��!F9�Iɠr����, ����w�|�%��7ow��c��?C~�kK�����cú^�_OCi���*�6u�\�g*�D:z��t{tM�zϖ����{��<�7lX2����m�b��q)���m�5̹z��W�)��!���8�1QnS��у�=�8��<b��`ۃ��k��m��0�=r	��enq�:�^׵[�Vۃ�F�9�ۨ��n<�ո�+C���Qq�K�"�4]>�{��{��-H?1�շEJ�j�ms� ����z�����v���n�5li���׊�`����?��X���������5<t]ULڻ*�`�w��DB��� s�Հy��?(��G�')]wrM�p	�&�[��@�z���� ��h�����㑨ےh���3�1W���7��`�w��$��o����K�T]Ъ�.�� �o�D�}�-��r�^����?d	��՜��L�۫�\]��6�v���[Mq��km��vdj�N́$_�;���t�?.� �Ϲh�U�"n<s$x�wPrjʪ�GՕH��s1�@��9DL�n˙*�\I3Wx��� :d��I��5�d̬�LO'�$��=]�@;�� �hW��.,�T/�H��s4|������ϫ �o��n���������X=7.:UwEtPݫ-izM��Q1�{NTIlu��-W��c��5 �9��*@9��
ˍ����M�4W��=m���f�w[7���H�_���4IrrV�݋ 5��I!LBIJ�B�y�H��"�,b�y����`,6А�l���B��D�  1d"0����-�]E��0��dE�A �j  �  �$�(���h�=_�X%1����
���]��)�o#�hT��"�� Dq�	͓PC�s�c�@<NH,
4j["�W��?J�SU�$0��`I%!H�2V��M@��ЊD�H:��y$��ӄ�.:�����Jֈ����Q�"���T�<�'��`��7�a�kP��@;v�W�E�nU�mPMZ���L�}x ���/]`=y���TH܀�qĞ'$���@��'\��y�, ׮�z]�z��TQ))b�J�{��U�,���G-(�v{9w܃I8�cn.���k������=x�^������N�T��!<��L@��@�빠z� �[x��Y�DL�)��tj䙛Wdլ ���@���& :H� �X�e�`�I��ۓ@;��+k�=oxrA���^nw��I=����"H7$�"I94Vנ�?���|�� �n�/;)��Ȧ�աg�Y9�oW�v�:���X�Un�����K/����H�$�70�Ǡz۹�r�� �h��@�ˋ�L��
�`-�Έ���׀9���<�������o�����Q0�
��m�����<��@�빠r�^��eb�"Ădb1'&��mz�]��Z�>_����^���_��4�IspL����g[� ׮�Kn��"	 �b�T{;�f}��Ͷ�ci4M���v��8�X���	�iz��4Y����S���� h�)�OJ�n�v�t<��mq�>��׋ȱ���]��k�٩.�RZ��Mv����y0`э�-���Xm�0��$���u��.M�bM��E���T��g0�x��ݰ�`�u�����-���w�1]��|S�:���mY5m/Tv�Vލ�M�썞2�ݢ�������|�c.噴$f��D�қXu�:u�Qf�����p��|��.�\���_qtm�y �8������z���z^��:�\Yd� �1����f���?�9}~z�ύ��z�k5r,nH�I7&��z��Ji�,Ī�z~�M�:�"i�a�@���g�� k�x�"v��`.Y�b�cq,Q���˺� ��h���zS@��B�#��O�j��Uz��m�Z��Q�g���<������6�픍U���M
G�z���Jh���=l�S&E�L�F&��?&�g�Z�"aR���"h�����Հz���w"���q�z�h�נz�����.+�R4��8���Z��Y�y[^�׮�բ��$�s��I�u�rL@8��& =Rl��.�vY
燢F��iGk�;H[sH���!�t�Ѱ�^sk$\�O-KZ����~�~ ㊐ܘ�sP�n�y�x��9�׮�˭z׬�<��jG*��������9�.��^��a$*_�TD�+3f�� |��~�W�H�l��z�٠~Vנu�s@��@�l�S&LI
db1G&��^�@�n���^�u�hz�dq�F'q(࣍�jx��A,=��ݫ:��Y��7Rq���i3����m``m��� ��PW��*ˊ�D�!)���9{�@I�\sH� �X��n���#RI&�u�hVנu�s@;����f�IȘ�rA$��?+k�<����w�I&�_��HY���h���!'��S�z�]��(��_�{� �[u�}���:�+�f�΍��;�;��^w[X &�K�a^U��4��v\E٣s1���m�??>������1��H�.U��������)&�w���mz�]� ��7���}>b�2!��#�h_wV��I)��׀_^�����X7�k�z��s@;�� �k����wu`+T��ws336��ͤ ��@ɨ\s$T��"����vgY.l���r��J�k���p�=��	��P��[�\��^����n����u��#ю���gn^��=��c�X��n��wn���1vܸ���7F��\��ơ���!\�Wlд�:D6ݶ��-M��Ѩ��d�p���0D<x �ci�d�r�X��ΰӺ��Ŕ���{o���|W��C���<n��m]���݆������hEO
�g�wvL�$�ݗ7.�fܵ�)�Y�8��g�OLn��I�כc9��e<d�D�A�����M�^��n��f~@^�M�~kq&�m'lI=��9��*@�� �M@{�u��	8<�9���s@;�f�B�Q	L�{� ����6vtjnl�����+s6��5 >�P�� :9���U�$�<Q�Ll#�@;����G �j ��3j�(�<4$�tڐ�[h�s4�a습m�IQ��X�]��1�剜]u�:�GpU�m�>�}~� o��(��@{�x�:�W+��.�.I�79$��{Ø�����!y(����o:����Kn��9����Jb����@;���׮�k�,&$����@���9��*@��u��I�i�ē�@�^���s@7�� o����Ұ�Qr�n
������I��s�L���mG&���/a�x���7u�pg��H��G�L#�����4�l��Y�y^�@�����9?�LfD� �j |�:㘀�qR �K��qńy	$��f��z�?����=T	���߿��� �����?[+�O呑���rh���>m��z��m���:�W���O'��۹�r�^�wu�+���y$?��I"�&
�E�Gk�jۜ��;=�+��vç�qt\��N#���75�G�Sng�*�����h�W�~��hG�XL��LM9$x��y�(IBQ29���=ϱ`/[�=�Y��N6��m%�+��6�a�._u`o� �켒K�	�s%�]��D%�V���� ��߫ 7}��K���������������b��(����Z���hVנ~�)�{��@M)�$rLi�`�=qgp�u��V+��<s�\Gs�\�+v�3����$(�x�G��f���z�^/�"?/Pt��Հ>��M�V�.��+3u �9�I �1 >sW𯪒<���dX6�1<�z����������9{��.,�.+��H1ͩ���_�!V���X�߯ ��u�~�ՠ_0�X�L��LM9z���	��u�[�'۵���
"?�**+�ʢ��������������EE�EE�QEO�TQQX(  ��
������**+�**+AQQ_ TTW�ਨ�������EE�
����**+��QQ_������(+$�k"����i[0
 ?��d��-a�   }  B�        
 � H   ��@���		BJ�JR�� 
P *H(���J�� "P(
� 
 �!@�I
�   ��     ��4�M4ـ4M4�L@ � ��Afh�wpPk4�@�` ;���I������� 3�/v���)`����z˓^�ﳥ\�R� ��}��|�r��:W6�6wjU�  �      @��+��g��y5K�[���\ zn^��Η|�=+���Z�β�����Tɯ��ͥ,YK� :v��oCswof�{���=��� �^�7T��.��������_ �� P  � )� ���[k�}iw���������w��{^ N�z����nv綞Z�{�r����ׯ0  f  �}���6|�� �{U�=�}<�WN�=�}o�wM8�=����{�^{u�ݼ۶��n��|�P( (�   � �}i�v�rj�n���n�N t��>�+͟Zriz��T��������Wy��  	��p���y� n��ͺ�n-�W�ܯ}�ŕ]���R�e��u���� 7�@��   P MPR�ﶮ-��qg�W>ܯ[ŕ, �����S���W�J综�yG A��s� q)@ �����)J0 �i�14PR���R�oYҔ (�i����Y�4cA�K0   ���U)   D�I�Oe)J� hǪ�*���@�  D�*�)� �OЕ<Ԥ��!����"�&RRSDɠ�ZL��w��+�W�M_��j�P���2r�6NNZ�L��+���
���DPT�eTW������
��DEO'�?����_�H��l��$`���M��$(ib@�JA"D�@�10:1�yM�$���h0$��g� jSR�zq��4cC���#��j*t�D�pr��DrH�)"BbP��H0�^h�`�bB!�`��B,B%H2$ P�D��`��J��$$�i#tR"�Ѡ�u���42l�D��`B�,Hh�*B ��I1�B��KT�4�a�$`AG��,�V���Hk$�p*ÚQ��H��;ݡ�R��&��$�,	.��Ԑ)��}H�b���B��,d�$��� Hj6�paM9!$������j���6p���H�Hs�tƌ����T�	Ma�Ã
��o
����M��P�XS0��#E��q>X3|>)"h2];�ڐ����
�!���'J0�����@�
�$�h�0�t�t��|��B�ԆMԲh��-&���T5���H0�K��8�)�6Q�B��XI	kv�!�6ER��bw1�DW"��h0�5�»��S�#$�i�j6�D$��.���2RXSK
+��SXh@�&��$`P�1�����SGXIxO��_��9B:�(?"0bE�@�D��0i�F�*%+��	B\vFA�ܦn0���&�l�����!@�I1�j!*0�)
D�H�iSA�J"�pm���[�Bu�))�aT�
D�V�+��`5 ��VWK��0Q����9E#�� �$�CK�"`U�HR�HрP�	0�#a@�H5�&i���.�w�7��vK��2g��_g�_a���;��2�?-hɒ?ERIk�p$J���<�~��xҀu6�O�Qu�q�]���{}�Z%?~����?m3)Pb&N�џ�)����ފ�fMa����\�ö�{��I�~C�P\��ǀ��E��?�6ف�QI"�����ަ#��ݭSl������{�M���~O2��[I�w�e��z
�;X#�~�}!k����NL��T�Jդw4���SPq���)�ɢ%,��"�bA`$@���R>P5� �"&-�OR �`1��SR����f�!���:�5*�4�PAb�S���$X"����A�+q"0 �`����:��
���]!)�IyZYI$7.�4͝%�8��3Zq��ڒ��*F�F(c�1h˗��͚c�>%u3��T�h̛xbϒ��d�L�0�*KIJ��)�_�]I0�фh�L!B#4$Z�`�$M��f����$�'97�S��&�5`B|n�Z����}�q#�$�I�	�x9#&��G:��c]M󐦶q�,,)"�@����Y���v|˟-��T���[�Lnh����鄸}�9�3	Y�g���]��]*�(��u��Ŧe�)����l��H�;6`E�R5*i���u�8��E�k��5�
h�FMl6]�T4,���I
��K�
B��-�2�P�%ф��ߍ5�`�XU�60�(��!B4H��9������ax1�jB�	M���9���*@�4hĠN��A����$B,Z�׸�#����!M1��ӛ����+9�J��k8�Ͼ�%�m�$Jo �B82��;�XK�ћ�A��8���`�4�`���L7u218�SF�6�b����x`}�'5�s����L6p��6c�� G�
�iH��t�
�D��Xi4u0��%4�)����Y�%��wM�vS43
�Yf���SG4o��/�5>�)�h�So>�\� #������B�$HĆ�c
�(C��)H�"Gi� %4f��P��D4fu&�z�R���!�lx�F�}����!M0ϙ���|M�fφ!s�%ޗ�9+��H��tx������(D�e.���MaV)����)�$���Ms����XB��f�ÇCE�Hң �����*(�E���e5xMݛ8t��]&��n����8B���+�WH��Ȧ� �|���c)��^�X;xa�$�Ƴx0�s|}}͜� f|�&�7���uܗ��:m���ą]$�A�i"��3��C�4�Dڒ�e4X.�[�g�~AHU���B,	H`�4}h�Ӵ�ƌ�4`xh�@��$C$ ��JjD�&�B@i��� 5�&�握�lRl�6E��kg ���9�]h��ƚÌ�ͨB��фn�HWC����4хt1)�"�e��%�laC���`�/�<� Ɖ�
*��i�%5K�ԛ��g�%u\�'�'Ȓ�	�8�D`EJZn]f�����a���]���	�%�vS���w���BVaaH�!H,"F$b������Nk3�WX��Z����ף��R��U��D��!B0!]@��4�
k����2]f�˨i�atB�i.�C7'h͜xH����L�}��8�亡�����<>�ܹ������|w�9�J�,w�H�v��]oP�q���5�ւ1��tA� �C��Sl��	RXa���q"$g����u��SL�h SK�6�c 8|� @�``�x����p�L���YX�ekW
d�b����4�HXQ1��]�����bF�q�kf�́����a@ц���H�8q"�фɢj��sW���Ħ��5����s�.^a5�̻u�4X@�b��5�� 0�HGp�"1
k79�e��Kxi!3V�������%�.�R�V��)�SP�aHV#F��#����v�:LM���4���C浙�L���^g>��@�`Ku��3{���n�e�ߧ�!Y�SD��H1��hA�SD�����]A 1����dv�G�_�vJv����!�Hq�0"M�g�4���WF�x}��}�C��W�_��A�"�H&�Hc3�#���fgR��s�~gTp7���'�	�/NF�&�s�4¤:¹�i�S�8;9�2�$ILܷVpv>%5�!
&�� I���2]���Y���48�� ��.+�Q�N���BWP���8j��.vw\M�����j�.��tdhu�ӾB�H�!cD�M|X���K���6��6��	lK��z,ۭ
	�$�=%u�a�Ҝ7��ӎ��u.��4��G`D�+�Ɣ����E���bB	 �$hB�,H��F�!tn��IB(B�x�Ѣ�4}5�Sif�.���|5�� |<H#d�o�``A� Catb�2m&h���	�K��.r6Y6Ma���heѽ��:�at0�B�0cF4�?���
Bᴅф����8�N�J��{;�l���vl����SY����)�6��h�h����f�:�����fd���4��6m��6B�t�8�.s�#])��d��@��*Ɇ�_�n�6���'&�aM!]0.�MNsz�i6�{�yM�k���Nk]QYxa��Չ�����N[��!5�ޱ�(�֎o�����a�_i�d0�aټ8��d�MC���(h01��f�7sFݛ1l
l!M�w��$4b;�����w�)�]H]g6��!e�2���
�ja�M~\������{)u1:;Lù��Ѱ�aIL�᧒A���j�Ć��׺�u�0��$\7�s���K���   �   ?�m��      p       �   � m�     %��65+����;�䛫��mqT(�[����<
�\�����6�������3$Gngcv6ܑ�3���YuŞZ�i���l��\�֊[������� ���J�6L0$v� Ft�� E��6�n��l�"�kl��m!��    �m8ïCq�ж�	 qm��   	J�T*��]�`�]�m�[D���5f��UU]��ԌlY�7h���n� �i�N%�ul��az8�lx�`�[�i � �37a�������k��, �WK*��k��JP[P�P;f���:t����B�ɭv�����^w�|��k�m۵�k��[jU�]�a�m�\��h��e��H�t9 ��2�N�����c� � ���e�����2'����}�8[\���pN���m�/2�]U+��4����ej��U����@h�h�@�-� -��pkkk�� 8   �eweV����{���8 ��$sm��������$�[��ր� �6��m���yknm� H "��	�6����ݍ��':�6�6�5&�U[U�nʪ��vڥ%�@
����jݥC�#i6o��a���ݺ��j��`�3��6�:���
��uSh
�.�N���i���e%��iV������>��[w� �h =zvF�{.��4�R��մ��;mղ�R�Kg@�S��Ӏ�$�� &�a�U�P6����VVU�*�M�����J�QU('[l�c$mɌhMm8�5u*�=m��e[e�H8�M���j�h���UR�K�*l<�UF�l�1��ق�:N8K�ٮm�lL�ʬ�ʷ]��N�e��@%�S��D�:��_�~G�K�ʦ-R�JB���� ��J�m�S��Z6�p$��n�0�95��E��@7m�����MK�W彴�����ŒJq���m�-�䜝 m�mٶ��e	V���U��G[����� e��L蕀Mw54��+m��I���'j�l��E�à�
�� 衲�n���Wluёc\�]R���k�*�  �ɬ� Y�Ā�l@K� l� ���k7Tn-ur��UM��]��H*�Z� �I���h���kd�ݺM�Z�  -�aͻb��l�M  �I{Vi-�6sm��am��v h۶ �`�fC���H8�c��k` 6� 3��o���k�$�v�H�X���m�2�n�� ൺ[G��|m]KC�����/7cT��v�ձ�� mY�lm��f�.��۵���m�m�q�j�u�֭��-�� ��Zm���[q�pZlrB@��m$m!S^lk5�Hf��ҭV��T��9��m�z�����^���@F�pA`gm«j��j��i�[lp �`88l  ��  8W4� pv�mm� 8mR��֤��m���$pm�C���ȗ^��kv[@8�	m� ��k5���f��]�@�� $m%�v�K���m�m�	A�Ͷr��$�j퍷�$��h[��m� ��m�Tu]����$$ p�Mn��i-	��KiqT�Uu9;BiU�Kh��{-��cjؕz�C�O���QJJ]:.����6ی��.�U�p�+֞J���6ݚ���Z�5m�V+hZݩ^ݬ�R�4uƞ��V�\�e�}��H�� ��JH^�n�i���l�^h��� ��%���6� ֜ ��uN$v�kbs��5��A�.�V���Uz�h$-�ɴ�﬙l�4��o� ����8�0�� 8���붓 /Y)m�[Nu��7j���	5([d�[�2��j@�v��vx8յ�m*�m��   6�&hՕmY!�)[l$�n:ԉ6����;[i$�6�X�� K(� 6Ƞ0  t�2M� m��ޤh�  p[m�:@�-�m-�U��mMR���١�m5n��Ā m�ӵI@m���g  n۳i6  ^�j� ְ 7m�/,���[��@����\k�lҶ-�kDd�!�e�l 6�m�:j*�m�PCf��U�����PAj��������U���\�l͒��l 		$�����pl�� �i6p�)m���������I�m$��5��
�U�����zT6kj��{=.�-�����YrM"@I%r�N���� �l�m��]n�HH )@-� $/m�6���m�l�v��m�( ,cm��AT����Í�Z�WfNN�\��Hճ��=(Er��]����}�>r�͸��uu*�r���+K��X�e��wE�!!��M�HmV~����Ntg2)s�u�z�n��a9��n�9Fwa��f{g�mͶO1v�]��ћ��T�}���k,� }%ׯM&��L�I�;v��� 
��Rv���`r��W@n�ۀR�,��k6�BKnCe�� ���d�D�[�vm�$��I& ��׭�-�% �/��d٭SU3#�#v�{I6i�	  ���m����,�c�١��5[J��R�U����}�Tl�`��	 z���h Y%�I���m��E��s���R��ۇ�d   6�T�Z���j�  ���Nk�ksv�`m�b�[�78�>Ԁ�ktڛkn @� p�f��;��:�v����\x�I�h�[l4�⸴�ܐ3��;: q	9��d��'@kX� �`[m�CE  �|���Ț����v�8H�h0 M�d�A�@�����K�u�  xm�icm�����ZN�l6�&�$���` qͨ��-�k�V��ٮ��oj�q��tV��c�m/�ͷv��9�>a6�Tn�[F���@8�[�&�gPIf��x�d�@u���#�ٺ�+g��jU�o^�g@?�SD��o��.N�Hݶ�u��� -�-�m� '@k�,8/i���:� E���m�I���x�Y0 m���|}\ Bm umT�U�Ľ��6�� mT�-�Ѷ�n�f )A'8[D��H��!��� !mZl�`�n�l	�`���`f�-i|�z��$	 ڤ�m�   l�^�:��d`�U��H��jVz  �`�[p�J�[���j�ځchUB�^�����H$m&�����J���s�N�dQ4���v�`	 m�8D�A�mm9n�L�����:[@   -�t$ 	l� $����m��@[�����@R��/�U],rFf   -���k��0���p۶5�{6�kx$ 8�	 6��6��v�|I�mض��� m�lIm-��v���×D7H k����6��p   � kX�  C��m���t�  l6[��M�z���t� �  m�@6�||l l m�-�$͛U�ui9.x�}�z�V�m��  �m    ���-��  �    մP����UR�P�+��z��!���-�μ8m���m�6� ����H�   � m�4�N[�Q�Z����0�]���"Ke���Ե��o�C��M���඀  m�N� ��� ��ŵ�_[r�pH�8I�l	h pH2� ��l [m�lVK�l8� &F]�hݶH � [@��[��H   	��� �c��yv�{t�AUUF�;u9ˠ��7 �����i/��n�8�m���>�� �C_V�	N�l�� Id�`J����]T�QH5T��w�^�l�U\�h 5Mw�+m�m� ��[@[A��׫r���h��m&�k"M�m�h V��&���v���-�n�(�'V m� -� m��x[B�Fe�i@ 6�n��m�Ӏ6���ݶm�B��bCZݻlɴ�$&����]��M+�*�mUmU�TUۓ��GAt�.�Ԫp�� m*��v�$�N�R�l`
��8�Uv�ݻ`�U�e\�H�)��1�L�-N�˲,$n�:W��[
� mmm�6� &�L�6���ݕ���U��2Dۢ�jU�*2� YT��:*�н���(��G�W˷l��n�V5u���X( m�Ϧ�~ݶ�I�tYZ��,@�K��
�m�(�bt$�	�V�2u�n�[Tm�ˌrs;�`wU���elv;�n�����2j�nM�""������ ���b 'P1��O�s� <�*@T�(P^��\򉀈q>`>Pꢟ"<Oh>��]'W�0T1�a�pT�6��8�uQ������#��2?��'�A=�A��
�v��*#���H�H�E��a��*<_�8 �o��(�i�
� J
� �< ����bU�*„���A4�����@�*�����\b����QBAA�~5툏*����	�E|���@>jQ��+���`�"t�(>�EFD^z�tO�(q'@I$ Ax�}P��ޢ��]���@�mP
ʁ�|-:)��uU{�7�I�2 lހ�E�&�
'�Q�Wh�U*l����G��0j������?�P  �,X�ޞ�t�5~�  -�i[US��,e�9Ƹ��C�sf��Ƚ[e��V����ET��6�;�W��AFA�.���;-�]�]ـ�U��ڸY8�� \�k�b���Mn{`瘻���A�Z�Pe=�I�M�tH�UKs���9��2����ڗ��r�8�{���x�dY,ܾY'!�
��'���ѻP;����{vp<��z�睱l˶��:L]6xf��Ƶ���u�C��Ӽ=��3���*dz���.�d�p�����Ʒ�� ^��q����70#��˟l�9�T�u�c�F�F� �T��l壷cVG���C��d��,��T9�6�b��U�8R�X��m�t� ��5m�m�d�Ӭ��(���m�;�����M�غ��ɭ��&���B�7b�v�MƷl쑦m��eՉ{v��*�u���v��e�j��g[vXGB<�s\�:�塓֠Nހ�Z
�BU��˓��{(¤�+��p�#��q�`7�tmˮ��
���c\C���R'H�����<ۗ�OE�I��.Wj#��N���qK˧�y7%�gvꬕ�+�[*L��l�It8�����.�gu�#j28�F�ވI�-J��v̕�<
�n�tv��f���U�Ŏ�\�7�6��I�O�d��,�u���;r�Pk�G'\���X2BVܡ��-���nh/$�ҝ��c�]ե 㗲p��j2j�By䢑[t��A������v��3F*����k��c:x%���m7g�m�l(����n�n�.kd&͒��]r�q@��֣d�t�MU*��-Uq�F%���
�-<������+5���K-����ٗ�W+��m*��m�vu�W�\�{�g�9��Y�x3��)D�u�.T%ێ(��m^Vx�䞑p�O9��vح��ղ�H=�Z]�]�۳����z�=6��-�ҽk�l�k[���mq�v�i��MkYf��� 'DW?(R$R`G�| q� �Dx�_�oN� �G��so�n]�=dtem�&:v�6��7EQb6���zL�]��\�ܶ�z՞�vz��<�u(f5� �5niآ
-8��ny�+�B㎹|-�nEr�8i[\"n�Ь<���uˮ�c��&k<�)���u��n��;��n�ĦR�zy	 �9�$p�/[�{#���L�Ƴ̓;�6k[��ۯ�z^��e;��=�plB	�[e�WZԥ�MY���Ǟ���g�9�c��p�E �D7@���NL��K ��ײ� �'9��n	 �}{�����MD�,N�߯6��bX�'}o�(LV��T{���{��7�����m9���]D�K޿�T�Kı;�~��r%�bX��k�U�8���-��&��J�:�\��ND�,K���Sq,K�����ӑ,KĿ{^ʛ�bX�'�{�6��bX�'{o���Y!�Eі3��bX�'��6��bX�%���T�Kı>�}�iȖ%�騞�kdMı,K�Ӿ�	�	rk0�eћND�,K��{*n%�bX�{���Kı;�kdMı,K�{��r%�bX��/��^�Թ�!5�I\�Ɥ��ѹ냒\=)۵�ӳ��ѹ�D�;�PV�1��A�k�É�L�gw��br%�bX�ﵲ&�X�%�߽�m9ı,K��쩸�%�b^���%��\�Ys�"X�%���["n E(ER�H��
�6��xZ����K��m9ı,K�k�Sq,K���{�ӑ,KǏ���rj�e�I�w��oq���~��ͧ"X�%�~���7ı,O���m9ı,N��eMı,K��z������Y%�8�L�g8_��eM��D�K����ӑ,K����7ı,K���m9ı���'�Bi��@���w��oq�X�}�p�r%�bX�v�eMı,K����ND�,K��{*n%�b�����F���F�B�H��Q3h!B,�mDtg:�Nւ�90�q=v+�+v:��ۖk.�Xq>�bX�'}l���%�b_���iȖ%�b_��eMı,K��ND�,K�m��Xk	��te&�
��bX�%��{6��bX�%���T�Kı>����Kı>��ʛ��5SQ,K��߭�fB\�̓.�Y�ND�,K����7ı,O���m9�
���^�W��Oe�ʛ�bX�%�{��rq3��L�~�6�KD�KQ-���,K��ND�,K���Sq,KĿ}�fӑ,KĿ{^ʛ�bX�%��:R_���%�0�r%�bX���ʛ�bX�%��{6��bX�%���T�Kı>����Kı?"w=�Y.�eˬ�E�)��̓��u�suOY����m�^J��ڜ��'���[�w�{��7�������m�"X�%�~���7ı,O���m9ı,N��eMı,K��ߐ�v�ZJ��[s����&q3��fڛ����j%�����iȖ%�b{ߵ�&�X�%�~��ͧ"X�%��g�Bi�0����w��oq���~���m9ı,N���q,KĿ}�fӑ,KĿ{^ʛ�bX�'�rI��멱Е�*�/�8���.���q,KĿ}�fӑ,Kľ7ıU�� ]�'�O `�o�3��M�"X�q3�����Uj
D�T��É�LK����ND�,K���T�Kı>����Kı=��7ĳ�oq���~l6�1�U�)R" ��7T�q�v��m#�	��xP�,:Kjݮj�I5���r%�bX��ײ��X�%�����"X�%���l���%�b_���iȖ%�b^�Zצk3T���&����7ı,O���m9ı,Ov�eMı,K����ND�,K���T�Kı/N�Ғ���Y-��ӑ,K��o�T�Kı/�{ٴ�Kı/��eMı,K��ND�,K�ޚ��3%ɬ�f�j]aSq,KĿ}�fӑ,Kľ7ı,O���m9ı,Ov�eMı,K����.d���al���r%�bX��k�Sq,K�����,K����7ı,K���m9ı,N��]��B$Y�ѥ�,*a!��*dY�h!)#��B� E�Db��M��L
k�k�������Th];��ʕH�$a�q��%I�H���΍�j�+oU���sp����n�8������#J�<�xٮS�tN̻uv�8Ҧ�\P{&��i�G�9yv��Е�G\�v4��
�=� ৎ9�z1y��b��3<svk�0��Q��:�dW8x�@h�[�(���-���=�QO�bTH���a��w�y���űiet�׭����c��e�ێ�鸻'=c4t�^|2�6Dm�Z٬�e�շe�ʝ�bX�';���"X�%���l���%�b_���iȖ%�b_��eMı,K����z˙�YrMe�k�"X�%���l��o��"X����6��bX�%���*n%�bX�}�p�r%�bX�;}���PX�Q-O�&q3��O�ݻND�,K��{*n%�bX�}�p�r%�bX���ʛ�bX�%�{|:�D;�]����q3��L�}ٶ��X�%�����"X�%���l���%�b_���iȖ%�b^�Zץ��l.L�j]feMı,K��ND�,K���Sq,KĿ}�fӑ,KĿ{^ʛ�bX�'�S~�~hJ��ۊ��X��m렴�ι�<qv2�2�fև���;D'<ɗ�^WFŹ��%�b{��ʛ�bX�%��{6��bX�%���T�Kı>���_�&q3��OwH�-��v�Y.����%�b_���i�p���>Cgț=�Ȗ%��o*n%�bX����6��bX�'{}���X�%��N���2k5sX[.�6��bX�%�u쩸�%�b}���iȖ%�b{��*n%�bX����r%�b���nZG8�ꅶ�,8��ψ������Kı?{��D�Kı/�{ٴ�Kı/��eMı�7�����i�j��w�{��ı=�kdMı,K� �{��m>�bX�%��~ʛ�bX�'�{�6��bX�'u�{VK�%����Kte����X���:�u`œ[�Ձst�n��E[+-�EX[QŇ8���'��iȖ%�b_w^ʛ�bX�'�{�6��bX�'��l���%�b_w��a1��d�s5���Kı/��eM��GQ5��~��Kı?{��D�Kı/�{ٴ�Kı/�H��c�ڊIm|Xq3��L�����"X�%���["n%�ɨy8�yS�Ñ>�y�s6��bX�%��쩸�%�b^��5��:Ѭ�[s�"X�%���["n%�bX����r%�bX��ײ��X�%�����"X�%�{�MY�3&h���3SZ�&�X�%�~��ͧ"X�%�}�{*n%�bX�}�p�r%�bX���ʛ�bX�'>=�d�5�Y�XM�@
=k��=u����!�]��_�cXK(�	[�74@WLc��׻�����ou��~ʛ�bX�'�{�6��bX�'�}���X�%�~��ͧ"X�%��nZp���#�����g8������!��D�K���7ı,K����ND�,K���T�O�"{��7����������"�j�߭�ı,O޿�T�Kı/�{ٴ�Kı/��eMı,K��NE3��L��=�B�P0��Ӗ�Ň���D�w��m9ı,K����7ı,O���m9İ3f�VH��0��XT����Sq,Kļ�o��c��\�35��m9ı,K���Sq,K���{�ӑ,K��o�T�Kı>������w���w�7��ǵ�e<�����@���{NIg,��]oK�.m�ɸ�39B��sjɱL�&k3*n%�bX�}�p�r%�bX���ʛ�bX�'����ӑ,Kľ7ı,K߻f�B�ƚ�I5na��Kı=��7ȠGQ5Ľ��ٴ�Kı/�k�T�Kı>����Kı/}�[tf��5s2�Ժ¦�X�%�~��ͧ"X�%�}�{*n%�bX�}�p�r%�bX���ʛ�bX�'}=�kY�u��\�Ym�fӑ,Kľ7ı,O���m9ı,Ov�eMı,K����ND�,K��[�.�32ۚ��jffT�Kı>����Kİ�޿�T�Kı/{��m9ı,K���Sq,K��{��3u�f
�,��Y]��M؇S��O����p�d�N���t��sgF�9���;#�p;�#����\E�\
��Ƹ�p���WnSg#V/GX����m��@��C�gՓs���:U��x3́i���H� /=D��V��[��O=�9����D=���GQk�s��@�9$�Y��^��wd�9�g%޳Q���A�	�ߗ\K�ė�~��P:�\��u��m�6�9�j$�c�-�9��y�j���Eh�t
5�ܩ��vzdT�7d�5�@nȩ���Bұ0�V"Z��ݸ���슐\T�#$�(�e^v�/3��k��ݑRk��였=����0t��K-�{�� ��q`{�p?$��m�w̑	�i���U���@rd���v~ �͚��ŀ{��56�h���܃�[::�m��v.9�ݳ�gC�K� T�6�KBAʰ�ݸ�����ŀo}��i��W��쩱�p{��H�D"ā"V �$�DdH�@"�u�95߽�rM�� w�� ��ܬpE��aP�1�"�� �1 F� $���m��e�ڥ�`��X��� �{n����7��j-�����N�R ݓF� 7dT�����������~��=9����
�$���qF�xv�S�m��@nby(^HF�Q�׮,�l;���d� 7dT��"��& o��]���������,��l��iP���k��l�^8�	�K:x�w�Tz� {ٓE���	��D�"$R0H��"#� �#"B��$$��l;u�M��h%@�#X��v�#cej��j�%!HBkB��Z�� H"�BD�㸙"�w�h.�*Ya1aR����2�mP�� �#J�O�+���x���z��Sx��: ��C�"�(!�"g�: ��(�b�o��'=�f䟻����;���[+
���J`|�����}�\��Ł��}����G���㴲[3��b �\���o���d��ݸ�\\I�~�?�J������k����N�^A��{�\����	ƹ�_��}}!�7i�*������`�� {ٓ���������3$�<�3+��H������{��@nȩ{��{]��mM�Vۖ� =ﾸ�����~����'L�9�u�̣�s��=w�{�ʐk� U*�u�"'�s=�ٹ$���~�3T�&��f 7dT����였>��<Oz�-PW����A[xH����nơm �ziϛ��
�箴{�ۋ�1�יH	� �7d����� ����V9jn� ;�ۀ��{�� ����=�f�,�һQUe�1���'���� &ȩ nɈ�l�ۃuYdr�In����?{�L �wn ~�����5�mr��̮�e >o �7d��s�*F���ww�����N�ԁB�Au:�36�t	���U��$��H��<]iŉ�f�y�θ�7�����q�\�=�S���@�γ�q���>M�0�]<q[������NN�pVh$͗.";�����v��w�^c��;+�(�c���@��A2
u�W�/mL��M���[YĶT,�D8w71�-Y8!11�<�����d9��`��J��9��fc��9u���\�R�stfw������܎NƗ6�T�n�S���,�B�N�{�}p�� 7dT��^A Jnv��U�w2���� ��@nȩ�y�6��͛U���Z�m�;��X��였>nb z;����ʰ�����)6EHvL@���1`�ѷ�§-C��`{�p71�"�� �uy*�xWq1Y�r�ζڀG�wU%�N�%�2bH�vr6�<�2��\�GhH���� }���7dT��"��& 5����/+;�9*�����$�9ĸٽ�ŀ�ۀ�m��6nϤ��J�ev�KU��J�>�ɣS2Ha2I'ss6h�����j�V4�%��j��& �n*@8��6N�Q��u�̢�31 8� qR� ۻp�O��~�,��;b D�G�tgmq�.��tu]<�v]s���Ɛ�V�2�RKo�7w�X�ۋ 7�� =�ۀ}�'��q��ʦ7,E�e|��6L@9��T�$q��§-M��X�ݸ��t8,���Q�@Ts=�sf�~�n,����;BJ:�n[��b7 $qR �& #�۝��v�]��T�ۀo�����9������}���m�;���T��EDu�]<��v� �ϵř����:!&囥�L��#J�v��$kd�`��X�ݸ���}�ŀoc��KF�Y,��2��1 8� #qR� �ݎ��9al� =�ۀo���o� own�{�ʋk	j}�@F��*@d��[\�̉m����D�T�J"�*�=��X6L@9��T�>��E�Qy��{/nɉ��ln�[hݛ��Ş,a�3�Ls�p,dm�eu�婵� 7�� s�� ㊐�vw�������w}�@9��T�q�Hl�:�fͱ��Yd��IT-� �{q qR �& ��܀^ee�E��Z�o� own {}��'��ߖ��{>�J�A$�Y-X�& �n*@8�ܮs�Ug;�� �<�ҕ^�{B�p���c��
��n3ۇHf녗˳tfݮK�1�Z��$�lunq��f���p�@�h�[��K3��y�ʭu;��ƌGc�n�c<�D?���w�i��0�:㶝�9T�\��'>^�9K۴k�u+�I�:)�Zo(�+�r���.҈{Ok�˩�f�֬��!㥷G>��$���׷Z��v�zѭ��p�:�6�<ݨød#zzk.�9�:l�9�GVX��Em��:UQ"n*��o@7�}p�T�q�Hl����ܣ:e;Y�U�s�� ㊐�1 8��ޞdc�S	(�\� ��q`�1 8� #qR q���S�yww)�CĪw�ݚ �͚.�y{� �f�,�БWX�-�o���� ㊐�1 ���x�yy-�Y��L�׵���	��z�Ѳso5<g�ǖUK���Ӫ�%n�J�m��ۋ q�H�& ��܀gr��w��3-��7$����\�0US�!4�D���@�	62d�L�k�������w��]��c���9+�KV ~�ۀ�b=U��]�<�=<� ��v�VWo�_k.���@9��T�q�H������j,*!�������@{�{���{�1 �[��;��f]qn��;�N&P��Sv���x)��\<��F��E)�jJ"Հ}����{�@������v� f�;��m�Sq�V w��?���q�����=�ŀ{��X�n�+�бWS��j �� 7dT���o+�g�� ߽���E��+vU-����}�`{~ŀ�������\�?�%�K%v�2빙H	�*@�b �� 7f��<��Aʉj���[b �I�6��Z��Gg����n^�����w��5���}��e| ߽��� 7dT�}���5��IJ��!�XK-����c~�sʐ였w$��ΙFv�2�/31�"��#�*�����;��p{���^5-�j��O}��-�v(켚d��P�e�֙�y'L�[���b�·x[11�2��}�R ݓ�9����H	�*@~�7rJ[�c*�'H��6�+A��� ꠆�v����}��J����>X��=<�����zh{2���p�_8{� ��H����[�r�Yn���ϒN�'J �ݚ �דZ�;����$M
Y"-�[j�;����?���K�߿����� ���69*J�PjL���f�=y�@{ٔ�;�2�߿�{��%*�8���,� ?w�4.Ifwyx͞(�̚��4��6BH@�!���M$h!��)���!�L*@���e4B�# SI
�bc��]2�bA�#�#Hj.�@�$�
1�A���BЛ"�T4����
�h����iф��#�� #
i����3
��"�$sI� ��M$+��M2�0q� 4��H��Q�خ�B]��:��^���SR��tB!vVjVjP�%e��B $H"F$HE"AXP� b��T��� 1GA�`�1b����K4Lp��0�HB!��atiKČXO� ��Gm�$!$� #�	 E"0#B1I��9;���&ۥ���d$� KE��S=�]}ϟ����!�8X0��j)B	�K�0�*b�BI�����:@�Ck�#��шY ���*��D��`ۮt����H  l$����.��&λ������L×�� U�����]�Z�-����+�7CU��P�:g5�M̊Үp�� ��I�Lh�����]� ��lc��W3[���"/^��F)�Q�x"�*�m$4;�2V6��«�V��9S+�Ci�NՄ��X�m��V��]�Ҷl��*�u��9�N�n]������Z8�{*���8�ez"3���ݲϛh\��w<���vB�;�����b��{C��sLmp�rg��˳�e6��KU��[g;����2���m��@-���F3Ik���f.�yi�06��!1֣��Z���+���
�ԁukv2�0��	��&�ę�����S��ܨJR$;B∄�f�lޮ_=qۓ8��\H)����=/�kU��.�qjpb��{Lng�m+8ùr�YQ/-���&ŋW��n�q��n)U��C��򛷓m�t�d�K*���˰��v1 픫�	�q�+� �ћl�8v��&�6�v��=t<p�푪�۪���vf��V���8��]�I�]���� =�:e���U����n�������bl�-�g#	�v��i�h�$�`8��ȑ��%qJ�25]��
��-�#�m�h�
EV�M��ƎGX�ld���'m7n-�qЖ�!⊫�k¶�/0*`����*�]�5!��v��z^�j�eƶ�Z�<Ҝ�a��U�̉C۵fCr]Z�(p#����6qj�UWm]Rd���ԅ0�f@�5Ӳ��:H��b�b9�:�Bz��e�����z����C����>�Xj6���S*P��C+U%�Ò�ѱl˜K#�^N��@���Y��I�����X��pD�n	��[q�<9D��yuGպ�� 9=�mAEB���B�[r���n�A��s땤2�x�;nm�2�gݴ�K��mQm<ۨ�!�N��ǎ��%�w�Q��U��/�^�����۟�P��@
��U�?�����v�������-h-��k��h��^��=^d���wq�-]r��
�պ�t۲U=����\�9y����Ժ�t0��.7=�s�6y�uڱ�P���Wz8�g)ch,)9"�J}�blUEq�\QP��Gnۚ��њ�8�srt�m�^^v�@ �"-m�cdԆ��X��u�Q�;���Gf����n�sr��[vM����$
�G�_�I��W��;�[B{9�N�{������4㛮2g؜§S��ĦL�B��)�\���z���p�{2u3|�z�f�Y��+�x1ڰ���>�I�����}�\��şq$�o���YrYP����vh켚?�&���@{��k����C�u:Il���;�=���H��{�o�������:�vU-�;��X˝����<��� ?w�p۵4��N1�а�r��j��:}�Nj�uh�VrX��;GXMa���̎�B�䈶�m���ߌ��� ?w�~����b�>^���IP�8놳Y7$���kx��yEt�G_h4� �R�y���vz��׻�TQ��V)e��o� �wq`�� w�� 7��ZVTH����n��T����& �+��ߟ���K;e���3���Hא@�b �f���ŀ{��56䵷[D���Z�v�,�n�y#���f�,3[�t�ī�
�%��ܖ���0�ݸ��� �wq|��n�� ���I,�T2ҧc���&Ɉ� 7^A nɋ��W=�؟ѱ��v�[�{�}� �qR%:��Ky1 Ms�Y���ے"�ն���߿, ������p:�wqP7��lrT1:�Nڰ�}���@M�R슐�n�v��2ˇU��+��zSl݂��sݸM���X�\iKR�V��\�a�t��m���~H� ȩ��u 8�Va�e+++vۀw���ww��ـ�_7Wй���3���H�*@u�v`w�p�w n�I$�]m�j�7*��?O}��}�\�wq`,��AdH�@��D3��|nI���k�VZT�rۀ�m�?ww) ��Hu�@����e�w�K�fFRv:�ܕ��yt&�$[�g�x������72'�i��v�W-����X��� ;�m���߮���VIQcr@���fU��p��M���4��4���>l�G���bvFKi���똀�fA�̂���3++q*Բ� �}� �ݺ`��L����|���ZVT)������p�7׵��y�@���&L�@�[�`iUUIB�Vܩ�T�9-�E 7nz�1��+�ò���sv�H�^�\1�a�l�@،���Ţ���q��Nwg#��Uq�jvv��9���-���}���Go� }U`�&��c����.�
�#�)�=���9�=���gS�,k��DOVh��3��q#@l�����[[NY�l�̡�s6�㨷-���[&��_� �P2I��&�l]���Z���ٕ�fUN\v�q]pO<ƭ�(��
+�y��2��p������� _�&�=��v�fK���<PwDC�q/.�2��y��/ٓ\̙�=����o���qg�f�����ʫ-2�;}��������� �� ��=�M�[�v��nϿn|`�� {�ہ�o�o� ���ܪX<D̼KĔ��˔noO�/���}t�=��*���G# �f�7A�nc�[������r�t�1$��ٿ��?e�E���-_�7���������0�oذ'����!�RYn }��P�6�A��Ҁ�ͥ@�ɮdˢO�ОT���!L�<���<Pl�#�ds؀��_k/�s��e�<IA����(/6h޼��h�߸�툇x�^]�"eC��% _�b �sG�@=qRIWW���y���k;9�˵�C��O�{r�s��,u���FH:i�BM���m��b3�dX��$��zh��
�yK[�{͊�	����`��n�}tϓf�~ŀk��0��n}�6y���nU,q�-�sʐ�Σ�k��7�؀ng�ݞ�G%Cc�4KV����~�����߿,��gŪ�����_s���� >� �z� �����5�����B��K+V�R]�s�Il;l��d�G;=�١yxn*����7\\9���b���*@\�}`o�� }��P�ք9L�v�&ᗛ4w�4�s�~2\� ;�"�Uu�%�1�L �~����n.&��ߌ���`�com-��k�m�p5����f����@}�(%%�&T�ˏ��J�3v`ٱ=�c�� �%r�7�@}� ���u n��ܪ�j.�*���U����,��*8� ��ӧ��Nuk��ŵm��U��p�Mѫ7"��3/�|�g��s�u�@}A��I���|,u�Ki�y��0������~��3��&�'�����/131@y�@}�8Q�̙�ۓ�����5>�\UXT)�C������ �@\�_murPr��v�;�\T�w�u }���� |U$�8��6�zG5���܌�h�ӹ-;maݯl���iy; �l[]n�9�8�L���6�c�7/%�6����N;�B���kn��H����ܿh��᧓ͼ������f����e��;����Kf�
��#�:{m�rZ�]mv���`5����$4���rU�ݭkS*��ͣ��@j׃���Ɨ��7cq�$�M!�P�w������y~����?�g�������ѽ�ѻ1�&�b�]9i�M��U�F�۩T+�k����� �� &��슐L�6�)S�V�0����O�/�7�}� ��~�}��1�[�����bk� >� ���u =s{��%V��mv�L���k�`����Lݞ�S��|,e��� 	�b z� &��슐I$����a%L��JW(�q��B�C�sq�M]�n�]�+C!���c��[�m]t��˼����{^A �EHo��O|lU[X)�ۀo}��VW+�]��EHI1 ls}�U��A˳���� �EHk��69p� n�H��]nIj�� Ms�15�H�*@93���[e*��F;n w}� ��q`��L ��n�����]�V�%�:K�t�X:�Wp�c��'�1�ɵ�g0��3k�,�\A�[����[�o}���� o}���~`o��y���$��9"-��m >� �&��똀���6g�9(7���m� }�����a����F2H@��
*�H�A1#@�!!� ĂFDH��$a{96}H3SC��{Jl(�� �H!F)<�!T�D���@�AaP�2��Κr7CD!���u��U�h�2$��`mJ(dP$a5��$#$dM�H��
+D
�
���jd��| �C>M=Pڎ!���V(EP4p S�a�Uw��ʃ�D؊��}߽͛�{��M�>/��������r���� ��@MqR슐��p'�6P��R+P�m�7��H�*@\���@;��D��6�3r���pQNf��u�,����)@�1�{5��/-�EZN�nYj����� 9�@�� 	{۹�fIj,� 7�ۀ�m�7��X��� ��I��k��ѷm�wۈ	�*G��W.��< 9�@8�9"��-n����n,����m��N.I��� ���Q�
����y���<� �� �bk� %����s���z��6,9�+����V�uȚ��r���2ݕ��=��l̤5�@�א@=�Ri�f���H���[n w}� ���~�]0{���n�;X)�C��א@=�R �� �b �������0r�'���� >��p����L ��l�DHKUq�r��1�~�π�� �EH&
`H���1 *�M�J
�ݝ�O[�I5l2�f���ERS�:3r�*��n��F�Ѹ��B�@\�쮬D�m�:�C�N,���OF�n���aSk�Mq��0�,��VL������(�ukr�Ϩ먔�̼�\V�E"�aP�@�s�ka.$Wv�%m�`��ѳx�R���VtVG	��mh����C \Vsx�ʥ���tޱ���X�ӳ�`3O����y,I(~FO�J[!S�$LEqѭs靎2� x#�.��E�'���GP-�0T�h��0�����?bk� ȩ M{p�l�VYkuWd� ���}A M��1��+:w;���o���ܾ���<� �& �b7t�?y�j$UC#��L ��� z� #y��{n^f�����.��������A�y7v��l�Z*�أj�����+*ඛx����tv��v���&{�������%t�e^f #y���1 =s0w��?i�nY)�~�]1���%Ba2CC�������zh����4v��	j�7*���w�p����� �}�,��9&�e��U�nہ��7~���� ��U@=���}���H���[��%���L슐�1 ls��ʮ�Յ�n�,k��A���W��[���U��x��&r�5l�Ӗ ��#����-�S��ŀ�ɠe����o'J�#6%
P�}2�̤5�@�א@=���<��m����ܶ� ��ےO}��ܻ���DV	�`�r��W-&�T���*\˾�egk0�15�\T�&����`�Sh~Ӏ9\LnS �}��u�@G15�eTe8������b7e��sƞ��lm̞�<#��TcX�,�္�ĶGe�t"���o���&�>�ɠ3�8wzsz���33-��J�ݷ ?o���]0wۋ���{~�w���UX��]��k��\T��g�� �� >�%ga�%ɇO<�&ePrd�˙����* �� �/&��2K̙�a�)PXM�A�P�&�	j����>�����ۿb�=��X�?F�D壖&\��u�c�������v���/,P��@�x�������I[nYo�}�\n�~̥�8{�@c>�I3#�aL�<��w��YrL� ��@��RI�����U�C��d�YtYn`���T�&Ɉc����HG}�%u�BZ�*��.s����� =���w��5��>^�ʀݍxٙ���w�fw�����@F�� 	��nI��gʦ� ���$��kF�s%:8�]�uֳa#e�OD�^W�Wduv�Y�c�����=�6�L������t8g���<�+p��@Ղ�c��XY�[�8�nηi��s= ��Ю�1�a�m�gCţd�ō�Qxe;3eH�[s��Ӭ\s��*��ֶӬ燓9z#�M���# ��`��U����������j���X�*��n{�޻����ߨ��Օ�R�kڹܾ�u���#И��h� ����М�N���{���/]-�Q�-����ŀ{���{�p�����]e�5!T-� �wqW�$�e�̢��h;zh��U�ɳ��C jж� ��}pc����H�*@;�d̺���{[nYn��M����n�� �wq`|�o�}��7�,U�b��p���� 	�b �� >�d�+���4�"�Y���k���۵��������Lt�)%��q���:�@IH�ݫ���T�̚ �^O3s7�;w�P.����Z$%��r� ����Ē]��fIb�	�ɠ>��T�2�k;���m��۔��Kn {����n,?��}�, ��}p�l5�EU��Q�. �������ʐ�1 ls�5���ƚ�U*�=��X�{��}�\}�ŀ~���dUH+	A�x�Y[���9���nD�[�K��$�*��#3-C���5h[W���� ێu��dT�w���8gK�����gsqΠ#qR슐�3 ��KUmX�;f����=��TrM�L�!$2VͿ|T����lP���ߖ�	)��`��, ��M��Ƞ��Ϲ��[���*]L��*�3ٓ@u����nfҠ/۸�ujs_��Z��)N9Ճ-�|����t�m`�z�G���o��C�Q1��e���34	����T�{"�;�p�l5�J�#�:��Y�o������T�<��@m�:�>r��V4ԥp����ŀ�ۇ����L�߱`�&�qPm	Ҳڰ>�;���o{�@e�R�d�3��̭�Iq~�+��� ����NW�����?�"��I��v�yx��T�̚�[~��~t�Tۥ�{my�⎖	���]���U������m4�9Y�{JR�7Q�Π#qRu�Hl����N�����-R&7j�;�n,�����f����Pw���;����y�.��&Q0DJ��٠>fE��s6�~߱`ݲM�WmnJ�v��%�$��݊o6��^R��I;������IQdr�T��0��������fElҥbW�@���R,X$�"F$�A��RB@`F� I1"1 "�`��#�B$H0�F$��I F#�H��:ѧI��i0�MH[$d��\F��FB1+��H�� �<0��R,'�Ҡ���I,",�(1E�hD�� m��y�L�Ru�ub�`Ab#BDZ b����B��D �$bFH�H� 6�P�*���B�Gw{��N�_{���~� 	 h[m�:r��$z�,��l��%EFő:��v0����P�T�N�m�R�V0I��#+�էU�*�ȴ��z �v�fAp��|9M� õۓ���&�ntɆva�J9�N!�습U�J��Nð��e����u9�]��N�ݤ��;����ɸ�ae5�i�-���فN��
`�ܰ����ٰ�ه[{<l�y�W/K�6v/vq��1v,�GKk�fWM�H��Zs#8㮀�C.��%\)�1X=q���z�xu��>Kn8�$ڸڝl������ˢj��2r-�MZ���q�X����Z�ƗaC�P�v���j;���J�l�#�`�$�n��۸8�Y�u�ҘSkl2�	�����q̬�.�)�����0O��6�ֲ`}=���Ev�$��ە����u�ԴȽ�H:4�����r�����h`8A�ڬ�0$b�4i�e��T]�HM�`l�Ǯ�8f�;�A��{	�-.���3M�n˻/k%�͊W�7��5/n�Jf����8����e�c�Z�ϯ\��Fy�vUY5���U�=������1\Y�����j��ڎ��;@��Q�ǎ*q�uHI]A���'6��)y"LM���D�v��l�Nԕ(�!m��H]�۶����6�e�ܐ�b����-�mx4i96z����1x6���(���L`zn^�A��%�H�t�ɫ������VV${u�/�	v��Þ�M�g:�[�l�:����l��h�uِ6��gB("�j5�2t�t �[:-U������.���̀��+T��J�]<��I�k�`J�fdu�e$	����̮�lŮК��R�0���ti,��ke�v�nt�A������8��$�:�e�K��n�P2[���I�ַ=p��]l�\Q�\j
��g��,��lͻC=�U;4豧IŎ\d�́Ƚt�Z��m��wV7����f��l�G����wwwn0��#�� 'x��Tx��l訟.��譜��ߡy��(UkNjg�#��OZ���[��»�0�5,���:��#ܐK�d���:�mn;M����2�i���q�:�H�T�V�"��+���d9	�.2&�x'[�7��Xx�M5R���b9d���uN���A���9�(�Ic�D,\���R�����PT���޼��>ܽ3�so��=
�G�y����z�޽�T��q�9�bNՠ*�&��:y���Tu��n�v9�ZPo�w��c�#����-n���߾ŀ�m�:��̙|ᷛJ��Dn̎�"!НD�fR �� 6�N�&���"����l���_	����~��MqRvEHk��udr򳹅�ީ�D���g���P{��=y4��=�� �����KUbnՀw� 	�bod�k�����S��z!Ϩ�����5a$Rє�P��X�1��XGN�;i�qŴ\v닿�Z~J�ʍm9�V�~������	�*@nȩ�Y#�-rZZ6�_wfb_��%���Tk��k�ٹ'��lܐ�����y%E��R�,�7�ܤ슑�<��@;~�P[��}���D�t����ŀ�ۀu�v`�n,�DݴnQF�MJ��`�1��=߀��T��H� Gc�fXܴj�l�U��=Sî�FƑV\t���[����N��:Yz�Ћ� S_m��w�@e�R�>��\�ɓ|�m����ߜVJ��V�,� �{qg�q6w�T�<��@;nu |iat�Qy��s�9�{f��{ٹ��  ��̚Lԓ$�U��E�yJ�2�!c̨u!)�%Pk2fe���@�� �{q`�w��$�am�KKK��b m�@{�{����� M���ܠ�v�-���EYyX���C�Y�'Ggk�d��v�� �/.����1�v��U���b7 >�*@d� ۘ����M�ʬm��mX��ŀ�b m�@F���ʻ�����+	�J��T��4��E˔Gn�,���ذ'�E��W�J�m� �Ƞ2�)Pfe*
fd�bd��7	2vI6�d�s4��]4��y�LD�v���u��I 	�b�{0�q.l��'*i�I#��D���n�i��l��½�&Ywn���ݚwﻹ���zUDĒ�w�^��� g�&���ɀo���}�{Q!-
��`{2k��7%k��Q�g~��T�v���"�krGm�ѷ-�<����J�fw��Ҡ�٠/.r\u(���镙��:�����Hk�������`��|�Ҷ�v�Kj�?o�) Ms�Π&��|��T�s�N? ?J�q&t��:k�kvEukM談��lq�;�9\�<�������H1UV�F�Wx�(���D���g[�g\u<��@4����&.��5̦Ʈ��6�^.unkg�7�8Gi)n(�6�S��M���51���ٍ��'9mg";t��V	���L$��S�Wgq�t��E�=��[]!>wW2���e ��\�Ce�Q�u'�/K�ɬpC��xуu�@%sb��sէ:�,ue��[hݢ#BjUl��o�\ �^M����%�̛��ԨO���g,RQ�e���n$�M�{~ŀ{siPz�k�&I��{�x�"S�aL�^f <� >�*G���$� =s(�Ã�h�P�w�!���?�y�	�{�1�����s(�;ӹ!)�%P{2hI&d�y�������ŀ~�n�*��B��--ok�u�A�ݝ��6oY3��o�!���P.c
�X�)�x�w���2�f�˼�@}���3/�d̒���4�wL)S3.J���b7&��s���d�R �� ��\�&d�(��;�u.J�wP�0�L� �~T�&Ɉ똀��H�K���B42:��`}�qs�o�}�����G ^ۗ�������:��� �^M���͹���nm* �����Z��أu��S���ѳso<6|���v�CJ�y)�Fn��[���f ^f #qR��6L�UW9����p��٬�B,�LnՀ}�����ovh/6h��U��rd�4@wlD����:w�T��4w��77�U��*qQo~�=�rN��ŀwv��5���ѷ-���s�N�y�@nfҠ>��Tﷻ4ln�D�IYUvKp����9�w��������������Q���ʶ��&�<<�	ۖ�h��<��.[pY�5vz�פ%Q�ʬr'mt����q`�vh�y:�&K���TZ6vdw�!7Vڰ{�s�$��Ü\�6�� �ͥ@}���Y�e��&Q���y�r���U�e���\}�ŀ~��X�ݸ�w�%Q�2�h��|�L��f��n�* �fM/32faRIs��g����k�=�KT#�`I =�W+��?{> �{��&��ͦ�qv���<���&�J�݇k��dٴ�U��:]�^ Uq[F{5���) M�nb7z������}�`������]��n[����w���2� g�&�332�d�$���"!L1.J�&&h��Tי� 7�� ;�m��=�5YU�D헒fU�L�$��ߕ m�� ]�M�Iq?�~��yY�UU����@�ɠ5&fnfI3(�ޟ۽J��3)P3%,�˒I���w���p�Il\�����@���8ga������n�n�u�n2����wp�oF.^7A�5Һ��5E�9�j���� y��'N�.���Ճ�Lt�'GX�-p ��v3::=uɱ˲l�N�Cp�gh���au$�����ɞ�i��^Q�Y`]�.�������ب;9�P�WU��[u��]���dU8�UP㩉��!�o=������~���ۛ�m�iw72�����'+үv�{n+�鵩����(���l)������w���2�$̙|�o���&{_Ҧ�b�Ze��ۋ92d�{wiP������&d���l���v��ݫ ��}� 7�� =�m�7��X��q=�YZ7r��1 6� #qRs�ʽ��� =���U[��KFܷ =�m�7����9�{f��{��A���ĸ���s����vU���#� �]n\+n��=/n	���L�G�շ7=:�w{�������kYfr�3b�A�A�A�A������A����߿p؃� � � � ����6 �6667���؃� � � � ߽=��2�3WZ.f\��lA�lll~����<��@O�b�*�A �>
���TyA���?f�A�������y���yO�A:���`���z���M�W��b �`�`�`�����y�{�lA�lP���y�~��b �`�`�`��]��u�X�D�Z�L��؃� � � � �{߳b �`�`�`�����b �`�`�`���߸lA�ll?������f�A���������-��4fI&k3b �`�`�`�����b �`�`�b���^�|lA�6667���ٱ�A�A�A�A���f�A��8�&�I_�(Q1.�.�Dʒx��v�<����:���y�3۔ͳ��ͷ^�^�{�~��5����55s�?A�������6 �6667�~͈<�������6 �666?���6 �6667������2�I��)na��A�A�A�A����lA�EK�{�lA�lll{߸lA�lll~����<����~ަ�j�r�̙�͈۬<�������6 �666?���6 �6 �v��"���$��ͤ�w;��w+aIeY�s�����$�i?dIIЌ�FB"� "A�� �R�A�=���&���^iC�� ��Ҍ&�
�A�D��E���5����CL"�
��+(�Դ����a�t����:�h�BqU_���� �!�EH���� �����y���؃� � � � �߽�6 �66q��s~�}a$V�(U]r�\K���ll_�X�������y�p؃� � � � ����6 �6667���؃� � � � ߽=���3WZ.f\��lA�lll~����<������]{��6 �����؃� � � � ���p؃� � � � ��~��h�Z���mpf�m%�8�%�#�^7l�nL�Ttg�q[g.5�9u[�2G9&�,���w���;�6667�~͈<�������6 �666?���6�����߿~��A�A�A�A������:�Y�d�fflA�lllo��ٱ�A�A�A�A��~��A�A�A�A����6 �6667�~͈<�-����S����fh��%�f�A��������A����߿p؃� ثl��߳rCw~� �uzDI��u@v��~���O���ܒw��nO����4(����z�wЉ���i�V Msnbk��I ?s�Uʿ|/�����X���J�E(B)%$��Y..��gTO&rt�,f�c?�k���uLV.���?~���� >�*@\�ٻa$V�+*��n����?n�, ��n {�۟���wM�����L�̼ʠ6�iPz�h���٠6�iP�2c*T����&ePs337.�� zObk��~�_��� ���xg�9��f&h.�hL�-�ߗ�m�Ҡ���ɓ;!$��8.�ԑQ+,��kDF:W��4�1�:���P�ۜi�/e�ۮ�4랧uN�;[`��%wI��g�ZO9NLn6�ҭ�Rx{�R��x�����=�"��U���ݡ�Znx^�����"�)4�v��z+�������ƀ�cck�����`�:�)�[kg���x��m9g��F��]���ѵ=�p9{{��������e�r�����xኸ#��̓#q�j�M�{f�s��R��;�����u�� ����ŀowq`���0>����ȉ>�+���`dT�&��715�K�\��Uv�`��.K�2�̪ �ޚ ���?�|�������ذl���U��d����3A�3;�f���J��fR����v�H�-�T겹n��Ҡ9%�̒����f��]���?���N'�l		
Ś���9���6�t��hu�v:ش6iM]���(�@M�R �� ��� 7h�mm�H�5%��`��s�\�8��}0T��QX�qU_�+�I�}�����X��ŀu�퓎&Ԋ���� ۘ���{�\�U���T�<�� ��������� r��?��~X�v� g�&��32g|�٠�Y
�M�*`�X��ŀ�m�{�p�������Mzvx����8e6 ��au[tv8#C�\�5�B�K
�nZ7j������ۋ�%�$�0��}� ߾����]v��﹈�15�H����1{�I.&��}�����T겹n���H	�*F��\��w�y1 F� �� ZG��v���.$����� 6�f�2�&��I�}�ߕv����R�4�[V o}� =�m�7��X��ŀ���V)��IYSJ\�f��[xg.�����s�ף�̚�Y��������&W8�mH�e��7w�o}��ۻ� 7�ۀo}��Abv�9�����s���پ�� 9�@���̙���d(Q!;�ħ�T�|� Ms���UU�$� <� 	����*��h4ݫ 7�ۀ�����ٹ<�r8 �⪾U^q$�}/���m��봴m�p[���U��y�}_��T�&��������IQN^�5q���1P��X��ٻvŝ{NO\��j��<�Nf��qt鯀�^R�>��T�̞L̙��������_}�������]� ���X6L@��n*S��*���J=��E �*����{�@�{�X�}���t~�M�(ղ� ���@e�R�>��T���/v(g���C�b��� �{q`�w��� =�m�3�f��z=�b�LNpk��!�D�<�5��mc�U�ŵvۄ�JF�q�ۮ����]P�6���&В��Oc��	�i��ے�����f���qշ���jՙ��Zʮ�6�n^MD^:I���۳h�oEg�3:PMzIK�M٦��i�`]�����$��2v���w�㍣�Bh��kay<����L/{[ݘ�;];^9��e՝�:��+�C5ːt��U�e[�<�z{bR�����=<���v(���+@o�T���u 6� &�� o|���*��h4ݫ 7�ۀ����n,���Ϲě7���[[��]��n[����7��X$����}� >��plݪJ�%�J�VW-����s&J;7����T�/"�.�&�?.�Nж8�k�`�w׷�@w�@_�)P��v���B�M���=jr/a�<k�۩:+�Hݶh]�N���}%T����TZ�T�X���m]_�~� m�@=�R�"�՚>�.jj�kY-����'{�f�O�P�fmL�5|m{�T��*ϗ�@bs�{*Ab���-�=��X��Ň�8ߟ���������E&�C����U�f\�&h���1�z(��h?$���, �x��YU��A��X�/"��I���fh�ޟ��J��3)`�܅R��X9"���7m�=�J�ɌY٭۲l��:�~���Ip�pR-a��2����;��؀{"��EH���=�v�+���*uY\� �wqg�2I���Ҡ-�6(��h��.���[]�Հowq`{�{�����M�E��O�;������:��#%�Jy��	�fU+}��P�� ȩ6EH�4�)Fڒ��ـ�m�>I%��������Ԩ>^E댇,RD��-�f;]u��Ӽ���N+�;m�N�+<`x�q��u5Ku��YSC����,=�J����k3$���l����
#�^e�X^e &ȩ�� ��@{����s�q&������Ucr�ls*���ؠ�ɣ�ffw�ݥ@m���=�f�h�u�mu�%�����̥@g�)P|ɗ���2mL�LN����~���%�J�VW-�=��X�w׾ـ�m�?vx�&�n0�U�eV���2�:��.�ӴF��k�-CK���dJZ�YdqY]�U�owq`{� ˼�L�8e�Ҡ.Ѳ��<ȉqW�`�/O����߮����7����6y3��PjJ6[f }�؀�ȩ6EH��P�n��(&ħC��&d��ߕ��J��߶`$�ۿ\ ]�lQI��;]M�@M�Rm����{"����Ȏ�.� ��D0
�1���JU��2Ť��0J�H$T# $c��Y�{��%;��w��7d��CV�ńHlD��4�,��>H��#ME����}�|j�E�0#��aD�w�'eCJ� ���������w��|p8 H [B�UHe{��7����6�p�}s<�:���N�`rI-��tUUϑ&U+Yu�d]j�cBȆJI9� ��Ԙ������1c6�ײ:�D���۶3�)
�{n�,��WdU��N
�۶��Y�pL��k���dF�n��c��i�u���.gq��[Lp������g���!pXW�se;����E��ٻ�#O$�v�u&�9n.�ɝ�<st�=��S�ps*�瞶KpŮ�Z��l҇3�[Y�E�y�=��Àǃ��լ6�Q�JF�s���e����l9�kbh���c���.ChRn���,l<����k9d{kmg���aMV�U�sH;n�Y�h�N*s�ا�}DK�RY-z�_H���:��w:5�\�Q���ѽdS�p�']5siWb����m��g�]�i��55�m�(S��4=u��0���@�j �W< �!0U�b�RUn���T^�Sn��Zbk�n��=�����1s�r�p�$a��,0�h䳴3�u�N��R���	�t���T&����;������geZ����[U�w;4�ɴq��]�(I��e�MUS�.��W'T�S���F�2�����s3�U��Z��ձ����5f\�۩*Y���ډ�fl�c"3�k�z�4�3Y{vxe�R�n¯m�iG[];[Xӎ{sG"�Ց5�]Ժ�(�[3�]r������i�2� ���-K�e��϶�f�q�nN�nV��eS���j���a��ѥ�nuV]�u�������z��,Q�=V���a��cvªƦ�]�JK]*Ľ��kq�NE�˓J���q�-��Q&C6{[g���`إz��Ige\N�A��-��yP9U��EU���/Ѳ�:X�rV�,c���Y*ڭ�i�l��=QTA���8GnT^g��۪�
��c�1�Ԣd7I���ѨqѮ]�*ǂ�3�1�cX�T��q+�Y,���D�sj�N/��EN :G7QN�l[��GA� ?�ݹ�vy��S�kt�l9z̜`�v*�;p�����ሲ�)�ZMέ�+�7`�&��5��#۵��9:�X�쨏6&��!Y2,���W�H������6u>�d�t�s\��i�.�ד[�d�f,1��F]6� +n$�h�t�,�N3�0;;M��Z�ݼ�Ep���<u��9�^���{ �*�Dp�ɸ����{Ͻ�>~�n��z	�\��3�6��n{ztN�����\rއ���`�8TH�t�]�������dP]����\����Ԩ���r�J���K0}���� ����:��3�6}�ߪn�Il��U������T��"��s�71 ��������X�����?�b�>�ɠ�nI%{�T�#6	O"�'+-�`{�������ŀ~����G�8��[vah�t<p�c*�Z�ܭ�{��s�ޝ1bMl4�wv�;}��m�(�m� ��\��ŀ~���&L��}͊S���(yA0�%:��b슓\�+���W9�I�on ~����l|�(��B��2�'� 	�b z� &�� I�ɥeV9-DC�`��p���{�Ł��~��� ߧ��-$�;%�]��1 6� &����R �� ?�\I�������a�[��q�D���m�ֹp��ɨ0.[(��qٸ����}}ج�G*uY\�����b�?n�, ����_����>{��7,vG�ܾ� >�*@d� ۘ���K�.�y��C�r�[V }ﾸ�9�\ʪ�2��\�Ԥϕ �Rj��=���%�[�����p�~ŀ}���5��;;�������y�Ʌ1*�� #qR�"�6L@���7j��%���媒��P��ͫ��v���'U=��ӊ�H���|)1E�!RՅ�W�o��Hl��s�� o�4���%��v� ����l7w�}��,����=�a���cn[www���1��ꪪ�*�}�*@{~���kR��r�U��p느I 	�b�ʯ���q󔕥.�wk�X�,�++�ʰ����	�b ���	�*@M�۬�����]��t��}C�뗍�F���U�d���p��,����]�r�7,%�`��p똀����H�FN��{v�$u334��Mjd�;�y��fm* ��n}�.q$��f���:��eM&h��T�yJ�fd�w6�f�2�n /���v��;Vˉ$�~��P�l���h5�>�oʀ7r��dV9-DC�`�v�.=����߱`�w ��Iqw��n֡ ��`�"�m�͌����"`���]t�Ŭ��iut���K��u��1;�Aб�3�˕�W�eEM��v.��ޖ�6�����Ͳ<pve{d�]v�����ۮۃ�6�jK�g����ҠfH�Q\U�n��Ny�`��l��g�l�B�r��e� /n˻s0��9l�����.gY0Cݴc��l��L����#���|}�o|���=[n�9V�7o�n����ɦ�m��p�恸[��:��cnZ67m���p���}��{�po���R��%N�W-�7�*@}T�&Ɉ�1~�����}���'ik�`��`�v����ۋ �Q7eM�B17,%�`�1 6� #qR�"�٣/i[R6���m��{n����?n�, ��n x=�jv�Kym����7�9���۟=e�ӦB��^aUt�8e/&��Ab��� ��q`�w o}� =�m���R�!�Sj�N{�ٽ���>CH�9'����7�ۀo}��w�9�dV9-DC̤6L@\�n*@}T�rX��Wlm�F�v� �}� �{q`�ۋ 7�� ��m��]v�h�%�� #qR��6L@\����X�F�hPrW�-��<�ι�z�:�mMü��.��u՚���x��}�@}T�&Ɉ똀��H�Ⱥ�C��r�[V own {�ۀo�����ŀ����i�ۢfb�/ד@_�)QJfL�̅*�Y{�����ـjg���X�ʚ;��� >�*@m�:����wS�s�[Հ~�n,�}� ?{�pww�5V�6���a"kkl��i}�G1��E��G\W �8��x	��qҩ�VEc��D;V׾ـ����,��q`ݱ�k�Xۖ��� }�buvl�X��޻�r�s��r����A�p��ذ����:��0�}� ��k�[$vG�[}�@}�*@m�:�7\�\��ʣ�� �M(	��͛�{�&z���v˼��s2�qΠ�1 �EH�ۋ 7_�0���Ғ�VBVܷ�ss�oY]��pѴԤ�
���W:k2�b(��]��� ��@=�R�����S7�]E�R+P�����$��H��P��_���V�U�/��.���;�H�ʐqΠ����wq`w�9�dV9-DC�`{������*A��9W�{�@Ow�.�Ĳ�ݴnI,������q`��ŀu��0.s��)���⥮��*Nh�g�7=���f��%͌�ݜM��ˈ�r%��
�f;\q�6����-�M<��*���8��>�1��Q��S0�\
	�68dgJ9x�N���� ru&1qW+^��pH�:�n9]+���C@pp	6�������KvjZ�-lC��L]�5��:�?�[��6�2����N�����y?��F���.�WW2L�հ��z������	����[m���V���6��V+NAeZ��Ih� �������X_�#�$��f�����L�C�C¾�w/�H�EH��P똀�ȫ ��.�SqPln��`~�� ��&�fI�K�I�E�u*� {���8���m���n�۸���ŀu��0L���� V+@�&h�2�̙.d̯;��>�E ~���udEN��!B
1ʬl�rk�:Kds�["��j�<�a��k��Sñ^���w2�k��mΠ�1�, Ｂqm"��j"� ���a�5N,F�� �8�������͚76��^R�I�2N��/L��m�K0}�\��qa�\\\M������;�����Ih�s3A���h���/��P{�� �^\ϻ�����'*�ʰ��ŀm�:������r]]_e{e`��^��n����փ�Bl����cX��n�cV�El�$�O1�T9D67lrڿ �Ou n�����l���	ܰ$i�
�[f w�ۀ~��,�wq`~����\\l�3u�꬈�;@q4�v���)Q-l̥2I!�A�!��'sp#[ִ�D�؀��� h2D��V�d҃�F�	�&�AB!R,�LʹM�+i,�
B��H�F=�o��P�@��R�,�)t�Ѧ5%aHQ# �֠F��A(��@�H����"ƌ*1J
�J�,�H��*�`A�6��B,�H�D�&��a0��JַMluд� 0�nB�� �q���2i`Ԕ�F3Z���E	mJ:��Ic`FV��++.�Ɖbq�5��5d
�,.��1�B$���		h�)�����1qD��|P�Y�.ϸ�A@�Y�G�S��U�E(�P��� S�"Uǀ�q:#&'�Ƞ��k��K�x�`D�*���Ҡ<�y�^M$�������n����*܅�c�`~�� �s9 >� ?s��UTeO}��f;n�d(#=�յ�@��1�g���ﯹ�u�t��g���$��Vx��>��T�̥��32f�>�E����Ɲ�rZ�U�ۀ~��,�wq`~�� �}� ��XKl���r�\� ���X_���\I��߮���Y��g�j/�T9D67lrڰ>fI3=�f� ]����R���fL�������t��Z����+m��^M�2d�ٻ��^�*�w�@{0�sߝ!3��v�&����oU�N$�Jvۜ��5��v���n���tg���p���ȩ�ȩ��� �s5��/��SY�Y���}�� �+&�1�z(szh�2�rd�xBxҸ�r��j�<�~���n�۸���ŀn�+�JK�ҹ$����U\�n{=�H�EH��P�ݮ6ZWe��X��n��?ww�Ƞz�h	��|�e����Kڳ$m�@R��!b�v�IJl�ڠ�Ȼ�n�(�h�bst�N:p�^�Π{tkxV�F�v�Yf��d�G]����v�/f ��b��qx:_l��áɱ������9#�7��Y�.����m7M9ڶݸص�շV�p�?���؛�j�X@燶�=�n9�#��E�g���;t�(8���v��2v:C�q��MnNC��{��b�9�ys^�q�E�d�\���4���j7�kf1K(Ua,�[$�ʥr��oذ=�E {ד�&I��f�*w;1P��v�-� ���`{��n��?ww w���TR4ԅb-� 7\��EH�Ur��z��Hr{�L�����,VVKp��ŀ~��,��ـ���~j)��5,B;�H�EHs��>��� ܯb�&,�{r��XI$`�%����[��ʽ�]��6JE7kF�2���<6��]�E��H��P멈���l�`��ɣ��촎I,���nbI&T�I$̵�U��*7v����=���%U�kuV:��?{w�ȩ��W.����{��Wo�و���%D�J��d�E�w����@����q`�E�h8�7ls3)��� �u1�R�R���ߗa� 'vz�����xn��:�soa�͙n��L��r�.��t??]�N9tfg~ nW��R�W�W����>L�:� �YSNEn�۸���3��ݥ@[�lP�k&���io�>��b-X}�ذ�{fI\�I�����n����2i]U��Yy���s��'�����R��ŀn�*�Imm�hܒY����EH�EH��P�s�o������b}\ҴU4�+m:��O5Ӈ3sm�95c��aS�]���"�K�����~��R�Rm����b޾��Y%�Aʥr��wqg��C_�L ��\��q`�ܒ�:�;����nu n���ܪ���*@k�� �Zsh�"jB�ف���I�n4�v���)P|��`�'�����8v� $FD��K�%�޷� �;箨�EeM7+�����*@m�:�5�x����ڙ
�g+��P�0]����mH�	�:���\e6���dW�^��n͔����s�[���EH��4��܅�mڰ�{f w��p��ŀw}���e[*���-c���@�� >r*G���*��yRܟL���U]����\��q`T��nu ks��v�e]�;��l�U+�`�n,��ـ��\	���7$���IE>�~�l�����Qc�E��觊
�]����+�c��.0��lY�H3����U���`xw�S�F<��ո;	��n��˵^��жvY��h6�n�뱥|�C�w;X�pW�a�<vr[�����5�p8;3����b*�٣�V���nIga2�a�u�cc(/��s������mgu��I9����q��բ���v�+�i<�n2��������o��v%+Y浌���^7h�mr���c����v���F�j�uT0�;��_�����~��_�w~�ߘ{�� {�4���F�#�Ffu ks��˳g�� �<������=���)*�rˀ~��,���s�[�����ٜ��(�e 68���� ��q�V {�q�H��Z�ݫ ���`�;����T�#�]_I_�K�|��ی�T��<yz��<�\v˱2��n@u=01��!4�րhČ�������o��9 68����gmΝ�;����eU�,��n��ܜK��.�=�ŀu��0��˟͚���r�$�H9T�ܤ�ʐmΠnw9 ���*j,+vڿ~m�M܆6�}��_ߛl��+���������~�i�N�5!b-���o�����m���q��w��~��~��m���o��v�X�:����yis���e�۳k������V3*��BR�����B����o�b��o����~m�M܇y�F���f6��?H���8X�;U����Y����d1���y�����n��m��q�aUoZ������^��7m���o���+�P�,��P:*s����3v���o���m��7��i[r��nXcm��ݾ�r�g}홻m��}Ü��Q׳�Cm�����d��%eU���6��U����n}_}wv�"����]���{�K���(Z�U8�݃V�+�#ܽm�R�p�u�Q3�@�Oa�Ѓv��q*�ʮ6���o���m�n�1���|����g�q\m������J�vʿ~m�M܆6�}��ߛl��+���{��~��~��Rm�R��cm��������n��o�����ͷ黐��{=���E���v���g�q\m������^��7m���"�X�1,`����}g9m����ʐ�b�Wm��������7r�m��{~m�۸�6���Z���p�����wC<��Xz�]��g�R)�[L'=/� �yؑ�Wc߯������6�~��ߛl��+���w��~��f��ZVܵ7[��m��{~m�۸�6���o���m�n�1�߶�=Q���YUvGo�Ͷ{w������~m�M܆6�~��ߛo�����,�U+�\m��{/ߛo�w!����^�ߛl��+�������%���e_�6�싢����.g�]ݎEX���[�W�]݈q>0�$ a ������~�|[��2����t�d>i��$QqM�4��K!a!A����6�$��!bR�c
J�!,���"��(N�20� �х"������! �T�*l�'ʞuR��TYФa�ʩ�1YlHVH�#$X��bD�A�H��E"�aP�X!)Si#��i4�CHH���m��m�@��hn�K�.c=����Y�n��vL��i�,�)��Kh��;9�% �Tt���w[Zm�+c���
'�n��}6��b}Jz�ËP�F�5V��;w�Xݫ��+�����u�u���U*N8g��v������W1���s�������%��*�ͽ���ݺ���������o;�݇�f��x)��c\�w'l��;(aP�є�9���r�Az����ݤ�ayx��"����(��U�!F�ؤ#n�9X.ֶ�m���䵘12���s��Z�j�%yw��+�+U���GH�]� �q=��i�^-cG���9Ɲ�yJr���j�W-:����"��&ӓRg���#��1��[���8HS�g>�> �vK,q5��):l�˨������[�}��};=U�ZWH�E\]/>2g?}7�t��F�jۣ�3�`g����;��k�J�j�7.� *�Vz\7N�h���0/Z�w.ڭ$<v��Ӈa㵵(m���97fY�ɦ˳h��N���@�)��]�^TsԔ99B����`D�FvwlqӔ�u��sn�k9�8��桔��b�+�D���q#ƨ�:-�R#�������`��v�'�ʟqAP�ɵ�lkg����u�>�o`z�ͮ�/bm��ԡn$K��һ����x�H[����p�����'��<��'N���a{p2q>:m��.�c�n;U�b�\l��k{#�60
�Y���F�!(MQ;]��&Ÿ�kxܭJ�*A����	U�ha:뜦۲����
��*�<�T��c���Y�l�R֦6��euMR�\�-\��v�v���+���t8�͛�*�mF����6m����1���md�C��y���`�3lʊ`a��A!�>��u��v�ajܴ��#<J�����q�6��m��gnuX��v����ע	t�qC�p�1��պ��u�X�eC�{N��fd�"���G@pE�O���tO�N�Q 4<?&*=��uT�^�'~�ɬ�f2f���m�Zu�23���].��Om�@κ�I�X���Ԥ�uצ��:�l�znp":���*���{n���!��:�u��{&���Wl��"5[�[!n�]�Uq<X+���[�ڹ^�x0�Q�u���i�-�pܳ�a4�tΦ�3�΄�<�nт����W;GM����R��v$;i���2>yćav�������s���~�e��;���k��ۓ��:�R_TH��M�q�b
�3h���}?Ys�N�m�����~m�۹La�{q`��L���,,*,u��� ��n*@}A/gf/�U~�w��C�t�����ay��3w�P��Tw9ē?}>����8�6V�3(��) �EHz�1 ls~�9W�oߖ }����KJܱ7�`}��@~�9o���� ȩ�ԋ2��-����]��r�EJ�Rp�;V�c�CT/N�[Kk&��d�A1,k�V� �� >� ȩ �_f 5�ȇ,�K$��J���qg�G8���$�ę�.fI��w{�T?ll���po�̪+kA`W,� �wq`��b �� >� �/�f]���b�fU�2L���@��@}��X��� �x���E�� � 69���H�*@;�و��k\]ۘO<XLUW7�Z�I�F�l
��Z]�q����k��&���<v*�m�� ȩ �\��+����~���8�q�[��v����y��n {�ۀw��Y��}����KJܱ62nI��k�nI;�}��+ "�0�� �?4��=�\�����~0=~�[��%e��[p?�r�w� �T��<�޾�@9.���,�U+����ŀ{���J��~���	n{1 =s[�WW�A��P;,fk���m��:dS���iE�]�Ƭ��߽����V��"�w����� ��@n�� �yp�V
�FX��<��?���p{~ŀ{���g�mq�TX��	31 ls�*G��s�q�ʐ��f�#�ڝ���u4;n���O�߿�{��lܒw��Y�0 M�D8(�{�n w��q�[��v����@~�r��| �=�� #*d��������];u��0��l�n�7Z�k��a�5̊��ֆ�T��g�w�1��H�*@m�}�-VZI+-,r[��m�?{ۋ �wq`}�۟qs�����vR�l�U2����<��y~�]�sو9�@{w^Z��8A�aKeX��� �3�1��H��켬�V�lΗ�� 6����r�9��'� =��X��I=�m����YZ#v�9"5:�2˛�g�n{C2�v���eV��z2X̷b���L�n��۲��1���Щ�l��WF�5b�7�o;{i͔�zl�iٖ7n���a�Y(@����.�3܅���/:k�`��xs��q��1��]N2�`u�����U:��a�w�a,Y�,�6�7-�m�Wd8�m�۩b�Ls��j;b����]���k�9맳Y�0��J]�V8�]F8膨Gm���gv��Jd�g�9��Yܫ�34�Ob[��dT���m����jv^��C����Ur����T�v��1 Mvw����Z�ݫ �wq`}�ۀ�m�;�n, ��oeRҹlRF�X�^D���h]�*�ffnL��F�u`����`Ui%��:� ;�ڀ��� �;��t\������y�+=rzomj�]g�uŷ�ޤ-g\A8$-(7e,�r���J�}��@=�R �s��69�$]̫�gn���kZə�7$���������_BE�� ~��� >o/�:b����	�V w��p��}�ŀ{���f���ꨱYSD�\��s����� �T�{"���q ��h�P�m�;�n,�}�ߗ�<��[��m�?xס2XH2%iE���M��W�#�֦�t����)���� W]U�P�j�=��X�}�h�y<������6�rI�;��:TL+��9� 7����������=��X_vCXG]rZݣ�Yp�wٹ'��n
�"Q~Q0�Y�{�X�nˀwwr�e����R�n�s��U�=� #�� �;�c�����9l�A�$�����ŀ�;�c������L���(˻��ڌr�+;�tj������F�.Iz�\���Gg˜��,�2©�I`��~ ���� �� 5�� �EH	d/*�,VT�%� ;�ۀw��X��� ;�l���I������}� �EH�r����终�{tz���Z�ݫ�%Ǿ��� =���ܒ}��7'�4'�� "� H���Q��ԢHB$���wC2t�Lʲ3mP�d9��`������r�����@kqR옰����s��)��R�&qXm���\Ct�ۢp��X��k�ҏ����|�.��+�K[�u�/�>���{q`��, �}���ܩ�G-��9T�[�kqR슐����_˲{޵�;i"��IKeX��`{��s�6{�������Y6�����\�7$�}�k78ؖ%���T�Kı>����Kı;�kdMı,S8�=���Qbv�Ie�/�8��%�u쩸�%�b}�}�iȖ%�b{��ț�bX�%����iȖ%�bT15��ݻ���e֊e�f`l��BSu�Wj^�k6�Qx-��qWi9��غ�����=p���<h�u�z�4��S�����>L�a˲Ͳu�(��T.�V�W�䕴b���	��U��
���e`�Br]��mbϞ���k��]v|�Qs��k������.���Hn����@�G�=�!�]�E�U�.w\�OX�b�y7h�Qc��>�鿿��{�{���߯���ݺ�	��۴��z�8�4=p�t*�Tv���=���m�2�ڑ�K����ʞ�bX�'��~��Kı=�kq7ı,K߻�f��'�5ı/�k�T�Kı/�ǵ'뫆[�L�Ys�"X�%���[��~:���%�}�Y��Kı/�k�T�Kı>����Kı/}�2�a\�F䒜Xq3��L�~�\��ı,K���Sq,K�����ӑ,K��}���Kı;�wZ��e˗Z̷2\��fӑ,K? ���M~��eMı,K���ND�,K���q,K�Q5����iȖ%��{�����i�T���Mﷸ��%��{�ND�,K���q,KĿ}�k6��bX�%�u쩸�%8��q-^���T��%�r�m|�R�^P�#�wDv��WF��\tM�����֝���V段�3XpI�=�hr	 ����͉"~���=ı>�}�i���&q3�W�{ �
HE`�V%�b_�ﵛNB��٧Q2%�}�{*n%�bX����iȖ%�b{�1Xq3��L��i�N���Z�fӑ,Kľ7ı,O��p�r%�bX�ﵲ&�X�%�~���m9ı,N���ug�1���CW3*n%�bX�}�p�r%�bX�ﵲ&�X�%�{�}��r%�bX��ײ��X�%�|t�髆[�L�Ys�"X�%���["n%�bX��w�ͧ"X�%�}�{*n%�bX�}�p�r%�bX�kޅ.������z3㭞�3`���ǎn)�ͫ��v&���i�.n��&�nl���{�[�oq������fӑ,KĿ{^ʛ�bX�'�w�6��bX�'{�l���%�bw��<~m�VZ�Y��~����{����{*n%�bX�}�p�r%�bX�z�Mı,K���Y��Kĳ���~?F�H8na�����oq��ND�,K���D�K��M$B�0���a��RwVs�\���$��[�Ѷ�U�$��
R�0p�LHA�*�H$SDC���1�!�� ��D4D!%�Zj,B0���T B�>ti!�@ڎ�!���䣠�SCP�H	�і�fj��oz��# ��d��6N���pC~w�a����R��+`5���L[� 4H@�PA�љP�<$��	������Tbc4J�t���@X�aK��,�`���P� �\(�G> C��+:�z�))���B�=����͇�O�j%�b_k�L�g8��?K-�qF�q�YM�"X�~Q j'��\"n%�bX����fӑ,KĿ{^ʛ�bX�'�w�6��bX�'N�ֽ��$�4]L��aq,KĽ���m9ı,K��쩸�%�b}�}�iȖ%�bw��ț�bX�%����2L�fh]WZH���s�eu"��3�b��LS��EnLdL�Ԓ7RI6g�����bX��k�Sq,K�����ӑ,K��}��?ND�Kľ��k6��b���-S�H��R�!����g�b}���iȖ%�bw��ț�bX�%�{�fӑ,KĿ{^ʛ��MT�K������-֦a,��ӑ,K���kdMı,K����iȖ%�b_��eMı,K����q3��L�{�FJJ�#���J��Kı/{�k6��bX�%���T�ʚ�bX����6��bX� �'H*�Z"VDB(�R!R%bЀ(`@������PbYA �g�}~{��P��N2q�^:�B&Ix��ySr�5�ND�,K���T�Kı>����Kı;�kdMı,K�w�4�ᓌ�d�.�D�$&T����]���,p1�D�5��N��`�g@�秲6��`�A�s����d�;�߸m9ı,N���q,KĽ�}��~Y�MD�,K����7�L�g�}��X��1�-�g�ı,N���q,KĿw��m9ı,K��쩸�%�b}���iȦq3��^^nͶ��c+�Xp�,K����iȖ%�b_��eMı,K��ND�,K���D��g8�Ű��n����.q~�bX�%���T�Kı>����Kı;�kdMı,K����i��g8���6¤5,B%��dKı>����Kı;�kdMı,K����ӑ,KĿ{^ʛ�bX�&�? @���O���kF�ubع�n��,�z�z�9�8�+;U���t'<�G���pʜA��M�O��rhY�N�]�rX5�o��_l{�j�m���Fzw-�㓎�-nN�[�������2�#M��I�oG;5�{r�nܗ]�f7[l��9�3�[�FqK�
=���� �t�h"��Dql����nt����u�󳊹�fu���<��]�7m��R+�x�k?~g��U&�)ʇ-�[;��}Y���x�c/+:u����B���c���ja��S0�\É�%�bX������7ı,K�{�ND�,K��{*n%�bX�{���Kı/��5��R;k,$��É�L�g����"X�%�~���7ı,O��p�r%�bX�ﵲ&�����'z�~աk�b�����{��7��_�&�X�%����ND�,K���D�Kı/{�\�r%�bX�v�y+v���J�&q3��]���iȖ%�bw��ț�bX�%���ͧ"X�%�~���7ı,O{�������GIeY���g8���n�D�Kı/��m9ı,K��쩸�%�b}���iȖ%�b}�a�&�t�Lf{O=[�����k�;8z���{N�u��Z��I�F��"n%�bX����6��bX�%���T�Kı>����Kı;ݘ�,8���&q=��n��GhW5�siȖ%�b_��eM�e���A���Ȗ'=��ND�,K����q,KĿ}�L�r%�bX�5�j-�HjX�Kk�É�L�g{��iȖ%�bw��ț�bX�%���fӑ,KĿ{^ʛ�bX�%�����n�3	e�6��bX�'{�l���%�b_��m9ı,K���Sq,K���{�ӑ,K��&��J�%���J�/�8���+�{�ͧ"X�%�}�{*n%�bX�}�p�r%�bX�ﵲ&�X�%��ջ��ܤ��F6��T"��m:&�ܾrv���T���[Sn-�2�աkZ�2fӑ,Kľ7ı,O���m9ı,Ow��q,K�>���q~8���&qw�r�º��kL�ʛ�bX�'�{�6��bX�'��l���%�b_��\�r%�bX��k�Sq<�j%��x߳�f]j[�5rk5�ӑ,K��}��7ı,K�{�ND��W�h�A�F�n%��~ʛ�bX�'����ӑ,K���n{Y��՗S,��D�Kı/��m9ı,K��쩸�%�b}���iȖ%�bw���Ň8���'�=��klj�B9-���Kı/�ײ��X�%�����,K���kdMı,K����ӑ,K����0��٫z��{v(���{W[����W
�[��F5�ϫ�R�ԇ�m|Xq3��L��w�6��bX�'{�l���%�b_��\�r%�bX��k�Sq,KĽ:wD=��[�L�,��ӑ,K��}��7ı,K߻�ND�,K��{*n%�bX�{���Kı.[GKe�����&q3��O�w�6��bX�%���T�Kı>�}�iȖ%�bw��ț�bX�'w�M��h�v�8�L�g8_��eMı,K�w�6��bX�'{�l���%����"�5�O���8�L�g8�_�`�]v�G%R�̩��%�b}���ӑ,K��}��7ı,K߻�ND�,K��{*n%�bX���~�J]~$�Ԗ�m&s�m����֍���YZ�L��U,:e�.B��[�I8�%������q���=���q,KĽ�����Kı/�ײ��r&�X�'{��"X��g�o앑��8V'mGL�q,K߻�ND�,K��{*n%�bX�}�p�r%�bX�ﵲ&�X��g��T��5]����_�&p�,K��쩸�%�b}���iȖ?�����~�ț�bX�%���ӑ��&qzl�IR,D��,8�K?@�N��"X�%��~�ț�bX�%���ͧ"X�%�~���7ı,Kӥ��	.�d���iȖ%�bw��ț�bX�%���ͧ"X�%�~���7ı,O���m9ı,N*����jr�p�m�XAj)�I��7i�3Q������m�e��;���<�G�,^)ա���.ۣ[��8�X�Y�G:;d2]�Wd{=����� ��r�=�@v�+�䵮Y�/0�'#�,�	�ն���x�yu�K"H�V��b��1f�s�]���63<˵�.#��C쯞+�xA&�ZѮѭ�,�Ƒ	cyk ��9YE�2��3����:h�Ho�d���]]]��άi�k�Y�v�����?�����nxgC�՞��=V,�u ݽߛ�oq��K�����ӑ,KĿ{^ʛ�bX�'�{�6��bX�'{�l���%��/i�z�-+��갲��_�&q3��~���7ı,O���m9ı,N���q,KĿw����K�q�߿���DS�K���}���,O��p�r%�bX�ﵲ&�X����MD���\�r%�bX����*nq3��L��ܒj��1�-�g�%�bw��ț�bX�%�{�ND�,K��{*n%�bX�{���Kı;�}��,���u���aq,KĽ�}siȖ%�b_��eMı,K�w�6��bX�'{�l��8���/i��UEmN����Xr.yQoTI�N�3�m�I8��nbx^�&[KFb��El�E�������oq��#��X�%����ND�,K���@��ND�Kľ��\�r%�bX�5�V��kX�.�K��7ı,O��p�r���k`%��B	V*'��+Ǒ>�bs��l���%�b_{��ND�,K���T�Kı/N�Ғ��K�2K.a��Kı;�kdMı,K���fӑ,KĿ{^ʛ�bX�'�{�6��g8���t��Z�%���J�,8X�%�~�����Kı/�ײ��X�%�����"X�%���["n%�bX����e��Y�.e̙��Kı/�ײ��X�%�����"X�%���["n%�bX���O�8���/�����Ild��y�8o����^x�-��.��:�Ў���bv�\��ִkXk.fT�Kı;�߸m9ı,N���q,KĿ}�L�r%�bX��k�Sq,K����k^%3&Ye�5�Y�6��bX�'{�l���%�b_��m9ı,K��쩸�%�b}���iȖ%�bw��[�Y�4]e���D�Kı/�w�6��bX�%���T�K�z�E?��A�)�O�o�>��Kı=�LGL�g8������������6��bX�%���T�Kı>����Kı;�kdMı,K��}3iȖ%�bt׵o�SZ�K��R\̩��%�b}���iȖ%�bw��ț�bX�%���fӑ,K�>�����g8���K�@�VH(�:��'S/d'"��֖�v��W\Ɛ2�8���e�).ۗ5%�0�r%�bX�ﵲ&�X�%�~�����Kı/�ײ��X�%�����"X�%��-���:G-E��QŇ8���'߻�NC�Pc���b^��쩸�%�bw��p�r%�bX�ﵲ&�X�%��N���Y�5���\ɛND�,K��{*n%�bX�}�p�r%���MD�{["n%�bX���ND��oq�߿���"+#��*=�ou�g�`j'{���ӑ,K���kdMı,K��}3iȖ%�T�dH�Q.�'3���7ĳ��_}�$�ZV1�J�g㉜N%���["n%�bX�}�Nm9ı,K��쩸�%�b}���iȖ%8���[�ڇ9YF�!�cD�9v'��q���kp���V��ݒ��k�Q�Af�۬�Ym.f7ı,O��6��bX�%���T�Kı>�����MD�,O{��D�Kı/�O~�k2�ܚ�3Y�L�r%�bX��k�Sp���MD�;�߸m9ı,O{��D�Kı>����r%�bX�5�[�Թ���.�3*n%�bX�}�p�r%�bX�ﵲ&�X�%�����ӑ,KĿ{^ʛ�bX�%��:R_ۗ5%�0�r%�g���_�*n%�bX��Nm9ı,K��쩸�%�b}���iȖ%�b_x��Ѭ�rkY�����*n%�bX�w���r%�bX@? �u����I�;�߱7�O�H$��(
���(
��� ����TQZ�*��� �+�
���*����� ����Dh$Q@!P E��E b)P(�AA�1E b$@�A�*���������(
�����PE~TQ_�PE�@U�uTW�Q_�PE�U�U���d�Mf��#���f�A@��̟\���  }@   � �      �    � ��@ IRAJ�      P
�!R���PER�IJ	@TR� �  ��%B�   Y%@  P(c ��6��rk�{�뷻x��� �T�ݔ��\���g��,�S� D� �  �� N� ::iK��� ]`��YA��(=�)JD����@����  6<�P   ( 9� �)�H� �@LMѧ��(�@�����%:1��=���i@���ޥɪ��}| g����6T��>Mo=)�ﲽz����u/g��e\ �畼q�d��ݼ�]�y5/x }�@      ,` <��m�[�[nm>Zrj���zz� =}�W�y������w�Խo{u*�� n���7Ͼ�����u�N� 9�  - 4�
���٪�ʫw+�y�{+��P�y���>��|��������m� ���P �@Q� S�O���{��_6��ݼە��{ʮ� zS/}�]��u���=v�o}�)\E�^�w}�^Mx �x����{ޕ}�}������^�p�n=�/-���oo} �{�K�t�����e�ۥ�כRp }�@  P*�Z@^��6���ۙ3����oMn ��mi�޼��w^��i�����&^�}ϯKşx ��z�-ͽ5� vOJd�ҹ��}�]>�zW�����n}���|Y�[������zt� =AO	R�  T��5=5JUM4�&C<z�R��  D�*�IJ� h �?Е<ҥ* �"Be%I�0��*����~������SF����$�30�����AТ�
��EE� ����*+T���O���Y�X\1�X�kZ�:aqaBZލh��1q֎nH\ѽ��6lމ�fMf��5vǜ�����u�M�R����gX�v$a�f�$$�o�B��])�ّώ#.&�\�#��6�Wo{"Q�0ӳr$(bivF�o��Xމ��̉�ѭ�r��a�s'2��� �y��@o�6v\BS|���Χa�X=c�gw�Yq��!C.�!���8c�"L�d`H����Sf����7D��)΄�h���I�G3���0"�v�"�_W��a�[�����^��!q��6j!H���NJ\�޻��M��oil6'��NX�ϊ�?���~D�3��~aCa�>X.nd���z)��H���k}4t��Ά�cH]�}zv����|I�ѭp�*�!��~���t���~5�G>ފ�fMe%�h�A.j\�H���5�$����p���)ao�B�L�RXKN�O#���MgA��*��i�h`rf�	�Vo7j*lW�S����W����U�/�`f������65�1HP ?�24Dы
���7�4�M�w��7�B�҇R��F�jh���	�a��h���`���j����)7��Lx�f�#�j.��cO�B�,����0�,k
щX.���h�f�bF���k� d �lB"Pd��)��I$��0����l��$�0btVcSyﵣN��XJ�đ�	2�)�2�;�J���`�	#\T؄�x��q��Ѓ�-J���a&L��B�d;��Ϧ<��M�2l$�|�$A��X���,*E��g0�|ɬ�aHf�o�O�4� ��4%B "�Z�3F�6� H�Z�XD P�a\��˦�RB���@��]Ç
t��%2�f��ӡ
q�o�,�9�sK���j�� F6kf�l���5��INi!L I���kP��!��$�hpI��3�2P�4aFm>g��J��%	P�#Qa,7�Z8�!$�)�B��Ʉ+��
33iU�@��@��Ar]F�s.���X`�N�	 �D�1b5ؐ�
EbHQ��e%�H��a
g8m�X�i۲%Cf� �P7ICz��Iv& i q�N�'5�gO�|�f�):JvR��HSƽ�q�D�)DJBBh��ʡa��<� �$�l.1��X]�6,J�vl!~�g�B�7rߛ��o7��R���+;`C|�:B��o%>:��w�Y~��M[J��b�a�s;�d�>��
��#B0di���)�6R��13gIIq��C�˜��m"��9��'��믲�s�o5����I�>^�O�Ʊ��a߾��ϵ�!.���[`�K��x��M5>�ٚa37�,k�B��.h޸ˁ)�ᡃ�X醖��ZsU��\�an ��v��������e29���A.��rl�sa7�4�%��S4B捇��{���Mf����sA���K�rSA��}��\��K��fM�.�6VR�\�%�e7.]lasL����v˛1&�	�E����.��5N8�!L5��1%1�0HS\4��h�nT�/���
�yR2~Y��4��"kD-ȴ��h�
m�B�2�XR�+HZbB�Yn��Gp%�oP�ZS�0�R����֒�kN\��C�Hݚ�.�$(���B�!J�hP�H�dPcR,x�p�kaǁ��k�"Ub!tn����X�<�7bB,H��h	��bE$0"Čc�V1`RA����!�Rh��"A ąYRP��&�h�GB��%V W��/�J�2Y�|˚�Á����2���R^�3(B���H�0�smI%��p6�!��51�6�[Ć��(˭�y���O�'/�	R/�R���
i�)C	G
������s�[M`�k�i�k��}�9��� �9��Z�A*B��G	����.���4�]�D���m�f��`�ы!�fdunBd�6���\5 �F-p�mt�B[�&�F�|K�l��6�1ѣdod�:�ݳT�)��HҸ1i�iV�f,(eaZ��0����e�M�70({���C�X�h`sĮk7�{�>v�`� qӱ�7���ƲoY9��e�E�v˝eIFP��?�a�j�١��!K�(�pK��N�B���p�;.���}��˚�Ir����7�5�|�H�
}���u^a��2��IL!@%!s�\���z	LtB����s5˭o����ᾬ	ߊ�]5�HS\p�X��yY4��&��k��F�sz��5��hރ��a�zS��S�1'YB3R$��`CF���>��a����w�y�9��$�F$ @�B���B�B���0�0�!C�}��)��U�\�aP�)����t���ǐ�hv�ǁ���ͼy����4�4��Z�kY��HP%p:�G>!aL������7�|s��*}I�DR����a	���B�HS%�(�.B�(���0��y��Hl�eÔ��BF�p���,��1���8�97f��Xh`KL�MB9a0e%���2�f���#Ie0��SO�
a���Jk:/�f�d�,I
��2L4n��,������1�)��@ �6�Fv�Ʀk+#�xs�~�W\�2d�	a�S ��q��p�p�%��aHXR�Xō0\!p�/�L�Ͼ"��0hiD������t���D2J3n)Ϯ2�E�ޏ�����9��p%��Fod�汲�L ��1"т�cC1�T0�FH`Q!cL�X�%��P!HS����cLHSxu�H��HW��Q�SF5�%��|� k)���Ʃ*��Z$H�X,V(@*��@
�!(A�B����"1 �!HЉV	% �"�XъF	!  "ĈU D�Ĉ�"	�E���T0�I�ĉFD0bE�A �X�,E�q��b@RHD  �����\։D�P�0�a\LH���_&�Bh6萍0�!�2�C2\!L�F��4o��La �7��k����1 Q�H�X�q�9��ᧉ�`jSLi�d)�R�˔��]m9trrp%%2�p�~�HD�`D�[ �"HJ�(
� u4
0����lv��ЛEڡ�`���a��D� mB\]H!��SjŮ	�� �@��`F�f�ŐJ�����A�b�\��`a��j�)�.�k��\tl�͚$�sF���ݼ$H��NÆݛ#Lѷa��p�CC�xJ�*l6;�L4�ٲ@ă\v���w�br��?s�y��*�ԟ�3�>���Gֈ�&�w@���Bz�	s�wN�H]t��l$�k�B�8q���s�!q�np��IsL�ą�
�H�1�B��H��P�t�����#$�@�B5�D"V41J�b�R1��o��w�i$�}�s��\�x1�ytn��)��P�9���YL4��epc\��0�Pav��H\W4`U�!�i��|We�%���]oq�捐���]��r�{�����>�r�V�m`C�.e0��y�2�7�B�¤�iơ����I���ޝ;���;��U� ��          �  h @��R���R۞�P 	-���`m[��l�eÅIZ��(��*�O����/�h�΀*��f� -�[�n��]�Ts0U-�;=W���M  ����,����,0�qB:4%��f7`�3<���-�]t�mm���e��m�� @|��l [@i�� r#[�K�    :� H ڶ�im    � 	 �m�� -�e��l�@�����.���UV�m�m�      m�  H�[@ ��  ��     � 	4T��l�sm���� �kh HH��ٶ-��P  8�۶�l �Az�  l�� m� ����`m���L����L�l  ����=%�$��m&�['B��6ۀ �� �f�	    � mH� [��ێU��Z���YR�d�N�  -�������d���6�M&m�$ֱ��$ H	6�#��m� @ H M��iUyv�I���V��z�9���a M�Iv����f��.ԫI��K�83��.��L  ��k�Z[vݭ�À �9�mgu$MH+�ڦ]�\��w������طM��m�kh-�AT�f���q�|Wk�m�v�7d�pH�&��CN�6�r��{^�H���n<B�G�$�g�P:XZ���9�n۠3i�� $� ):�%�<^�fٶ MP���]{SE�
�$��9y� �l km�m�� I׬�.���ݦ]�Fu�!"en�	�e���ϕ�9��j�m[G.�E�mmm�h��6�jy��2UV��`5�Y%].���VZVW�&�A�'���+T�����kj$d��[�i;m�-� ��8��)��ksi6� ��&�5�����/^�6B@m6/V�m� �O���-� i�I��$I6����H     ��� � �m��e0��-�   -�H6�6�^-�i��70�ܶ��-� m�  ͫ�Y�r��r����ڶ[o���.�l [x�6�j�-��� ��I/ l ��lm��[@�[@�m�� [B�$  [@�$��� [@  m���  ���Ͷ jڶ��I[ myձme3N���&[@ �-]�-���vm�MdPѷl8 ��$t�m���4��   lm�[@��    	�m�� 8 -�m� H    l  � m�m  �m�  $8�qmn۩�lm��F�v �[\����6�m2��e�vt�L�	$���4�m�- [F�� -�l �m�6� � l 6�  �      m� H��p$�� m 6�f�ip6��h;��r�2ܛ�l]6$�`$ H   �� �����$-��$� qm[@8{moIm��%��-���'��-�( ��h3M5�l Y@ߓ}A�V���]�Q�)������[� p���[�I��l#�  [C�� Eнn�m�l�\�$	/i�@  6��m��  -��R��6���O�kX$�n�-K(�nm�sr �[M�I6t�{)Y,uB.n��u�h�Uz��!��Ϧ��GN�\� UR��:��X�r��Tl:��55m�u�![�si�R�;��l!V�:tp���Ѯ�ɍp[kpC��(�J�@�m�2��\�D�ۨ�c�]���m8�s<]t�ev�a�,Mtl�fi����K���[��|�SV�5ѷb�K�J�	kc2�܎m�	��h	<�ҼS�U�7kl�Uۭ]�am�͐�������U�)м�m����e$	Z��@e~g|.wew��m��N�ۼ��:m�MT$p��Կ}�ײַH�Ak�6:�z�[�p�b�Fb��-�X�l,��ĥ��	v���Îѹ��z2�f��
�u;�ЈX­UU�h���g�[[m 8�%� ��[&l�_Z���h*k36�YFN �- �l+�ׅ��[%�d���$��X�m�	�Ö����o�:�\�(n'R�b�m�$��΋z��[d8 ��9z��Z� �h�w���ӁK#�p9�lC� �� �vt���ʻ��u�i�t�-��	�Z�:ᶾ�rvF�-\ۇ;u�r�,髫016!g+[��l  �I:��cm��I�G   mm�b�t��%�Ͱ $m�� �\�p.�0�N��
�Vʝ�0��Uuܼ�zڶ�9֦�8���A��r�h i6�[R H �4U�z��@N�����>|햃:���R�Ļl;Z	y���"P탵+��.��;Q4�K����Nvz����rJ%�� �> �e� [E�knʝ`Wj���1B��,�ne�t%�bږ�����E@m]+���T,��U@h6ӥ�i�T��pT�A��m[��s�b.̘U���
�#m���5�JSm�N��g�a�J�:Yy�]��x��UURc=�!k*s�lڵh�^Vv<6q�m
�6�n4�3����&�s��؝�zYx�^i�.��f�pbG �i5�/T� z�@�[D� ���� ����\[	g8�8m���N�$ �γ�� �e�O.������r�ݺYw�,��!x������lk��p6ەv��$
ۓp=�Z���� �:Me���)r���h�[L8�6�j��.�|n�-���kX	 N��[w��L�v�s��i���m�_mYh8��  m���[�)B�U%ڕ@�8���m:�kn�ꪮ��"p��A#:���Hqi�����H�� &�\;i��Rԫu[4�m���yd�:;\H i�kH[dK/ګ�)iYZU��'������m���s  ��m�-�	 [v�PrN	9�gSzT�kM���oZ���
�H��@����^�d�e�(P+m��=��	�m �@���X�l=)�{D9&qZ,5��Y;^/�ѰWUT�*�YM�hU+3Iv\������v���9�`����P <�F�p��`0p�ϳ5*[e��+v�X\UQ@���@S�s�B���[\��@U��v�$ l�����eP3����.�jp'E� ���9:��7Z��m[]nI69�v����� ޠFn�V��v��\�k�q�h֖պ���ta��k��/c��%$�jR@�&ٴQUU��+el��mm  7$���� ��@��$�be�����&]�v��kmm� ������H�m��$  ԣm,�K؍w` �� [@ �m�4P8 �f�I�#�jͰ6�8����@m������k㉵Ź6F�խ�%� [�� 	 � H �Js��ۭlH��`
�Uka�m����	��caV�������� �:�U]mʲ���U�;/UԼ:��wg{;]*����V�v�.���n�g���V�YK9,��0$���@�n͖�q��$�ۜ&� [Q-��  	�Y|�X�mU[��l�\;E
� WR�U��  � ڐm���mpm�-�hn�$�0 I$� 6���tSm������[��v�E	$M��  [Z*�Z� -�ci$�7l [D�w[�  ڶ$  � �������[QB�m  	$P�` � A�� 9�Z�6� [@  ���iɵ"���� �d� ���H �p�f�]�$Zl[�ܐkZ@��  H�Z����������Q�m�Am6�  t�N ���	 mm���	8m�l�-[���|lm�H���l�dۤ[GI� �]��m� ֶ�A����Y5��n� 'YKJ�V��x �VGUt�T����Pm�h�m�a�H5�m�hԙ-Ml0��u) �&�g����T�N��n[R�l��m��彮l ?C��h � �	 �%�,��d�m"AU�p�b� �[^p鴆�"իx���cj  u�ya�Q]ɩ��Of�ggv����U�Z;ᴮ��n��ڰ o���@��W� >m̨l6�]�m���@  ��h1m Y` �e�u���¶�.�� 8 $ ��YxMR���� e��� �-�l  ?ӽ��{����~N�����{�)�"!���Q��"�O��8*�(	�:E QS��誴z�\ ",D�ľ
��P�oVb(`�z��t�(�&*��j; M,����� bt �>D���_(�� �C������!��
�ت!��:�p)�(|�"0Z�v <v(p8���u#�h>�"`�"�Ȧ*�
|�Q?H�(Ez"� *�� <��T���|��X�q]���4(���qU��/���t;CN��j�U�t:"��j��D/�R<TP�Ӏ���!��C�)���@\�O���P��Ub��Q��C������ j�t	��P��V
|��s�Q�y�]��mGI�hTΠ��_� ���v�/ʃ�i�T|�/D" /���T]+�Q4��G��EEx#�?�	3��w��| � ��5���i�l��[�j��j4�>D� �z��M���K\�d�]�@ٵ� �浀m��E�E�	8ZT�*+�58A�[t�j���=g1F�p��3l
uL����K��Ѐ��]���<�D������Mu�x���U��Nb�Nڍ�.�i��l�v���mc����"�#3� 8Մ��4cv�N��̷U��;X�|� T�4�:�t+-$M]Q��&��Y%Uu�Z�s�%vGB�Y�Sn=
N沲�4C�y$"���b�	�rҝLMl��[A�;	TR���KvNeU���
�L�h�gg�����^0`J%N�ݐe��Uu�*q�	֭&cfP�
N<���+s�-%���e�(VXFG:�6�\�B�fw���o`�.���t���M�6�w�Gkri#���������flq͌���f����{WbF<�� I�|��;n�N6��)���v�8�p�f8[-:�z;M+<�(m��P+����bM��N 1a��2���i�[.���N��-�c�¡���y�����7�a�Vʹ�p�k7�lԘꝱ�����
����-�ò'a�f�ܴ��6�x����(*h��ԑ�K!�:7�Q�c<��!:�`���tu��j�M��Z��Ssu��>[n�[2��4:l���DE�v�F�n��� �r�O=�V��G�c��8���]��tont;qt�@�wc9�v��ڍ�o�wa��c�V��CZm����;;��  ��:�ۜ�l�Z��Iï^sdb���7]'v�^ݽ8��6�9�1FE���Wv��cNhN�-�i�s��q����a�W]MJ�ڔ]V0΋����u�_ YM�N��{�����%��.��]�7�F̨�5�p�<eHD��6pe����N�ڶXl�ŧG]�3���9�M� Ƽ��U�\Yv�rK�Ε�%˱%s���������O���F���
��SN��x���
�<��.��Y,�։�L�&�r�Ƹ�n'��'�Z��v'�+�1���n��"s��@�˩�I��,�ʂ��UwQ�Һz�@���Tѩיp�k�cqy����:�G!�#����ä���ݷ����#�۰�����M�n��mv3�\��r;"�	��
U�#ŘsŶ5�6}����@K+H��':���3��u�q��Fݷ$l����`�a�v��UNAvy�p���T��T �e�D̴�^m*��y���?zL����T﬎yK\��Y]� ���3�|������@N�*@yȩ q%4�2�L�7so7�L@s��"��ـs�c�SQ7]u�J�y��@yȩ�1 ����Y�4(�ksov�ݤ������L@w;� n�M
CX�r���j`ݠ�������Yy7`("^�0��z�Z���� �tۙ�[[���v�b��}1R�w w��ݥ���%��0>wf��#��<@�Z*�Fڪ�U�=�T��"�������"v��e�yݘ���Ň����`}�L��ۚ7I��m�ʐr*@;}1 ���>���7#��$�XG,�Հq�0>wf�wf,�7q`�>u�B���ڤ-Uhz�]s���sB��ے랢��Kn��(����,#����埀���`�vb�?sw����9ݱ��J�N�y���� <�T�v�b���͆���"U�j-�`ｋ ����� "�~b#�+�e﷘{ݘ�۵ɵ�[uY,U[j����v�b�LT��R ��.�Ktn�Ke�`|�����X�nҠ-�6(L̛zNg~O2K�L�K�'�l�0묲nޝ�LpqHR�[g�:�+���5	knP�NZ����ŀ~��,��ـq�0oknhڭ�cNn�nm <�T�v�b��}1R��#��%�ZG,�Հq�0;͊9$��sz)P�ԨK��Lf�vn��n =o� 9��H>��~P(� ��A��@��-�~�ɀw}c�SQ*�N��0}1RϢ����5��߫�n�ߩ�\��;��m�b3d\������zn��^.�,���];vv�5]�ͯ�� ���I�}1R�k�kj��X��Հq�0�ݸyݘ�ww w���R���w7w�5Ϧ*@>�R���{��X��
R�n��'��O��� ���I�;n�!w[w-�9m�U�s���|����~ ���rN��f��>1�8�B��@�`u �q�� %�d-bB�$�5{$׮[[k4�sb��hW\#ڶ��8�a#+u��7��m�>��@݈��`���U�,>;�b0pl��[�\f�.:�u�䛑�X-�r[V
��P���swl�i�,d�]e����5�-Ʒ/�W�m���U��#/by{��ck!չ7Tj���.{N�,�<5�Ů�nwv^t��5p3Vݣy��W2 �!��.L�L`�+�Y§<�I.�6���S\U��Q9�����h�nE��2�sw6�_O� >�P�b���, ӛ5HQ�[+�`����LT�}�R���r��]e���W�f�9��H� ���?wv�Wv3`"U��Y*�9�����M@s銐ͼɷtVUd�Um� ��v`������X;�ŀ$�I.C}$g�7B��7��X�����"�\n�$i1R\�y{F��N���dr��Il����z��vb�9��,��ـq�u�+]qГSW5��;�}�7�3�uD>P<�����?�� ���=�j�ۻ�����-�ʰw�� ��v`������X�l�j��E��V�}1��1Ϧ*@>� A�3"�$�l�W,�?>���|��ow���w}� ��v`�ݑ�$EURvǞ�\�M�gpsizν2sOK�ל�ض�J��SQ"�:��`�vb�9��,��ـ~}ݘ�݌�Ue�"Uy�J��;�����E���sk�h�YU��U����ـ~y�&mdڙ632��ڊT�m* �͕�-Q��RKe�`�wf�wf,�EHo� Ηw�m���f��n 9��H�*@;}1 ���M�_�ڂBDK(V[Rl�ۍ�f�c��eW��a:�ݹ���K]�ذ��si �EHo� ����� 7{dsSn�-r�eX;�=����g^�� ��,��ŞI6��ny6Q�[+�`{�L���X;�� ��v`��ɵ	�Ⲵ�ف�>��|���T�������	"*HQ@�>S;��䓇v'�۪�ڋ%X;�� ���gw��{�L���X�U�E%G=Cd9s�����%�l�y9朹����/F��L�VJKh�UU��U����ـ;�1Ϧ*@>�R ��6�svͭґ�e�`;�s��I�{���ｋ ��v`��[v�+�:R�nϦ*@>�R�����s��惣�li�l����ŀq�0�ݸyݘ���9�I-r�f�������� H��]��{�����>�Շ�K�����9�j�C�P�h�xX⺆�P=	�4�zyl���+�i����镥PѮŊ���G<�@g۱��	9*��qn:�f��U��Վ&�gr��:uKI�rk�C��ZH<��jC]�WǵmȮH�j�f�."L���sXф�*m;W-�Nϣ�rrc'�n��x��k�kv:z�B�tVQo�����׽�}��-f�X��۹���}`m�dĽ4���c��앺zw6!�hA���j�\�{�,Kĳ�����Kı;�}�6��bX�'}}���X�%��}�fӑ,K�����ֈS.Z�֦kZ�n%�bX����ND�,K���Sq,K��>�iȖ%�bY�{ZMı,K�ﰾ�K-ѫ5�Y�6��bX�'}}���X�%��}�fӑ,Kĳ�����bX�'~ﳆӑ,K���{Z��F�fk�h���%�b}�wٴ�Kı,ｭ&�X�%�߻���Kı;��7ı,K߻�ֳY��F�52浚ֳiȖ%�bY�{ZMı,K��}�>6�D�,K߯�7ı,O���6��bX�'�N��Y���]2nM�oF��ga�u��@qs+	�B���ގ�.f�.(
؂R��*��7�ı;�}�6��bX�'}}���X�%��}�f��ϢdKĳ߿k^��oq���~~����W���L�ӑ,K�ﯶT�6��`E�Đ�Ab$���\W�K��}�fӑ,Kĳ�����bX�'~ﳆӑ,K��v��n[��2�Z�7ı,O���6��bX�%�����Kı;�}�6��bX�'}}���X�%�}��[�%&f��kY��ͧ"X�%�g}�i7ı,N��g�"X�%��_l���%�b}�wٴ�Kı>�s5�˅֡u��ִ��bX�'~ﳆӑ,K�ﯶT�Kı>ϻ��r%�bX�w�֓q,K����>��oإ�yE�ͭ�9�k����eݎ�v��3Ʈ�n�+cO-8���x���tkZ&�4q>�bX�'�_�*n%�bX�g��m9ı,K;�kI��%�bw��8m9ı,�R�Z��F�\�35���X�%��}�fӑ,Kĳ�����bX�'~ﳆӑ,K�ﯶT�Kı;�w�ֳY��F�j��kZֳiȖ%�bY�{ZMı,K�w��iȖ5'�U+�ύ!��<T�!�i�C�6 i�d^���$,�| n#�I�樲��$R-�
�:k��{������t��&�2�q&����&���D� �|��(1�aq�p�rItR�Q���"Ѕp�H��3Q�V3	R$	Yp����}q�c �
B�$1�hZ���H��H� " ,)0�R%e	�Q�E��*Ċˌ!.����$�W�=�\Ѯg�RҤJ�`0B��:,tj�-K
��D�;P:��P <W��Q؂��M�iU�(t<�m
�S��z'y}���X�%����>_��>L�3�ɳ[v���,RMf���&�X�%�߻���Kı;��7ı,O���6��bX�%�����Kı>�wm�Ku��ֲ�5�f�Fӑ,K�ﯶT�Kı>ϻ��r%�bX�w�֓q,K����p�r%�bX��������kM���Û��AyN�*�BE��nIdݎ���lƖ)�krB����,K��~ͧ"X�%�g}�i7ı,N��g���L�bX��l���%�b_ݿ���JL�Klֲk5v��bX�%�����?#��,Ow߳�ӑ,K����eMı,K��]�"~L��,N�_�]h�2�u�]jf��&�X�%����p�r%�bX���ʛ�bX�'�k��ND�,K����n%�bX��}��%��֮�L�h�r%�bX���ʛ�bX�'�k��ND�,K����n%�`T*�
"��*��D�=���r%�bX?t���I�F�k��Mı,K��]�"X�%�B}�M�$�wٳbH$��obj	 �s������$�k��FՎ���;��{;uy�E	��V�H����ԍ=�*p�3$k��kZ�OD�,K����n%�bX����ND�,K���Mı,K��ן/�ɟ&|���٬���W,RMf���&�X�%�߻���Kı;����Kı>�]��r%�bX�w�֓q,K���ݷ=-�fZ�\ֵ��ND�,K���Mı,K��]�"X�%�g}�i7ı,N��g�"X�%���s�e�sZ�]\��Mı,K���ͧ"X�%�g}�i7ı,N��g�"X�%��_n��X�%�}��K�&3R�5��ֳiȖ%�bY�{ZMı,K�ﳆӑ,K�ﯷSq,K��>�iȖ%�`?@ ޽=,�4.��&�url:7ے���9Sqv���1I�a���2\���k���(� �\��.єDIu�̣j�VBDv��b�q�صΆ��5	�޸c�ð�lF��O\���p��i�]�֝���^��v2Q!��{G�|a��g��K�t�/i�
ki#����^֎�b��5�ۧH�d�r9�k3�[��9�shΚl=�~{�y���c9b�S���[��,��!]`���6�/:J�j�o`�dh�D��r<V�U����{��7�����6��bX�'}}���X�%��}�fӑ,Kĳ�����bX�%��ao�e�F�5��4m9ı,N��eMı,K���ͧ"X�%�g}�i7ı,N��g�"X�%�.���F����*��?�&|��b}�wٴ�Kı,ｭ&�X�%�߻���Kı;��7ı.�~?�ϵ3$k��������ou�g}�i7ı,N��g�"X�%��_l���%�b}�wٴ�KǍ���_�k��l̾��oq�����p�r%�bX�v�eMı,K��]�"X�%��^�17Ļ�ow߿@}_�S�ݐ8d��z�3��F�!Գ��ۮ+�WeR�@m����5�f�Fӑ,K����*n%�bX�}���9ı,O��ف�9"X�'����iȖ%�bzg�?�-�jus3EMı,K��]�!� #�2%��^�17ı,N}�g�"X�%��o�T�OÕ2%�u�y8�(�-������gɟ&|�/�f&�X�%�߻���K����;��eMı,K��~ͧ"X�{������]��x�š���{��"X����ND�,K��l���%�b}�wٴ�Kı,ｭ&�X�%�zw�e�2[4kSZ�.�Fӑ,K�ﯶT�Kı>ϻ��r%�bX�w�֓q,K����p�r%��{��?��~� ݤ�6��7m�6�wf����%��'���-��5c��ֳXh�kEMı,K���ͧ"X�%�g}�i7ı,N��g�"X�%��_l���%�bw>ﵭf�Yuufj��kZֳiȖ%�bY��ZMı,K�w��iȖ%�b}��7ı,O���6��bX�'�����K��Y���k5sZ�n%�bX����ND�,K�_l���<x
��1)
�S��k� a�����ͧ"X�%�g��i7ı,O���s�k2a��asZ�k4m9ı,��Mı,K���ͧ"X�%�g{�i7ı,N��g�"X�%���s�e�sZ�]K��I��%�b}�wٴ�Kİ�*��~֓�,K��}�8m9ı,��Mı,K�w�۾��]Uh���a����1����9"Iv^�OV]أR؜VF�j�\�m9ı,K;�kI��%�bw��8m9ı,��Mı,K���ͧ"X�%���ٗZ�S.Z�֦f���Kı;�}�6��bX����&�X�%��}�fӑ,K�s3fYP��N2q��݀}D䩒fIu�6��bX����&�X�%��}�fӑ,Kĳ�����bX�'~ﳆӑ,K���W=�J�5���ZѤ�Kı>ϻ��r%�bX�w�֓q,K����p�r%�`u�����|4��bX�'�����Ya3�S�����{��7�ߟ�kݸ�%�bw��8m9ı,��Mı,K���ͧ"X�%��=�s�8����X�<.5�X���仗��儶m�/����Ɇ��1�t���mi9ı,Ow߳�ӑ,K���٤�Kı>ϻ��r%�bX�w��w��7���{��>��\t��Sf��"X�%����I��%�b}�wٴ�Kı,�}�&�X�%�߻���Kı=3�nx�̳5�eԹ�4��bX�'{���9ı,N��q,K���{8m9ı,��W�ɟ&|��zs`��)%q��Y���Kı;���Mı,K����Kİ~��i7ı,N�]��r%�bX�w^�th�˅֡uusY���%�b}���6��bX����&�X�%��뾻ND�,K�{���Kı:*�����M�}>d����	Fn���s
m�c�h�9�Z�;���v3r�s�4c��oC��n�p��\�&D.�:/I��ӣ�M�)�ɧlZ��"k>�kū<1c�r�Z���W�moc�97`q�W������";&������Qn�.鼚|�i�nN0��̜K�I�,{hŜ��bi�RwK�-��nHB6�r3Xu����.u�J����Z�2��uӓ�ٮ�M�`\���Mm��rG�9��;:�Kb՞X�@�J�&e1*�`��N2q6wQ��Kı;�w�iȖ%�bw/}�ӑ2%�bw��g�"X�%����;k�tf��|��{��7���]��r�c�2%������bX�'{��p�r%�bX?{�4��bX��~?��bs,&`[U=���7��,N��q,K���{8m9ı,��Mı,K��}v��bX�����u����3/����d�>�}�6��bX����&�X�%���~�ND�,K�{���K�q��~�|�и闆�n���oq��%����I��%�b{�ߦӑ,K��^�17ı,O��g�"X����ߟTq�N�s�yX�t]\���������1m���v�P�Z�BpܪgZ�]K��I��%�b{�ߦӑ,K��^�17ı,O��g�"X�%����I��%�b^Ͻ��S2ff�[5��Z�ND�,K�{���8��0�(P�@�E�! ��05@l��i
)���Q�ț�bo��p�r%�bX?w�4��bX�'���m9ı,O��T��r=1�C/����oq��߿�^ND�,K�{6D�K����?{^�v��bX�'���bn%�bX���/��٣Z�֌��ND�,K�{6D�Kı=�w�iȖ%�bw/}���bX�'�ﳆӑ,K=��~�;k�u�]��7���%��뾻ND�,K����f'"X�%�����6��bX�'޾�Sq,x��{�������ڲ�p�:�n� m���r��[b�%l(u�<��X�c���\Kfj��MkZ�ND�,K�{���Kı>�}�6��bX�'޾�Sq,K��u�]�"X�%��{=uuuu��[�s4f�Y���%�b}��8m9ȡ��,N���T�Kı?{^�v��bX�'r�ى��%�b{��n��L�4Sw�w�{��7������7ı,Ow]��r%��""w/}���bX�'=�g�"X�{�����>�T�nHV���{��2X����Kı;���Mı,K�w��iȖ%�b}��7Ļ�oq���\?yr����|�7���%�ܾ�bn%�bX�{��ND�,K���Sq,K��u�]�"X���~w��4nKe��\�sX���9�:ݵn�^`�(�^��&Ţ氉u��{Y�]]]k17ı,O��g�"X�%��_l���%�b{��ӑ,K��_{17ı,K��d���lѬ�֍]f��"X�%��_l���%�b{��ӑ,K��_{17ı,O��g�"X�%���\��)5f�.kF��h���%�b{��ӑ,K��_{17ı,O��g�"X�%��_l���%�b{;�M]Y��r�\�Mf�6��bX�'r�ى��%�b}��8m9ı,N��eMı,dX�@�'�uȚ�s�������ow���%�<Y,��Y���%�b}��8m9ı,?�߯�9ı,O���M�"X�%�ܽ�bn%�bX�����5��֤3"�g6ٹ�]ѻ67s�b,�3�7A�\�]כ�{�ڀ���L�4Sw�w�{��7���}���X�%���~�ND�,K�{���NDȖ%�����6��b�ow���~�f�$+q�����,Ow���r%�bX���f&�X�%������Kı>��ʛ�b3�ϓ�̓��$���H�3���3�bX���f&�X�%������Kı>��ʛ�bX�'���m9Ǎ�7���}�������o%������Kı>��ʛ�bX�'���m9ı,N��q,KĿ�I}$�&�f��j�4m9ı,O�}���X�%��U����m>�bX�'���bn%�bX�{��ND�,K!�� �V�0!	�VG���|z"�HoP%�_^�!���aZ@5����P##!@�e�����?�<E�F� |��HG��h��P�Ě�{U� �v.��M# p)	�a�hF$X�����bh�p�Q$��n����K�#���FB0�B,"�bF		��#	��́��R+ ��X�%:IB�R@֚=1F�S�K���H�C����ȫD6�"�g��H�A��Ct�A_B2�HMx �#�H$CP�I$	�I�Џ��1 ��d�o�m��lT�zz�G��)Í�B�Z��8����t��C\�b#��MuU����m�@�ז�X`jۢ�,0I�i�٭6�	N����P;��Q٘V_='q).Z̪��1v6D���3�*�b+���tر���IqvAYb����t�˃sӳ�2Z�`s,��؂�T�r���4m�Ӵ��:N�$�ml`5�m��@z8���vf�-ˋwnӛJ-��Z3a���S2�����n��"m�����':0p����3����
�I��7v�rem΁]����g�٩V�)��h	ZX*�m*���vP�]�&��4���B��e�2-Tݝm�*�\����)C��I��m��<��nnK���˷S�ڔ��j�2���=v8g���v��KL�NP��l�����r�{�>7�"p���rl�˹hj1|���~d���=�ۋ��1�:��]��#=���T Pm������L��e� �	��
6��=`L�=��s|�˨x��&��vG�'d^y#M���r�(m��f�N�[eL�v�#l=l�;V��60g��0].�W��!/nN+��^M�ݱ�W\����<q]��]�5l	�]��0q�/����$D@pY��nF�;b'<��U�41��ٖ]N{X����C.�at��Χc��$�\�J���K0�r:Բ[����e����.�k.	���-m�Q�qm�I���:7;�rvX-'E���k.� z��.����3���p&L��^I%��pI�.: 'DX�rl�v"E�by����ɛi�s\A�)��.2��2cb,�kCW$T� ;-�H���:�#!��ۓ�y�=���Ҕ�B� ˢ�f�@m�Us���k���v�:ʴ� ���|���X7[s��q�fڥZqvh�j'l�6!A0�oZ�ki�r����u�rqs[����3�v���;UŞ`wS�\����LV��� :G�(�>Q�4�;@���ŉ���D�@x��Q5�X��"9T��ؚ7�!�R�`�.��togFL��^�;��sucK���d�l�֕���J��Wܑ<kn1�굎-g7Hy�q�c���g���zN6=j4i�����R�t��d,�ٖ7WL�����{ �]���s��1�˱n)�kѳ����x�Z^�df����[��Л8A�b�nڝ�����b5ױ�9�#^���=��s���^nx2۫t���'.�ñ���t����-0�Վѫu�\{�w���{����~�ND�,K�{���Kı>�}�6��bX�'޾�Sq,K�w���aR�ڨ���oq���X���f&���ș���~�ND�,K���7ı,Ow]��r%��ow���%�<Y,�������K����p�r%�bX�z�eMı���?{^�v��bX�'���bn)�&|����6��dm�9k�U�/�X�%����T�Kı=�w�iȖ%�bw/}���bX�'�ﳆӛ�oq���}�gl��[��n=�"X�%��뾻ND�,K�{���Kı>�}�6��bX�'޾�S���oq���}��s�i�el��릩]pmvv%�$+�LsXvJ�=;��d���^K�j\�ճZ����r%�bX���f&�X�%������Kı>�������,K����iȖ%�bw��R�e�"}�7���{��������rw�V
� � tw�,M��eMı,K�׽v��bX�'r�ى���r�D�:{�忬�dѣ5u�WY�iȖ%�bw�����X�%��뾻ND�,K�{���Kı>�}�6��bX�'ݺ���)2�j\֍��Sq,K��u�]�"X�%�ܽ�bn%�bX�{��ND�,�L����
��bX�'j����Bu��Q�����{��7��?>�&�X�%������Kı>��ʛ�bX�'����9ı,OL����]r�Rnx�:vP#;tnv��qn���M�t�q7iqD��fU��f&�X�%������Kı>��ʛ�bX�'����?(�&D�,Oe����Kı?~��۫MkY��j�Y�iȖ%�b}��7ı,Ow]��r%�bX���f&�X�%������O�&TȖ'��Y/�L�	��2�Z�7ı,O�׿]�"X�%�ܽ�bn%�C�R�ȝ﹜6��bX�'޾�Sq,Kľ�x��a���l֦\�ӑ,K?*�2&O{����bX�'{��p�r%�bX�z�eMı,��;��I����ٮ;A���;I-���/߻٤�E�H���?D�,K���m9ı,K;�kI��%�bt����Z'�[N��Í�z�.�Å�3۞.�=!κcO-8������ɵ�1]w�%�bw�����X�%����6��bX�'�{����DȖ%���������3�ϓ>]�zѢ2��URkEMı,K��m9��"dK������bX�'����iȖ%�b}��7�2%��ھ�5ue�n�j[�˚�r%�bX�wߵ��Kı;�}�6��c�"w��ʛ�bX�'{���r%�bX�g��Y���<�&""bb&e��d缙��#.��t�r%�bX���T�Kı>���ӑ,Kc$X2 *�����������kI��%�O��q��d�D��V|�&|��b}��7ı,?Ǻ�f��%�bY�~֓q,K����p�r!������O\E�17+��Y��.�l�ZKpl�=�n��&4���ww8����3Z�\�kY��"X�%���fӑ,Kĳ��ZMı,K�w��a�E�DȖ%��_�*n%�bX�N�G�E\�l�Wlϗ��ϓ>L�9�}�&����MD�?{��p�r%�bX���T�Kı>ϻ��r=�����;�ow���K�8��+i7ı,Ow߳�ӑ,K����*n%��dL���fӑ,K�9��,�d�'8�����A3�W3Fӑ,K?)"w��
��bX�'s���ND�,Kϻ�i7Ģ\�-��L�8��N2�y����kR�h�֊��bX�'��}�ND�,K�溞���'�,K������iȖ%�b}��7ı,O����;��~n�'X;Qi�ʇU+4q�9I��������N�H;6*�v�:;sN�ӑ��MͶ�if6�����]�[��k�]��8�����nۛ�ܼ>���:黆C�\��n
<����hm�	g��+#���lQ��OZ q�u�L��K��;�-����d�nF)��'j��#��1��d�7
�3s�����cojDg@��{��=�r|����g�2Vv��,uF��e�ˮq��/g���⃱綍0�X��̗��!s
�6u?D�,K��ߵ��Kı;�}�6��bX�'ݾ�C� ���&�X�'�߿�iȖ%�b{?�����5.5����f���Kı;�}�6����"dK���T�Kı;����r%�bX�}�kI��%�bs�ݷ�.�d4f�.kWZ�ND�,K��l���%�b}�wٴ�K�dL�g}�ZMı,K�����Kı;=��ڙn5�e�f��*n%�bX�g��m9ı,K>ﵤ�Kı;��8m9İ?L��_�*n%�bX����~DU�D�l�ٟ/�ɟ&|��g7mMı,K����߿��ӱ,K����l���%�b}�{ٴ�Kı<���뜱t��l,��p�N�v�����Ԓn]�E^RN��;H~��o�ۯ7*�%ֵ��Kı=�~�ND�,K���Sq,K��>��a�'�2%�bY�ߵ��Kı/���e�,�5�\ԙ�Ѵ�Kı;��7��� �����,Ng��6��bX�%���i7ı,N���ND�D_��������X우�\�ǻ��,K�����r%�bX7�{4��c�!�2'����iȖ%�b{��ʛ��{��7����tk����g绑,K?$����4��bX�'����iȖ%�bw��*n%�bX�g�������{��7���~��{2�M��n%�bX��}�6��bX��}���ND�,K��߳iȖ%�`߽��n%�bX��m����I���k0.��0��ޝt#v%����m��.Jt.�����pJ�ԫS7=���7���x���7ı,O��{6��bX����ᜉ�,K�����KǍ��߷'�{5�����{��7����ͧ!���-uQ,K=���&�X�%�������Kı;��0�y(�P�3���(�������]��,Kĳ��kI��%�bw��p�r%�	���6r&�{��ʛ�bX�'s���ND�,K���5�k]R�R�Z�n%�g������r%�bX������X�%��}�fӑ,K���:���i7ıL�yo�7��B�(K*ϗ��ϓ��o�T�Kİ��1���m>�bX���٤�Kı>����x��{��>���~�^�ӏ1<�r�m��lU��&7PDsp�u���;��3U��f�35��h���%�b}�{ٴ�Kİo��i7ı,O���l?
�>��,K޿�T�Kı;�_~���.�-3?=���7���w��߮�p�*���,N���ND�,K޿�T�Kı>Ͻ��r'�@9=�������f�؅ji��2X�%�����iȖ%�bw��*n%��Ta�2's��fӑ,K�����a�gɟ&|�oq��;$j�d�ǚѴ�K��@Ȟ��¦�X�%����ٴ�Kİo��i7İ>Ch	�(Q«9����i��7���{�7���h�nJf�{�d�,K���ͧ"X�%�~��I��%�b}���iȖ%�bw��*n)�N2q��$�Y�\�`reD0��=�G^H�{^�X: �ݸE���tv�h]�F
�����Ɋ<Q��i��]��.�&|��b����4��bX�'�{�6��bX�'{���2%�bw;��m9ı.�~}�]Z玛��M������D��{�Ӑ��r&D�=�ٲ&�X�%����ٴ�Kİo��i7��P�3嫾���J�*�U�/��ı,O{�l���%�b}�{ٴ�K��R���7��٤�Kı=����>_��>L�3��d�m+-$��5���X�~RD���m9ı,�߳I��%�b}���iȖ%�bw��*n%�bX�wW����ɗF���k5�ͧ"X�%�~��I��%�a�F=���O�X�%��_�*n%�bX�g��m9ı,N ����$�ޚ��vGʈ�r
[��q��q>6���[G�X���N��f����պ��ۭ���ʪ������ʘ�-��Ӊg`�!cJ�Y&�UFd�NV��i0�Rۏ$�d-�'�9��團�����u�ɱ��l��<7(\XI;n�[s\�v2�������ls�=����H�]���h���ۭ�s��l�q&$�4�&D�����aHNK�����U��c�ƺ]),pz�ݮ�b}s�+3���ɸ��z�Q�5�.Jpa�����>_>�8,�Mf��,K������ӑ,K��o�T�Kı>Ͻ��~Q'�2%�`����Mı,K��ݷ����M���eִm9ı,N��eM����,O���fӑ,K����4��Ͼ���9ͪ=�n"Z(�ڰϛ� ��أ�3'|��Tgu* ��拓�\M������O����;��,��J��$���4d�?��T'O2�0�T��Py��L�fw|��;������?�_s�o�,mUlm[�U���� �m��zU�Z]& �Q��s�sK5p�9���k�Gj�{�b�?>n�������ý�b��I=h�Yi%�Yj�>{݊�I�O���2dA���P��X9��=��6k���@�R��>wEw�J�2e�IDn�Ԩ}�����J���7I%�[0s�� �ݥ@|����3�(�w�*a8�vG,vՀs��X�ܝ���8��L����9޽pk �EuDȤ��,\ە���r;��W��#.��Y�'*Ժ]�}�|Z�WGS��;e���q�ޘ��ـs��_�K���{�ŀy���Y�e{����1 �EH�*@zܘ��%���*��kv'Uv���b�9��,�:'�Fh`|FL�X'���A�c8�V���l� �HN��G���F��"��D�IB,F$����$t��B 0! ���m.�p�HeH�ظ��L�a1P�REH�F��`IC���#c4s(���0�l���4E�@�E�f�+
$�A#`@Ƙb*�!)R!`!�`��4�a$bD�X)RVA�*R�� � ��.�<�]� �p Ҩ@S�
`U�#�/�;QjiLQ����#�� |�|����'o��܇;�r7T�v��U]� �7q`�6bۓ�T�;�fM���7L�ݭ��@zܘ�v��} �R��{������Um�D�@�����s;T���̖�+�8y;F��N�UfeM$D�LL|>wEw�J��ݥ�ɒ�Ï���8��d�q*���-�wEH�T���1 �Ɉ�K���8�vG,vՀs����wfI|��7��z`��X�ڍ���墎f&fU���P��fm*a&ho�sw��5�a&�B�2Ym� �䘀�� ܊��& ��,�)���)J�竗7&�1͔v��6�;�b����ibҺ�C�v�&�U֥U�0����nEH\�ܘ���F^���e�[{��nEH\�ܘ��{����&��VZYmVڰ�wq�rb���} 9�7w.�v�$V�,���>N�� ��b�9��X绳 ����8�����f��R� =rL@;rb���Ur�1U@�j/u$ߪ�P`��VoH�$5��9��N=���iJ��j*;�3ٱ;����6�6oTpf�M>;�����=����z;�Km����#r<�B>S�����Q�m�M��q�Ѫ�u��|��#ki��ju�n�:��'C���9�~����[z�ϤE�׉��@�jqX�1ʙD����^5�1N�r��-��ѪG��2溟�S���kP�˭HfL�3�6�uz����\g��n\M]+�E�F�s�շJ�v��UX�U�7,vՠo{�X绳 ����;��,��F���r�Gl�� =rL@;rb���r*@K�	5	���e����� �{��sw����:����'u�Uwq��R� =rL@;rb����C�%r��X9�� �9=�O�u�ޘ{�ŀo7�ω(�#��ol콋�e�V�0�̯G.�DA���7K`�٣KMT�YZ
�K-��V����8��0����~a��ذ�������I�����>�{ٺ�J��0h�L�o���R�/7Ԩ�wb���5�eޢ��9-�ـw��X9��|����0��� �v���⬱�c���&���H�����k'���P�U�,���E��V��v`|݈} �R ��]a[fn��ne�ܟ�`eo*	Pʜ��b���ͬ܈�/N�s���)-����E�d��g ׿�� �3iP{�����~ފ_��S�;�nm���� 9�T�nEH\�ovg�I6ot�A��t�Հw��lܓ���nm��)P� �I��\ɒ����(��Tf�Dl��e�����`������ �{��=�����ߖ s}=%�:ݕ�"��fo{�@s$ۻ�/���@|���o���.n��F��ج8)���'"N'Yo,�'n����.N[)��#4�S]���v&&b��ͥ@]�Ҡ>}ݏļ��+�׿�� ￨���⬱�e�����\ɒw-��(|�36���y�GS��;e����ـq�va�����b�;�{ n�6�&�,C%����fo&L�6wފ��J��ݥA��*���:� :�����}���k#��Ԫ�f��q`�/����~����8��0\҆�k���lF^y�SgZ�q"v	ݹ5�wWHs������}�K�ir��괤����w��R�$��& ;�*@wM̼��l�&&T���@|���$��L�4A���P��T��*�I�L����^&b���[]� ��0��� �7q`�������K����-�L�ɒ}����J���v(9�$��#���9���*�8�vG,�Հs���$�;�>;���ͥ@:d�J���7	�c�V5a�n�:UFm�X�h5�n�Xr�k�. n��u��6w�U\V\��ۭ2����T4�3���S���z𛱛��v�"q��nF��]v9��╸.3����Us6
ː�+�.�'F���5��ud��H6�'k���7�Ύ`H�cܼb��V�C-+6�F'sq�9�q����ns�@�i�uW+i������sb5g����{�ލ���>:��L���2��@uI��Y�9�V�ݎ�3ۦ�.�$lg��w��þ�J�����￱ �Ɉ} �R �,ٗxR�Ș�����b�$�y�2h���J����P>��s&L�^�?<���ejU]� ��`��,����8��0���Q��iITv�$����*߷����ؠ�o$�;{֨{�����Yie��-X�ـq�L@s� ܊�ߪ��g���̺��Xմ�@���r���٭��7C�c͸�x ���e�B4�6�z��������h��T��/%���1�ފ}�^d��\��&f&b��ͥV�L�k&I,ff�����T������W3�{�?B��n��ڰ�}� ���0�o����7��X�ڵ�(ʥ���e����;z(|�/6�3�o|���z�1�]M��e���ـowߗ�;��,����5�t�Q�k%���:�a8[ۇ+E���p�sa�#ţ��q��lՂ����ejU]� �7q`�wǽـ~|ݘ{�qGP�����76��T�w:b���9 ;�a&���Z��Հq�v`�7fLD} � ���w~ٹ'>�`9�\��[v�H��ـ~|ݘ^�*�6�$��;z(|�&"TL,��K�����9 � �t���ـo��ٌ��l�[�p	oi�;�V��2V�f�O@6���f��W7G�{�y�y�H�*@;�1�rb��ŀo6�r�[���v�-X�q]���;� � G,��Yy[�]�����[��T�o���f��z�cqYZ�Wl�;��T�m*�sb�R_JHdÉK2gd6'��!�J����ܓ���̺"u0L�D���@]�Ҡ<���%����}���n����h��N����O3�g��lW[&�Pj��:�R}��e3�*�)e��mX�f��v`��/��;��,���X嬡(��KlP=��rw7;�P�Ԩ}͊�L��}���u�r[e� ��ذs6�d�;���P��ٲlCʘO;�;���ʠ�&fO���1�z(��f��$�����w�y�n�kU�7wi �t��& 9�T�nEH�S�����j0$�eS���� �a��'�#�Gf(q�u!!$�!��1 Ē��D�@�B饬M28 �!��c�*�  �� `�1�BDFE�>%b�!FB0KhT:VAbAXD�֝ O!����"���	��G�$���� �`���O@��`֮�p�< ����!���4��~�mi�K%�H���M��Iq��@��c�v��;#�DYv��wF����ۄ���t�NKn� -��m��`N����m,BJ��:�5��C�yyƻt���UTS�
̽M�bN��V�s;s�cYȼH���d�5.y��WC6�PP�uHۨ^B�;2�c�pt�g��W��f��.Z�ۍs�k�Y=;`"�i���J��<��G��Ҷ�F�a�-*�ү[��#U+͗m���s���b$�$��� �A�V� @�W�Gl������l쭝�m��㠐*R�����@� 2�JK@J��rݝ(	��e��m���6����-ʵW6�niS)h6n��)C��Ϛ�/l:����M;	���sjYX���p[H�[��s���7�	�G� qIb�s�����nq�c�ƈ�̔�ڴ�.^����9�	�\"�<�=dOI��bM�v�sO</g!:����v��%�r�����v�k+�l��T)��vGk�6�ܕTGcY�n-�;Sd�u�xzò��
�2�e(-�� Wm����y7n��cS�;��*�;V�8�3�KW *�Le�:�ј�K��l���	��C���i�vy�d|ݍ��IŞr����]�Tt���X-�5ܰ@�ڳg����۷-��Ps�v67N�mX9qb:"���N��V�im���#��b��u�;ظ�5���#���^{\vu���,��[;���
�ݣI����V�V^�d��r�b��٩�� 9"�� ^͑gZ٠Û�y��M����p�n#:{=�{�5���9�6� ��x�s���VNd�����;b�Uv��P�)��L�j�FU� ��Uv��������g�0�㱦�FD�j�Y��We�U�������ӭl	y�mp��\�Ln�L s�g\���:�]����]!����8esN�u�u��[u�Y�Y���@M
��p"�/��)�v�� �ۣ���o>�,�L��0���h�'=\�u�v:��4oF�#��;T���ut���t8�ԅ͘��\]����9�ۻm�%�[����F�tv�m�C�v5��+A%�oF���=*���%�x�q�6�c<l��Sv6.�9]�<;ց7]�çq��m�n$���:�Rm�(;N�j.��؉��j�Vz;u�;u:{	����6�:�K<���6��R�����q�;���9�jrR&�i�m:;r<��<��]�j�[���ש��Ӂ�������7�1�U�7,�Y�y�0� �7qy%�_�q�}0=��l#��)Uv�/6�w�J���6({݊�32�_|�7��P�����;V���� �Θ�v��>��M��~���M��*bePs2I�;z(|�/6������{��<�vz�-e	D�Q�f �Ɉ} �R�:bX���~��t�H5÷n����<f&��
�����尼�u%ݚ0a�{���ϟ06���՛��'O� �R�:bۓ���I[v7,vՀs����KA�$̟̐����;�@[�tP{���&��~<�"��]��V����-�v(�$��J���@z�̸���ڻ3sw7ܘ��"�r*A���=����8��;��f�nҠ9�;�_���@[��Pl-؈s�:�C�ћ{v.�(n�m��̠�q�V.��v��tn���,��P���W*�U�s���}͊��cɒf^W��R�=�K�}F�V�VZ�=����� �7q`��,�l�{��9k(J'"��Y�'o~��;���s��Ġ��X��XP���z�훐��v`�7F�u�r[e��/���v�֨�z�o��@[��Pfɲ:�RV;#�9j�9��X�=�����0�w���<���'+�n�u�NOM�gp�ٸ�lp�n��E�_���|�\+�|Elv�m_����`|ݘy������ŀ��F�j,�����b�;��Ԩ��T���~2M�{��TDV�R����ŀ]�ң�N���>wEy���'��4��si ܊��L@;rb�"��BBFŁ,"�D ���Ty��nI�{E��ӊ�b��V�{� ����7{��sw����wI$����〪�����"�1�	���Ax��v2�������ݪq�lBQ9v��5����7{��sw�{� ���9+,Q�Q�m�1@n�ү$�gs3�����@[��`���V)+���`��,^�f���ޘ��ŀǺܷ�+a[{���H	s� �1'EH�K ;α���,�Y�q�v`���36h}͊Y��3!�����q�ɨ-������;�$�Aj����LDl݁nw5
+Wn�.�u[b��L�nmX���@���F��W:�n0vPl1���\v��
��1�K8Zer���t���@s�ny�#ÑŖ���"C�e����q�x���y|mOHc c�il�"�
F���Yt˩�囊��Yt��ݸƌV���p٣[`�C�n�f��f��'?8s|�&���\뗋v�q+v�1͝à�R��+N�U9��1t▷eD%n�*���w}� 33f�����^fW��z(�ީ"	�ejXYV w�۟��l���`~�w6�y�3��ҝ���LDy�@}O��rb;���k@���8�C�$M��y$��7f��b�s�p{ݘ7G%e�:�I-�ـn�q`K��w��~�L����7��2�`�AXح	@��W�����<�=;]���t�:��7�"k��-�ӢQ���Tw�4������y3%�2�{�J�=��;���`R�*&&h}͊�d�RI%[���m* �͚�_���@�������XG,�Y�u��� $� 7�P�L@;�MͣDK���&"b��&f~�� foM�{� ���0p��MD겵,,��.�f���$�;z>�;���ͥF�{����}��^��gb�����h�C�^s���H��-�f�,a� =,������@|���m.fL��;���l�$�G\$M�f��vW�2N�v�* �ޚ_sb����2M׿�Ò��U$��l�?���� 9�}��pX�E����8��k�l�:�v`���J�,����L�fI3�f�����{�@n�����]�B;`��K-�5�v`�̕�wG�woR��٠1nk�>��K<'��#��>Y.$9}�+J�vu��Kaӛ���LR+���4�f��m����E��J�.�g�&e�?oE��tʈ
J�NR�f��ş�_|�a�呂���>{݊��ɼ�I��ީ����VV���`￮�{� ���0��,��c�~u�k�Z�m��L�'���-�(��T�bd$��*�X�D���	�k�r�ܞQ�*b"������P��ɻ�ߗ�;��,^�f��V¦�R��ӵ��I�29����zglM��un8�8m�8�y�-���+���$�Kf��ŀs���}͎I���p���/zNO�K+n��rZ�s�� ׽ـ~|ݘ�m*�$�/2d�(����L�"e�/3*�����{�G�d�ݽJ���`|�Ѧ�d�r�e��}�I��gtP�Ԩ��Td̟����Ǿ󲢂r��)d� ����=��|��$�[��V���>{݊�5�% ��W߉�^je��hִf���v3���Zz��:¬ܦ�ػ���㤝y5�9̻.F�d"�C��goT�;��I���.��ۨy�s��Kv٥�cvnN���ڃIv���E�l�;)c�ke���c�N�M��z��Z�r���7qFs��\g��%��#���TnSi��L�����nMq�����C�{��ƥ8y�P�lE��͞F���{����w������["��r�g��I��5��B.ld��Ș���en�,4�V�+�x��uĬs�����@|��d�&����b�;���{�[v�ը��^��y&d�[�tP�Ԩ��U�ɓ;����%�Q�$M�f��z`��H�*@;�1 ��y��w�w{Z^f��� 9ȩ �EHs� ���U��z`�S�ʝ�Xݍ�$�`�w)�:b���N���{w+rvz�.7)�vn�Ҁ�<MR�n�$�n�NZ�i#mO��ޕZ�Y:2�S1ߒIO��rb�EH�*@K}��K�f\�sY�f�rN_���)�Т@� �EW�%�ək73$���w�P�Ԩ}͊�K�g^��ʬB��Ӕ�Y�o�ذ��Ty�N����wE�nҘ�'N�+R�eX9�ŀu�v`�7f��&�&��z��z^#�'!ɘ�S(��@c��PL����J��ͥA������N��vi�Vk�6�n�����\�:�%�Ҽ�v<ۊa,���u��Ͳ&�fU�n�w�}�:*@7�R�͘7\���c��Kl�`��,�fK���z�Ͼ�P=�����J����nY%� �;���n�?}��R!��"v X��4�B�����ǂ�� �� @J�4X�Rх�����/b��#�k�5쩝D"|t��R,J&1XX� ���h�1H}������E���_���6�m�8qv�
�2d�Uʰ�ejf���Eă b$4�yD>��yW�)� �U:��!6� �? ���:*:ɗ]�nI�}훒O}}�.��u/3*��ɓ7�QӾ�Ps��tT�o����^J�/v��!�b^f(��b��d��f�w�X��� ����8-�J�K��	F���^yn�F�[�:��H�-ۏs�Vhj�
��NR�f����9��,����%��}�oO{)"N�+R�f����ܘ���1 ܊�������$�+-��Q-X_}�~|����6=���6 �666=�p؃� � � � ��{%�f�ˬ�u��[��lA�lll~����y���y�߸lA�ll"q�"(�`����.���g��6 �666?g�~����̲����k3Z͈<����{���<����{��6 �666=����y���f�A����w����������m%,T�#�̄id�0�]u8�nd���S�v�h~{���vhֵ3Yn���\֍�?A�������b �`�`�`����ٱ�A�A�A�A�;��lA�lll{�߸lA�l=��w��n�w����ߴm���L�|y�~͈<�-�����߳b �`�`�`�����b �`�`�`�����<���0r9���K��-ֳ.f\�j�Y��A�A�A�A�{��6 �666=���6 �6
66=�p؃� � � � �;��lA�lllzg�~���5isSY�͈<���� Q2>�����A�������b �`�`�`����ٱ�A�A��A�;��lA�lll}���p�!�Ѭ�3F��6 �666=�p؃� � � ء���_k��ٱ� � � � �=���y���y��h"�)c'����r��ꛚ�C������3���i�Ɲ!���k�H�7G��j�NK�9:��M����q�« �hh�ձ�ϧd@��d:�-1q]:v#�!�tv�s�t����V���+u�Xm�Ո7 ���9���-��<m�-n�d��t:K=y�[��:rN��C�4�q%��m��	�g�N)B��j�r�57���k����d��lPk�4Y��L�F�jR�M3V���g�u.�n���r�=z<��wkj���5.oP�VkW)�Zѱ�A�A�A�A�;���y���f�A��������A������ywx�����������3�H����<������߳b �`�`�`�����b �`�`�`�����<����s��f�@S� �����}~���$�b�+KO��w����������A�A�A�A�}���A�� �r>���ٱ�A�A�A�A�{��6 �666?{���f�f��[��5�5�b �`�b�X ����b �`�`�`����ٱ�A�A�A�A�;��lA�lll}�߸lA�lX�K�/��������ڎ�e��<����s��f�A���U�;��lA�lll}�߸lA�lll{�~��A�A�A�A�C��3~�<h�p^t�S��8y��z��vkr���oS�E�����8n8)ʃ4���w�$�&I�L�8��;��7;�Py��=������P���Yd� �����AF|"�Q�"�? ̏��T�oE���Pf�R�Dʘ�Q*f%P{��{݊9�3'|~�� �}�X:mrm#-q�Q-X|��;���ݥA�&|���ݍ�J�!c�[0>n���gw��3;�P�����#\�1��n�p\;]N�^��"4B³Ɗ�^ c���&�уUL
b�+KOͷ��������*��c̙$�p���/:C������ܱ�V�n��8��0>n���Ş_%�M����e���v��ʠ1�({݊&d�����*��ŀk���M7l$��+�`y%��>FwE��J��ݥA�&O���@q�\��	��%�K0sw�Lٝ�/����-�v(L��V�D8��#p۰�F�^�Ȇ�	�]�OC��t���;�l�S����F~?9{;Lsu7pI��� �ɈnL@7"�pM��Zdv�ը�����<�K�g_}�3;�P{��ɓ3;�����$%��Ɉ�N�3>wEw�J�3&I;�wb�:��L����܍�D�Kfw�J��ݥ@[��P[4$ɡ�fd�D>U�� y��w���o;CШ�K[��c����ŀ%�M��������*��������F����q�&�睞����ʸ�d�g=Z��E���.L�en�m v���[j����`����/&ff_��5�n�Ԩ>�7?�c��F��0>n���ŀ]�Ҡ-�v*ٹ&ewC�A
"<e�f���ʐ�ց��v >�& 9����`겵*�U�s���>n�����|�{�~X�o��Z���U�3v�ܘ�v��r*@7"�}��﷚7��v,����B(!q��p{@p[��7�z�%N�y�ӝg#�&My�z�+=WI ps��̘ڬ���!5zc��j�����&j���H� i��t�v��\�KVdླྀU�I�*+�.��n� ��>��Pk;��=xE�sz�m�p�����[�\[)����񙓃�ݑzzt�kt��X��lm���㭭q�9.���8�e_����D�+*=vN�l�����NF�n�Iш9)��}���!�h��/a����}�b� � �ɈnL�sn�,�ҳ3w3wȩ �EHnL@~|ݙ��&�w�=
�T�u�,rʠ37�P��y�'{|�3�� }��1.̻�y���T��y��(ݟ�؀�?�� ܊�ȩ-̻�FU�闖f��� �1 ܊�ȫ �����wc
�bVV
;��� ����q�T��O\�huZ\߽����f;kn�[\%�K?��ذsw��ـq�v`���\M��aIU��rO���o���W�#�w�^g��}�s����7�͵�Gn��h��@;rb���r*@7ҕ�y�D�3�D!�f(<�ɼ���;�E��R�.�iP�������̊"&b&b��ݥ@y�fo2Lͻ޵`k��{�@nn��K��ΐ�Y�&�^rj-�x�"�.$����:ۣ��+�ۛ�v"k����ͳp25�6�����HnL@zܘ�nEH;�w��kj;e���{�<�K�8��L{�b�9��X�lnj"v�8�e���>�{ٹ'~��n(t#� 8����1A��~Uy���6��z�o��P۰l̎����&&"b�����*3��o��@[�v`���\M��aIU����ŀs3$�d�6ϻ�`k�^�*Z����rW*�Wd(\k�p\C6��ќ.��\u�[�h��,
5�٥P�������K�&K���T�v?BP��Y#��l�8��3�|����Tgu*��b�2L��oB���v�Il�����`��,?�_|�}}����z`���,T�*nX�2���T���o{�AlɢS	E!��	Ah�C��ߺ��zܞV(�ڰ>n�ۓȩ ܊���eR�sk3p�	�7|��	����獰�l�����u����і3��vx��������??_�k��T�m/$�|Ꮭ�@��x�����������T�o���& ?>n��_6oM�*�n�:J��`���& =nL@7"�v]̹�0΢G�2��T���3�(|��w�����,ϻ=	(7a,������Ɉ�T�o���& 5��hO���`��*��m	u�D2U"V)UF-"	�<��D$�I1C�E:l@ٶ� ��ǊaE Nw���(��)F)��@�+ƽV	^I�B2d��h`E)������4F��0`D"�Z�$9,������B �*w1RDp"X@bXXP 0!eWr�¸�1�Bh�Sh� ��̈́a!1VY"w��O��kZִj�:���N�q��3�إg�c,�RU�k�����%��$�n�₭�ڭ����Y�nt]�� �%Z���j��^ZUPx��*��Oi{i��5l�s�5;+ZUUp����'���hBQѦ�M�N�݂NQ7\N�XL����ӻR�L�8����Clh��K�������n�H��]�3)q��\9��{=���.�c����7W"����X��u+iUR@�,�ڐm��cM";�Ʉu�v�Yp2O �N�T l��A�������<���gێ�*U��g���� 4ږ
VvS��scu����ʛE<A��e�V���k��d1b�i���Nƹ�*�Yn6����p���9�VO]�2S��7k�yɮ�w]�f�P6�wOLg��x�М�LY��F8��<��m�(��b�=;O�q�F`��mzs=��7�-
h���:K^��)��ҝ[�#�K���
nmp{wK���k0ݢś�Z�nԍ=�m��N:��mO:��qXl�(�VMڋ��e��N*P��HlKv�Bݭ/.���ptq��k�jx{= �mAMY�n^�˶�\����.�l�(ݜK�3Q1�5���J�۴��G�����Wp�S4guJ�n{����k�4T]� �.6.Er�'dݪi�v-�tȷ����� �����.��6p��<Cs��9�i ���m�I���sϭ�s�g�0a�-�s������ɶ۴��k��=��e�`����dIY�&Nk��e�mTU�³�h:M���:ۇ^Y��lٲZ�iWn���[al�����s��^��z��34�ع��nL6%Hb�R���em]�Sm�!���j�ֲ� u�l�8�cm�g��݌Ҧ(x�g���Kָ��v�!#���)�uɸ�D�wl��+�]�acWe�Xk6�r��]86�z���U{tLB�X-��u���h!����h+�eS��=(�E�B	�v��Q��1�<�7��"��a�2V���f�I��fۛq�A;vベ�\�\¼�����l�l�u�cg�;z�˚LQ���s�x88���3�ɑ8&lؼ9�#��`�7m"�rlX[���ަ��v��@�v�J\U�;s��3d6�v��G����`g+�b��G�&�w%�V��=�5��#��QG�T�mf�v��{3]N�r�6�bٕ}��&\��Ej���Y&��ɣ�rd�Y�]���t7I���&Ƅ�q�d�۬a�T������;E$�Kf�wq`y��{ݏ7�5�c�o�=�5ET��c����ŀq�v`|ݘ9��<�{���������V����& �R� %��y(�ڬ��ev��ϳ���;�{�ݥA�L�� ����f^����r*@7"��& �1+�:ݾ�3�<��'5��=�O�2����9������en��ز���+�U��&n�"W�fwR�-�v({ݏ$�7��԰�ߣ��|ԣ��KV��ً~��؜A��Cs��{7$�훒}�����$��ݞ�����n[0���@7"�r*@;rb�:en����{�ff�f� �R���ܘ����|�������aj��Sr�-H�*@;rb���r*@W�߿%�	��YYm���#"�*���:�)��̹��6���\t݂$�ҥ���@�6�
�����`K��؀��1 ܊��ŀk���'jv�+�`�7f ܊��T�v���밮�fiwy�f^����3��w�J�fI8�	�*�	�_��ܓ���nI�z]#�i�Ib�[*����O��~X���ؠ���;�T���3�%��F�� nM@zܘ�nEH�b�;��ƫY�-�}[e�4!�x3��kY]�yz3jD��y���,�����.io(����Ɉ�T�o���W�X���:����c���I-�ـs����$�foR���>{݊���p�!J�N�0�2���Tw�4rL���}�w��, �=nMV(�L���b���v(��T�2_33%�#�6>���9~�[�&Z.�[��{����1 ܊�ȩ �Ɉ�}ߟN�sr�p��f�����-��]�m�ٍ�<2<�zZ�h�K�S`T9���@7"�} �1�rb���:�C��)U������|�:���wEw�J�&L��sz:&fS�%*e2�|��أ�&I�3���`ν�Z�,$�H����ؠ.�iPy��9�&|����+
�c�RKd�`��,�����c�tP=��)�S2Q��,��
�Y�y$�UH��zu,�r�uN��H�K0Νͳ�tݹ�f<�Ս�
�m���2�(Hi�f�f�/U�xϱ����v��gk�����O�l�g�w%�rlp��������gB\w����w�$�.:�� o7s�h�n;q�GGm�D���Wf��0�H����-x㹳��۰���[&�z�rՖGr�T���#H6���z,��j)b�Ӈ ʱ�v$��.t���<�;-��O<�왅v����S��c����{ذ>n�����9��X�z����Ym �1�rb� �-�nj"r���ev�����9��X9�ŀq�v`�V5>��K,� �R���ܘ���1 ���h4;Ib�[*�9��,��g���}���n��;�ulM��9T��c	Aͥ���(M�˻��&#B����;�8�Ev$�[jh��QmX�f��v`{���p�ޥ@vk�2��Q2��ֳrN_����*��1T�����*@;�1 �t�ܻ��(���l�;��X9�Ň�_7����8��L�v���'J�M��`�T�w:b���9 �^f@@� ��bbeP��33\gt|��ŀs��X�\ֈjJ����s-:;u�������6�:�7H�f��8��nYl� ���0�w�wq`{ݘúm�N��K,�P{�������ޥ@c��P=��ޮ���K��V�wq`{��͛"�GB�0H�>��3p;��,��f�mQ�Uj-��%��>�b�}� 9ȩ �EH�{r�ʤ��� ���0�w�wq`{ݘ����dC�Tu�H�wcg\]���b�9n71��أXu���h����|�s���C�RKd�~{�b�9��,�{� ���0��+�U:��&Uw�J�s&�މ�;����W���=�M�Q�,�`���zܘ��"�} %���*�M��bf&(937�'}�;}�T�m*_Pg�`  ���s7$��׶8
��,�Y�w���s�� ��ؠ>{݊���һ�!�!��/.r��ۡ�ն���c�Xۜuu��Vܽ/8�"򥦿�}��`X�X�Vʸ￱`���& 9ȩ��2nn�^�����Hs� =nL@s�R�����=���ڣ��Z�C������9ȩ �EHs� Ι�Y�nQy�ff�f� 9ȩ �EHs� ���/�'}�s}OI`5b��ܱ�V ܊��L@;rb�������o���"��yR�a����md��g^{6�F�2�\8�V���=q������j�s�v�N�k��v�ulr�Q��۲�:�b1s-���m����6�����⧀5���#���ͬ���N�Lt��w,�Z�n:��l�u�6y��s�j��d[�9B�����W,�1��O;\��y�wl��'	���&)����O���v>(����=���{�?!�8m����M�]"��=n3�Zn)x�ju�b8Y��E�*��2e��$��X(�ڿ����@[��P{��Fd�/ђMp��*����8���nYl� ����;��X9�� �����k����K&"b��ݥ@]�ң̙$�̙�F��рk���w��B�hv��*�U�qȩ �t��& 9ȩ��2nnʅ)�T�"eP������fKg}�;}�T��*mF���.<Jx y݇l/\՝�%A=J�\��B�'kKѬ�h�ө�]v��$��� ����;͊�ȩ �t��tͭ��2��+35��k7$�����vE����@ę&V̓%R�s34a��R�-�(|ݙ��K����=%�ՔM��`�Ԩ}͊9���w���7;�P��j\�Q�-�`/�ϳ���:�� ܊�ȩ-̼�W�y��e�����nL@7�R� =nI�\�ѫJEVV
V;Y�n 1Ѻ�m��sG�O^sC�����wx��|]9M[\%�K?��`��,����8��0uv�X�+R��X9���rbۓ�T������/���mD*r�Q-X}�q�va��s��T�Ǥ�H��G-֘B]&.���A�����`�B�(ݚ��Rakd
3�Քs�|e |���05)j؄`����	�n��̡C�)(����l�(J� Im�Kj7�\�IL���8� ���L��"b�MemaB1��#B%�\�pd@��������&�y�j����IBRRV%Xā�C2��*J��j�	-��H{*8Ё665��Z��Y�� �\���F	H(��$� �"���|&���$P>b�tD�(�O���ffi�ϩP����u��T<��y&"G�����b��ͥ@]�Ҡ�ə����8���Y)"��[%� �;����T�{�@[��PI3%����ۋ�6�M��Z���Ppsn�C��X�f؞�:�t��sq*�6&4��7%]��Ԩ��b�����ffe�f�* �}$~�Er�Gl�Հ~|ݘ$�} �R_L��W����ydLK��o{�@]�ң�32N��Ԩ>�� :sv�ZDյ�Yd��%�g���P�Ԩ��b�Z3!�JY��_oٿ��L�Wn���uWZ�Wj�.�iP����d����@]�Ҡ�}��X�i�ʫgE
c5ӌ��wT��8��\u�;RF��,lc6\:gnћ����1 �Ɉ�*@7"��n�2��$-nV�`|ݙ��_|�L�Mn��P��*�ؠ>}͉N��M�)%�[0s�� �7qa���&���L����;��n��UJ��fU�fL���*�;����ؠ.�q`ͮ9���Q�-�`�7f�l��ޥ@]�Ҡei��3;����nz�L�u�2�f��˗E�.5g���M�ݳ�{n�����t���5�J��;m�Y��Zxۇ1�uQ��Kcu�Xzsq���;��2�5;^ms���\唅YΧ���u#��t���ǎ�Z�3œbq�<�p煽��3��<�����R@ �=h��
���2�z�Ӯ5+��Ns��k��2�Y�oo��
��Ut�$���-�+��Ē��,��|��>ǻ���k���U�u����e.9�V�᧫`�ۧ�UΘ��Qn5"fbf4}ފ�6�w�K�f_8[�t`����&���%�9�ŀq�T���1�rb�v������u��Uw�J���v(䙒w���;��, �vk����QmX��}o;� ���T�o���%b�;	�r�0ϛ� ��%��wߗ�;��,����7���G+ Z��ɱYx��th�)۷&�G#�T��ӻ6�h��hi�eM�8��RKd�`�w�wq`�7g��}������+,MU*nYu��}�}�t�A*�<
��$��c�tP���m*oeȍ7���e� ���0ϛ���7��`������Z됖Wl��əy$ѓ��P��T�m*�ـ7V�%U5mp�Y,�9��,����& =nL@J�(�m�f�s�I���M><#��y/<t�vb��Y[�-����W0,��v)Uv��w��X�{�@|��f��3z� f�s���.�(�S(��@|���̙;���f�*�6�rL�fh�7ǔT�b �x�&f(}����ͥD��ؓ�$��Ҋ�����{���;}�ٹ'���hn��ܢ�[%� �;��s�� ���0ϛ� �7q�+,MU*nX��ͥ@y��;��-�(��T�w���7��'�LN����њ\�e%kM=��y*��3Ze[n���Kssv����@zܘ�o��} 5�c�\q�,q�����ٞ�$��Q�z��ޥ@m�kגfw;�<�UN��K,�`���wq`��x��ـoWn���v��*�Ձ�̒e��ѻ޵@{c���{�AL�(�PH� �U�ލ ���D��5�rI�w=sZֵlyDJ�D̪n3^��%q����Ԩs�� �{�#���-�
���c�n���]2��ח�4J���65�D����W�~H�9�������7��X9�ŀo'u�{ݕ���ܤ$�KfEH�*@G�-�rb���ee���M��`��,y;��L��(�}������Pq��]���� #Ζ�v��} ����>����=�~����+�W�q�v(d�y&^���wޥ@m�k��j$A� �
"���|b��*�P�V7,E��4�=��>65�H�A�$�W:D#�r-Y�D"�lީ^4������Cx9ώ7T�8*�b�#����@�=Nͳ�7'3ś��9J{*��`��Y2%6
W� z�lsټ-�V.���^1�mj%�(=u��^�tUp�L�c�y�f��I=q�\ۜl<��ې�{��>�}�׮�:�6Y������#^�o{���r���nQ�];S*��.�m*J��t����Iu��g^ޔ35���-lZ�3,��~}��|��v����fK�|��l�LC��)Uv���ş�M�}����z`�w s�5�j����j%� ��1 �Ɉ� �R9R̨�9$���0>n�����9��,����8��+���\$�Kb�EH�*@z�L@zܘ�#%���4��NQ�]�G���H��4�VV,��<�\W���3KD�������@7�R��b��Ϫ��'ʐ��h��	�e������W�I2��|���ͥ@]�ү$�;��ѿRBJ�q���}�s��X|�}��Ǿ���]�,��[!,���$���*3z����Prf{��L���,�i,R�ڰs�� ��v(��b��ͥ@rfI6���C��-tk\e��t��&{����v��\��^�L�=SU?w�7��+�q�w�$�o���@zܘ�}�S�X>�Zr��h�9$���0ϝt��q`��,����/�l���V;GTN�%�[0��T�m*5��	$$�̄�	E\C�GYo��ܓ��{7$����,,MU*nYe� �;��ϻ� ���L�M�Q�޵@{}.?���%��3*���v(3+��ޥ@s��X�s\�B�FB�@�W��D[�&G��)�t�����Ok5�56��e˷�yfnm�����} � ~�����%vV�%q;,�`�wy�L�foR���>{݊�d���S|���K��V��`�n�����9��, �vm��jn���Y�A�fg{��-�(��Td��b@�� �E�� *`�W�E�I$�w�X���2���9jy�����1 �EH�*@rj ���f�!Ъ0�%R1�T�3k V��Ʋ!g���^y{\h��`���`]���@7�R�������ꪪx���`���vKUJ��;j�9��R �P�& �K��v��M�,�`�n�������}����`�`��I+q�Kk���& � �EH�M@.\ܬݻ�/o*�73q �EH�*@rkrN_��ܓ�bp��ŨJ�1�)�C�"@�YD��X��
��� ��	P��@�@�P�5� 1��"bȐ�0�##b�`�A`E�%��%Xҕ"��!P�V0%���XQ�0$�!�0���+
�"@�"ƌ��1!V6��<��
�
+���I�5��!�Th�4X� �a
@"T��$A$BxH�+d�{��}:wߧ��[y�.�*�$�|�mt���-] �t��$6��nSs{vi"@9�wp����$7!�ֵ�l�f�U�XamQ��U��@�	��#҇R�WPs�������Z���V�هnj��iϧ��C��A	�U��r��<�r��o�_#�܂=��fF�ٝ�Ŕr9�6{]�=sۛ]�)����Nq;+'6�l��<��ҧ�=��uMj����m��i����iٕRUl�R�F4O%�f�����`vLٮ��(#Y��W�*������J������鮰BqIwPZ-�v����鴈,@P������4�Ϝ�ϐܦԝ�lm0P
�U�[P
�qc�8�����2�@��
�v ��d�\a�uU�m�z��'��s���~z>|��m�\۷P��Ku��X:H�c�k���Їc�M�W�C����sq�FO*\�K��P��rE���5N{ ִ�S%Pö��Gj��5�eN7]���;i�1"��gO+]	�V��Rqڲ�n�g^ƫ���ˇ�
���p����V%T 8�nu�\ϟ+��1C�pv l���y-��6���Y�=���+�r#��:�Y�Ogs[t��<�j0p�ymʆpiC90Hs��]JY=�uP���t�YD��:�KU7=����2lr��:8�,���Y�K&�.	 ���ڲ)�e|�s�Oo������X�g��"�+um�K�Ѹ�q� 1�gJ)���vI� f��7`�@�(td��Z��Z�ٶ�<�<Hl+�M6�:k���n���s��(�u�tF�r�Y6��.^�-����[�������1�L:_Q��@�˫�#�n�&�օB�+km�1��Jm�� &�� ����dl��>6������ �D�1Td�S&���IH[Pclޛ���2\�\�v�An�@/Y-P�q[�^J;Y���-�F.zh)v�vu��nEHX�[������������_/� ����\*��G�T?/���@�./Q������p%�V�y�lUz��I�4ӳ��^:�[X�z\hy��<:{+�QMv��7e��	UkJَձ˳Am9#x܃�=�Z����]�=�S�W']��q5F�C�n�6H�"��$�e�ҕ�@~�nv��KC&廛�H�rƊ�x��qmպqH1P+k�&�v��˛�n��Hn|��皜��7P<^��]�{��=�wx^�++��j�{`ޮ7V��ugv3�^7V�;\nkĽ�n��fP�����1e�X�X�Uڼ���ʐ�����c�=뻷}b����6K�q��ڿ~m���Sm����r�~���ݶ߾�s��� ֵ}��]Qi"�����o����ͷ������_)'{���~m���Sm�ov[-��T��m��ߛo�w��|�w�����{�Lm�/��r�ޟ�6޿{���J��9j��o���_�6���/��S�m�N��������1���u���P$Y5ͺ�8ٷ���8���%�b8N��E�/��|~Z�(6\N�k�����ߖ� '7g�ͷǻ�cm�s��~��{'a&���[�2f���jn�o3�{9����� �D�?�T~Ϯ���f������9m�����?��@��~����<L��� u�ئ6��;���Ͷ���cm�ӛ������u}4�8+3���������������}��z��ww�/v>���̚2;�QN�ow�zK�������ߛm������7g�ͷǻ�cm�s��~��{�TG�0�Ü�5�.����ˮV�g��0�C�=/F��u��B^�0�	���g��s�����f���}��('{����� _�������0-M?������3�䔑��}�~��{7�m��sv~��}{��0��r�-Sm��r�{���nއ�ax1@+"DFʰx*h ������8�|~�)����F���7l����o�%����Lm���z~��|{��6��;���ͷ�vj��W$���i���N{��[o��s���m��p�-���ާ� ���ϯZ�#ӛc�.s9� �Gn��8��N��vJ�=y�h�7��	�O���d��g8�}~�)��������m��r��o��������n��4ݤ�J���]��}=^��~�̻���}� �& s��b�n"�j,� ���,�����|����`��6T�l�$Lʉ��A�d�q��@[��Py��J�;R"�G_{��ܓ���kZִ5UR�%�[0Ͻـ}�{�����b�?>n���oe��%alq�+>s�\p=oZ^�rDʃ`����okA�
qD�nXnE���� ����rL ����7�[�@$�n�e� �3iW�ܷ����.�iW����	<�r��[]� ��0�{���{�ŀswذu�Gc�6K.f� �t�} =� =nL@:٬؄�v��*�Y�s��X��sw�_o��@|���d�,fZH��"�53���r=�\��hf�pmѩM�=S�.���]��n�l���v<��y\�{dN.LfͶ�
!4ݤ�i�&����1SJl���]��;V�6,6��+�Ǘs�8-�q�lllE�;3X#6�ͥ�e�4g�`�1�dܲ�^VS\��/#�ۮ��H��dv��񙓷N�d9����y���4�1�&�.�0���u�S�Snh�3�˭K���D.{E#��\�7�7G+vr�k]�:䭤{bkm�Ge�Jۨ�Z�*�����1�o��t�ɛW[��i�2�feP=��~3/��c�z(��*�{���}�ɳ���-�UT��m��ܟb����& �K�,,aaP�[0s�� ���,���Prd�&^I��'��@{c�<��7l�Հ~�w��v`�{� �;��[�ϵ����[Z�YVVT.�e�ͺ�����2�]�z�C�4�Y�+��f���x}�؀��L@7�R��ŀײ=�I[l�Y,�?>�f`(�xD?�G{���lܓ�{���~|ݘ�f�&���)U����Ҡ>��T~&ffw������b6!���(�3(��A�3=��ʀ����ݸ9�ŀw�d�SR�%-�f�� =nL@o�������8�s�%�.��\�H,�d۞�.۶ʹ�I�.�ٷ�V�䉫5.:�`bfbf(�͚�6��f���fk�ǿ�� ��;%�",*������@{�*@;rb �t�y33 U޹`��[j�?w�� ���¥��H��^�� �<��J/�7�]��s�� ����QIk#���j��_'��}�Ͼ�r*@>� t��%]�y�wvf��n t���"�{ݘW"[����U$��B�S=�t���#�`)Nx�M�/�+x:F����޻���4ݤ�KKm��}� �{���{� ?wv�zl�#L"���Հw�*@z�L@�5Ϣ�t�ɛV�d���m�`��f ~���;��,����8��촃UU+r[m� >�٠2�iPy��)�0�d$7̝�c!#*2�,�d!!"�$ T�*"xA������ٹ'�}��
DXT9[������7��X��ـk�v`�}�xl~�� �V˹�gF�����ڛ�:{6��]s�p�V�FI(1�,v�-_��wذϛ� ����9��,�����%��BY]�@zܘ���b����T�����'�h���K,�`}�L����7��X��ـqvk6!4;[�;6�q �EH�*@zܘ���b ��li�U�ڰ�w��v %���o�����`K����`^h���yճ�T��=�ݣ,m�wlg��E�Tr<�8l7:��xB�n�l[6�-�ڍ�rΫ�kͮK/�7u��"v��X�1m��J�&wcH��v�Z����mûmֲR�`���˿̡F��o$,���*ʱ��7Q�l�u��gnX�� �џ5�kWv�c�MY�kiڮ��a��k��7i����*����{�{��/�,	�;7j��m����������nxW\Z��J�wc͍�v,.��-SrZ䤲��?>�� ����9��,y�ŀq�u�i*�V��f��1W볺|��O� =nL@;�/o76��ۼۼ��} #��rL_;� �M�M7ebn�e��3&~��o��@k�lPs2|�����RGj�HK+�`�7f����o��} 2�;���ݫ�];Vab2e�9��v��ttAœi�<n%ޔ�l��݄��uV�-�K?����s����T�ـj٬�C��;���ܓ���<P⮲g�훒v�0�wf wuǶ4�*�����Ӣ��t�[�} 'M�ͭ�Yj�ڰ�{� ��v`�w����8��촍�U+r[m�-��>���T��Θ�鄠>�:&�_��a�Yl��4�9���*��<��T��@ih�u���(} #��1-��yْh1�+v�-X� ���0������;����v�T���U��lPq��Y��Ha�t��p2�5��j�c��'S�p��n��CdFb{�ޞ��ZJ��4�>��ӳ����Al!"B$ H��aXW��c��*�i����D�H����,p�,L&r���O��
���XD�R$ �! �h@)) �Xń��C�>��%�t ��� D�ɠ�!�`C���>"��>b� �	`4�(��0 �@:FI��Y�q4��6$�	��D�a$ʖR��tӢ���AS���h<3a D��DR#�&�h�����6.�W���� �Ut��N�E� ��6������{{X������MM��m��\��ϝ����J��ݥA�̓=�oEճ���v�bt�� �;���w��v`����#Sj�au��u��2��`N�M���Cav�a׃��,OH�����TU-E�`��� ���0rw_�_�owذ{�����:����wi�1 �t�>��r*_~�_/�:��vZFʪ��-�ـw�|�} <�T��Θ��yy�nٶf��n�f��EH9 =s� ��,c��RH�BRA�H�VP���`[LDKsUv#�Y�_k�rO�g�3?Im���]���� <�T��Θ�o:Z�LX����_�e
U
��+��-ɑ�f��z��ݎKgu=�.���'��f�a��{���>�y���*@{�����Saa[l�W,�9��t^m*�ݥ@|��̙�ű�thv�bt,� ��`��� ���0rw^ wu�m>U�ڰ�ة�1 �t�>���o2m�UW%��j�?=����׀w��XIϽ훒mU��O{�H{/�V]h�(����2�@��6˭��P\���p�V�m���Mh�����i�Z��5��CiwZ�֔�6��݆,C�5K�ϴ�۶�y��7��Ŵ%ح����nv�����b��5
�Tݦ��&͵�c���|~,�˻C;����E���u�c���r�&a����!�6�n22�۰���M��-�]��	�&�ں�ZEG/�Is䕫�?Xȝ
��,�Z�Añۭ��qN�[WC��.�#<���c����%�6UT��m������w��X�n��?=�� ��Y%e�,*��^Ϣ�������K@G�����A7l�Հ~��,�����|�}��<{�ŀw�a&��ʬ%�ݤ�t�y���T��R �}���\u��er���׀w�����ŀq�v`���,�!T���Ym׬���u���5�W�z^��&ŵZyP��;�exy�� ���X�f�N���͢*�Q-XIϽ���(� ��&]�:��0�w�v�6��ʫ�������o� 9ȩ�"���%Q���nKm�`|����ŀ~��,�{� 9��䬱�¢K�����"�����L@;}1��F9���Id�[YmI�f�7=c4q�#
gr0�]nλK������l Z76�׀}�ʐ�L@;}1�EH�SrX�r��X�f����;��X�n����&��#��[-�f�_��ܓ�w�7:�:H1:5,���ŀu���8�5� i�c�:[��>��r*@z�L@;}1 v�"� ����E�`��� ��|�f���z,}�E��J���B����r�2�;���̅��NJ��ں[O! i;F��j�o����v�b�EH9 :ffmmٵ��w�����o� 9�T��R����|����nб7YQ%��0��R�EH\�o� #�̼��n���e���7q`��f�����_!	!�L�6�ճ�j��ق#S��Ii\��V��v`�.���7��X� :��"��XZ��n����l���]`��k��0VN�[��sb!갏-Q�Gcl�W,�5�0� ���_��?o�ݞq���q�Zt�X���R�EH�K@;}1~�Uv�2/QeU�j-� �}�X97^����9��X����+*��T�ݤy%����nEH9 ovI*�UU+rR�^����=�K3����Ԩ��z I3/�sG6!�pA\���W6�[�ŎX/\VΓ���ص�sy�zOkuL6X�[��݃�D3���yn�[Q�h�ձ�ilq&���5r�it3��(o;c�qv�Mx��X9۠;p�Z��F����W6�-ٳ�����CGb���FS��%�s�V�n����3�4�q���7H��I�����G�۰@q�OLL�� ��iUֳ3V��u��5�y�.�.�YH��X�ֲ$�a�=R��dt!2����ގ�-n�;[v����	-vY�9�{�"�y%�����72�{���W{���H9 �- ���rb��M����ɹ,r�9ev�������~&L��J���@���Va���wf雛ho� �R�D�rn����ڄ�q�Zt�Y�]�Ҡ<̯;�_��@]�k�תvs��K(�[j�c5m���*���6{%	�\�M֚V��7���u:@}{����z�3_�3/�3;�P��s�5[uRKU�Հs�u�I/���!*P���;�����ـ~��, ��d��5UR�%��0�9�T�ꪻ}�ʐ��b s��V1�XIm������?sw��v`|����ۚ7c��n�e���R�:b��} :�����u�1�c�U,˅���*�D���5ۧ�:cK������;CY�ݦ_��؀v�b�EH9 ���#��[+�`|������?sw��v`��&�&���Ӥ�LPy���v���d��I%��>�2=��`|�� ��"�"���F���EH\�o� 9�T���nm�V�T��m�`��f���2�iP^�*�vI��)O1��]qm������6N��b�&K���Ѝ�T��6�2t2��:�����������s��"��t� �K����*�5�"e�&(��U�̙����T�oE����9����쐴M�,�`�"��t����*@wM�2QrZ�r��X��'�� ���`�}�r`�_�Q@d>	3�����T�q��-��0>wfϢ��������R�Vfh������M'n©���]�.��7^m-���[��\�Z��u�Zt�Y�w��X׻J���69�������B� ��+�Հ~��,��6q�}0���wq`�kslj��X��Հ~���L@s��"� �L�ͫ��\��m�;� �;����Ł�O������T��XIk����J��fL��Ձ������Q'�@EE� ����@EE�EEh�*+����� "���EE�PP����Db� ł((�X"�0 ���1 �(B(��PTS�B������� "���QZ ���@EE��tTW�PQ_�@EE��(������LPVI��_��" �X�` �����[�� ��*Q !�b	@���( ((����VlT�UA �8��(�* P� UD��E(U
$  (��U% � *���P��D�*�T��J 
D�   @@   
Uc kN�����{���|� 0�x9FN��p;���K���� �n<����{���{Ӈ{�g�|��r>��
<=3��y���#���Up׀  }  B�����(��mK���v���P;�Vm�3�;n�v�X{��޼ ��P O��  H� D� =YҔ�� � l�8� @��ݸ    �K   v(( P (P �"�� g` 3` >�� 0 ���G  ��1  �� w�O�c� oO,�g>�� �+��      �{���^ í��f����}8� �� �   P�1 p�A��c��2t z`z�t94���@��r}�� e�p�7�Tw �Gv})��r�o->��}�� �ﴮfN�c���t����� x  >� �� ����)ɮ�_}�Kۉ��T�ˉ��y��x��gҜ ��q��$ ����n�d, =8����`y3�l`р�v;(���<��=!T��R�  4��*�@ Ǫ�(ʦL  Ob�Rm��F�T��%OmR�* �"$�JR�D 4x��������?�?���}����/{����TW�������*���������E�D���*���!��k?�5aL-��]p!pRB-q4�"�]B% Ԅ $_�%15�:�R�p?�R4�����o��~<cBVT�ͽ�������50�P�@��O�?�f~�<�cE�!Y]W\La��`L��!!,�$��沷&KS2꤃֬S�79CSp9�v���9�b2��ҶdI�!@�MH�6k'=������L��(˅�ˤ�j�{Н��I'<HWkԪ�sYT�9t�]i�����U��&�R�!�9���`�Qs�dT�ZS�5ުؤA�b{u9(�y��W��&v$�K�ҧ���N�H�R'+�Y�EȥPuNŬD508C�')}]���<+�N7^jQ�Jm��:J���^�mnצ���)0%I�(F��6%-hi줘L3�^���A����(E ��E�R�(�*�ӯ�A(�j�G%0�Ё@ 0p5W�%{{�{��)
A�	JU�,R
A`���@� ��X�U�D@��g�G)d!�3Y��p S�_#Ǆ0����.i�č]8�h�B8��)� ���0c\H��o�?&��]��+�T��mT��߇%�s�(�q�IW0\�8i	ʨWw�����%���U��+D!��E�$�*KR,�I��4)VRwV��S��PI#'�&[	��$��fL܅���K��*K.k)��+d+�&�\�\4��n�J�!
bJa�x�l.�a)�3���5Б�3bHk���(a���[�j�@��O�zjdB	�if�8t)
S0S��o^o=V3|��k=�[5)�J�
�U5,�C�j���MvH�X���F���JIswҁ
�FJT�.�	���qR�ܝ6jcՋ�e��H�{5m<��ʮr��S��B �C�+ p4�Yaw	LL�2��B�.hB1�p�hK
�%ͅap� SH��p%I4!Ёt<�
f���(@��0�H�����B����������<?5�xx+�e�a&9s�`�:�h��q����U�R4$�B\B\
ٺS$�09㬸l�$��#sN2�/%�y��jJ�ی�Ǿ����5aILӄ�+Ra�ӹ�K�9��uzOSuZ��M�9)4�)�%�nϵ�ċ.��F^��S���s&�FN���{�^^���������}�^~�*f|��P��Z����O~]��^ك��Ä�Мb̼�/
�؛�V�}WR;�eM
�jb���$�i�&���cE5����ߖ(��4���Y��lySD�;�t�<�ݩ���6��"zh���B�u=6)VD�W�BV1!��U������\td!5W厼z�NoG4��2�ٻ��ܒs��"�=^@��+�Y^RRN1{oջ�u��=�?FZ�w���կF('�-$,��R'7J�MM�$;�J���Ŕ��H H�}!��}��)3������ٹ����P�9��
�C!IM�O�7N��D�O�eC�f�v���I(J�#�.�,+���!d��U!!a=�3Ą!x�+���B��¸@��$*��F��b���e/9�DevB,O�,�
E��.,�$H�,VF	 LGy2�Os|<O��Hzq�`�L5 ��H1� �q+P! ��A�7=�D��}8G44ĎT��"a��d��#	��LXE��q#��k��R�L!9W��5��֭��n����zu�wt������;��z_�w�33ww@��p�.����B�.�8p��d1`<����9/��;���	L�Bf��B󛁹�������4#z�Gs�Ǚ��n�夌$-�%2$	H�e�	e'#�6P��,�X��c�*�9hE7�SQ;;�5�T���$����!���Ja��������X� �F%ЍR&s�~')�H2�<��#Bm!i#!'&&I�L))LWA�XA�-1Yp��4�{����ǕŬE{ٻ�X�v�Z6�jb#���ہ��u��8����7��K�f$/���K��ap�\��WWp�]{j��50J���%ʸ!�*|չ�M�'
��A�����0C��5W>�^�x����!0��.���kLc �����g	YHKp%&�7��4%3}\4�K���j�nX�����Yp�sV���U�RP��7NK�� \#L`S$
�.,+�nk��ILB5!y���Fp$�R��bo�)�4cja>����(k�o���?0�� J�\&��L׀pb�� "<@�\焾±�33Y�JFRVRYt�4!wp�H1jD��K��i�
2鰦@�*Jp�\�|4笸s�%���$p� �L�!1p���~���aX%%�%�fl4�1��cHU�)B	X�'���������r�'i�͟%k,PC�5qhP�!!@$Pԍ �H���s��$.�'Î��0Ӛxq�Æ�)����ĀG��y��	�1 wg��N,u����|5aR,�0ӆ��\B���`��\	L!pe%!�!�!ϣZ��i�p;sH�*k6gF-cB%]B,@�W����jũ��˚M2ˤ+��LB0�!C�$ �bS�B�.��OJƨsB2$�$$BX� A1!$Jxk
a�1 ,Va7Q�=�=��W��m��R����'ʖg�� �
�JS��m����]�
W5s;�]]LZ�g��u3z�ij���<�����e3V7�	sxp#s���k������YL�4\v7�8��i�4�<��B@�	Ϧ6 [�B��x���y$��ɻ��W�5O!9m8c�isVTL
�0��x��W\� �HM]:�ir���4��z��9���7�sL\�qe��B�hhB����paU�u�p�Nn��ʜ�o�	�	r�Niz��U��3xi.q%��i�Á.k��7�	sx��(ơ��Ǆ)�翿p# @	<(����A�sv��Y���k�VV�d&�jjӾJ�Q����p����-`��0�������|5����(�F��*�t�kʇ(R�D�X閶5��1��c��HH
�K��i����B���hB�@��s��H��~$�a��/��!��!0�
�1�ab�j1H �ѐ 0"����`��m����4 H-YR5$
B��"�~�2:��I
8�Ь$�#��� ����H	=�CAjc�8���J���e!��y�$�@�b!�ܿ�������ݜ5�{Tf�-��	k.ː�ǽ?v��H��^���~��$삤r9�sP�j4^�2�ka�3 a,��o�f<����9���x�HR4�@��,���&'@�+��ץ��Mc�A;�U��5j=��|�O�<7�B~�4��B���#M�[����.9�'ols���V�r��K�1RDkGA���{���c��nG��6ok�������������L F!�H��< �5��K�AZ�7�!�I�J��cבSw���@TB�N��o�D7t���x�=>�'���0��;�(����b��78�p%q��9�$Jl�ϔځ1���O\��^��)T�1!H@!H��Ny�D�|�{��'L�#su!X��Ș���b�<U~��}T�VfD5 3u��ŌՄ48= �%e8x�L��RIG�IP����eP���oԦ)��7MC���������k2i���!ŌXR'
�ZHM{V!M�Xd8�HMJlXHB��aL+'�Hs�)��-"	 IV���<�	31;�~揟��)��XI��*8P�)��������Hhۚ��$!"$B �2�֖�h P$(������꽆�MBd7>���xn`�Q��p�D�S&��ZO��Z��B@�Ay���^r�	��D�B�������%��@��ƒ��x\皝���m��.�ґ� �	f�w�Kٳ�,��2sOiM$ۮŹ�X�!�f��6H�hS��%��y��<8���Q"I3�o�̼�
H�H����8�<9đ����a�\!L�9t�?R��K��5��i(K��D�	#.lk��p�%Д�hL����2T��<��l�oA�%.B�\����rid�n�.xi��P�B�� d�H]���n���8э0"4���i�C1
���'�]��f`! P(@��!9Fϯ�p_���Fա�W$S�U^�><�i9I�$�&���x�2���g��@�p�!�*V��Q�dR=�!�B��w��&��r�XQ�YY���*F)��m"BZP�]`1~q4�GWucS�,X@�]MdB#Q�SH514tH��P�BD����u��!�P�R5\:sv<8l�h�n&��L{nn��=/nwN��������	 @   m�  $<b�l�f�^�6�Ls��Oѧa�/[�N�>h���m$!�w]`αu$خ���r}�`�c���9�{��sr U*�#���ʅIIpm�uܑ�q�-	6�;R�BM�*ڶ����m�\�ps'-�%.�u5.��PU�T��l�uU�U��&����*� mu���8���,s6�;aRԉ���;]�@����D�,�,�Hd��m���]�:9� �h�Kit�Y@4�؛�"�#���P��]���I:�+UE�*���l�j��m[-�u�[% -� 	&�KQ�`l�[I6 ݶ�^�nٖ��Z����=U.�Q�5<�Qڕ^�Ji@�����m��Ͷ������[*�����$�I��k��[D���� �-�.�j��m �8-��g 4�M.\�Jql���-׮�)C�m�	��4k��n���>.�    ���4PH��m�� Kr�Z�� � ��vky  �z��7K]�I��������'����ņ�m��  m���>  -�h��Ѷ����t�V�� $m� �`6�;B��V��*����km���  $���Ӓ��z�msi6�m�Q ��Z����l�ܲm���m���l��U�n�%U��-+k���oN�U�N �fV_4F��9�V�h[@ �k ����v;m��8J� H���W��෮�m� w-������Z�j�i��p�� kk��:C�뮀�����R˴�N�m� m��m���lj�ɗ60sѵ���z���m�l �Nl�  p ���nH)B�5�2�3մ9U@��T��<��.�{k1l.H���l�ˁڀ�ÊVUm�d��t���N��$��i8�i�Sm���鮒�["X�M�����>�흚�
�e��Ll� �kv:�ȭ�˳.� [Fܴ �L�%3����ĭ٭ۡI��"�a�yU��Ѩu�6�c�[:0� �\�$��-�:�q��t��;^*-HU@��8*�
G���8�� �� l���`-�LS���:�{ *����o������*�j��-m��J��Ԯ��U����eUT	�$���p5�"/v��,��� �����@�����`eݖ��/#{
�{6�U	˹�V�����k��T��^�]T��m�����hC��+rUݜ�l�-RUhmyI�eM��f6ZH
�9^�RP"�]i��sI���
���3�z)n��ƚ�U�%Ir��)�	����	7���N¢l�sm���@[@,nB�Z^��bͷ^�V�+n� ���eӥ�V�
I��uCb����2�U��U��1�cz�WkaQ�en5z�z^Z�\v*��Jғ$���������l�2[U*�);5U/��f�iY[Η��Z�
�J��a���⺥PR�� ڶ��Ym6� p [@��N�u���9�ԯ`��.��5J�YNW8 ��!fnY��A�z� ݵ���j^뜴1�Eu]O0��S�Irl��-�\L��+j��g���ƪ��U��+nN�v0�bR�����ƺUv3�Wk��ܚ���퍕���f��[(�̼pt�ӮvA���we�����x�R���L��f=�ɷ��*��7*�U*ʵ�q��lc0Y�K�p�m�n�#�i�+)��+�(j�:���]��;tuۨ�یă-g6�d���r�@n��ڐ<�0���:֝���
q�����˒�藍jV��Uڪ��ٰ8����>�����m�i��Ћf�n�;�P��4�BTn��ү@uU��V�6N��H��ٖ�;�n�0�@��i7m�  � e����WT��.��d�MZ1`�*�WQ��m�ݠ��Q!7m��N6�t �m�f�nDY��)�7Pp�I!�r ����t�˳�Vy��e�\�*^��;j�Mz��N�mv�b�S�d����mv� �[��   qt�t4��oa#�l��jN�)��cZ��A������Nζ�KC�m�EYbYB@j�=vP*�l.v���R۶ �!t݂Cm�@ �ز*�T��mt�d��ST<��X�ʀvz�������m��P�$��ζ��v�ٽ��e��Wj�w|������.�m��]�1�f��uN��Ѷ�[%{m���m�8   $m� �E�Nq�l�#���߾�8&� n����,��5��9�]�	�����]�?a8)�/m��Q/Yr�7/n�� �i��v�6���l��b|�m5V���5$�%�KoۖZI� pm�oie��[@8 ��   6ͳ��h ]���i�@.�h��lc�rL����+��U����Y�nIl��9r�m�`[@�(�^����ҍ�I��HHt��6֭��R�o6�rGK�5�޲�����k�K\	��)���HG6ؐ��-�.�i�'1ݓ�m��s )I��bFt�e���A�-��l�襴8 H ߛ���mUA�l*ԩd��UO,��Y�H�On�'mװݻaŴ/Z	8:�Jp���,U��[N]�d!z��&۰m� �im� $ �U�n�4��aum��U�+��rM#��f� ���i��H������a&6� ^�� %�'u6� ۗ��/Y�koP^��i2�+[U~����e�ꃍm�� �l[l�b,�ڪ������G/h�; 6Z �� I��mu��PR�� )�UN�Zqr��V�m*��5mvWZ��T
C�+@9�5[v2G+�mv�m:���6p�$$ ��&�J�J���TPR�X�]�-�`$m�˴'n��=�'W=�ɳ�F�;m���ͳl�J^�tPK;w[��h�����հs����&�t�uUM�c>"�^ZڕҀp�����8�Z;[.%�Yz�7R֭�BI�a��uX���&;]5a�DLA��UZBh�(j�����r��Ӹ�eZ��G�3@WX)��C� *�Gm�-�UUS��ʠ�R�9������˻=U u���^6j� �@t	 ���N֣��)��p�@��K�tXb�썶�c�k6��@����`�Am�P�ml�v�A��&�iL�`��{e����V���]n݌�*�!5�����sV��yyW�����26�m�F�H��O�}}_e���UJ��[��m��6�l .6�s��Vۮ�Lp����lh H mZ� ��d��c$$[EҶs�����H�8q'8I��s��l*�Ժ�)�6 ��[@     hq�I� �C��˵AN�>�}�T���� �d� L"�!�J���˷Uc'�]l	�k�-�H��p$m�%���n$ �  �h���`rÔ�0�W	��QKp\�J��$vOi+f���:@  v뚼6��'-���on���
����	V�A�#Yy�ۖ��-����[@�     �;l6� H ��� ��7Y�vH�B�T�i8�� 	��#8����4J�Vڕv�K,[��tH	m�iŖ�Z�v :�؆�� ���[@Um*�TK���\������Pq��)[����	 �e�v	 N�5�Unpj�����Y�P[@8�t�� ��������R���ZڍH �UJ��3�kռmɶ���̭$�.��.�'L��� ����al�pM��K&E	 :��f�#H���uN���NCY���n�v�f��lE�%�+Y9�MW��Fu�����X�q<�[7�9�A	x2����T�+�x�I$;i6�ދպ[Km���ﾕj�Z
U/gu���[Vզ���`AmZv��(j�*�PneUUj*�H 8q� @ �m�@�u��f� �ml��� ���h   m&� %���n�l �lH���	 6� �h -��n�L!#6�ڐHH�-�l#}�o�U�:�$�8�K��&�M+��   m�KE�l��l�a� =�=� $8ڐ�A����6ش�5uUuP��J���    �Yv[��D6�lh � �[@ ��`   �n�$��oP  � � 6���� $[N��� -�N��X�Zm�}l66����f٪���R����ݺ^�N�l	$�Kmi&�l����m ��  	o}��߾��Bɹ�qѦ���
�||t��S+ -�(D��U�Px�*��[FE��%�3�#jd��QEKp9��Z�d� ,�mZL6ͤ�m�bI  �lh�� �`-���A#Z�   �[I� p�-,�N$�EP��[�S6Hi$��s��nIN�o-1jг���y�\s�]�"d;l�ve�r�.K����"
���	�?��H_�R��j��Ă�'�ؠ`	��x�T�Z,<�N��k��x������+���WQ�N(��/�C� ���q?% 	��P�#�@���O<�x����5"B ��q�
��G�Eq����?==�_�>�|3���~L;L ���@Qz����? �R����P�|D^	���"��GШ�^��x�T�U�P?1D�AC�+���'D��U�'�� pE_�+��}A
k��>�A�(���?*UG�b���*T<  <@uG��pCA� �"� �*�UT:��l<�pE?*#�T�xP��
�P��@����O�� ������ �����"%4���A�",T�ō������ݲ���]3��ڷD�]u��T u�\��f�{kjy�HU���Ѹj��7h�ѭ����s��i�\T��Q��1+]nE�vr2�)>�����8@^G):Q�Yt�q���Ҧ���4N�r袇[R�U��]�����Tz�e�Ո)���]>;cp�:��8��)����"M���Γ�f��
���:
��q�$&�I�Yv��:�vô9@5k�]g����%�<�8n��=��v�l
�G�g�y��1��9���3�떊^ɻ�l�w[d�D��]�K�]{Km��3��B��/=I���Sm�-)72B���d����U� >���C��<�����]m��{=@6۝�sk��]G�[�{kS�֠n1�`T���N��}m��8��7Q�ER�l�	�S�BZ��g�0͜p�`����X�I�6�v���B��*��퍷N�mWmv5lv�r��.V�Kd嬢��2�23��6�d�ۄ{=Y�hDzMn���.��p[�u�m��U�z�K��]k��d^�:υ��v\�Q�yt�x�km+��nJ2�%��4Y\9ɮ��%�xrK{xuE�OR���Q��4!�A�h7ap��\�ZM�d�=ăq�\c;��Ѻ�byz��v��ɦ6�&���:��ږ�a�ɲ�����g���P!Ժ�H�x�v�8N�܏Cfγ��.ݲ�����-U���qvCex�c�]��"��U�\ɹm�x�Ɓ��[G	�g!��#=z�ij��غԀM+���dM�<;�b�ѯ�ò�Y�Z2޷Z�]�i\�J��l�p��bv܈�@b���mUҷ-��9��e�\��&�p�7-�2'���Ga4C� QڸnZ&x�ڭj.�nRt��ͅ�n��B�8����<�	�U_nʹN���U]�Ѐ� �8Κ�8�v��U�f��h�ζXкt�."C���ug8�Y�y�L��4u�i�6n >:�ꢸ�F���⇊*)�?�T8%Dz"�⿳۹�vI&n�.]�L��=��<��h1�N� (�� �q.σ"���1����5vwm�p�sJ8�7Y��I=��\D�Ml��F򜻤��h+�&�ڗ�+ݎ�ٞ��`hM��^Gl�
�3�,��<v�٣!���9cl��v�튺޻���nA�|u��kdh�"�茜�6�H�Y�9);Q�tF	�@��-���@8�|�x#w��fZ[G�n��`����<9}�g��;�Ó+�w.���8�9��F��;siP�6�Iy���U����}�
Dń�I�^�h^�@/[4_U�\�x�+��I�2I4
��@/[4]�@/[4.\�6�q7�@/[4]�@/[4
��@�4ew$����rI�Z�Zz٠Umzz٠��<,ƱLPh�H�O1c��W:��J�ʮUa�H[�=H�D1D��1)�ȴ��@��zz٠Z���U'�y&$�ƛrf�u�6g�yDX�+�T�c��(R]�`gN�/[��~���iLq`�ԓ@/[4_U�^�s@-�4��tɒ%�֘-Y���7�k��Drup�o ^�h�*��`�I$Zz٠��z٠Z�����>x���/9`����uv:[rF^���ej�u��#�vΌ�u���� ~I'��������h�f�g\;Ɗ�q8��I�������� ��߳�3�=l��G 9&6ә��'�g~��N���'��� 0B
0��IB�d(�;�u`��`fI���lY�܋@/[4޳@=m����?p��?���Ʊ�&�_[4�٠^}V��n��q׶;z%�#��Wt[k�ѐv��w;�I�Q���4�ɸ���9��[f�y�Zu��}l�:���&B%1D�rM���w4�٠������)<XI$�h�}\_��WuUiG�.{\�ǋ�P��D�1�3@��^���o$����rD��F����j�uY�:o T�(�1�՚�7ws��]�@��M �h{��{q���sb�[/��&�8z+��2;�����g����v��=�e�6m#,c��/��������uz��h̫
�$Di)�Hhu�@��^���Z�Jh�|RO�D�1<mɠU�@�v���Z�l�?W��������[��]��R��=�. �[4���:���dB��L�h���w���z���vDzBH�[t@��$�ܺ)�RdʪhU$dN5�e5.�4i�[\nz�4��̵�k�3͗�.bޡ�#W���ۍ��k|�O2����ae;lb�=s'n�B$��K���Kͽ0��`�}�..��q���8h�s��������%�+:�gs{v�9|c�N�]�gt��[[��4�gq�������u���Yų��V����������������a.F��۶*�it��M՛v'\h�c2p��MC'<xI$�p}~�}�h�ՠ_>�@���X����M ��4Wj�/�U��� �;�h/���M�ڴ��hu�@/�� �ݏ+�8�̓rG�|�� �h�Y�z�V��ʲ�#K#���Hhu��;7��Ξ�`vmq`~
!(Q����S�l��7Z���9q��n(��Ѳ%j�H`������0��<��V���o��k���J���@��p�;2�Uma��������J�
�����b `VP@�&	���#$��-	eQ�Ot>ѻU�ɛ�p{a�5��:RC���F�2`�܋@���h�S@��^���Zz�i��<$�H�>V��˯�@�v���Zp?��X��y��C@��^��fu�|��;��=�S@3��q�Ȇ�� /�q�j�x�q�:�k	kf����=���}1��FL>L����$z�ڴ��h�)�U�@�{&V���d�ے8���h�)�U�@�;V��U�+Y$m0nE�{���_u�o��3|��B���;6w���'y��9SL�1Dۆ�W����Z��u��?W��2c2bc�M��Z���)��f�U�I��I`�gr�rN�dW]����dx ���}u�zػ��n"�q��F�2`�܋@�_U�wYM �u���h��qj�چ,xH��\���.�!�I��H���].\՟5��PD�܆���z��h�U�wYM֑��:�q7#�@�v����)�~����X��M��2�&70s$�ܑŠ_g��%����s��^�8�\�����uU�<s�Nݮ�c�Gx�{j�U�ݝ��N��;x�Л;	�Jumxmt�@^���ՠ^}V����H���Q
&�4���/;V�|�����?W���̘����@��Z���S@/���]j(�FLiȴ��h���_u��j�:��J6��&I$Z��%��9��G�.��5�]�]S������f�p�m@�{WOm�0��Pxyxō�۷[s��g.ݻ 	�]f�99�ֹ���6�=m�C�qp�Y	�;�����?5�����↲u�m�֜lG=�0�e3�MVư���gy��60��*fg��ͦ^�G�n^*3�g�����,�rr/]un�Q�mlX��h@k��ZU�Q�ۧ�p���[^�AΩ�Ĳͻw3r曲���)���͓9�\շf�A�n]�&(�nG�����vW*�Ӧx���p�A��[������^v���Z�)�Z�9������nI�yڴ��h���W���vL�ȦD�c��r8���h���Wuz�j�9T��f(���m�r-���*�@��Z�h���i<���m�@�������ՠ^��^�D�s�k��f�giZr��E���m�a͝�Wk�:#� ��q�4A 2m7�WZ��mp�Y�]U �ɜ��b�[�6�L����I;�w���Ĭ*��I+H�볺��7����`~�u�R��cɃ�I�z�h^�@��z���.v?�ت��DY&G!�U�^�yڴW�h����s�Y8�M���/;V������� ���,��8_%����d^s!]�SH��;uj�]�Jc��s=�n�与L�ȦD�B&��~���@�e4�٠^v��h���k�Y������T�OI�y"�>�@�}T&<m�q%n^�������
m�92Ԫ�εb��MBW�S4��ӹr)�Is�uhUH��)<!/9��`d�+��c  ���$X�@�s�mA�I3ysX��n��*�-/�x�=?3IO4	=e�!o����f�M�C
@��d	m�F�R�YsH����O��ČZ@��b,ᐌ ���a����������<�� ���D 0|ǰ����c
a�c���s�c��Z,"j�	�g�`���v�[�Y�FD���/�aS�fg�a	�0	�X1C�C j��q�e�|
��	!��*¸�h��Xs��-�7);H�^�HQ�2��B&��cL�aM.00YR- �n@.������0`�U��1�e��B~/���<ᎇ�+�HG!X�$�i��r���5"���%R��A��{���S�z������"+�)"���(=S�:�����~*�(_��=���h��y����D2D��J��ȸ���6��]�W�wY���p�v-�nR��3qf����\��'C���p�k�o)��Y��:�W>�n�D0P�ܺp��og����M��sƵ�gm���{�O���:`/�����8�y���Ϯ����<�.ꕔ�_%K6��[��Ӏk��t�HjI��8�7����%}��+�V�������"�ﳀ��q.�'&À���z���4�lrH�>�_t�pM� ׼�k�W�QW��Z���TW�Y�����E��Vf*[��3upoY�~�s\_�9�.߳Ɓ�ޥ��:K+/Ts��^^�e�E�������jkr]:�';=I�j���>o���>�5�3���� �g���$��'ؚ �(�	ǠZ�[�bG��ˀ�l8�y�KH���3i���#7n�{\oYĺJ/9��"�=o�8Y[���7wwupK�$�py�����=�.0�C��,6�U�K7N��y�J�d_�Oc��o���'�b�Sޒ�̎m��n��gQ�l5�+�n`�:Wh�zvC���܍�8��s�p��=;��	1��v3��7�%Ӟ"GM�����s�ڸ6�C�l=��l�=��v��c��#���utݞ\$��d�4v�
sՑ���cڱ�gl[x0�ö�t�3'<$�Z��g]�r,N�o2):��:pÝb�f�۞۲���k��q(@U�r~���w~G��������ݦ����:e���m�=�N7bSn<�#y䱒K��M�5��Mq��RG�>���@�}V�m��*�W�{��v9��qD�c�E�_>�@��h{��-v���;1F�'�7"�-��}�h�V�|���U\Br(���� ��4�ՠ_>�@�e4��H���b�������=�/�#���y���ߟ��حm��x����
�.UOOG9�-��j�N�8�(P;��mN*�^�7K�dwW �g�����k��K�AH��;ತ��aH����`v�q~Q�]�]�8�\��k����Da��Q*Xn��v�7N/9��6�WI_>�@�e4W`��<��E#����@�}V�z�hwW�wc��Y����=�ڴ�S@������bϻ�j`�L���9a�v0ʦm�hŝ�Kvt���:Ԅڪ�0�1I�6�8����>�O��uz]k�/�U�}���O��L����Fۇ�>]~z]k�/�U�^��yۉ≤@q`�z]k�/���J��Ԑ�, ����#�1F5�J�,!D�F� �Q�K�κ��3w���**\FF�m����h���_u�]k�;��I$@�rI"�=l� ?�{�{�����\���%*&�so]I=�TX�"�-�b��ƹ��MN�V��M���:2r�bŽt'^;b~I'��@��Z���S@:����	���)�@��Z���S@/���vL���țM7#�@�}V�z�h�Y�^v��2�LJ3�o�h���_u��j��T�^f�{y$�{{�f�Hbf���f�yڴ��h����z̿`,�&�cjc�p̝�l�\s3�:�Z��$�7vKf�-��ja�Xnch���b�O�}_�-��Z�)�U�@��.�?���F�iȴ��h��@��^�yڴ�u�T#p@��I"�/;V�W���hϪ�.sز�!�$�$Z_��~�� �g���=�p��.*��+Vnn� כ�]�Ok���~��f�X(��9�534�̹h�e��Mͩ
]L��U]��{H]�z�JX@R�����NCçW%�����%����<:���^�z��Okם��9�#��VC�1���@9�f5x��#W.�Mqn�`ۉOn�)uc�H�>ݦo�����n]3�Cӎɹ��㔳�Ց��ˀݷ�ˮ-^0|����ժׅ�I`*F�a��%�w�����\v�l~���G[.úK���L�Ҝ�c]�����u�|�ۓ��v�V�@Z�h�hQ��;�Z�j�*�W�Uֽ��e�Q�cx܋@�e4
�����@�}V�|ʛV4܆Fa�4
�����@�}V���h�n�iY���j�R����*��<�g9ߖ���h�Y�w����)��q7#�/�U�u��}�h��v���߿�`n��;�i��\�����an�Hٱ�P^Kt�$��n$d�8��k%�$�E�u��}�h]�@�}V�s�sU��	�4�����â, �@����K�:��"!dP��S�vl�;{�� �˰��!��)�@��Z���?��}>4�M�ΙS�E�64ێ=��Z[)�������R��D���o�hl������~�����U�~�5�XGp�E��:a����D�ǋͻF�i��.���i�Ԍ���p�33NZ���i��Ϫ�?[)�w��$0m�!R���<��#��M� ?��׿�pAL����y�Z[)b�IE�$�:�{�V<�5p�'�c@��I"�:�M ��h��@����0�W����D9 ��h��@������<�.7����F獺zp�Ŵ���!�'6��;(Z��3�닳����j�m�Vנ_t����h�Y�~��*n(�rFƛqǠ_>�@�e4���9[^���_�ȓxbq��r-��8��x�5$�{$\��*1��7
�(�34��RQ��RL���o$�� )���_�����=ҌX�4�Xfn����UU�\�ȿ�rl8�y�����V�R��e ��wh���FѲ� mV��n�y��^j�H�G��2n&�z]������}���I��9AY��*�������"���yI3�k�yҒ%<��T��J�Ջt�"���y[^�Wuzu��P�O��,XnV������L�"�g�=g ;�h�%QG�F�m��k����������}>��m���v		�"��Lg��!�������x%�c	 Aw���k��'�<��RFR~T�q�I`�cXB�!A!=(V�`Fb/!'"#�#�fb�"A�E2~���Oށ�@ &�?P$!BH"� L (؀O���%��2X�����K�
wh�Sa�Gy�
I�ME�{<�@)A�Іg�bIw0��	�fh��Mu@U�[#;m��=v�3�j.�[�;�i�����m���V N�/Y^�<<g�8���clr�pv�V(	��ʜm>����{&��zy�{\�2=&������UN6�Jq�Uٴ�i��vŷQF��F��� �Wf�N̦:gY{Ogd�ZTқ��'1���:Ìʁ�1�o��YWv��i�P36"�H]�nY]<+[U�`7n"^���E!�o=S�J	r+JѸZ�\dwt�1�&��mۘ^QC���EB�KN��7��͂�q8G]v(ݳ�b����#�ȏ0gk��X\Ξ��7'C���$�$�K�l�\nn��dRp*Ge2еxͺ��/\Z㣝;N�{ZRI2:�G�lu���@��#;�L��GC�W�Mtתé}�;Q�֭=�\g6��՜�˔��u���z�rj_8	fV�:�в���%�>2�^�W7fj�]�x�����:�R�B���c?-V�CNZ�'�y�I�h�� fxk9;\����۔�f��u�`���!����x.�s���^	���&��b�mK�.�J���˺1����j�W&����9ę
��^Θ��;�6��;5!�G`��'��	sU�GE��7Of�Nz�,����s��X�Q7����zۇ��ۨ��s	���\u�t��@uִ�
��Ƿ1�㋮�⚇����v��MkS�ZU]���!p�pu�}���[<ä�\F��Er�%4T:'3i��&��s�h�iZDM�Wnvv66 6B�7m񢙵��ESi^j��A�w�6
�l�֬�jM3������iM�<u��k�!¹�9N]*��q۴sH�ئ)9�Jj!��1|�ξ��pv�9�C�v��]�����.%�j�z�.x��v,��8�	��^����ۺ:Lr�&�1U��R�r�m�TXP�H���N�bM�Np�rl'h[��%�붹b�I����-�꥗�V�n�=�lۆl�sdۛ��P��=Q^Tc |���t@� j�q�'�?�".��a+ݔ���ۭ	�m��(ݥ*�[��ֻe5<b�s��8�z�	�l֗��;���cV�S�'V�b9�zg:��O9�啯T:�D��9%�V�\]b]*����6�n��g��t��hx.^5��hLY"�7 �_2#z1�p�n)�.��6�뇄c9��������k��]�6��)	�a�|�ګ! �����M�����x���K�i/m�v�u7���ۀӫ>���)��l4��D-�[��t� �ō�7�ȿ�z�?ƀ[�h�y?�E�{�d��n�Q�fi���D�2E�E���:RG�$$���`�ܓ@�?�ZW���e$��p�o�~z�	j�����n����pM� 7�9�.�,39jT 7w3w8<mp��O�_��-����. �-m!��"����������I m����k�8�&U��M=�Ly�&8�$D�~ ����:�W ��Ϯ����������|���6����I�s���u�1�� BP>ݟ_��r�w�Uz��1#�R|6��7Q7�������y�k�t�Q������*�x����I����>�h�o獮	T�G3���,2Q�n�Q�,��4��T�ȿ��9�Wj�=�Y�� �4�i)q����By�]�sӰ���dW];q��	��w�|�Sx�A�6ӑ����h��@��_UU��wu����8�|�a�Un#3un���5��(�px��WWi�9a��R�wVn�ɰ�~yû����UuWY�rE�I�.׫+�*)�H7Q���Wu_]��Ug���8	�}���5��UWUy>߈����1Ȝ#�G�r�PWWWuM��I��~y�~=B����[�-��c������zZ��c1/j�&اy�\kS�v���������b��B�f���c���z��������"�<��fn�p��2�7W ��t����H�9��"��5����'�%Y3w3A�����8<mq*��)2E�96�o����X�b������������w�.��{��g$�������C�QF���W���O��D�ȓr)"�-u�]U�ۓ��Q��<��?m=��N%z�:�t���\���%�m�Ȗ��;l��GBj�����wڽ��� ��u ��p?<�<�.�������%<�e*Xn�7Q�� 7��]��WUW�E��g��>\��t�����:,��b��3M�����g ��k�uUwI96=&��SŌ�պjՙ�f�����Q닀rl8�ox%]]�sd\W%L��me7����7��>����ꪫ>}������-������r�31�
Nzv��(Mg���9L��n�K��.,g����gwSm���Y��d�ӝe��R�]gwjӤ� �N�:,�=��ƻf�d��np�]��X�p:6y�@��Ӏ�t�mm�S ږ��ݧN;;-��Z�Ƀ���I'kǢ�������2q�9ex+��`q��θ�Ӷ.dk����[����1Y����#TR�H�Ig�wwwu���n�4���8upq�]f�lk�%�&roi��k�#�g�9�U}��0o���L���}��6���R�_����1�э��ccC�M�6���\��p�����H�����Օ��7V�<qpoYĺ������I�.��>)nn�I7Vn�	UWJI��	�7�i������_��r�W>x�8�A"��_[��WUw��U��}�~���6���[�q�4�ᛐ[��2dљ#��!���vHmѻ�n.�byzK��M������o�y{�:qm����>�����poY*���=��@��>i�L�B(�d�E�^}V�������>�~��O���䓽����U�������ݹp�w-�sup}��p���*��"I7��\��5�Z�p�Q�fi���WwY�?���� ��k�U��)'C��2A��&2�9$�:�V�y�Z[)�����ꍱ� ��,qqq���'r����k�N�g=�vPc;��mN*�w�����4B�<�7"�/�}]�hl��?�컻��@�H�N+7�ͤ���7W���*��	�7��$\�y��uUi��:�J�jԃu�t���ﳒN�;�Ɋ.���򣚭w�{�����<i�LX�&�����Q싀�\��p}�]Ww������m�����/����
��l��k��uWuQ·����5�o8��~� "�	.��l�3ܠ��]������J�����LMv�t�x�F�7W ��� ߞ�z��uuWW��LqpW�
fmj��44Y�p~{��ꪪ�BM�$� �����UWWy��σ>*���qfa��� �>�x��q*��Ҏl8G7�����In��Ջsp��	uWWt��$�9$���I�Ip�:�ʪ�r}��=�|}�H9$����ȴl��7�x7�y���������E�q�^�:�W2m��J�o%�;z��������tq�n�o�{����ݏ��(�j3[��}��x<M� �y�wuu_�$� �����T�������<�7�*���$�$�p~{����"3*�k2�MZ�0�ջ����z�%�]�$OI�D�x{-����3ws3+supJ���NN� OI�������
���XDA� ��x	UWuiԓ��\��p
��	 ��_s����f�[e�Oe�Y7�]�f	�G�yp�^[��]��pۆAV[��u�Ja��6ɣB�����l��a��7lΊ��M#c<mٗ����{WC�� ��k�m��@`cdssk����<�0p��x���έ��һe���p;���ò�G�ѭ�@������#�I9������$7T=����U$	*�����w���ތ�����
���.]��in���蓦8�[.��7���������BM�ڲR�[�����o ��k��z�uwwU��}��;���Q�&BGjI�_g��WWUt�$��W������U"�V%��﷉�Kı:OoNMٛ��[.n�ݺ��bX�'{�vq<�bX�'r����K�UHdL�{����yı,��]ND�,K�=%����rɻfn�'�,K>A��>�߳�,KĽ>���yı,罺��bXȏ�
�b}����q<�bX�%���)��2l���ND�,K�w��'�,K��@`}���yı,N��>�O"X�%����aY	��	��c��t�ə��j��=�#���`�m��r��?߯�˾�A����C:�ֹ�Nz�J�z����7���{�?g~���bX�'��;8�D�,K�}�`*�<��,K��﷉�K���������j٤^�/w��bX�'��;8�C��7�㦀�!�!'��G��,O�~����bX�'�=���yı,罺����2%����$���m�dٙ�8�D�,K��19ı,Orw��'�,�G����?�����Kı>�����yı,O}�ܷr�1���K����bX�'�;��Ȗ%�`�=���Kı=�y���%�`| L�������bX�'����3.�tٻ��3wx�D�,K��n�"X�%��G�}�Ӊ�%�bX�e�ىȖ%�bzw{���%�bX��٦�@y�rXؘt��nX=�(qPm�y6,���l�N��t$Č���/}>1��..��,K���s���%�bX���s�,K��'{��|?DȖ%��qm�H�E�.�c��1�KR7l����%�bX���s�,K��'{��yı,罺��bX�'��;8�D�@��M�`ߋ�e��?�a�7ws�,K��'����<�bX�s��ND��b����H��iU�Vx���`��~�O��)zR��T����(�#�G��P��T�XA��@=�1c�h%��Wu�sa@�YMU4$$HXFXOɊ`H�4]RD�c"45�BR�6?�V4�#e!T!x����"�`�2[��#<�B�$���$້P.�֤�A�JR#�JZ�
�$	,^J�s%"	s�$rV6�j��`�#�!r"��M�S8����Q
�����9�TW���O?�PP�8���|��M��?N'�,K��/�f'"X�%��}�;36����˗&��Ȗ%�@�?o~���bX�'~��N'�,K��_{���bX�'�;��Ȗ%�w���;���Ӝ�/M���7�������O"X�%�����1<�bX�'L�ﳉ�Kİ{���r%��ow��ߟ�ޝ\M����9j20��\1ph���=���'l=q�Yn�=�Go�|<���6ff��Kı,��n�"X�%���s��Kİ{��� ��
��6%�b}������%�bX�}w�6�X\f�e-��ND�,K�;��Ȗ%�`�=���Kı=�y���%�bX�w��"|9S"X��w���Y�l��͙��O"X�%��w�Ȗ%�b{���K�D?�lM�g��۩Ȗ%�b}����x�D�,K��ӓM�wp�.��ݺ��bX�'��;8�D�,K�����Kı=���x�D�,���*݃��n�"X�%�ܝ/rw).�lݳ7gȖ%�bY�{���bX��Ͼ�x��X�%��w�Ȗ%�b{���Kı=��2N�7t��g��#��O%msoQF�9����ҙź`.s:�a��9�Ω��}����d�'{��yı,罺��bX�'��;8O�2%�bY�~�ND�,K��I����.�fS778�D�,K��n�"X�%��{��'�,Kĳ��u9ı,OL�{�O"X�<ow��q�3]���/M���7��b{���Kı,��ND�,K�;��Ȗ%�`�=���K�L�ث�:TҐ��(��.�L���D��~�ND�,K�}����%�bX=�{u9ı,N����yı,O�;���&�k3&f��r%�bX�3��8�D�,K����Ͽ���%�b}��׉�Kı,��ND�,K����;)>�r�.nf�ɛ��q7k�n�y.��0a�6��C\�d�%KSm��ۜ���q��[y��ĩl;��kC�Wu;��힛b���8z.�dݽ0����������l����Lc&����rݲ���ۃk��f)ǎn�&ֺw�^�]���ܾS��'k���v�]�l9�"awl�S^�ج]Fa�n�h�h�n��{s���{��wy�www~}߆����W�=&��c�A���f;hݑ�ݺ�V
Ν;nr�ac$�%٧L�͸nn�Ȗ%�`�>����bX�'}���<�bX�%����Ȗ%�b�N�M��	��	��ֹYH�*�K��ݺ��bX�'}���<�bX�%����Ȗ%�bt�{��yı(��y�+!2!2)�l�-i�ٺf��'�,Kĳ��u9ı,N����'�,K��{۩Ȗ%�d-�.�L��LQ��%4��%
J�����Kı=���x�D�,K��n�"X�%��{��'�,K�goUB�!2!{9Z�T�H�&�e�ɹ���%�bX=�{u9ı,?�=��>�O�,Kĳ�����bX�'�;��Ȗ%�bzzl��m˘n�8�[��:.�+v|�W�<O����ۗ�V]sV��]�^�^�/w��oq��O{�vq<�bX�%����Ȗ%�bzg{��|O�2%�`����r%�bX�g���.�K�l�͜O"X�%�g}��r.����a�*��9������yı,�߮�"X�%��{��'�,K��3�ۓͻ+s377S�,K�������%�bX=�{u9��"w���yı,��59ı,Oߏ{�3L�u�˴���'�,K 2��`�	߾ߧ�I���l@�O�wg�}�O"X�%��߰�3m���0��sv�r%�bX�����yı,��jr%�bX�ӽ��<�bX�s��ND�,K�?t�B����H��Y�;4��i�Me:x�=��1'b�)�.8.B����_�ww�]�~^��k���Kİ���"X�%�};��Ȗ%�`�=���Fy"X�'~��N'�,K��&v�K�\�$ɹs7S�,Kľ��w��Kİ{���r%�bX���vq<�bX�}�59�S*dK�~8_��4��73.f��O"X�%��w�Ȗ%�b{���Kp�BB�
`&)����0�6%�w���Kı/���x�D�,K��Zvf�̥�7�۩Ȗ%�b{���Kı,��ND�,K�w��'�,K�����S�,K��=>��f�ivM�����Kı/o��ND�,K�V=7��'�%�`����r%�bX�����yı,H����)�4�ˮ��Jm��E��ݍv<��bMt�p��yۉ���t�f��e̗7w�,K�������%�bX=�{u9ı,O{�vp>D�&D�,K�s�Ȗ%�b{��|K��L�����7w��Kİ{���r�r&D�;���q<�bX�%�����Kı/�{��yı,O}��!�r��&wnn�ND�,K����O"X�%�{�wjr%����/O��x�D�,K���S�,K�\��T���r2��T\/�	�2&}��jr%�bX���}�O"X�%����S�,K�EPT��y���%�bX��)�)s�fY2n��ڜ�bX�%��{�O"X�%�ʌ��]O"X�%��~�Ӊ�Kı/}��ND�,K��I^�O1=n�[]n8;sD��!ǰ�ͦP�.�tcZ�K���{��W�7�mv�ʈ�׏�,K��;���Kı?{�vq<�bX�%�݉Ȗ%�b~3��8�D�,Kޚ�m�I���]�wv�r%�bX���;8�C��D
�M�b_￷br%�bX�3����yı,罺���«����Ο���4�n�v�͜O"X�%���݉Ȗ%�b~3��8�D�,K��n�"X�%�����Kı=��L�p�n��˄�݉Ȗ%� �������<�bX��߮�"X�%�����K�� �>�۱9ı,O�N����,��˻�n�Ȗ%�`�=���Kİ�@�{��N'�%�b_���ND�,K�;��Ȗ%�bt��!���^]ٷ)�1�6펽+t�(Os��3�v��m������>n�3���bִ��V8����Ҫ���n���QN���&�<�V/'#دgF1�V�W��=\�r�`-�Y�
�X����;��p�������u�bS�;p@q�eƶZ�,�.ݪ�w1�\j�w`��0q�v�������r;���zguY\����>�κ�rNtl��I�;��9���nlɆd�nɹ��5�{�r�nL���ۅ��@��GBj�����is6�i7v����ı,O��s�q<�bX�%�݉Ȗ%�b_�{��yı,罺��bX�'L�����\��v�ݜO"X�%�{�wbr��؛Ľ?�����Kİ���Ȗ%�b{���O�2�D�;��s�3,�7nf�ND�,K�>���yı,罺��bX�'��;8�D�,K�����K���ȵ��S	�jf\�*j��L�ϔ d��]ND�,K�}ϧȖ%�b^��؜�bX�؟����'�,K����'��i���m������Kı=�y���%�bX���v'"X�%��N����%�bX=;ΡY	��	��N��Y5@�&e�m�v̧m����7/V�˺�F��Ns����q�b|��Sj]0�Sn�3G�a	��	�~�۱9ı,K��{�O"X�%����C���&ı,O�����yı,O���e��[t͔�M�؜�bX�%�w��'��@�B�⏀�^DȖs��ND�,K�{��'�,KĽ���9ı,O2~����[t72�᛻��%�bX=�{u9ı,O}�;8�D��PdL�~�۱9ı,K���oȖ%�b{�:�˦l.�wnn�ND�,���;߼�q<�bX�%�����Kı/���<�bX ����r%�bX��tϳ$��m�v�ݜO"X�%�{�wjr%�bX����x�D�,K��n�"X�%���gȖ%�bt��Y�4�&;f�M���1r]l��]V��{9%����%��6�����&Mۛ�S�,KĿ�����%�bX=�{u9ı,O}�;8�D�,K�����Kı<��p���3ne��sw��Kİ{���r%�bX���vq<�bX�%����Ȗ%�b_�{��yı,Ozi�����.ٸnn�ND�,K�{��'�,Kĳ��u9��`��������K�|��<�bX�s��ND�,K�~;a:e�2Ͷ칛8�D�,K�����Kı/���<�bX�s��ND�,K�{��'�,K��۽2�̖]ݲwwS�,KĿ�����%�bX=�{u9ı,O}���<�bX�%����Ȗ%�bw���Zn�]7l��g<���{���C�r����c��o3��8�ť�2�t�ff���O"X�%����S�,K����oȖ%�bY�{�3șı/��}�O"X�%��۳�vm��&�wnn�ND�,K�w��O"X�%�g}��r%�bX����x�D�,K��n�"}�2%�񝓦}�-�ɶ�ۛ�x�D�,Kϻ��r%�bX���{�O"X�%����S�,K����oȖ%�bz-e0}N��UT�UB�!2!<;��Ȗ%�`�=���Kı=����yİ=W�E}NC� �	G��1 '"d�n�"�	��;B�754�әs2�j��X�%����S�,K���+��^'�,Kĳ�����Kı..�!2!3;�ˢ���353"��^�mfr���:���W1���8�jvJ���u���x�;M���7���{��{���%�bX�w��"X�%��w��?DȖ%��w�Ȗ%�b|{����l�m�e����Kı,��NC��L�b_O��x�D�,K���S�,K����oȟ�+�2%�����w2Y��m.��"X�%�}>���yı,罺��c�"C"dN��}8�D�,Kϻ��r%�bX�d��Km̒��37p���yĳ�Q��~��u9ı,N��}8�D�,K�����K�� I�3���'�,K��n��K�i4��sv�r%�bX���vq<�bX����"X�%��'{��yı,s��ND�,K��"L�V�YA�ICzEd5H*�O1j�!V��`P�E�FIA#$�yZL�{Cr�n˛/�an~W�F+�� X 8�`@��cZ�D��>y�."hr$<B"T��%ĉ�
�� �"���@dV�JQ��$H�	�ؗ�!$.��Ȅ$4I�@a�+#$��."E�$ Ą�gwM���ҙsww�n�#�D���:�L�;9(��ۃ��u����ڷh!�]g�sjg`�bm�{#���/UBnCQ7.�	,�t�s7a�ݧPEGt88�BЩ�4�A�`X6��n'��m�v�K�\���&`�P	֜v2;1n93��ݲJ�Lv648�a��UZ���K[%I,��n��vʽ��f�Mv�۳.���s=�Jmֶܲs�(��ճ�8L^|�&U��i�M��5�pն���
bt2�$��mPh���Vٯ;.���Vݭ\�Ҙ���i;G2��{bwmvh��
��D������[�iTH�%�n�my��iɃ� ��������F�X#`z�Y�I=bz��,���l!wX�g4t�
lnB����ܡv" �ˤ�^Ʒ;u��m����GC;��60'E���vsu�o6��RS�ţ�e�S�'��;��%X��m�u��#���痒+Be��<��ѷ[���#\��=1���6�uG��ktRRv��͊�����8ȝ)��%�g�:���8]�����H��S��f�W=	m���m��<I)���VS��6$�8�v�A�J��Qj�	$�$L�s7���4��p�=���D�݋X���q���.5ȮC�Î�� �v��L7m���˴2˲��[$�꧂�L�g4v�M1Y���ݝ���v���O5������b�ݮ�=[ꬔ�ܺ�ظ�T�&q�y�6�"՝ˢ�.D�V�VҼ�J^vT�{qsv�=np�%�c�-Ճ�hu���ms�]�\r�ͮ�w;vhNI�M���]zGi�:�b�X�=n�qi;r)2��� קhw(���]��&�.�R�����1�4٨��ʭ���G�7n:C�gV�(���vd�\v�V��W[�;TuԻ����m�SN�+U���b�S��\��/\,���m����J�oj����rf�ny�i^�q���: TC��R�@W�O5@� Pᩡ�~N�����ej�wu����L�ɃqUgi붰V�<l�x[v���ۈm��ϳFU�{k{$;a���QH�L�.��m�uO0��1��1�����ql��m�P�K��6ӉzvYDGh����)B�0oI�=nI����uݷH��z��s��;Qv�3<�O1!Y�3���g����c<�m�2�W8ɲ]���f6�h.�U#� +���o�!�����&f���4s��(���뛛¯l�i���m���ݦ����s	̜�-�3m7n]��?D�,K�����Kı?��8�D�,K���C�'�2%�bw�s���%�b����˶�6��:������ou�������%�bX>罺��bX�'����O"X�%�g��u9�Q_�7bX������i�v�\�77x�D�,K�o���Kı=����yı,K?{���Kı/���<�bX�'���{�m��훒f��ND�,�RD�y�׉�Kı,��n�"X�%�������%�`|	2{Ϧ�"X�%���>,�v��d�r��'�,Kĳ�{���bX��}>��^'�%�`�����K��v����	��	��S���*�k��D󰤃�8�F3�3F�,��	Ӓѳq�n�����!.5�GF�j�~���bX��o�^'�,K������Kı=�{���g�ı,��S�,K�����[nd�v36�wgȖ%�`���jr@j�=Q?�1�M�bow�Ȗ%�bY߾�ND�,K����Kı;'�z�ٙ��wn��ND�,K�w��O"X�%�g��u9��"z}�>�O"X�%����S�,K�釧�wr[�d�n�����%�bX�~�wS�,K��w���yı,}��ND�,��;߼�q<�bX�'r���}5N\��������	��u�q<�bX���f�"X�%���gȖ%�bY���ND�,K�ﹷ~ k��u�p��I�������!�N9i��^�I��٥Ĝ�&ˣ�T�r���Kİ}�{59ı,O}�;8�D�,K����_�6%�bt�����yı,O����l�s0�f䛻�S�,K�����?��2%�g�}���bX�'��s���%�bX>�����bX�'oKl�i�K�36q<�bX���ND�,K����KV�&A�٩Ȗ%�bw���KİgKos-6�]�&f��r%�bX�����O"X�%���٩Ȗ%�b{�y���%�bX�{�wS�,K��'�z[-�f�2fm.��'�,K��٩Ȗ%�a���>�O�,Kĳ�����bX�'��gȖ%�b{��t�dr��8&9�jf�[mo0��\�/M`�h=9��\H�˳�v-��G�D�,K�{��'�,Kĳ��u9ı,O�{��'�,K��٩Ȗ%�bt���;�%�n�v�ݜO"X�%�g}��rG"dK����yı,��MND�,K�{��'�?��D�;��I����nHf����r%�bX��}ϧȖ%�bv{����c�ș���N'�,Kĳ�����bX�'�:p�̷f�mٙ����KϘ���Ȗ%�bw�s���%�bX�w��"X�'�"!�ڡEX�0H1�B��)0�A�`E�dH�����W�$�$@���"D��$� H1$!��I"�"�����Cr'{���yı,O�����6�/PM�ϻ��7���{�����yı,K;�wS�,K��w���yı,�����bX�%e���$Cx�G��4�29 _c]��(�&�Ll��А;�%���o�wy���Ggk��͞'�%�bY�~�ND�,K����Kİ{��jr%�b2�_�&Bd&(��'�7D�B�2fn�"X�%���y�����)]��,��jr%��!�2'�o���yı,K>�۩Ȗ%�by��zM�2L۵˴��8�D�,K��f�"X�%���oȖ?���,��n�"X�%����}8�D�,K�=��e�ݔ�]ݻ�59ı,O}�{x�D�,K�����Kı<;�vq<�bX�?w�MND�,K�N��l�5��ۛ��O"X�%�g}��r%�bXG���}8��X�%��w�Ȗ%�b{����yı,M���߿����{T�3�uuk��@�C��v��vx:�n�D,��8��Mn�q��v7!�g�Z�h�L��i�q�p'V��pݥ����l�+nq��;l\�Z���w��lc��-�:�� n�uK�vUN��e㮮�ݹF�孳ی��:�l��%��ƷW��V����+<��n�38wF�]t����51�Q�DT���w~{����}�����d�9:���ۓ��JА�n6��;
�@�m��<�ϣ6�nwwwwS�Kı:{߼�yı,�����bX�'������_blKĳ�����Kı>��N�2��.۲�6��<�bX�}��ND�,K����'�,Kĳ��u9ı,O�}�O"��lK��5���7.d�����S�,K�����O"X�%�g}��r%�-�����!��<TB!n��C	ə��O�}'��u9ı,O����'�,K��٩Ȗ%�b{���q<�bX���˙�fa�d���ND�,Kþ��'�,K��w�MO"X�%����'�,Kĳ��u9ı,O}=�rMm0�m7f���2�^�1t��gn��ݭ۩78t^��˽��uS�Gn��i�iw7��Kİ{��jr%�bX���|8�D�,K�����'�2%�b~>��8�D�,K���ܹ�m%�wn��ND�,K�}��xTA�dKĽ�;�9ı,O����Kİ{��jr'���;��,O��'�?���ɻw3N'�,KĿ�g���Kı<;�vq<�bX�}��ND�,K�}�Ȗ%�b{���ܻv�n�n�ND�,� dO��y��yı,��MND�,K�}�gȖ%�b^��ڜ�HL��Y�����47D�r*uE��	ı,�����bX�1�y߯�Kı/�϶�"X�%�����Kı==$�z]��ni�L�C7PnGT�F�a�gb�6Ϯ�{v�{ue�5`����\&�����Kı=�}��yı,K�s�S�,K���y���'�ı>�ߦ'"X�%���岟f�.I��n]���%�bX���v�!�G"dK����q<�bX�'ӻ���Kı=�}��y���M�`�?��˙��a�d���9ı,OO��N'�,K���{19�N���"A$@��H$"  #$`�@$�"��h	�D)��y�Ϸ�/Ȗ%�b_���ND�,K�OyғvI�v�v�wgȖ%�� ��}59ı,N�~�8�D�,K�����Kı?�;8�D�,Kܞλ33fRYwv����Kı=����yı,K�s�S�,K�����yı,������L��^���d�UDˤ*D3s���M���z�r�=9��kC�р�iz���츎.m�ɻr��Ȗ%�b^��ڜ�bX�'�}�gȖ%�bv{����bX�'��{�O"X�%��S�{sr�d�n�n�ND�,KӾ��Kı;=��ND�,K���'�,KĽ�;�9쩑,O}�NL�0�6fېۻ8�D�,K���br%�bX��}�q<�bX�%�ݩȖ%�bz~�;8�D�,K��;2iԎYU.f��&��	��'w��yı,K�s�S�,K������yİ?��� `�����H�"��1ܑ;7����bX�'{�e;���m��fn�Ȗ%�b^��؜�bX�'���gȖ%�bv{����bX�'����Ȗ%�b{�M���h��+ƹ����b��!�g�����p^kkɮ��Z�Sڍ"��6��&����7��bx{�vq<�bX�'g�ىȖ%�b~���8O�2%�b_���ND�,Kޛ߈L�L�l2�77gȖ%�bv{����bX�'���É�Kı/}��ND�,K��y���'�eL�`�'g�ɗ7v�˻7wf'"X�%���É�Kı/}��ND�,K��y���%�bX���f'"X�%�ܝ-��Rnm�dݶ�O"X�%�{�wbr%�bX�����'�,K���{19İ>&D�}��yı,N�;�a��۹��7s3v'"X�%�����yı,N�w��,K���{���%�bX��{��,K��PA�'�B�S�	'���S�s$v�4����ɱ�Ƣ�r�he:O+�iYN
b����8��ë<e䲪nۋ��6�t��[u�z6��f�Y�Z6]�l6�I��K�ю1�T��vݥ�ώ<�M�ٴ��gGgt6��$�0��'9g\�g�\�D�ۦ��v�^�1�v�<lz�=�ֻ�Y�hʝ㙊L�4�ݹn�rG�n�2�D�=�}>�|���r2m�G���i�ɱ��qq�W+���ڹ���֧��7A�(=ΰ�n��yı,N����,K���{���%�bX��{��y"X�'���Ӊ�Kı>�fW�͹�囹s6n���Kı=����y�#�2%�}��؜�bX�'���Ӊ�Kı=��f'"X�%����,���\6�ݳss��Kı/��v'"X�%�����yı,Og�ىȖ%�b{����yı,O�:e�e��*d�rT�Q
�L��LKm��76S@��^��/}~��;�9��$X�X�����M��z�������������m=�Џt�6Dvc�'1��l�z�.Ё��nNl���.����'	$4^����h�Қ{�4��vX�'����_u���Wn���VU�T+f���p_��˳��ʤ����4e�M��4�*����_��z�\7�ˊ&A3"��;�)�r�W��Y�������}��h �|���&4���9{�8��������6�{Y�J����s��؍F�P;s9ݮ�6�j ͮ8xW�<ޔ�T���RsZ+��c�����jG��}������;�)�ywW�{Ϯ6�$x��Ȥ���)�$^��@�gƀ~�f�ݝ. ��"E��T���n��5%��@�D����H	i����CI�mz"�hd���@�G|TLL<�&��a ����)��8�"�*�`���P-Y1�U�aI%�c���R)
i)�J���?~:��?��$�/�x���C�i��#0��(�h���e��O�q "'2�	!xJ��V�H̭��K����̓cHЍ�H��HYhB�5ME���[x� �D0 �!1S�:�#C�_A�x~�z��Ti��� �����4�YM�Η�c��`��$��u_d�����}��7��=��� ��vX�7�(�� �z��[)�wt����s@�n=����/�9�9�Ǵ�q�KY���g6ktv6sD+�{Y�K-�`L���b��7'�=�}>4��\�����y��)&fV"Vf�,+V��?����Hm�8y��?��M��9'dcxH�dNE�r�@/���[)�_>�@��F�/RKQ����S�o���p�y�"���T�$Q�uQ����ݯ@�}q�y�I�~�S@����uz}l�?�w�~��dEhܻ�9ՁW��\�ك�$b�D/'[���;y�͍(s:H䊼���I��o����uz��4��h��Xd��0Y����<���A�I��6��k�����H%:MZ�77A�7w8��x���|�x��ng�z��ef=�kUn����~���7�.��y��S�o 9I33�fn��5l4Ϫ�9wW���������~ >Ѫ��
� Ζ�0$�H�#�g2w6m�tg&�B�83=����4�c�\c�UջvU�2�󼳶̑�a*�t���xNk����O]�]N�m�y�5�.��#<�R�j���h܍v�ϬU�M��,îv�6�v8w�h'���[tQ�X�=[����h�Q���s�{tni͹��&ފ;n^����Ş�.h`�.�	� �٩ݸ��R�J�"%�;�����{��5����#��Mqk���E��nP�2�ٱ�0u;iK��w��^�'�D5m�'"�<����������h������R- ��h���/>�@�}V��?�٘�k������� ��I4����/>���&�À'��ޯk�m�Y�Aj[�p}Uj=qp����{�7��w�Xdb�@B��E�w��h믮�>}������<����T��I��+u��l�7ZW$m����uԝ�,Mۂ`K��M���C�w�o�r��~�x �~��|�������x #?A �`�`����8 ������&iK3w3wx �~��|��7Ơ<N�*q2>A��o߯ �`�`�`��=�����lllo����A�6667�Ž��-������ۚpA�666?w{����lll{���pA�6 ����߾�>A���߻�� �`�`�`���{�>�ɘm��ɷ7o �`�b� �D� ����8 ��������lll}߼8 ����~�|����ޛ�	����l�����lllo����A�666((E_���A��������A�666=������llla�ϯ�2��6�v�ו�\�����U���p�:���6�n���f�2nL�2�7wx ��}�� �`�`�`��w�^>A�������E �`�`�`�~�ﷂ�A�A�A�A�M���ɦ�tͷ3N>A�����~�|����s��8 ���}�|������Â�,lloN��l�]��,��sv�A�666=������lllo������lA���¡Pr9w�8 ����x ���t�n�ۛ�d͹���� � ؊� ��w����lll}��|����}��x ��{�pA�666>�gL0ˇ�쥙�s7x ��}�� �`�`�b��
�W������lll~Ͽ����A�A�A�A������ � � �'x��?<��v�j�ź��`�����k+�-���ݸ�~�����Y�q�uĥ�_��w��|��Λ�sni��lll~���x ��~�8 �����|�����}�� �`�`�`��f��>۶e۹��nn�>A����߾�>@@�A�A�A�������lll}��8 �}��x �O� �r6>���}��6�\���pA�6667��o �`�`�`�������lll}�{����lll{����,������%#�F��=��nh��]��z����a�"x!Qrx�UbN��@��>��̊
$���~k����s?�=�7��m�p]U�����q�����Jæ�P��͹�mkĈv�qkk�2q:�\H�/�F��:��$�V�p���o���@��. ��u5��CNH�׬�?[w4���zob>S'>M45���3@g�}��r�P/{��ww�@�9�bI�9�����/��@��^�_u��n�|?�J�j(�dNE�r��v�X��V��;R��(Q�����߳�%�[k�ٹl.\�z���v4s۱&ɖ�%ݷ=t��\cZB�Ö���ZM�V�K6�ɞ���6� �`��ڰq�����V�=�훦�l�S�Qu�@��M���6�ȳj�nk�؎��r��=T��;Z88��!���ۮs�8�8��Pi-Վ�뒳J �j,�nV�]�M]Bf�t蜣�҉ IWW����'PY��{6�n�.��e;tK�E���2�g�N���K�	&�SP*��R��(�T�v�X��h��h���=������1ō<�ɠ~��h��h���׬�;������5nf��}V�˺� �z���s@?_���G�R����O�����6��~�5�Tv�!H6�b���~�f��޵`nN�5���BI���?D�T�1ф��ӎ��5H�[��ZΤ�r�=�xp\W��F���ƞL�!Dܟ���}��w�U�r�@?^�@�4sn�M(�ITS�V��;�)(Ja �u΀~�f���M���F�Q$i�f��<������wT��6�8�&��$jb����M���`{���3'y�tD>���="}#j��4D��?[)�{Ϫ�9wW��/�߿����ꋶan��Sj����N�=��1녓et^�rF�K{s,�bNC@��U�r�@=�f���M �����L��#�h���z٠~�S@���@��e�Nbj6(����3;���uqgB����MB��(J"�$��o�`y�}6l��J&W%!�7&���M��Z.��׬�;+nȄҎc$"s4�h����f��۹�{;��,���m�x�J3f���T-�puU�km�ض��۫.��\���5emQ���~�u��Y�~��hϪ�/���+�e�-Fn� ?�{����#��{�@�ֽ�?�#������F24�rh���@�}V�˭z���{:\Qq��hry�Z.�����䘆��`"�EL�����';)�u���D7$&!HG"�9u�@?^�@���y�Z�Q^��:��t�d��Y%ey��LxF�<V��pvx
F��Mk�Q�72b���l�=l���>�@��^��gc��h���f�.�I����˺� ��f�n9��#���4y�Z.�������Z�en���m�H�>U���w�M�v��}V�}��Lb��D9�{���v��v��uz�U�`��bBR,m�"�>�A �=�E�!�B$ 20�$"���`B���T� �.w�a���%!m<2�� ��I0�!	$ �P$B��ċBuH���-%��34��R��X��'��1�*��%2\Օ�D4��`8�����	Q���Tɰ�!Z��wA���D�)�yi'���DL�R$"E� @b�#$c#��c!3���H1!X�@[{{��3ws3͓`\ɲZO=b:.��<� r�����z^�
�F�n�,g6�Sh�i�)�Ū�p���CV��vx��|��qI:�*Ƣ����ȏݥyzvV�,;;sq��PnD΄%a�0�kv���'Lcfr��Tn�ݞ���j1�һ�k;�����u�QcC����5-�=*�-!��xN^Z6c�n��m�
��3�`,'&���<;V��@$����r
��M�L�M�IlL�'��a��K�]�v�=[����wk����r�l=x�n����|iMh͸��yt�Kz9����;M�Ù��&;�n�c�6��v�vQ�{�C�0�R��1�!��j�c&��\h�n��M�p�E�Xp�s��1��5j��u��Zݼ��^�F�]n��<��7\��qX��X��s�ե��P�}�����s�1�n����2�����#s��1�6���mMI��jQ�!��-v6�^��6�*�y�(E�*:y.N�m�%��;b�Lj%:��X��^}uA��Q�l�-Bc�[K��8���M)�vm8��gڃU�]�]���P��rn��uѤ.ųA��.x^7�9�.p:픠����ң=�0�8-� ʢ���t;v���!㋘灹��n�q���cm[��d��lz26�l�㩍N�<�J�����m+�#�yMhm������w=i��\t+q]�����v�$���l�j��g�r�nκ��(ت���2�T� avQ�[T�����9A�`iU@X�x�r����K����걵Z�C�9A�+�W��	��:�94��, 덇��T��u�td7a-���=N��j�c���v��;e�T�2��[�г[ԽS��&P�6�Er8s��{�n��<s�q!��=���z�Gָ�n#���%B N��,t�팱B�	R[�^����:�Z�#5�=�m��4�*�׉:�.v�6��͛��J �{��@��OU8��O U�U㠡z���=P�_����~�Ynن͢A���v��;��P�b ݛ��3�#+�:�f-����8'��cS�Ŵ��4ն�ۦ�&佻r�)=`@n��Z�u)\��[���Ҁe��ml\v�q[�/%��ь��4k���/��������uy��q�^aMw��)�8��2nz8tқ�"[r��0��)�{b��$:N�	���5�gn׽���ﮰ�.:�#tq����n�:m��N�o<�yn��ٹ4�sn���3Ky�Ja��h�h���z٠{��Q1LfH�Dqh�h�k�z٠z��@���rD���#�h����l�?W�h�h<��b9��ID�@=�f����@���A�.~������ʌx!ȓ�@�_U�{Ϫ�9zנ�l�?qؑC[o!��GG���9����[,�7X|���,�'��O%�m��֭����	$Z�����z�����x��86�1�	"�9z׸�$������`nN�7'y���fA�����@?^�@�zS@�>�@��@���+i(451G&�����/�U�r�W��Y�{=��q�8��hNf��}V���^�~�f�����?u�����Ȣ�$�v睧vك<��Xf��svFƄ�Ѽ�9�ڪ�RdnHLB��E�r�W��Y�~�w>���-�]���
D������~�f�����;Ϫ�9{��-�\lȌ���7&�����;Ϫ�R��"!�I(��oM�fwU��)�'���Xn�������^���
�������Jh���86�1�	"�*�W��l�/�U�{Ϫ�;�;FѓD��EX�i,stk��Q����&Q^��.�s��kEt�݆$Ϭ(�#�޶hϪ�=��h{��?.�ڬiD� &D��/�U�g��(lݞ��=��=��`by���s.3N<MŠ{Ϫ�*�W��ﾚ�w�~�������#�h��l��V�w���	+�J!)ݫ�`\]��RE�9#�޶hϪ�{��*�W�z������c�3o��GF�6�u�ݸ��SKm�ʘ�L��X3�e�TQ51�"2!8������@���@�}V�z��W�rn�1�s�n���y�]ZC�8������[�bGZLϓ���܊G�}������/�U�U�@��C�n����(��h��hϪ�9{����3���w}>M�ƔI2Ȥ�y�Z/uz��� �z��(��b�ƜK&���b�n���(�K�w[�(h�oU,;��`�����gt�Y6v�M����E��ae�KB���m")�9�v�v�mj8ѹ<\���O$�^*;U����[<����g7i��9����m�{<��Rŷ��筍�v/y�m�0I]s��t� \/
C��P<�I�΃��<몳�ΰftv��;�[�"��K"KGa�t���_A��EU��^����nt�-N)�I��8�7�*���?^��׬�;�)�~��t���@BpRG�_t��~�f�}n���^��.+���%#X<��9 ���_[��r�W�^�M���N$��q���/���9{��/t��~�f�ʉv%��H�D������Jh��h��hg���ϑ��	%	#����ePs�y�F�3�U�4���7��.(��t90X�F�R?�}l��^�@��s@��^��Ǘ��<O!��� �ޫ���B��E%
��\Xy�:��h�F4�M��I4�)�r��@��� ��f���j6��')!�y{��*�@?z٠_YM���6'���ए@��� ��f�}e4/uz^S*�&t�����8��Y�m�x3�jx��`��K�vΌ�\[MznX�o�����h�S@��W�U�^�yܸق��ē�7&�}e4��hwW��Y�r�.Ʊ؄�x�"RٽV=ޛ):��%p�$�!Q�ޫ����ɘW�3�dnE#�*�@?^�@���/uzy�����#�׬�/���9{��*�@����U�Xbr)�8䄐�r6L�*HƮ�%��X�Sf�z�q�ݞc�H��47E$�/���9{��*�@?^�@�zʚ��)�rb�/uw����v�X������4�R��ए@��� �z���h{��;#�ē�""�C@?^�@����77�ð��(�/j��;z���P��C�7&�}e4^���\X�z�ݱ2C�UHj�Iȉ�K��ѡ�h���u���O�d�n��k�ͮ.��j��5�D%#�I��W~Z���l�~A�}>4\y������dl����)��Y�_[��r�W�r�`�Zx��p�޶h��h^���)�{���F8�&@X�@��s@���@�}V�z����V�m�O�7&&�h�k�=_U��f�޷s@����<�	�4�n玬��ʑ�]����!�v�8�����L� �i��t�^ήYfI�mC[� ��aۀ�m�X6J�zkl���s�83��e�S�r1F�R�;Y�t�x��i㵚4۞Ul�Z������]<��ص��s���3�lb�[����c;���;h���;c3��;�>/G6تn
��Pꎱ�w�h�F���3�����;���z/��c]���gYrv�+5f�I��u9D�X��3����]� �㍓s�Q��� ���v�X�ֿJB�
�qT\�$�F��rE��f�޷s@��^�������ț$ ,q���;��h^��W�h��h^�嘔�$I��9{��=_U��Y�w���?s�n�����G#�=_U��Y�w����Y�r-����1�<1��L�WZ����vP���rz��;7�̭�c��p��4�Z���z�������Z��kdoi@y�@�[��H�H�x�)������w�w�@?^�~H�_}�(�Ʀd�<M��*���=_U��Y�w���?_�F��d'$z��׮�޷s@��@�\��R0�`�rE�~�w4���/uz�����V���/n��Z�է�S���ֹ!n3&��nL�0�\�\�뎬�m�廚/uz���׮�qe�i�ʈF�#Nf���^��z��빠w���?s�v&�HF��@���I<��ɅCA��_)�8Tt"A� B+�A#!		 �ܹx/Ie�� $'I(/�
��A����B�A�BP��P�$��F�f��9��{��8���y'��1�#�ѣ��$	m�@F�B�d!$c ��%�!
�.D-YA�$$HCVRc
�!��( �MQ�����x��������D�s��#�1UG�t��
����K<�}j�7���׋��������b���]��n���^����ץO$j7��@qI3@��`k��3�y���V���Pvۧ1�I�١�k����������Q�[!��7��K�譺�q�����r���=_U�{��h�w4��n����8)#�=_U�{��h�w4/Z����5#�
G$Z�[��w���<������/\��IST*�*�uJ��
}�}�`k��l'�罼�򮂱P��D � 
� A`,�H�D"��,�.,�<x�#L��9�/s�zk���sx~o���<�K��f9vf0ֵ�6��ˇ�f���9���H�5���g�J~�����׬�;��h����w0��̬�V��[��?��������:����^�߱#����GlmƓȤ��N����q*���{ ���>�5�L�x���r�W�z���~�f�����?_�F�S#ı8��h��?^��z�� �u��@��Bb	�=���ٙ�wm�7E�Y�4nۍɲU�����%E�hM������CJ���N�O��q���&��9�p��]���ͱť7�u�m���l`��lr!�u��R3�t��.�:죾��g�N�W ׵�oVL�.�D^ش�ن5����[/�󺼆-�D.Cu�M��\n�vm�[��ͭv�s���<��.�Rv�vR+�EYJ�f�{���_F�M�ۖ�\qt���%�GCְ�I���;<
�Ӧ��ɨJz:�Q��^����n�w��ץ4�"��y$Y ���w����Y�z��@�z�h^�<U�C$i��9{��<�W�~�w4���~�C�Ֆ�4���Ż�]�ݯds8}~��;��h����1������b���]��n���^��z������`�4�0D��\ݎ���:�=c�GL�&������T�Y���<�ɠw���{��<�W�~@{��h\w�	Ħc�,M��{��5��)a3;��=��`nwZ�<�qtcsx�'$z���빠u빠~^��#�E�nG� �rEa��Ｌ���`y���Ӽ�nEq$�dxd���]���@��� ��f���uf�$�G��\Vk
��y���!D�9R�_:�%�3�v�q1F�i
1�873@��)�u}W {�g���'���n��F�nff��8<�].��� ����:��}��|����O��3�Lͭ����I'�������O��	$`E��#'SH&(�F$��)�,��E D�����ԔDU�z�,���ܕE6�h�ɡ��߳@�gƁ����[��^�h1L�Y#��f�q`gN�=�֬��V��|''��f�1;�f��N^C���[ �	Q&��rto2p�l�v�oLrp٫~�ߧ�v�zՁ��j���q`k4�X��x�G$Z�빿g�ffbE�W������WWuIJ�)!f���
�ͮ�N����q.��g�~��-x�bhh�Dj4�h�k�oM�{w���%.!Fo��/�#��ń�nE!�y^�@?wY�w���?wJh�v�$fX�.�AoC9���tt�;/����bѵ26�v9�w5��w��᷂qO�m�����;��h��4+����TQ�mA����z���t���z� ��f�y���Fd"���tg�?<�U���G����up�OL��1�NHhW��?w]��7��.���~o��41�jA5SUN���Z�>��.����gu|X������,!#Q~��}g9r�J�l��Շ<�.ݰ\�s+nݕ�ۿ����g\l���;*0%��6wV���%�������4�iy@�2�k[�Hs�"[8�t\��۫��J�����Nظ�u�A�;K�{�+= ���M�FoE{]v�g#sG�2����a7J�׶��/�.Ue�)���F��sn5ϵ�-� f5t��f�u�wn��N-��][�����rWг���������;#l��l�u�;��$nv�6y,�j�rX����@�9�}����������ޛ	WUU�?7:���FT��Tә�`{v���6f�_w}j��۹���+���I���R�YK ��U���j���q`b|��y̧4Ct檨�n�X�֬n���h����Pi�E$�=�w������=��`fw\PӑU6ؼ�6��f�H,�����A/\D�c(�na8��RI	 �ƅ?�QcRf���U�~�)����;�w4��LX�Ɍh�&j�����z�B��d2����oZ�=����%��9?�K�J�L��$Z�~�{����U�~W��-������P	RM��s@�Ϫ�?���	wuuT�7?����x`���"5�����>�@��W�~{ϫ��uwKީH�^R�[����1u�5�籺�W�r��Ȓqp�mfx����R鶺��Ō$��rG�<��=�u��;�w;? ����YdI��Dӑ��� ��s@�_U�~Vנ~^�t�rQ.GEM+wzՁ��fDB�"P�DB'ú��j���l*F2���C�V�w�����`{w�X|�!�~���~Ջ!���r-��.��~ro����~�y��{�m�~F"�u]�Bf�n�Zt����x��{s��z��e��6td讧kI`�� �����s@��@��S@�ܸ���F�H�rh�]��uz�X� �m�K���H��т�J`�0܉��V��޲���4{��k俫����n8��?z�h�n�I�����>Au ( ���{�rIؽ�V}M'�j'$��~�����׻�`{:��<���p�2J�i��S��1`�s���n.�eMS�*�Cvy�8��#�cDnM�빠r�@���������I��&%B��zn�%�\���$~�a����{�]����Q̂�A9�����~����s@��^�����$	I���٠w��hwY�~�)�Z�V?�ƑH�rh��V�k� �wU��)�P�	 K��JD�S�@�0P���$��D��NR(�p����T�# � `�R1L!H0�����ol�/��r����M�I�/	t��"%$��`���b�.(p�H� A���P�j�!	e�4�`�N�ָ�+��`�,"HT�� �jK+���$��h2�A.)$�2�p0��u�E�e��)BN*oU��8p �#�0�BYP� G��"đ������?n+S����/7�Fg�WD>^��X/O��(5q�UX�]�;�	�e�j�����e�h�����W���8�uȽ����!�4�@�j�d�[�$�ed���@��u���Bh��m?X��ȦD��(
���x#(��Z1���dz�F]�r[G��\����9��9�v�(��=��R���R�������5�$���չ�n���q2�;��v��0��E�Zٺ嶴�@������α���M��T��1��)�7��r��jF�kY��nz�*�&얘ٝm�1��)p!8ú�;b�T۳������Bu�m{R�ƥH���|�����*�<��s�d0�TD�tE��9,���Ԝ{{h�����E6 N�9��6:wj�:z�a���7h��N���g�[.wGwV�V^qm�,����my��vݽtrӹ�'���ʦ��W��`��lfsOeZ�tpA)j�<X%�հ����ɗ��i��-*���^%��l'a�����kOXs�A竨5��A�s���ɝ��*3�9�8:0�5��>f�1�nV��7��67�����l��ۛn\/�.��!�K3��]x�g!�$����%ΗF��c.M��ڸ�.ml)���e9�m֡�u���͝�*�ф� �cYq����	��n�ɲNz��ұ�Ƭq.\��=U���ώ�J�3es�&��@�<�ij�줹�헡h���)�U�4'n1-� ��t��*��7:�'�<�1r���5i:閤@H�M{=N݈�Z�8ۅp�k��aL�w���Zș�i�`�΍����!=",�n̑O<��ʰWhme퍓2��ۅ�#�����K��&�R��*̑RJ�!kPF�I�c�'1��Vy|{XNۣb�m˩P�̈́���粼Wkv���`�����]d��,N�vI����Jq8v��pܵ�:g��4ݫ�����T*�V4�I���3L�7)4�Y�OC��/ȩT�ǅE��g�0S����s��~���nX��l���nV���]q#�\�b{v�gE�5����l��[;Y��Mq��疔��1�n&��*�,6�4�/p�tle��H�WR��N�O/X�p��m�Z1�� \��ՏZvj�[M�dk&5aOmr>�v�����>�����w\�MU壠��rf��Lh����?x�{���d6�f5�ⱝUk�+#t��w��^��uGm�W�k�^�g�9TЌ�O��n��[�D\>�u\�d�)G� ��Ng _��@��M �m�z������@�<��G$z�Jh�l�;��h����bG����7������8��x~o��uiUo�@���?yгX�4,���@��s@��^�ץ4��4
�Ԗ%1���E���/uz^��׬�:���9g����iF%$�xl��p�m�72�n��2vB3n���b孪�n�dx��1a ��@�YM �z�׮���^�����$$�i�l�y�{���"�'���\��䇗�<�=��:U��D�I�ZU���cNI�w�������e4��4��CI��&A��9�/uzz�8����������pb��ZI����@�YM �z�׮���^��[Ii7M�cM����c:9����t�<�#�,�m��v��<Z���@prHh��h�w4��}������^�|h��}1sLl�I�~~}].��!�9���p�����	
'�$Y��r�W�w���~T�@��ݞ����'�w��~��.C��NG�w���~�f���s@;�f���4��Ȟ$�jj� �oU��#��X��X�\X�j�c�	�7���H�:T�^zt�L��ѥ���=�Ɣ:t��s�9��urM׮�W���e4��4
��n��D��r�W�$[6bI~�o��I���K���eI�6�$��䒵�-I$���ߒH��MI$���ߒH�Yl��7���䔬̞s��H�uo$�y��?��]p������6�RI4�I�����$[w&�����ߒJ�(�$����~�???>�[C�s�l�L�Ved�7-�񍌢����t�k���AWb��]#$2)2jHJ�Y��I[%KRI+�g��H�w&���E��P1�c�D����~�b�uu��)�7��$��i�$���~��]�t����$�iȖ��_���$�~}�%*�1?9���%�K�I[tU�b�"���$��$��5$��u��$�](�$��z�ߒH�7^<L�#�s&��]�!*�Q�M�OoO��goZ�m��%��dFmʷ�m�*�y��v4v+��*�δv��4�Ξ���+k�1��>;V�] ;*@=������W�֖,۳��1���@�\�ݠ]�GA�%��928�th[%��dy9��Yxģ��
�qٜ�q��=��]ۛ��\��ݸ�,q�˅����K��Gku��^��sWS�9ZI'ms�����v�z�����t�H�_�w��{��wY�W�^^��ݤ���Dt^�v�nn�v{p��W�MqԩqU�tʓ s$m�I'�$��χ�$��g��$^��RBW���	s��X��@[���p�I����ꫫ��J9�rI%$���$׵�Ү���3���n�Żc2b��?~I%��a�$���ߒJ���I$��~����P���ɑ����m��wu{ͷ�k����ou{Ϳ�P�!L��z�o�W$�$U��檽�ګ���W���$�z�MI^�~��?o�����&��y��v��g��F�����{Qmʝ���{GJEӪ���<��#�-I$�[?~I%z�5$��l��$�IE�$��.,1ȱC$n9?~I"�Z�H��B�6�ou{ͷ�5ö�o����T�4��6A��94���~�5Ļ���H�M�	�7�i�J֜�dm�I$�/>�@-�h��@-�h��RF��r8�6��	jzM� rM���p���|�6�ӓngl!�q6�gI��we4L�t17��9�b�u=2����oxͽ���O�I���v�&H��A��h�f�� 9&�����@/�����1d�d�xH)���w��owU�)P$��
	$(��(��;z��7������7��3R4�Z�l��f�z�4Ϫ�-u	\Xc� ���M ��h��@��� �h������d��r�����ݗx�m��r뭣k���ݦ�J4�ˬ���[f����@;����4��V�Lj6�rh���٠�@=m�,�b�Io )�ȴ�٠�@=m�������`܊�6����~��}�Оw=�䞃��A\�"!�9��}>���6%1�#ı�&�u�h�)�m�}�h�O�0r4�]�˪�vW��yݝ1�9�h�v- <uoS;"���9�]��B�>�~���M �l��@:�4�Uq=5&1�#�C@:�4���������]]�CC��*�����f�����@:�4^��:۹��\�v<x�G$���ץ4m�pJ�����sx͛ji���-�Q�#�@�Қ[w4�Y�m����ʴM��#Ia ��ƃz��O
 p ���c�z�&�%�hզی��ݰ�e$:���I����lu��>e�sзj���;[n<Ě��ض]��������������ڃ��rrF��nD�v��s�к;{��"^�"qtTZ���e��������r��n-M�����rbH�]�hV�ع���wZ9�U@�j^d�vnP�yX5�)�N��k��:7Vx�#K0V�;:q�C��bd���$<��ۚ׬�����~A~��@��H��#�i�&h^�@:�4zS@�n�{�M�O�1H�,nI�m��)�m�׬�=__�16�,$I�4�)�m�׬����j��cƤ�4�q�h[f�u�4��@�Қν��2�7���U�j��@�����4�q�l��a�(hh���G ����Ăb�g�/�8��wL�{��4���i�1�d2\˻��O{��<G"UP<�;�of�}n�[�h��W�&5�Mޔ�:۹����٠U��,m�h�(
Hhm��z� �l�-�M����rI� �b�� o�x��?�q�8ͽ��~~�� ]���Wg�y��l���O�Z�a� (s
�5.��Q���+k�:���u�}��~�M����c?�	���)�m�׬�9[^��\[1�I�iUMMQ`��`��g�.�q�sH[lP���5ҋ�� !��r����"�%%��&S4x��V$���DB[	i@�����$$�?$�D߿$1�"')mR��JW�"��K,�1M��&	)
X�v���J �u�K1�F��	$	DX�c��i,b��	Ȥ�b�)�E�u����sGyLc ��� �~� B@�� 4.OR���z���)����5��<b�'�$ehR1�3"��6��{�0�*�Oʶ!T�%��M�z�p��A��xNO߉e��]9��x������!����0BM����as32�%�)i*�dV��L�1�D=ˁ*`�<��j>"����?@���=G� �q�G�f���'�Қ#�.�V$�0d�rM��}7��x7���uWuI9&�	��S6A�Ȥ��٠[e4��@-�h{�gM��P#�<�;"s�4�M]�ո�N�k���@���=�%�j���9�&5�M�)�m� �{*��5$�&*����6��RC@�n�[l�9[^�m�ߒ=G~R17"�21�&h�_���ڴzS@�n�޷Zĉ�"$X�sUV��;�k�{�Հ�ED$���D�E!�,�s�o$���z��S�`�NI�[Қ[w4޳@<��]UU)����YH�AX-����q%�;qnY��F�ݟMxzuƆ�s[M�kX���s$HrG!���nh�f�y������a�4:IҊ��En����������R@��H��٠r�`ݍ���D��9[^�oJh[f�[�h�WS�1�ƣdrG�[Қ�٠��+k����&�c��$4�{��� y��~�pwVy����ߙ���=q��� 89s�xM+�wڅ�����ܣ������F���k2cn�c����%y�x��묣�K�n��5����=���u��s�,�}WcEն����]���9�d�c�F�.�`y����<��Kˊ��X��]*=���q���`8��9<��9���S�7�.���v)����D�e:˺��gtb��(�J��P�<	ܞ�0u(t詪wC�"sd�'c��nF,0@nܭ�B�v�'�NIK#1�&�~��4��@��4��@�[�X��ȌNI�m��)�m�oY��H�Ϗ��,mFc�D��@��>4��@-�h[f��-W�mID���h[f�[l�9[^�m��9�v*����d�rM �٠r���)�m����]��I,�t;��
4�s�n�gvF�c���}�q��1p�u�tœ�6A�Ȝ��/�}4zS@:�4޳@��ز��SL�fnnnrI�����P_��Q�l��٠��+k��E�-�6�q
��٠��+k�-�M����$Ȍiɠ��+k�-�M �h�F,U��D ��h�ՠ[Қ�l�z�6��w��~ Ɲ�3Đ 6��N��%��Z�l���v��Ȝn�q;-�u�Tr���܋�}gƀw[4޳@�v��j��cjH2`�C@;��oY�z�V�oJo���9���W$��J�iXv�X��l�U*P�&f~iޔ�:����s�l,ęG"rhVנ[Қu��oY�~��eq̒Gn8��-�M]URrM� ���<�y�~���7w.���*�F씌�z;a��x�s�6�Mn�u{ve���S,�`�1�)�Hh[f�[�h[f�oJh�}T�H�)�Qӓ@-�4Vנ[Қ�٠~�0xV��LjI�r��ޔ��� ���=��t�&23
	��zS@�n�[l���#�p�%bB ��@ ���HH������6��}��vw��[1�L�<��hm��m�+k�-����}�dpc���c�Vۧy����6;(�O(l�ӻZ���8�f���[B��kM�[�_�I��o8޲]]_�$��
�)ѕ�D�29�@:�4]�@�n�[m�����o���v��r�
Q,����L�pm�q)"I7�jI��~�i�����7"��� �٠r���j�?p��$�LQ��Ɯ�oY�uv���h[f�s�3�;��)�i�g��\ݕ;��,��^},�2Gd;qs�t�۲Wv^]�w^�&m�78�b��b���n{��COt�v�u��3�5�;&���v�L�x"�bv㝛�m+��X흅��FY�S�g66��ʖ=pa��N�{T�< rGFm�� ���L�`���;up��i�Oܚ|mNӼ�V�d�T�ދ���R���s.�ܔ��$\<��&�]ܵ�瞶9���sVZ�޸䳍�U�O�rN�z�DqPU��=�;F��W�m��������@:�4޳@����<D�<�h���u�h�f����e-�c2I<��h[f�[�h��@��4�ǋ��H��	�oY�m��)�m��.v*I�q9�@-�h���m��oY�~�B��?�Ēa��Ct0Tr����VV�s�pIذJ���crjD�N94zS@��� o���@I&�Q��Kp�VKt�ݜ�w��x���y8�O���@>���-�M�U$���Q���@-�4�f�ץ4�f���`�`O�LjI��4�)��4�Y�{�˦9�D�<M�4zS@-�h�� �ٻo�w��{�����kT��쨷&��m�Ts�����iό�9�Ӫ�Yv�t�g�n���	$� m�����mp;.���ㄌrM �٠Umz�ՠ�4.\�6T� �f�����p�k��UUW_UU�-�}��}���=�����H�crG�uv��w4�Y��4.������LnE�^�s@��z �����>�����(��B�3��ܕ�؛̳[7��;N�)�M{vF݈H��<S"������|��= �l�-}V�z���|
��	��zz٠[Қz٠Uz��L�d�(��h���^�h^�@/[4e.\،RG����8%Z�O��"�g ?7�n����R!- �@$ ���)D  B�
�D$UR�V�T��,i�#7�ϧ$�g��}�< �<p�#s4
�W�Uֽޔ�/[��{���� ���0nZ�*�ճ����s������kd��nK-�m�b�"KN&����@��8�o~���As8<EL�����ubŻ��~�t���7��9� �l�<��X�����LrC@/[4
��@/[4l������!!0��orh[^�^�h�M���������6��@/[4.��G��G6�/~�p�uuWv+�؈*+��"
���"
��TW��AQ_�QE�E�E�� 	P*1E b� D�0E b�Q@�TBE�E `1T ����*+���*+�* ��� ��E|DAQ_�QE�D��TW�TAQ_�QEЈ*+�D���d�MgX���Paf�A@��̟\��|=  �f $��  @ P �vd �`�  f�+� $�� P)J�I*�I  *  	
$�J(*�*B��R*U*� �R��*I(�I@PG�   @     @1� i�@͸�s%�L�=N��o��g��}����y=u�x޺\���{ye�総�����z}��}{�=��/vt\`����}| >�#��}��:��k�_ ��P P 
 
����S�ݤ�W��Ǘ��g����Qxt��A���ŕ���wD������}}y��� 9���Y�W� �3��N�}����۔�������w�o7��{�|�o��s������  �  }P   }�L�����������n�|n���C� ���/=����Ϧ�{�^������}�>����R�wn� N-)CB���uH�&����P�� @n� �   @p  ( 4    3�*]l�Nvu�bj�@  :       b 0�K;r�S��H\J�!�S 5B��hue�)X��V6�C  ��V|�jse� ���=�u/x�n:s�Ԝ��{�t��A�p ���܏n.v[����/���� D�    ��я��9r�k�}�zy5N��n-Ʈ{k��t�����s�V����,�w�|  |�|�u=��}|� }����o3�{/�{���l{����}��^}Ǿǽc�}�ﯞ�����(0� '��JT @�=U)R?$�  "{R��&� @
����ڕ%H�� �B����5��O�?��?�����������n��g���їD�{?�PU�a�2��PU�"�
��TE�*�����+*(�������HN�}�۷��/�1֟�?����������9�><�<{���{��kІ0�!���h�m6>��>M.1���ٵ�tAbV�{gbT(;��\(P�.*r5�U��d�G�35���ޅ���&r0$������$�L8;C�A����>�ʳ[�x�>�xx��F:6p�������8����N��Rѷ������8i��������[7�3��➉:�<0Ӵ$��o04�'�b�bC6�I:<	�[��X�zY��<Bs\#���l�>�	�{<���;s�d�LT�N�疝y���<�Eo3=��H��5f�5�f��p�X���Vb0bhcY��F�XF6F:n��Ij�#{���4i���ְ�Fh�3F�58�Vh,tAa�Ѭ����Ͱ��N*4r}d�� ���6�g�~zC���t3�xk�|�D�x#��vk4,2"¸��n��l��q��L���2bA��0�f�U�,d1v�h��4@c�|���pѱ��s�4�h��O�c5��&�<��3DE�8m��h�pp4m���e�O�h�љ�灡=�zٹĝl�+U�5q��v�D
W�Åp��Z��H���5�����K5E �%��\dN�^��bQ)yQ��WX�D]���3r�WDr�@��ݐ�E�FYH:D���L�,:#l3�-A����p��1���i)��qH!!���I�iCiŘ�4l�8i������Kl�=7>⢁�����
b�E�h�ݐH"6�Z1�`���1�h��5f�ϼr��M�k\�Y���	��YBB������F6���#��IK228�i#\ב�Ç�0CA�l�f����s���Dfh�����?���h�߾9���������`,�c�$�Ŀ��8ﶁI�B��ū�F���U�n����B��������P��?
�i;�l1�|�~���������|@�ྀS����c���H-o�|�N\`���P!9o�|' o���r�	�m��r��U����8��0�sO�$s��z>�c�s9�C�41a�a��_B3[.s^�����Kc�lT ���6�w��KV
b���U. m��(����f���qto�p��Dkg9�q�|�!r�@�����`�r�T��#o�tS� �ɋ_>��pc�����y�	��u&$a��o�p�M����e�cxFǁ����.xg9�rќ���sFLo$5�	�a��3V��5�xFl��Ahǋ�2�x|���������G�"�˜��S�.���*t����q���٠�ӨsZ�k��Y143����&��׉SU����| /<���w�������
s��P��8�d�u�ļ5�Lf�,�\�3N�p�A�N0Վ�0c�q��L��f���ic1��	Á�l�1�i#�ki#�0�����<8h�4&�����1]�L2b��		���K&�����ib0`&�"	�6�M�d�2ãf�q�mtœH0|04�	#�A���HL H�����)%R�)"IK����M @��,8L2bh(!ȗBm�Px��{�M�� �H`F��"y��6qd٠�4����荕!	��tZ7�Fh��'a�$���l�8�a��#zJ �A:۾PA�i,59��4��7�051k|���0�kf�%Q��g#s�i���k{80Ff�6�4�h�D�7�㱰�p#'z4�f�����[6N�ұ�-�4Q��qѲ޴�E���1���gc�#Z �og#)"ӷ�oFju8�kTƶ�,l���6���kKa�(�F:��{������XX&.QA����+4A��,_��8���3���n&wl�#>r�iG3��A���LzTNk|�c!��xxp�7��ou�Ìf�q8��z�����g����,�|��	$�&���{���'�4����`�i#1���6h٧�a�z�6a�5n"��Q�l��F��<7�y��oi��	�f�l0ӽ��D�4��F:�	�`����Y���������FÈxXk{�A�Tkg)O6|l�[��xI��6�a����c�$��D�4�$#
�.�N�[_~��3G�{�3^��������p٩�^�P��̄�}p؊�:I���&��\'[G��u���,t�,a��\j���1��y��F����4�
f�q�0��;<|Gc4)��:mo�#>͟sZ�{�<o5�4�p��>������]Èˁ�i����#.筚�Ͷ�nsA����ۯ\!�0�0�����`K������sE���l,I��1�f����햶�=<ݚ�If�4FB�S�8�ŭdё��!��ai��0�Z�ݚvHfG���<�o��3K�DVkk��8f��yz�a��l��f�Č6�ko�������}��<9��
c3Z�N��2�,�c����ێG=��>�<��������ը'��4�$z�F�����n|���+�dfdy!Ek�ON�a�<�yf��k|֋�F&π�<C[�<����sÞ{�<gI���I�����;b�Ś�)1.EO�E�Y�lǱ]�f\{x��N�T(��RH�I���Y��c���15}��0c�1В���I( *���8��b�D�_�A��T�@ݏ�\
�
�^��f&���7�D��k��p�
�[4p�)���2�f�s��^�il�bX�v��}4FZ�8�f��-��'CfG����]<<,�Vl�f�a��՜�F3��"��x��m�$��¬Չf����k|ץ��h�=�VzA�O���yHF���4��'��^�8�b�����I�0'�łM�'�>����Z�a���Bl���ѡ�4j8@na�$�~M�< ���������c�ϸz����z���]c���y�>�ݷ���%�L�BFϏ@�4l8����ls����O��͘��JC�4b���C����w|�wa�}�c�/�k�Z,޵����A�O�d&�6p�gƹ�d��5�K6aa��=���~���	#@m��FMĒ�%��tl���6fkiFX��<�_g4�s4��6kFw�7��76r��TRe��3��@�ʀ(�D���D�ض$l�ӔP|!1F��9V�`�����`'�YV�1 )������ 催_b��.�O��ӀP5�>ᇆ���� �F�Fyf�pk7��$�0�9�f�0���&�r��Ί�EELN�T`��"SK#5�������Ӷa�pO�&ki��)k��ѷI�I�E���u��q�k���xo�]�7�q�<,��A��\�R��5��=>K��F��mk|��0��Ϲ�m��DQ�!�l|*�
�F�W��
"�����@�N#q|	;�yM����s5ɵ�`lьf����#	A�ٻ�O���G=Hg���7�ޘY����m�a����K��s9��0#�oLt(�>��`�8��83��a�#A�F2Ӛ6H0`$��0]X�����1��FBP6�58ht����#4naǉ Hx0�����R����SB��K�@Ę�v��yă&�HX1HŁ1FFLA��!1q`h0�I0��q!�' ��l��p��f�D��H�p�#^�O���p#�N��4��6�4N�63A��1���<�s�XxY��x�0����x�8�ێ{q���{pv���Ï�_��]�������r|Ā��� iA��L��������Vv�¼�^��;���zk�c�I��L�:�v"=3�.`��'��T�@��uM�*���U>R^^�lc�*5��;�=]7�(�!T+�qeFE���+�MU���Ny�x�Eu{�X�=��)��"�y��@�����U��/ Ɉʨ��L�+���25Fv�]D��"�}鬂r���6H��U�\
�6:k�&A_U��&�^WY�T�:c�IxY�:�K &�VO�M_�вP��wM�v���tGR�#�S����^G)š�{kv�FT�¨yYx�l���ɕ���*����\)�b�|��j ,����c��W���al��"ȟ,S���MN�P��  ��       �x�g4�h��;w'C���n��x2f]����J ���g�N»sV�5�.����G.��"������l�g[:�2�iڂ��p&bl�y����roF�i��i�bpvc�T$J�jV�!�Z��^ا�[���D������ճ<]��鸉��W��ɰrndw��)
Rf�zA�o)Ҥa� ^�:u�Y.D�^h�� ��U�X6Œ������1)/O#��<g&���7�h�Iu{\8��寧 ��$-�l-������\��m[ �`wF�9t�2���Η�r�ݔ8�q'6[mmP��PeRX���Gi�Uk<�r]����x'RL�K�@V� ���m&9��8��n�94�Rj�j�U�e٨
y�ùm�]��(g�U[prA�5^�q\��f×�!�K�n��u��+����/=T���(�&�U��3OG,X¯R�ѷ�����k�띭�.0�qU�n����W [�+� ��r�:*���C�^��շV�e���E�����z��%�8;f�s(捹��[p�V��촤փv8�`� �T��g�z^���'+�v�7+�|�IP�r�Y�m�tj[U�l��up]�v6j�r��<5WA��N�����E���l�j�ϥ9���h�%��N�oc�z��u�>2��6[A���&�8[eM+Q�/+�aG�F��c��nj�<\:�󗏊��:|%�/N�pu��ڶ��zÍ�kiV� :�V�LDZ9��  6�۩�*���!��&��S�]ú3�h\yb�[���̽=!��B�:%$ݭ�@im ��m[��3��I�kXm�N���ݭ�Ёu�J�]*����kQ<�������� p[m�5�q��@m }��i;�n�ۯ��F��;�[Gn�mr�˔�tU,�!;J�W,R�UJ sm�YoA�uj��	 �a� ���^�ɧ�g�  	��-���"M�p ��W�n��( m��$V�@`|�,�iV��w\�V�^�5�j՛��vѶ���D�1��<�'[m8 ���۶�� 	Ͼ��l �D��H[[l Ѷ��|�H�x7m]yql��lt�i3�Hx������H�m�sm���i+`rP�m� �ۀ� tAF�Wg�Wey`�ݍ�"�J�̽+��-U@(���&u����6�4�.������f��,�.Z/r�����l�Xၮvٔ���m9n�ض��	Ӛ�hM��	m�    ��6-�@�  �hH �H 8  �8lְ m  ��� A���  @���6}�)l����K@ f�e��}�Kl�1�j^��p �-�   M�m[��]x��		K�8 [@  �����m�     ��m�[dl|��]K9�I�a��l`����m��m�	 �nP�sN^�d�lez�����u5��@� �	ݭP[>� ȰP^������v�lh� 8�e��� H    m����f�� i!��� m� l	    �`   l � �@ �6�[@ p �HѶm�h_^*M���*]��m�� �[���8���o�|�6� [%�-��ke� h��  ��h��l ���i8I�m��YR�N��rH�v�IY��8 کF)P%eKn����gZÌ�UJ�]��R�kԝkrI�� �`m�m��� �`�����n�ۀ � m���Y�� �r�dݵ�U��+�U �Ԡi� -�m $ �I6-��i9�!"ڷ[l�sETLʝ�
y�UMSt���EM��*��6�Ǥm�a�ܶ!�!�lpH඀�m��@�Na}��, �l��J�t �R�-!*���mR 3��cV�5��V��V�)�+�JJ��Q��qT����ڔ�V;l��q�c��8L[
�9���U��F��]���HvvǬ9WE�����n7Y��$�!��6Žy��z��@ Y4���Fѻ U^N,���7eS����� G;4ײ� p��ܗE��� 6Z����nAn�����F�8�(U��� F�  I"6�k֚sv�`�	y$�m��oE�%ۖ�(e�@  ��\N���K �-�$�մ�L]�u�	zjM�[I��i�Gnj�P]UJK�&��#bH��ѩ��B Ns����/I�����	Вs��� 6����6�qd���� &u�Aٶk�����ev���Wnv�ӭ��Z���rJ? ���+VI�h�Y�n�I Nj�,��mml�2�*�{aj����Z��J�-B�u�A��*�WK�:zky�k��76  �Z~[��:�l C�knR��:^�Kd��e�&��@-��l��צ�g^��]�  p�"�՛r�7H[�F麧.�%���Cf� 9z��4�&��̲�m�
���8ݺy��'�1�VK+]J��U��R��oӝ[m��V���^�ld�ۣ)]�I0VP9�@�i9�ĭP�+k�����[on��P�a�K!Ëi$�2��f�p ڷn 5M;.�z��� m�^�I�p�[/�j�n��ڪ�6%�ȡ�X8��L���;q��t=v���  %Y2n�ۥk�lX��&L=m�TJ�˱-*q���5��)��ɇ����Hc��mR��q�V�ۊk�pv���� �o�l[A���h-����ZA��	2]6��v��i�em�	}u�:����vv�� ��!V�R��� 2�fz�A���>k�<�\[d l  ��+�K�U,�V��K��ieUj��ZX*��jYXv޶�q �l��uʵ�^�ykgf
��z��� 8I�U+$	s� F���s�+-P
���<�- 8-��M6�U��`   �����sY�]m�[%m� � U�[���"�΢��']V�9$�_9W���R���3sE+�4�u����8*��2�b&�m��Ė�����O�Vԡa�5m�e�uJjj��mz-�cD���Q����5�d�ڪ���]��qL�Rv�����k�9�,��t���8�b[#�E�EtJ���W�50b@  h��%��+6�mU�[2��@ �m��X��#����ce��i�n�֎9%��B���H �F� q�V�E���HR��۶�pHm�k�A#n�A��!�d[R�ݶ� ����j� �nE�I#m��շ�� $9��v�� 	88/J��� �� �	 8 �Ͷ��A������j�R�H�� �a�ݱ��ۮyz�@ �i��WnH -⪗�UT=Iە��tF�����B��}���mn�$����M�cYS3�p[Tm�����5 $sm��n�f��mI(W]J���J�(s��][\��\�P�@J⫩l��p��K�p����;e�]��f-�4�wm�$ [d��;�b�3v���D��/-U<�M: S#Tm����LHH$mY�au �^��a����j����)N�l�H��(/WM@�m���ݾ�}R�4�.U��gM���P�X U�Vj�n� 3l��d� Y�F�H�� ���;_/���[@mS����Y�cjV�YZ�}����i  ��m�U�d�#�IR۴�mr�>�oIL�/h� m��Ѷ�Գ�m�n�H�AT�UuJ�O>�)eU]5��4ky�,�� )W/�j5c *��xU��JCڪ����J�;��-��N�I������vc�$[8E���m�Ȇ���q�I� S(4�]uuP�z�m���ذ�C�8�J� ե� ,���A �m6v�x � Hn@�ݳvΛ��imԑ�ж����NF�*�j��ٶU��HM[5
Ղ�٭�5��x�n���D�*�u�U@v.�gn`�ԶU���R��[@��9�Ӛ�m-��Ǡ��*�z�evl�5Ulr8�v�V�U�zt*�u ��j�a]��WS۲���Z���[\�V�v�I�H}�|��GK�n�H  �rcSUյu���y��N�� �i���Z����j����Q�M�j 	T	V�Su4UT�J�`�$N�m�6�Ӥ�6Zm%�-��� I�ه-�3;�� ��L�K��pp��H �~���U�-��N�)��8�ڻm-����� ��W�]�m�[m�Um'�0�Bҫv`����Z��ݰN�`�-��)*�*��ؙ@:��ZGg�j�Y.�\mRl �vB�cZ�MT$[v����m�   	�Hۤ݋E6$ ݻku����u\/Oo\����r���ٲ]��=� ӟA�o�n�Rq���s�M�;��g�oXoZ?�@D_�*���S���~�q�H�h�&��HpK�D<DRHE�@�A���Ȇq�����YN��#�A ��OO�趇��>�|���@ ��AF8��� C�<D�E%YP�A�����OF=TG�	�T>3`�(��&��Mx
q��8��*mW������Q@ү��' ��y�x�x�£�<P4�? HiUU����@6z*�P!@:���t�( @�D$�
�(( '��@�W�]��C��c
iw��� ' � ͫ�W����DOSb�P�U��
�D^�^*|
�>ǉ�C���О|��|��*L�@�)�v�i��@D� �_OD=Z�
�&f)���D���@�AD���,I�P�"h�� z*:@S=N��E@` C!q��O�T��>�p��331��� �~Sa��k`���}%�.�z.�Q����C�nڇ�uS@�eATWb?��	��HE�0��r�U[!H.ی����)��]�sه�/�	�s�	P��Y��Ѐ��5S�a|m�P��`�2�;��S�챹���<l`�{g��!�ۻ�����Ycl̨'v�ƌA�SM�M��p�\�.v6��牰���r�KZ;A�7f�c�k��v6�7v�W��])������+,[�#u�ex���N��m=�8ek<�ѓ<��k ���ή	��l��wVZ�fǝϗ"���-�F����ආy�ܻ.ͪ���(�AS��p�xgs�nI�j�k�-�;BFV9ЫU[R���Lv�;�
5q�q45UH��ͻh��.���l��d�S�zPйC�	��������v���lV��W-�٪w�.�*��dƮ8��p<͹�db)I�.�%�,W�q&��Һ��`��b���w`L��WL��[��7;���FQ�\lY��W�Y�ogt�R`�l����sԬ�s<330=�)�v��v:Z	]n���]'�݄�R�\��k���ΝnW94���E;=k��غWU��g:6�ʵvƷl\���W��Mݚ+\���\]k���v7h�Ɗ�=i�7[<�)y�Iщbݺ�<�/<��v����%��ZE�s����K��@Vő�Xϡ[n�؀|c  :8���]e��r�n�l�=Z�g�rZ���W1AqsTg8�5Ɣ�k^v�pB��O;��ή{��pU�:^�ݥ��^��5�m�;r/F�'�x]k�Mp�Mv�}c۰�ۧx;8N��8J�[�@�l^j�Ʀ�x�r�S@����hZ�糊 X���h��4:�d�N� ��t���8/l����]U��]��EW�v�y\ܸp���ѭ���, N(�1��aVЭ���X�#�K.���<�Z$ˉ���+��{-ڙs�.C��{7"��s�\a�mrk�	����8&����Oa�;��j5�6Z�3y�5��iE=Q>a�?�� ���� ~WA��|'�|*���B$X�*� �5>BF܌�*BJ ��s�Cj��������ua�܀T�Ɏ72�m��t��m�U�z����Ys��]"�9U���ˬ��d�yF2�kv�]�E�zy�iq�n2mӶ�8��d\�1hU�ۭ��ej��P����%�75׶}���Ϧţ>�D�;	��.cU��S�M���!��[� e�G�����o-�f�QN|���)���_� p��<�TP�d�s�W����<s�)�>2��	��M�O�9 ^�0�� ����uB�|����d�t����FdI0Vמ�j�� �����l�
]dI��8&���-��V׀nـj��嫗�����$���V׀|�k����uۏ ��֣�l�n>!��ݯ 6�0��x�k�=����#�Ț�6�L�'J]��3�{p�����=٣)k�f����-�����i��I�{��>[���� �n׀]z���܈����f���y�}�s�S	�h�4B�@�8
`��">hz
b?���x[k���v�;ț|RA)rG�j���^ m�`-�������rRGx�v�������0�|��ڰ�����p��~� �ݯ �n׀}�Հ|�k�N�+�s~F���`��q$A�C�]��rz.-��-Dn��x�w7F��ӳc�4<�G�?��� �]� �n׀un׀|��|u�69$h�ǀ}�Հ|�k�:�k�>[�������J����+s�Ws�6=^���D{}�(���ɰ;e�`c��9V�aIO��'�j�� �n׀}�Հnـo]UH�nDG#m�#�>[���ڰ�u`j�s`�N%*�T��j���al�']��6[��ڬ�6
c�K���`+nl��^*�����>��� �v�U��-���ͣ����Iq�۶g�?$U�y�V���� �x�k��9$$I0V׀nـj�� �v� �*ȓ��8(���۶`�� �nו���LA���jA<T�� �(P�a7�o���]G�k�M�9$j&��>�j�>[��[��۶`-��F��crp;nY��{6w7hznwf����>�v&�M$���Lld�>.E�|�k�:�k��l�>�j�>���?�&�$�>)SS�ro��u`gKj�����$o]UH�ډG#m�#�>[��k�`-������x�"bc��Hܑ�>�U@.d�VI���d�.��~[��S�q
4����<�]�t :�5�I���d��s�{ʮP4h
 C�<2>d[aTH�j4�=�K���x���ңKj�m�����R���㈍��ɸ�]�۵ʞ)�������-q�����j��:k	�݄2�2d����{��v�<O.v:����'n6�v�X�t���.��F���:B�6�#�%��봊��<�2gգ.l;q�͇ۚ��/op�;%ˮz+r���s:�����qr��݆�VoZ��5��sy��v���Z�*�ʻ���j8���p](�L�qx��iu�$HU����j�n��ؑ��$�<��<�^��^ }�f nԫ"S��(�d��-����:�����`[����pT/�9$h�ǀ|�׀nـun׀|�k�-��M���$|\jG�nـj�s`b�s`b����7?�eZ�T��>6����<�^��^ }��O�C4n�%F��*4�dV��\�:��4���W.|G��T����ѹ(�p�(�m�$�o���^ }�g��V���q?1�IRD� �m��@>��Q:�� <#��z"b#h*v��ռ�������G\IN6��"�RG�nـun׀|�k�>[k�;�5U��Qp��E)Ua������`jo�1ss`���9�Qy#r�8(���-��s�:����}>U�xy�;��i�9��o4�9eEt����pV-�0�]�]b���,�!�pL'rH�� �m� >ݳ �ݯ �n׀[�ͼ����$� Ԏ�'��%�
G�3]�x�5�-��R�O�1���>&�����U�}�u��f#Uʞ8 ���T��M��ý�-5U"�`�$m�$x�v�嶼�^ջ^���o��H��7$x�mx��V�x�v� ݮ�p"mz��wa[�2�zy��G�	��b�Uf+����s��(�mG E �� >ݳ �ݯ �n׀|�׀w�V�r6@|�T��<]�;�
A#ř��<Y��}�f{��m�{�7 H���I���`gKj�3�Ձ��̀�E	8W�Fܒ4F���9��=��� �������߀��.��)��y^{��bM4��>.E�nـ}��o��K�X�ڰ3���vpJP�:a.����c|��{2:5b��\�L[�Z��7?���_��yF��o�￞�{V��V }v�z�I��2�m��{��W��RG��U�O6�`[����0w�P��$�H��mX>u`j�s`v�5`d2yЛC�0�B9 }v��v�z���v��b�����$$I0]�l�=���s���1�z=��7{����7�1of�6��,K��v-�{�&���۠1���cd8:㋧�tx��l��2؎C�6vݏ	u	V�)�'�9B�8.�=�9.�'N�7]oF�I[����qmۭɦ��q�v�z�����wb���|���{Z�<���˚.���Q����AzoRK�n�4��mt�7�W\Wgu:�Wns��8q��C��fđ��h"V
�t
�`P�|�w{����f�K;�F�]��J�s[%�,S�io;s�	������p���	l�8(���;��`k�`�l�:�k�/X���1�ܒ4�q`k�`�l�:�k�5wk�-��&�i�H��9 }v��v�z���v���������O��'�j��;g��3��a����Vl��R6�1�m��{��VI�Us&���y��un׀v�]�����G�����6c���t�%Qdw��]�ա��k��f~J8��I��V }v��v����9ך������E�1Hc�Y:�76X X�X � qL�d��`k�`tb҂�@|�pRKWs��y�:[V��Xo0��9�ERH��ڰ�ڰ�`[���H��mF��4E$��ڰ:t��5w9�1ks`}����߿�H!Ò�6g�L�g���U�YƶK̎�嵊�������޽����L(&�`s��]�lZ���ڲO3�G�6���ӓ�OVf��H�wu�'��U���{�/�H�Y�6�`�dm�$vI���O�y��ô>�� ��"0x�3A��0���I �h�5�FP�%�iF�A�h�:�&�A�g����v#p�i��a�M�
k�@�����~1�e� � K
���Iv���KE�6�0m1��C��xy{�v}��{����<r6�����05���y��I����Xa��a.��V�Zӆ`9�h��bH�f��و��h���xq���|[�����͑�oq�:0Č[#�17x�d�Ϫ���)�٢O3)#j(@k�= W`���~@\P_EUC0`+��~@v ����~��;�x�����j�$qIn<~�s&�I�se�x��vO�T)�g���羆8�q�LR�VI<�rY'h]y��$�wu�'��d�W;�_��-*��t��m���� ���Hj�cj�CWG_߽�l�T�J��p�J?�����6-nl�m}�F ;��`�����pQI#�>]��q#���	'�͖I<�r_��儥��Ȝm�DR<|��� w�f����`[�<x���|M��G�X��U��w|�����+� t�,Dʡ.�
��*�Ù/�VI�x-���g8�i����o?�_/��~������"m8F����|8���/����.���� �+M�%,�h]ι�mZn���ܑ�V��}�Հ�ـun׀n�����	RFۏ �]� ;ݳ �ݯ �v׀}G��8�$��RȰ�8�o��j�� �v׀}�ՀwF*PR.�BN
I�un�`b���ΖՁ�ỳF��EMn8(���.��v�y|�}0{��?B���xӒܑ�P���#����\�lJ����s�z�\nma�g	���ef�g��'t�+V�l�6�P�x��f���sֶu��^r�]�7$�K�^-�P��y�Ű��	&����P�wj@%��on[]S��0�=��%��N9����v���Y5�rmsvñ�7VDNu �u���*����K�s��(v��\��NT�;B���߾�q�߽پ��ك�Lnƀ�)ڗ�ڷJ��9���k�$��u`mڳ��1�Fڒ6��z��, �v��v���^�\ڕ�m�I#₎, ��V��6-nl�mX�9�������q>6����<����v� �m���(&�FH�nH�������k�� n�� �ݯ ޺�����G����>�j�=���>U�xWmx�]����B|j9��M��G<���ru���]6u�R�@1��MN)Ԑ��B9 w���v���Ǣ��O1�$�3�i*(�bHdMU������z"���́�-� ��0�P�.G���pMǀuv׀}�Շ�?~l�����V�V��mIDR<�v� �m�V�xWmx�o-���H�F��q`�u`j�s`j���ΖՁ�G�9�����T��R��]�
�6%�լ�۶��E�LS��)l�9��g�|'uf^R���������3��`�Ձ�#��W�PI�FH�nH�V�� �]� ;�fջ^�u5%�)#m�d����O9�,�@v�|: ����9�~��7��[��퉗�Ě��Nǀ� �ݯ �� �m� �e|�L��䐐��:�k�NЮ�<Y��y��d���( 9��`��:�=[�;�"��g��踶�<�aw`릓p��������գ���A��V�� �m� ;�fջ^u�V�"�1�h�G�|�׀� �ݯ �� �o7�~i��F��q�{l�:�k�:�k�>[k�-������3�7��$�V��]���sa�����z*�Ձ�<Ԫ��H���ܑ�]��+k��ف=]�;$�P��m9L8Ȉ�HHڑ�g�iڷ]óC\�Z��Ă����8�Vk��N8�r6���y�{l�5n׀uv׀w��V86I	ȧ���u`r�s`�Ձ��7�	�Ҙ�.D�2@� ջ^ w��<�W�����*)�ؗq�47�n�V&���ua���N[�l������F5#mD�����qn�ω8�5�$��.���"� � "@E+J��Hd��� �e����)E-�w�lk���H�w]d1���z3��<�dř쩃!�7k��� �@�l��I�"@n��`��a�:t����k�ј{�'nmK5s�8�ų�U_�;�o��ӑ-�"^��Tp��&�[�<�F�����)�<�{F�r�K[�Z�P�������V�n0붝/59�{�]\�.!�e�5of��������{�����;�Ա����p�S�tp���T�ͅ�������6(fiQ]]aΪhq��}0[��{l�>V׀[�W��̃��1I>�|�������{l��F��
���ܑ���x�����`�k�7��N�q�����>V׀� ջ^���������8���S�q�{l�5n׀uv׀|���������t*�8`;l)I@�\)s\p۞ܺ캇;!
�vr��V~�~���ʽ$$�rO��o���^��W�@n�� �+H�����pMǀuv���g �C�D��SZPv�`nڀF@��X�<O<��� ;�fջ^y#ʇ�<�r1�h�G�v�y`{l����Z���5o��l/��D�$h��%��L�M��[�76q�O�Y5�t(���5[�uv׀|�׀�Ͷ���~�[���/;��2�uƷWVu֦�q�v᫭�9��ؖ����ݩ֦��ܑ�I�<��Ğ,�vI<�d�Ov��u�uI�NFۏ �]�=@��we�z�5�'������^����F8 ��VI=��O{�͆*�Q���U��W���d���$�,K0\'$��NI�un׀uv׀}�Հ� �֑]�$qĘ7��^��=���0�����:�/S՟0F%96�\��Ά�Ol�-\㧳��3lћg�iw�)SE?ͷ��y`{l�:���]��m�)j&I#@9 w���F��x����]� ��x��a'�q(���5w5�'������}��+$��zY'�̴I9$�#$m��x�8������O9�,�eUP�"����B^k��N��?�����O�y��>����߫@i��lZ���mT��7��
�"�C�{=����'W+�����塺1_��q��ǐ�H��N	���0[�lZ���A������
T�NI	 �� �ݯ=���F������'�̗� �ѭ#�B)#�$�N<V�� �]�~��$n�� ��<	��q��)H�F)��  }����Ng�,����}^��y3�vI���	N9��#@� ;�f�s�9]�z������d�%:�(pD E!&Y  �(��@���4)E�R�f*_�1%�Aa`XF66�fXX����`�����c��`I�acb���E@X��c`�`��� �d�BIe�i%��I�&B�%�RZ~E�HLK2�C,�����/6T�������_u�3z����%;tuv�h��J���fb�~R^ȥ����6�%�GXX�1���Ɂ���`�����f>>܃a���oN����$۶ �Y����𻋮D6]�wg�m��n��HF�,aY�Y��g������%�n�\�t`����8�]���c�ej�tm�[�:���v�'����m�����q�ptT������O/���[y][v8�J&��Y:��Mн3��(뎑]�g7�W�m���u���&�v:�ɱ��$�{1E�@��н h�	=mq�`�5 !�Z�HL4V���dku���|�z|<|��Oaf��T]qP;=�x���bvx�ɳ��6)n���i�yہ�[y.ѹ���$�0C:II��;$����W��^2��S�:	x
ZB�C���ҫe��k�8��ᮄ�1�2Nѵ�Ni��嚺� �$$�c���d 놷6�l�]�m���iv�Wh	n�7�6y�e]j�Kfs�u�ۆ�J�n�ڗ� t�j��Z�8 #��^�{t,jy�z�C@E�3��g`�Z=	��q�bs��k����s�Ѹ��V��#�Eix 6l�f�֦W�Zn״㬕R��b�3���^J���;q;mqln�^u�[�'"Q������9V#�0�Η�yhG��狩�h�VS�[q�g�N��ݖu��b��+���R�	b��1��$[�g͟Y�In��Ӣ�$k;1�&�t�s�b�۶��52�J��n��lV���
d�
�e٬�<۴��7<���t���)�n����?1���ٳÝ�P�'��������l��7//zG�c�):�oZ�iY������7<s���sx
V0s��NMu����c+�v���uu��|ƛ�ݲ��r1`���Va�8v��8r:ۓ�	�0���k��p�q$�O+����6�I'E�^I�M0�I�:5�mڴ�7nX��$�H��٩�/\ ���ttv��r�y�E]%�nu���@�]��1����i\h�fqWq�����hg=���:�0�̎�ñ��yvN3;�k�Sc�vx�.Ӷ��]��N�zv�Y�e�7;{���Fkykq�[���i����0x��� �L8�(�b��|S%uӛ�a��ܝ杙Nn����~��1�#k�ף2���ue��8G[�N';��[MR��a��ְh{	�C�v��s�θ:^��3�u�����Z���d�&v�N�e�u3��./4��w���έ��ɢ��s�(޵�^E��d�Ѻm�qӬ�^�+��I�B%��kl�i^���6m��k�1	��tg����횜����<a����=�������wy�}_���^�6��'v�6K�������1n�Y
�.iGkz���:�����O���>CJ7��$��^����^����*�ȓ���$��6ČI
	m��x���hP���$��vY'���z*�	f��nGNFێ�<[��y��gj��fk�OWw]�yǍ�Ȅ�!9��x���KwޘV��$��ڪ�w]�z��LIB`�A9&�v�߿~�����u_y�{l�>��^I�AHD�'R� ۭ��g�W^�㫂n^�D��0��n�Y�	q.6���ـ|�׀����|�*l=�! ����� �>�u͂B�aW��y����߿K$�wu�$���*��>�����#��#@� ��<V�x{�H���Ż��9��p�q(�A���k��I�we�~Y���C��g�쓙�둲(�)�i�& w�������wޘ��0��m���	�"qi�mn��I�l�֘���cr�h�5h`�Ń��������6��^�x��0yܞ�@ <8�9���N��o�FR-�9��x��3��� 7}�|��~�*����y/xĊ��$2B���'7},�y��g�U��UC@ :���� �ԕV\R5 �ܘ���^y���OV���'�̖OF��5�
�䌐RFӍ�0��?z�u����w�X	�JR"D��0p��=j6㧬�!�v'�*��چ��"Y�O�wv�}�4�f�����By��d���%�O9ܛB�D�f�N��иB�Tl&T��I�f��'�͖I���d��3%�
#��Yr7	i�& n�L�^���8�����o���pt ܎(���&������d����$��ܖO�*�� �UQ!�����9�￵ʻ���w7�Cs��NG�[f�|��|�����ʞ!����pj.C� 6�r�������ʼM\�Ie���s�����_!rrrNI"RG����7^Հ|�׀|�� �ԕN��H.6�Oz��� G�7]�x�u�'���d����HH)#i�$X�mx������׵`m�H9$Q��#\jG�|�� �ݯ �{V����쓛�Y��2�5#���3]�{��7O�j����ۛ���*�Wk�usv����@��cp-l���9۶��RZ�7M[�=�-V��i0��df�������n����e�3ҹ�%\�Vœ�I�����%8��<�s�ݸNy��T�{��8��r�6��A����ˮ�RݞoH赮5��}��� ׅ7�;<�K�9œ��s�u��s�<׆��I����F�;~�绻�x��?��NS�z����z�����G�㘺E玝4tG��X�B�Y�;�������!m���W��X�������9���Uo�w�p���QD�H����q#����*�� �{V�+98��|�Ĝ� �[^��́�<Ձ��6B乔�EEETI"Qǀjݯ ޽� �[^�^QR��4HԂ�n<z��nlO�����kIQ*�v0�AЩmKň�+v%��p$�k�R�y��6ڂ�`H�HF)�$m6� �[^�^�v�z���9$Q8$�vI�gq��T��(�����9ט�����{@P $swK_����F��ӏ�<���o^Հ|�� �]� ��`�S����qǁ�C�[/���y��l��?*���-�\=8A9�8�,�mx��0[��׵`�|��q�1�C�Rfs+^ş�Vpy��p��B�r�nl��Yg*��Gs��8����l�5n׀o^Հ|�� ������''$�r%�����ڰ����l�/+U����F�I����ڰ�������tz���k{V-�6��&B�RF�nH�����l�5nׁ����v_,����'M9�#\qǀV�������j��ۛj9��s�.�t7P�bR1�\+��c;m�ca�t��t��M��Ó���k|�/�m�����y�nl:�5à��q�Gm���^� �������?q"�E�ӄ�Hӎ9#�5}��`b|���������Ů	���$�x��0[�����r�� 4���D0@��7�r���h�i��r9�LV�x��vI�fc�I�;��:( 3�w�`Q��@�Z,Ym�y^��/6a73h��t�7ssv��&7)pֳ�%e�����������6��X���g8��B�U#|M�#�>V׀]� ջ^���{UU�����I&�F��;$��{�`�k��U�� �����x���Br	�br|����x[|�����l�;]I;��q�Gm����N�q����y���=]�;$�
U\�HN�lC$���0�j	Kd+�6%^;���Z^�m�O;�=m3&�̫���:�:8ոvR��@C�P��t�뎓m07�l���\6#C�Nn�N+ek�:6/��2i�['{m�M�b!٬�j6�Ȟ�fnTaB�s�������2�n1^f.̆�u�<	�n�8��Q�3Ɲx���������\rl�h6ԉQaH̐&�9�T��WD�8u�'��4.�4ۙ�6��0^��֎���Z�:���|��.�)��ݷ������}v�V�~�[|��^��S�8�Ĝ��'��K�IY��
��:�|��{� ����ț�d�|�D�� ��q�'���g� K�w]�O76Y$�8���4H����=�~����u{��~��d����@
{7|�Fj�~fB�RF�nI�~Y�쓴 �7v|Iř��=]�;$�P8pl1�n����\ӇIknoi��L�	������k%-.A�r
�Rs3��O����'���d����UP"x�u�'74~���26jG�'f�U}�XP68���P��_�T>��sx�ՙ��?,�w�U$z�gAMIn6ێ;$���d��f;?���
��W��d�[�vI�B��IN'qɪ��16���ۛ�s��=��<�W�Ȥ#�|�Ĝ� �[^��������7���s`j|�h�p]���
���R�-7&�n��!Dr�tr�%�$�����ϟi�6�9���H�$���d����~Y�~@z����'���I�>�S�4dJD�n;$�w9�1>s`bḿ�y�����脂6��y�����nI���|����.C�20�J���! �1�B��D��p�/��A�%1���a�ADELL2I%1EAQ0�0L�+e��$�wJ�D���	$��Y�XChL�(�pTغB7�6$���F @蘂�Bj!�]p�B�9�P�6�$Q-(��!��*�6�:���"p�c�DIQ��4Z��b"a�)(�	ih(X�I v�j�5��3���r~OA8�>��A �!�0I�`&��'TE_AA��>�M�����*�z�����':������w�vI��k�Nf�"Q��rH�rGd�
�w]�qw5�'�}ŀ|�׀m���r�R7�Ƥ����>��( 3&j��Ź��������o��}��v=]��W�]��e=c+�K-g�'a-`Kt�Q������{����ͧ�A����O�f�|I���d��fM��UP�8�՛�d���R~$��j'$�E�|�׀[f��^����
�T��Z[�)
��`���vI<��d��w�UUU
����+$�{|���e�o��H"I0=�s�{|�]��>Wk�I}m�Au��H�$JD��x�ڰ~�ο_?�;�za'���d�
�f�М�jD�&'V�pV��Zūh�q��X�똇^̭�ͳ��.S��8���&ܑt_��x��`������{�9��@�rH���+k�5n׀n�� �m�<�}t~�ꉋ-H�A�Ĝ[�vI�_qY�����ޘʚ�a�|i��jGd��C�v���=[�;$��2Y'��ǀ}���@7Q9$�,嶼�o�}X.M��<Հ���B�yG����6�X��f!q����Us�#v�7<d��!�<�	+@���Zs"u��^��n�X�ˊ�u��z�;�@� E<G���g8�#gY��	�m�����烧v�q��.�;����9ݜTY��6�D�S�p��`����.Ѷ�Ή���m�;l���m�ɶ{e�c3p��т��#l&�i�5��a��ng7c.�-�{��{�����%�#�u��q�$<pLQ�����^��m�3VA�)�4���qv���0HɎ?�'w=0��x�ڰ����TUD�#$h�AI�j�מ��k�XW�� }m���A�Ɵ��h�)q���|�ׇ��#���V�< ����mI#�m�� ��0[��{����`��O��6ܒ5�x��`��Wo��j��|�����>���Mp���6��K�?���|7�L�y��Y�*���UNƸ�i��}����ۓ*I�N��;$�s������P"O;����"LRN$�m���:���s@���0,
� � s��< �_�un׀oy`7P��9r<嶼 ���=�s�Z���5w5�'�c��I����#%��T o��z�5�$�θNP��1�'��/(��d���L�v� �v�嶼 �����]�/p�E	P��ʩMy&�7Ks����s��V^��4P��܏�UP��a�a�ё)-��I9��`b���3[���bM�6�"pM�$|N7$�>[k��l�:���y�佪�B�;�D�	�&ӒF�R;$�wvY'���f
A�F���&`iQN�
(���(
@((_se�z�5�';ܳ���O�5#|LRO��o� w�f��]��*�\��N-KF��r0�����'��K$�PC�7_ē���$�w���|~����8�ҐL�dn4�ΰD���������m:�-4Lh��u��:��@n&�r&��v� ����v�ޠ ��I��K$�1�H�a����n;$���/@$z�5�$����>D�_y���G����$�V�vI���Ϗ�
�Iuo�����d�D�XP���Sq�;@P�;�,�ş�k�y���r�T�d%"��u���@sz��d��RH��nI�|�� ��G�����o��u`d9l�R���j4�k'gz2�M�����=�T�5s���ym�{���'���%QZ���5s�l]�l7�~����M��͸�H�CR6i��'�3]��($O;�,�ś��?.w��PT:���|m��8�n8�o����^��׀un׀n��t��I�"nI��*��7]�x������}ꪪ�s},���������##%����q�'�UP����$��?.�;$� 
� 9���hE���]�z�u��V�2�=J��ٜuk�էZM��[N��8x����9,�Y�X�k�)g����+j��w.���릅[���,Z�&vv�<b٬�;j9uպʝ[��^v�ЧYwl=��#z�\�:-M����M83Ɖ��gӮA��̛]x�[׉ԧkS�ax̛��7�4r��8�Z�f��j�-�9⼛p��� ����{��,1�㇬�u���g.��윋���;p�$�tV��蓍�����wwvM��U����QǠy< ��f��^��׀TZW�P$JF�Mɀs�/�UW�P���{��=Y�;$���/G��x6�O��7�O�|�O����ż��;�Հf��P�j��M�#h8�t
�w]�Nfl�I�;���
��B�g��d�k�����I3
%UN 6�� ��V'�lZ���}��5�nn.u���hw�'O����=��sv��N������-�~��z����̩t�̩�����V'�lZ���z1v�`y��Hl��q�����4 �)"��uM�o��|����:����$n�����H�)&�7�����X����9�1����%#ℂ$�߹Į�LV�<�v�s���� �V/q��H�I�0��x��x�m���|�~w{���b�n=����;r�fp�h6�摪�k�2�y��Ͷ���%�V�RH���G�^�x�m���0��x���cmI\rG�w2^�$Nw6Y'����?,�;�	ǚ=nݦT��ʒ|I;��d�.w��M4R��*D&c�
F��6ݒO;�,��3��	n6ӎK'�.��$�nk�I������L�=����6܏ �]s`~�-ﾬ�M��ỳ�a�JUIN^g��H5r�q�yq�9�V0�h,Z��,���N��}ӝ�=/aa�f��O��}V��6��6-nl�t4�H%#℉I&�ݯ?�$j��uo����0
�u���Ĥm���;��?,�;;�l�=�d�Y�vI#�XU#n4���5�ߗ_�� w}�}���r��Z��y�z���UW�N�O;� ���ԑ���$���d�P� x�7τ�Y�vI�fc�m�;��}5�u��z����j��9�ͺ7��q�\]zz]k������w��s|�a0�UU�4��`j�s`bm������Lw���E�"�n6ێ<��^z�����d����$�w���URG:6�D�qE��#�O�$���,���䪷� շ� �_
��䈑�q�>  �;�,��3]�x��vO� �����ǡ�FD���E$���6��6.nl5��7޼����� @�"���2�eELL�A$�AIL+,�A DLAE�3,�LL0A�DD�L��A2TC0LLEDT1w1)�
X �"a�$��Y$��$%�HH�T�Y$Ie�a�$! I @��&!����_��N x�z����a�fYaNI��q�s���<����ab��HL��QLa`A$�A1LE��L3�0I����0H�%0��JB�BHB�K$�$���D�	M�M�#"<�6No[��b�z03,��(��o���UQY�lA�K��0\�i�#=��YR��^�nv2:����Wl<C�	�zы<�,��Gzn�wj�.��K��y���9�6�n޺ù�2�v���#kKۓ`�5X�
��7m�j0�Lt��콜&;��q���F�[{\qv��a�lga��:��i�h�z���ɍN:+;lv���Ԩ��$��g���t�c&�3ӵ�+[_8����pu�W��θ)�Y�T�js��h��@3���nqE7`i��U�Nm)�XF�L��j���tsi^i]�kUT`9��<�����t�Vԫ ��o$�^���/]��� ��V��e���[���k��,޶�C;�kc�j]��ihrl��6��e�n7^���s�*��VВ�b��9'���`�P1=m����F�ۇl�'f��N4Ϥu�;s��]-�5��"�����פ�����\�X2jJ84n�,��ɺ�cv�L���;1t�-�zZ/�gj�'F��ۥ�2��ɯo9�j7� �&L����%�n��d�����z�0�X�q��gRۈv0�Hv�T
���v�S��#]������i%��q���ٶ��_dc
=�Y�8Z����n*����H���olUN�K�]�����O"��qt$pARl�;f۞���୷��`ݐdӈ,n�����ӓq�غ�7<�Q�o���v{d�Z�g�`�ݧ9I�;�&[]�f2��/p5��	�R���<�θN��ڝq��k��f�],�e�u�9�OvH�s������F���O���ƭ���L9wN�^3K��m��N���!1�����3r�����u-�I�&�@l�����'Oj�R�6[Ol׫���r�7 d\K��zP��M'@q���)�ݵ��L���/UGi�Q]�8�dk��u��5X�y'�s���vH��f�nz�[f�!�d��8���7�`y�BuDO��Eܪ�ǈ����]�������(;&p��%6a�(\N֢��@x���ŧ[�Z�+a�4:�kѧ�α�m�m��\v��bz^��+>C�I�q���
��� �汇z^e�u�N�lc<Woj�z���X�k�7v{[�<���ۋa��Ӻ���f�)�h��-����T�����m94Ҙ��OS�x��i��N��S,cS�f�v��]�]n�W���+�����$�vN���ؒ.H�����]ul&X+z,��r�n��u���{�Z>?Cl�����zI���O�;��'�fOx
��՛�d�3W����ҒFQ��'�l5��9o9��u�?G�������4�FH�8�{���OWv� �v��mx���3�GL�'�� (�w��'�͖I�fc�v��\��Ow�b!$P��m���u`bm̀f�V.�6�ƒ6Օ��Y����j��n�×�͊�؆�(�*/h�����w{�|��vUvdܓ�:��< �����{�`�	�(��0H�N;$���.��!���T��3]�N��I�̖C���Q��I��"��L�k��l�߹����0��L�U]B��dRF��x��m� >������ڼy8�✑���rL ��,��;�>$���d��w%�~�`oܨ��=���2�.-�׊��+��R��7n{f��t�.�S��v���9���?s2Y'���d��w'����{��>�3�ݲ�H�	�$���3]�  �=��u{�x�m�n��r8�ۍ���'��K$�ט��BR�*����ꂗ/~�wʼ�~�Wޝ�XE��D�n&����=��z`[��{�`��B�~��iŀ�Ձ��̀n�:[V�we\b��jەCR �����.�Z�9��)f�-���ä�sW!�ێ�J��6�ά�mXku`4rn�D�2)#bn< �v��Gk��<��O{��A#�f�u8�
	aD��I���d��3%���6sw��'3}0�A7A!4I\jG���wޘ�{�|��߻�W�8���m�I���$��H����; ]����6I�MDB�}{TPb������'�����̴��a2�� 9���7yՁ��� �n�������[��k��Y���Wu�E�6�e+�7����Dm�_]�׎-s���m\r|�}0�����0��`�XU\M�I��jI�|�מ�9���՞�ʠ9��d���$�'������8��mx��0��x��X�V��ENN)�`wl�:���k�`qu��r�?!D�2)#iǀuwk�?�g�� ��ӕ{�}�r�/� 'P$A�p����|.Ӛ�<�U��=r�b���b�һ�h�Ͷ�\C�0�*��6�qp[v擫j�5J�(�����#�&OD �1�,:��3ڭ���ۜ�-z9{RFNø܌���CvШӷg�d�.�5&�6=�N9�9"����Z�;�Z�0�rZG�6�2�[t7X]s��@ݶ-v����k=1��km�k#n��X-���=�ņ.���n�Qnꦤprb��L��e;rt��I�bݣ���4Ȝm�rI��;^Հvـun���[|��(/IĒO�F�%UM�f�W��	��l\��77���xPl�|���IZ��*I�'W��ɰ5o9���jmPku`orU$61��M7�����׀u_y�ݶ`[���X�M�I��jG�}�ڰ>��{� ���`j�s`>im٥�ME�L^(rX;N��=9�=���歑����'En���Gk��$��d�O{��<\�?�@q��~�OF�7��Q��	�
�K$�w�> 6Z�q�'����'�fKڪ�:�-zm��RD�ܘ��x��X�m���0
��r�8�D�>"'EPq��Ow]�O;ܖI��q�'0dK�F�jGd��3�%�@PY���'o��~]�vI��� �2�d(k�׸J�h���|爷RG,��	M�DY�k��!�
|�㒟��}���/�5o9�1ss��DDb]��`?���H$��N90��y��s�H���8�����㽡U@z�����'�B�)q�#�OV���?.f;9_�@z�i�� �%	%�: (
��w��?,�vI��N	a����VO� ).wvY'�3]�x���s����;A��E��N.�d�.��|*�����$�^�I�������ߟy���tg�iݑvsFI��7' ޽v���7b�Z�h6�k���D�P��TT�3S`j�s`=�Հf�_{��A�o�����'h��G�D��/^b�[A�{�e�ufk�O;��
�
 6w��/8
%$��c��'��K$ջ^�ݯ �v���/?��'#y$a� ���|�s���9ǘ��	*����ֻ�uʾ�l���X�9n8�{��O�
�^���	=_��x[���V��6��k�II*�:s���Z�l4���ii�cEL�v��!��JN7RL��`+��nע��';�,�ޱ��0Î"I�,O��w9��u`=t��舏z�Pl�I~o�Ƣ)����O�� ov���`+��GS�m(b��In;'EP�����;׺�����|[ٙ��:�52�Ě0I#
$�O˹��:*��T ��>qn��5��w|�� VP� k�����~ۏgY�c �m�vM�����#͒J[S��=q�y1�G*h{xz(�<{0��-��S�4/�c��U�M�e��u͇�n�C���h�2s����a��z�@��k{��ى��;v�sȾ��������#^��t�/oh�$�K�ZR�+����-���5hyn.F�bԛOi�u�E�P=�q,�%���bA����w����y�7�+�#�m��nQ6�
v�]��v��m��sM�\%����;�����#k�H���<�v� ��|��=�d��=��#w$az�5��T 	�͖I�=�d��w�  9�z)5N6ێ;$��}Vt��O�������qSJ%Ȕ����Y$}ט��T	����r�������?"C߻�c�Jhw���ԀȋN+��h|s���R��>��┥��ݏ%)L�m_��@z1�:ET�����P�E�� �OU۔�g��]�D�h��k�g�:������w�DS�')�+�T	�Y��)JP�����R���w��)J��Y���^ф��2Kqڔ���ݏ#��C��C�N�מ��(~���<��=���UA*�M#u�Ț0I+y��ǒ�������)JO.��$?�H�O����)JP�����R��X��H�$m�WT	����1���������(}���y)A� �*�Wv��u@��Mo�~��n���f���R��;��┥�}��%)O{�߳�R��^��JUP�T �:w��P�Q$R��|�o�h�ͷ���V�<��&�;A&԰�n�����Y��)�R6�R>�j�"�}�
�T	�{��8�)I��{���JS�����	��΅�Dq2�I��MIY��y���������~���)�}�����w�ǒ��~�~/��Ѭ��{�Y���(|����R��>��│���AǦ���2D$�8Je�(z�P��a S� z)����I�D�T$02�P�@c�N��9���O��%�����8D,��`�D0KC0Dc���vgo5��D�s33*�,�� �jF���t�`�R�$H �B@��iX�(>DF�q�@	6��'E =Q�N��B��PT�
|�i�{�wc�JSϵ���)<���vkzԍ) N"܂��v�  �(d��)J���ǒ���k��)JRy�df�T0.�xDAR�-�uE)I�����R���L~����┥'�����R��>��┥'n���ܶ��G]��������V��g�u��c��Fm�lp�)��TX���R���w��)JO=�v<��=����R5@�=�b��j��խ���Z7��XZ��R��{��y�!��g{�\R������<��<�]�q�ꠕP&��Ѳ(��$af��>�����)I�����R���w��)JO=�v<��>�۳]7Y�f���m�㺠MV�Q=�b��j�1���R�����c�J�@%��*�-���qJR����z�j����������<��<>�{�R�����c�JS����R�����%)O��߽�w��	3�8rA�iڹyn+������}D�S�6�5ɆY+�[s�wwf��u���[�F�[�T�)>���ǒ�������)=���JR�k��)JU�V,�'mIq�f�T8��� ��9)I��hy)Jzw_�g�)<����R��ֻ�t���v�{�����R�����%)O�����I�߿ly)J}���qJR�a�����$�#�U��O�Bӻ��8�)I�߿ly)J{�}�qA"���F�OsX�5@���7Sv���7��X���R��{��y)J{�}�qJR��߻��)����┥'�È)�1����o[-Zw��<��0���l*�u��n�װGe�kָ�]\���	�g�.V]����"�4X�VN�Y�S9��&wId(D}���=�)n2�u�4i�}`��'V�W'7Av�����>z�$[�̥�v�b�ػ1�un1[uǎu�v�g�������1�z�z��%H$������t�i-�m��Hp�ɵj�-ڞ�=��{�����b��caۣt�8DX�X|��������K�j�-45��vy�|�9Y$a�T	��|�T	����%)O�����%)=���%)���=6�p�#m�㺠MP&�;�%)O����)<����R�qw��h�� ���gѨ�r&�j6�b��j�F�y]P&�C�fA�/�A����┥'�����)ﺎ��m���������R�
d����ǒ�������)=���5@�����WT	����b�"q6ԛ3[�Z�ǒ�������(�P�@1����e)O�����)JRy�{����o{������#�g��n΋jZ����e�h�p�7tY����9��5�La$�&�ݼ���kz┥'��wC�JS��w��)JO=�v��*�������wT	���3[GdF#�0�N1VT�<>�{��B��Ǥ�
��D�e);���y)J{���qJR��߻��)ޝ��l֣2ѽ�Z����R�����c�JS����S� ��>���%)ON���┥'z}�Y�7f���{х�ly)J{�}�qJR��߻��)�����(h�
49��U��MP�Ȟ�i�����k[���)JO�~���>�����)JOw�ǒ��������"��'��	�	HA*9-���:���q���ԉ�-�Q�b����72�+v�y���<��<>�{�R���wc�JS������K��=���<���z�Ѱ�SH���WT	����ݏ%)Osﻮ)JP�����R��u�+�UT�P&�0�[$N$ْ�Z��<��>�����)C�wc���0ԧ�����)=���y)��/��"b��In;��h� �~���<��=;���)JRy�{���K���┥/����~6o-��vkz����)����qJR��>�����JS��k�R�>��v6j�5C��: L6c0�(��m�к��u�b�Rz�Ve��n�vJ�[�����p�*ְ�ѽ�Z�ַ�)JR{���JR�g�w\R���߻��)����qJR��>�6ky��o{ތ-�c�JS����~I�J���%)ON뿳�T	��3 �4<*�R5C7bzm��F�q�u@��H��6
�T	����R��`2O~��c�JS��k��(H��(J���(J��"��(J3�-��ݷ{��~��D�Jܐ�w��P�%	By�%	BP�$BP�%	Bfb����(J!(J��>?s����(J��J��(L���(J!(J��30J��(O~����(J��0J��(H��(J���(J��"��(J�w���P�%	BD%	BP�&f	BP�%	�%	@H���
��?�_�T�J��(J��-}���%	BP�'��P�%	BP�%	BP��%	BP�%	B			3a=	�1$�H�i���P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B{�����%	BP�f	BP�%	BP�%	Bf`�%	BP�% P�%	������(J��(J��(L���(J��(J���(J��/����J��(O3�(J��(J��30J��(J��(Jӻ��<�J��(J��(J3�(J��(J��30J����*�3�L��@� 
8Hn(��	�,h˺q{�7��f��!�Yi�J�6.��kyk[߂P�%	B{�%	BP�%	BP�%	��P�%	BP�%	BP�������(J��(J��(L���(J��(J���(J��/����J��(O3�(J��(J��30J��(J��(Jӻ��<�J�����J��(Jy�P�%	BP�%	BP��%	BP�'�����(J��0J��(J��(J3�(J�$P$P$P$P$P����&���1խo^x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�%����	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bzw}��x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'�~��	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B{�����J��(J��(J	%r~��?ek-kZњ�ֶ �N뿳��@�B���y '�J3�(J��(J��=�{�^x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�%����	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B~�~�~��z�5���kZ�y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP����8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�����(J��(J��(L���(J��(J���(J��/����J��(O3�(J��(J��30J��
��(J�����<�J��(J��(J3�(J��(J��30BEEEE�:ڶaQ�$a�(J��<���(J��(J���(J��(J��(L����<��(J��(J���(J��(J��(L���(J�����(J��0J��(J��(J3�(J��(J��=;���<��(J��(J���(J��(J��(L���(J����	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%H���3���H����@�E�cl�N�t����X-�����\�8���eힺ�������)���d���d�xώSm05�6�7REN���p�ܮu�-���])�^�rE���\��f:�]������%��3���m���Z�
���1�:���nk���轁7�ư��mM�T���V6�&t�닃�9���wB	�0������:�әM���j�x��n�=r�3�8}��5j8�V���wo�!�̨����;ݷx�(J!(J��30J��(H��(J���(J��/߻�g�(J��0J��(H��(J���(J��"��(Jӻ����(J��"��(J3�(J��J��(L���(J���ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�����(J��"��(J3�(J��J��(L���6�v������֙3Bܐ�w��m�(J��0J��(H��(J���(J��"��(Jӻ����(J��"��(J3�(J��J��(L���(J߿~��(J��<���(J!(J��30J��(H��(J��{����(J��"��(J3�(J��J��(L���(J�����(J��<���(J�J��(L���(J!(JH�H���41�$Ē"!��
�BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B{���8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP����<��(J!(J��30J��Ud�J!(J��5�%	BP�%�����(J��<���(J!(J��30J��(H��(J�������P�%	BD%	BP�&f	BP�%	�%	BP�� �@�@�@�C:�b�B\&8�����P�%	By�%	BP�$BP�%	Bfb�"�	BP�$BP�%	B}�߿��P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�%�����(J��<���(J!(J��30J��(H��(J����~�<��(J!(J��30J��(H��(J���(J��=�����(J��(J��"��(J3�(J��J��(O�ퟭ~3Y7o7�z-kz��(J��"��(J3�(J��J��(L�B��(J�����(J��<���(J!(J��30J��(H��(J����~�<��(J!(J��30J��(H��(J���(J��=�����(J��(J��"��(J3�(J��J��(O���מ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP�������-�m��Ll��l�5�͠�����{u���D=vK-��ߞ�n�co��7����%	BP��	BP�%	�%	BP��%	BP�$BP�%	B|~���y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�߿p��%	BP�f	BP�%	�%��g{�\R���s`�5@���2,�Ɓm#j���┥'���Gv���]��Mg���R�>���JR��{�Uj�43:q��F���"pU��J���w\R���߻���d��w��r�T	��͂��j�s�<6q��m�㺠MV������AVj�5C�~����)<����R��K���k�m�v�����}i��rBU�������w�┥�?�8����c�)�w��5@�]�r
�T	��ǅ�DVԉ���v�5E����.�W[=����\B�b�X�rtV���[����پ��O%'���JR���w\R���߻��)�w�┥'��{������zٚ�F���%)Osﻮ�rR������R���~�)JRy�{��U]8�B�Fb��q�P&�C�߻��)���������>
��CC#�K�(ZS��8�����s��JR�g���┥/�aK0bIMG#f�� "��m���)I�߿ly)Jw>��┥#���U��MP̧�)��2F�!Hx�)I��ǒ��������)JRv�������};��R����>�zDL�]E���jaϞ)86I�,���
�ݼ̬�SL��qv5�Z��璔�sﻮ)JR{{��y)Jwӻ���˒��}��ǒ���tޯ��K�6�m�㺠MP&�3�#ƀR��?o��)JO���c�JS�����{����v������n���.IJ{ܔ�?|~��R�����y!��d���k�R��_~���)ﺎ�:n�޶f��k[��)I��ǒ��sﻮ)JR{{��y)A�Bp�a�"�H&.��!�#-�H�,�%212M0�I$�I* �(]R��麠MP&��f����{3v�k{JR�Ͼ)I�����R���u�R�����c�JS����6z��ټ�ȁ�2M�ݎNU���:�0S�\��qڅ��+�/��5ΊŶ��qJR��߻��)������)<���~/%)O����┥/�	�LE�$a5�U��H���L��R�����ǒ�����\R��p��Y���H������aI7�-k{��)=���JR��{�qJR��߻��)������);߱7#@Ȕ���N
�T	�
�(u��┥'o��C�JSϵ��\R��
E��*�P&�nb3I�$-����z┥'׿wC�JSϵ��\R���wc�JS��{�)JR@p0ٽx�Q�M@��L��dH$�u�б��4bJ�1�����o�6p�lpq�0�`�F�`L��{Ѱ ޝ�ڒ�%�݁6��,t���1 w�Fc!�g8#/#B�66X�6XXa��@a�aaa��X��c`XI$�9�acb�&����$DY3f0VA��#3,� �0�0
�C= >$ z����z`���f�3L`A6�>���kq����v&cca��f��҆�X� {�Ǉ�����CkFj��Y�$��f��F���4$͆h�jı�Fa�-hBWd�`|n�����ָ*P�͓k`H��rg9�͛��:�sHi�&
L��&�,,,,�qb&�gk�d�;"��l�q��	�����q1ŜhE1İ����5���Y�h�a��Ao�@A}�M�l�:˻�lf
��g������ݿ��UWRӞj4puŷn�k�0񹽆s�F���۪��.�L���v��Cmf���bd�.�t��m�멗h�(���Wkm��M�nv��n��]�/G�:�w3�͏[�M�<pFU����<[v��ۊ�Hv�yn��qWb����p���6:��6�L�<�͗;��cj^��Ђ�]v4^]�{[x��TX�ޡ�6)ѳ��(9/d���M�7m�qc$ �
��x��rͪ�r�v�Y��gT�bW�[Pm�^�F����s+l/h��dƮ�� 3ZX9�"���� �4���p-E�T��]���-�����%	�����1�m׎��� x� #V��Xt*�UV��*�ѓ��p��xnZ��iT�7e+u��\:)獏k�+b� ��q0R�i �T�p�)yvBT����m���O�{;N.��.��N������뗶�Z��Ͷ�^癜��F:��c��#������-���F���`�Kˎ�[���mYF�a�qN�V�\��m������޽a�Cb�̑�c��+N��W�=�,��|����W�trq>zR|;��C�n����Z˲q[q�tˢW� 6)���HodM�l��U�a��x�v��mk�����Q����9�0)۟+�x��v�@h
�9"�YU\���[X3��u�;;�:�͗��O$�1�\s�
��>��)yU��j�yV�ouȹĶE�ܝ+�l�lXG�K�l�4�՛S��v�d�"$Jȹ:�6P��ڜ��s��L�qٶwm��ֳBr㳽]0�p��J�۵��\��&e{�Zcجlh���$un�K�g�&��1��T7Uö[��$�fܰ\��v+�=<�:7���ݑ���r�Oe�puu<�*��v �횔�M�u/X�JH�[l��/g�`������A�&`,�͡����!�眀s��'�Ksq��Ez�&v;v�Y�{�֜ݪ��C�M�DM|>��OP�������
��=��G=�{�q��ƹ��)u�f�-�-���3�p�9�oj�v�����c��ή͵�8�۶1SD6:�m')ҀI;"� ��'\�%<u�`��ulg�#�m�P���Wn	2;>�!�n��M��c�	�5���[����as���P��r�U��W1ȳ�<N�NƽN�n6v���t�Y0W=6�c=�v$�����FӒ�`.��^�wwv��YӮ�Ϯ{:��!�.ݶ��Z8}u-��9{S��j�\7���5�W�)O{�����ￏ��\R���wc�JS��{��Ȉb�R�����JR�������޶f��oz┥���JR�g{�qJR��߻��)���w�)����43�F�#�c�C)�*�P2��߿k�R��^��%)O���)JP�߻��)�wOMh�f���f�Z޸�)C��wc�JSϵ��\R���wc�J�A1{�߿k�F�C�n���bI�$aD����j��y��P&�<@���_�MPŻ��)J���JR�w�y�oq��Y�#�V��C
�U\���81��Y'5]��+s�ԗ�5�������,�Pצ���<��߻�C�JS��{�)JP����z��ƨT9�v;��hn��bm\���r
��j�-�v � 
4�%��ݏ%)O{���qJR���ݍ����"�����D&H[r6�qڔ�{��JR�}��z┥�̂��j�Vf;��hg3#q�Z;ٙ�Y�����%)O���)JP��{��)�w���? ��������j�zΔ��(H��F���P&�|����R���]�u�)J~��JR�g{�\R���_v���{�f��iv̘��U�������e��ܤ�k�g�w;w��w}���ƒ�3�d��)J~����qJR�߾�ǒ��������%(}���JR�����7�-���o3m�o|R���ﻱ�)�w�5�)J��v<��/���IUha��5�bIQ7 �5E)����)JR}{��y!��z�����")���9��R�>w��Vj�5C2�������\��P&��ha��f�Tn캠MP$W3�Y���CWv���T	���2��l��#����.�T>���y)Jy����R��^��^�m�w�����,�:�M��!�:H�Vw�ݳ5�2&����\�R�8od
޹x���Y��{┥���JR�}��z┥���JR���w�)JN��ᬉ��䄫��{ݷ�߇߿y��u)C��ǒ���{��JR��{݊�T	��'c(��Cru@�J=�v<��>������$C���Vj�5C��c��MP&�x�f@�E�l��*ַ��)�w���(}���y)Jy����P����U�C�o�JR��_i�[-�{��6V��qJR��~�ǒ���k�޸�)I��{��)�w���)<�;�/l18��g9š:��E�y�F,ce��:����\���27 =T���%)O>�{�qJR����C�JS��{�)JP��{��)Ӯ����,���z����qJR����C���!���߿k�R�?}��ǒ���w��uCEP	Uhn���dȕ��E��)J~����qJR��{ݏ$?�ɡ��v.�T	����*�P&�gz��uaFdm�㺠MP$W9�Y����uÊR�>{��y)A�Ue�~��T	��ѮF�jFJ����
�IJy�{�R����~���R��~��\R���߻����N������:����a/U�^��'�v��G�۪` ��xA&F!%�.3j�Lm=���S'WI&�ˇ��P6��Z8����y�Iv�c�<f�]�[:�n6am�G���]���#�"��"�۹�w]�dݙ_柜|�2<��\�S�6�Ǟz���A�XpZ�<;��7X��s=Z���=��3ʰ˝PY��H��ɢعKc^X8�I(�i"x���ݶ�73��bպZ e��۞�={����Z޶x�)C�߿ly)J_w���(}���y)Jy�{�R����8�	h8�R"�q��T	���.��)=��t<��<���)JR{��B���H�k�Z�"̎%-�qJR���ߴ<��>�{�┥'��{��JS��{�)JR}wY�Z�a�7�oF[�oC�JSϻ�p┥'��{��JS��{�)JR{{��yUj���	l�˒F���u@��J{�w�<��>���┥'������y\R������~?�j�[��x���lE*+�t��dae-v�3�V!�\PM�����u������S�k�R�����JR�w��qJR��s���)߾���vkFoV��k[���)JOo{�%^T5)�w��)JR}}�t<��>������o{��>���%�TD$�=���y\R�������R��;��R�����JR��h�Z:�kf�o[ַ���)=��t<��>���┥'������y\R���#�$1���"e8�Y����u�)JOo{�%)O���(Mf1Vj�5C��0�[l�C�ơ3���K��r��F�܄\֐��Δӱ�d� 1dq(	n;��hp�1��JSϻ�p┥'�������u@��M��m��8�18�rR����\8�)I��{��)�w���)=��t<��;�5��ѭfj����z��)JRy{��y)J_w���J��J��K�Ё��<�e����)�~�b�5@��p)���X�5#�)�߿s�R�����%)O��y\R�������R��~˺�;7��1��r�5@�<�1Vj�5C�̲x�)I��{��)���8�)K���o�n ���i븶U�n0yێ+��3�bknFj<ڐ��銊E�m%)O~�y\R�������R�����R������y)J}�ٚ:�kf�o[�����)<�;�D	����}����߾6��"��)=*��[)
Er!Vj�5C��wT	R��ﻡ�)���+�R��}��f�T>��N��#�B��T	���ﻱ�)�����)JO������?&%�:B� mmI��5@�#��)�H&$q�r�����w��)>��t<��<\�;��Es;�U��MP�u��6X=1�zɗ�^	Yv�tΈt��gt�]7n�u9K-��Pv�G�5I�7|��o%'׽�������(}���h�T	�ݱu@��M�:��b9��Fj��c�)�w���)J~��JR�w�8�)I��{���
5C;�͆��(̍�wT	���g�%)O��R�������R�]�;��h}�x���8[�ǽ�%)O��R�������R��>���'�!�����)�ƿY�?��of��Z��)JRy�w�<��=Ͼ)C��wc�JS�������{�ߟ>��<��;�'�ڇk�Pa��gG<��s�W��4�s�:3\vu�H��خ���ܩ�M6�V�]�vʥ�qh�h�U�u��Eۥ^7�Λ<����ۇ�ܗi��c���e�1�ˎ�z�V�k��yy���m�8�	�z^0G��m�V�d2t��յ��i8x�,�ջbp���r�Ε:�0g������K���<l�3;��'T��vL��z}�{Sqk��s���V�q�u��2�;��Ɔ��mfj���F
��خW'3qDM�)�w���)J~��JR�w�8�)I��{��)�릎��yn���͕�o\R����wc�JS�����)>��t<��>�_w8�(&�H��x	�aD܂��j��{�R�������C�Q?�J~���MP$V{}Y���#&�i;[���m�g�)>��t<��>�_w8�)C�~�ǒ���{�R��f`��K�,I�#��ǚ��)G�/������e)O����R��4:y��Y���N8�i[��6UwR����&)�a
ɮN3]�K3L[�Н\���H(��8��l�>�9�j� ջ^{e�)$�pn'�o|�ý�p}C`b��������'z�U�O3�/�T=��zI(8$�ܐ�'w]�qfc��URG}}0���`q�xؗs�E"r;'G�?z��d���K$����z������|���E�' v��܆����j�>�r%���'�n�;Q��&��KM��3�8v��76�DWl�Z�3{@Ap��RLI#	�$�y�������j�ݳ ��ȅ�I�� om��Հ�f����RGwF�j|	HX�6JI�'k��r������j|�ކ0$�I�O� �E����}`���H	�H&d�a�I ���F�PIQ,��L����(�F!�� �IWĒ$/4�\`�|��$�������F5Iac�fIF�F�`3��h�@9�<�7��ce�����޷(��6h�NF6���
ׂŀ����dD��,��36�
���^Tν�n��6̱x/����E�>E��@=D�~T��N�2!��:�	P[�<꽾>�9U����9�~��#�C�����#� 7�� �ې����s�����o��Q�"n�� �ې�� �ڰ�lͷ�����������@�����K����F4�e��.��`WI�uI(F:ܝ�l�e�05rC�'�7]�sb�I�{�| �O}�\6I�D��m �H�RGd��j�y ���~�����́����rH���ŀun׀}m�a��UIqf�N��W�	:1i+B)�$�&���?
�7w�d�,�vI�_qY,4*���X ��3]�~:v�*YrH��O˹��:�����.qn��'ᙖ,��K̂4��d�')�OTAyvߓ������Vƴ!;m���P�L��n�����9��7�Ƥ}�~�XV�x�܆��^�[��3��RF�,�����*�=��p�'�}�d���%� 9���Dj7pn7xｐ�>[k��
�9���=Y��ތ��Q"���Ԧ�O����d����$�w���v���mj�㈑Ĥ� ;����������,\���yǢ=��۸����˹�K��-Nz���v*���^�k�n�D3<�b[/n,�/L��1�^1�찤�$�]&@d�g�)M4�;�ծ���>����PK����p4�@Jh$�H8a+��&݂DWd�5(޸���Y�Y�ɔ���1vn���;��ͷ��O0�u�\�U��k��6��v�;F�-B�	��jq7g:���k���3$�c�[^�Üݶvλ9u��z�'��Z�
��z��ث��k��`lkw.nF ��}6�����Dr>&����m�`�f��^������Ŝ�9$k�� m�`]�����������3�O��,I	�$���@U�=�d�^���v�� m�`i�G����x�k�;�ۜ�������m���}L�U���J�h�H1mrlZ�6��6��:zVh�Ch�tg^9ke��� �;ns �mxWm~��|��{� ����8��!8��rC �s���@_E
��vI��c�O9���>��+ƒ㌜�H� ջ^z�1��(%���6I9���?*��I0LE`���K�$����6�0[��6��"@����5$� �m�`�f�v�U������kr�u�,v94D`��
��eoH�hx��v[;��{d�t��1=4�#��5[^�v�U����|�w��Y'sN���%!bH�E�ĜY���U
H���d���زOVf;$��ܲ㈃JH�i�d���vI��e�?Ui� 5F��*�P�@ާ�;$�su�':��"Q�����q�:P]��Y'����U������hP��jzf�,�mX���5w9�65�����������ԋ�VW��h)*T�+�p���m��Y�^��!Դ�e�;s�qr�%p�E���z`[���m�`k�`~���|D�E)&ջ^y#���I�=�d��fKڪ"Gst�#���$x�}����V�������� ��-�
I��I�G���R�M�d���$�w�,�gj
�pF٥[7���]����򄳄�>.E���x��0��0�ڰ�)r&�ۑ�q�\9�V?O����Ψ�+�3["gŬ==�4e(Фj�j�V�#�RF�N?�6�L����v����z�,�J7pn'�y�s��k�:�k���w�7c��O���U��]����q"�ޘｐ�>��W��Ƥ�	#�;$�w��{���<�e�d�
c��d�*��E0��`��Os2Y'@(w��C�'�$�w�쓢�W(@�ID�F�~;%IIds��z�^�:ۻ]�$n��<������6�=G7A�=c��ͭp��;n��y;*������Ӹ�ѡr�Y��mu&ܷ��x2'�(������b�W��`%��xrYy���!�͸��u�\��9��&�����h敺�Z���ɉ�ћ=��]��d�XF&���V�i�Csse���(�f-j����3��{�|���6�V<V�*2�vn71�|]tl�5�@뒻j�7]9���f��[��0�nN�s���d�
�d�_qfk�wl�/;�I7�$�p�C �]�=Ċ����� �m�f���5>%�$��pr/���< ��n܆��V�6"��i��m��� ��V��q`gKj�;[��_,�J6D�'�yv�0�ڰ{l��ـ]z+��� G���r�/=L�ifs��˪���[�K��J�7nl�������S�rs �]� 7�� ��V��q`d(�Lp�D��(��������2=��U7�`tw;����~���h��Q�
I�m�yv�0V׀�f sn�FH�	$|Q7&�]�� �l����Y���::6��qIU��=M�����9�V��q`}�D{g��g�l���n^5�+�5v�;�͔�V�W-e��B�C��3��/��|ڥ�	�Z����{�X��F �ڠ>�b�CI��m���V�}Ϸs��j��ـo]�圉FȜR$�vI��e�$�ט��P�D"�'��g�p��u`b�s`wC��R�)�T�%W��E���� �n�]�l?{�@
�s~I�C�%2�R�I om������_g0������!W�$��2mg�.���7e�#����Mǝ75���nfӱ�u^�ke���L�v��nC �m� .�\�g�HH���x{nC �]��'��K$�w��h@$w�e=%Ȥ*H�������fջ^�ې�.����pa$o���|���{�}�r�;��w+a���Ĝ�{�%P s'oU�{ӱ�&�I�q�S`j�s`cn�3��`4ۛ ��ߟs1玸�n���!�r��<m�\v��YN݉������f���%���3�m�t���s��؃�M��HףQ'"�q�����V{��Am��5[�w��0���tԜ!!� ջ^ջ^۷9�}�ՀU�[9�qG#�:�k�;�s��k�:�k�>\�gd�@�G�F��;�s��k�:�k�5^�\��X���KT:C,�S�D J�8���,8H��!#LDDDEA1A0�0S�4�!2�3#���Ye`�H&e��) �Y�d��#H	�0AF��!�FpD�3�OB���F$�$��[py����l�C#���!�q���'����f�I��.�0��4DDMAI0A�N��ְ��r8ˇ9���A��Y�H� �Hp5j;�>��u��i!EO�>�'w����f�
�Uθ�8J�ޯh��om0�ݸ��Zr��u�GWnM�.����	9xy��Lݫs���U*�7"�r[Z3�K�Y�Wx�d�{{-��t8m���ez����ֶ����:�筇���ß�\�N|��Da���e-F�;�=i����n��]���q�.�궴e�{._i���;!�n�`6t���cGKp��jŒ^[b�eD���s�2�;V��]�,8ݛ6��sqq:L�T!y1��V����K����e��.�G=M���Ȭg��4$�l�5U�T�L�`Ӭۮ��VUU��T���U#���9Q8FݷH.�ӻ8�F��}��z�Ks�z��c�㊵/l�;�-� ,����[j�( ^��l(MONݻp1f^-���vUr�I�VQ��a"H�T��m��}�k]'={4DqKg#NR5=۵]�^.5�`��W���/"��\�����A���qJ�ȴez��ɠ�Vz�'ř�U]��em۶�-\2&�M>�'\q�{:�f�9N���!�]����j0R�p\�Cb놵u2�$u�O螧��=u�����˾!�<����$<l�ûX��ݫH��u�N�؃�O��6`��-َr1� ���e���K�ݛ�d�x�"�OgkKf�Gu�Ҹ�ᛨ����R�Ma�fGp��vKlܠ���%.����t��ݺ!�
\q.��Ƙ#m�%�u�u�k����:y�5�4Kk0��kq��@���ٴ�����u��5<|���,m������6���9��H�IuX��n�ظ��=���Q�2(������m
��pn�j�U��q������-6U�k:�F��NB�*�]�X��y��۝�h�ͅ��ζ3�űi�ɴ��Ә�U�W�q˺
�2��早x�ga�r�����۲�h�n�D6;8�c�vlnCm�i��l�4�UN��q�y��$jᮝw��Y�f;͘彿�N�q+@���(��Q�<U�Tt��W ��%C@��=�&��T{��}ONmŹ�P1#�x�^7\���h7�][���5�����=�BYKTQ��;�ت.D���7���6��c6�l�ev��$�)�s�&8�G��g���{Mp�z��E�/2����^z��Z-)����ō�5�N��s���p\�f��<%�u�v`9�Q����<W\Wnrj������{v��(;H��[ׯ{����|��˻M����9!	qՋ�sk���X�:�mWo�K�����q�5#mp�s ��<���U�����y���h�7�9#�[�<U����U���9���;OD?A4�M��m8�
��<	�3,Y� �n�OWw]�y����%'M�� �m�`�� �� �mx�#v5rN58ܜ�5[^�s���W��w��0ݸ�Xwql�C�ۡ��n������gM%M����퐸���J�i~`խ́ɷ6�w&��G�D4a1�`��Os2Y �s_����w�,�����<\�vI?�oN79$��Dܘ{ns �mx��0m� �圳����r6��0=�Z�w}�X�:�7[��n?����cD��.E!���x��`���e0��\�!1(��$�+m����<�;&u9�T�v1���4ż��̚�'81�&�m��x��`���� �q��=�d��B��1E'"rId�s2��UP��7f�$�wu�$���#�IHE8��rs ��NU�{��S���
	�D?�
�\�D<<������s ��7�uDRS��l� _w]�qfk����I���d���WȈ�|� ջ^�߹�}��o�WŁ�[�;��*�g��m�F�vpcN������n`N��K�nbX�ݝ���,�}��@n��~@����X���9w9�éi5#�nF��Ns ��L����E[�<�|�ݹ��/�)08�$��r)��}�jݯ��_g0�����E����m������� �]�d��&&� .���  ��1�'��7ʈ���Ȝ�`�s���`�k�ݳ >�H�c�0L\�i*+�y�c\m��kA[�죙�	m��n�DiI���S����e0]���ـv��`tg7�m�HN&�OW3�UP�A"s3e�{��I�,�W4��q�r7#�ݲ�<�e�;@
K��M�z���p���V|rH��nL��9�}l���^ n��,j����\��`�2����p��l|�,=��w}����V�3���uױے�j�q���nM�68�=8�ʁ�ī��F���v����%�-�g@��k�z��n]�lh{c��Q���n�]���i��{۶`m���v����Uo�ɝ���`��N������' n�@��9�i�oOY�t���w.0��&L[e.
�k*t�Xݵ�����H�C@<O�x�x"�C����>ߝ-���H��#K�7���i0����>������ɰN��aj5�����nST�tV���������s�_;��X��0꒡A��ӏ ջ^۷9�}l������?$n���%'NF� �_g0���5v׀jݯ ݤiY���S����e0]���k�� ����Y'�dn��-��&FBn��6.�6�w7L�1l7���YA���f�cfReN����m��\�����X�چ��`S��ŵ�t�ajl]�l|�,n�`r����6p4�rH�1����X�ŁT�Dwޞ0/{� ջ^GyTU8�'����x�K�r�|�B�bI-{���Ijۜx�J�o�'08�$��r*�u$��}5i$�{��$�t��i$����$�^�68Aq��N9�$��9�I.�w
�Icv�Ē�5i$����K�����O+&�)hҘ�uf�q5�:;EĴA�w:��M�V�;.6���I.�w
�Icv�Ē�5�ɔ�~�����ʟ��8����.K���	-����I!ksV�K���bIwK�V�K��,�Po�H3��}�I%�dř���������P�D4i@�CA�V}B�� +rgm�´�[��7�I.-Ko"p���nI�$�����K����Icv�Ē�Ui$�!���i�H��츌K�r�|�Iv�1$�����$�]�� ��"�Îǌ[r� ^;fd���1㙌%We�-'�P��ћ�mqP�i�� >���|�B�`�Z�k��ݗ�$����y�8�$��r)��B�y�I^�|�[��1$���3������!���SUV$�Os�Ē�p�$�7l�I!v�1$�{pN�RF8����$���{��}���[���IkuV%�?x͑�M�Щ�rS�ߨ�<���;�$��&VH���j�E���홈HZ�դ����1$��� ����~����߲������H�����E._\��뗒���ӚXlc�%��S�p��H3��w�$-��ĒZ�k���h��Xݳ1$��G8��PTMJ��L�U�����1$���+I%��3 1����~�����y��T�B�bI7?\+K�f$�Z�U��]��>I#��\�"��&��$���^bI%��ZI%�γ_{�-��
�I}���Ѽ�MF�����sI-�u��]���X���8�G����==����e�q��nշB�[v�sѭ��fY�Sn���[[l9�W,�c
6�Ȉ�\]�q����Aca5�
g��9��8�u�e��qW�K@�u�=	U����mft���Z���B4��@���c4˓�|�.�l]��,��5s�m{v.�i�v�y����
�H�N���[��`z�h-�~�=_��f�mdL�\��$��U�C�����Ld6��\c���u��|>|xn��gvÓqkOAv�K]9�����b	�Dg�m����&޽� �m���|��}�]�Oѹ�1��NI0��X�mx˶� ���X�$B�58��r,�́�[� ��V��V촥��o�H1�#��^�� /��w�j�tUP�$�cZ�D���#2D�� �mxz��U��ݶ`����~�v8��M�e�X�1q'a��!F�g���:駍1�狛�.ɸ����^"7�umP��x�u�:�u���2a�9`��z�1�(U*�5T;B���~�*�9��O3]�yǵ`Z���>�!����8� ��� �mxWv�U����7ǜ$L$���r`�� ��׀}�ՀvـolT��''��ܑ�]��M������ۛ �p�J���*���bvnxl��v��Ӝ��˦J\\�i85#�r!H��jq9���˶�V�xWv��tN�1�5 E?&�vّ#V�x�����Ƒ�5���
p���A7 ov�+���뗾�������3$$��A$a�4�H���bK1�\�HX�%�������j��H`�`��h
"$���G�IB�#4��	-)$��,��= ��1|cҠ��'Č��BO�q� �e�u���zy�����ͮ�w���3�$���&BB�")�{��'�׺B}<CC(@� da�D��DU��J"�		�(B"6Z�74�AE$2 �z���}�rm�s�'���م�f��j5��P����C��U*#�W�U����CR>�'��D� ��qS����WFB��ۚ|�����t���z#I�#aDܖN�Au�5�'��M�������� ;O&�@��r&�R����Z��w:�5o9������n]jBi[!�u��ݨ�2�b�!��g���iN�K�p����v}�f�m
�Q�jﾛ ��V��?���F ߽<`��m��"a$m�ӏ 7v�V��X�����H����QQ(��nD� շ� ��L ��� ��0�l�nD)�jq9�d�d��3&��'36Y:A�*�W(J�P��BXg@��b2$� �U_����]�}�=*0�jBb�)�,5��9w9�5o9�1�e����k�Wg9�=���cd]bF�e��һf�:��srV��ٗk��7&�v���^����m�KSc�b|�GF��:����?s���� ��� ջ^ }�I:
�ț\�ǀ}l� }�f�v���^�����߅�����8� ��� �mxWv�U�����|$���r`�� ��׀mv� ����X(���+ b	���3{��;m��;��n��O��'0�@����&��Q�ge��̭ݭ"����y�b�8����$��D��@�Smu��c�����97]�bh��Lu�Փ�.h�蛃Om�<')A��<���S���Z�z[���Cm��N�j�ܮ|��:Y'\�PZ��v���X��xT��x�
��K�vy����1�e��I��`mA��d?pI-�\;�@r���p��q����F6���#��]�GC5y�7%�Hm
���v����?���j��l�5[^�퓊Hڊ8���`]� >� �mxz���t\|��\j@�q�"�>]���� �^Հmv��j���8NH�9�x�k�;׵`]� �v׀|���yO�$pDn<�{U�ܶ�Z��mՁ�ΥJ|�����k�=]Y&;��,��OWmSdVp�\�cxhS��ͷ߯ߧ�1ks`�V��V7��%VxT�������{�~��x��zt^��@�2n��Nc�VI�y��?��Б�#����M8� ���w�j�-v���^�ͪ'�M��Kvy��mX���۫�o���NF�Q�58܋�=��,��^9���<��+$�UU�����,ǡ�Yg`��i�oZ=�b��0��CtQ�]�>.>Hq.5'N&�_վ��m�z���j�/lMUȸN�1�
�l���ݞj�n[V-no� |�M�i���
&��;׵`��s���(8���A�P�� *Uqo��{��d��N�"�Br&���-v���^ [l�;׵`����߉��(���:�u�'�UU
[���Oz�U�sb�OÙ1�d8v���2k�]h� �;a�/6��Wd�h�b�ZE�ѕ&W��xFl���ݞj�n[V-nl]�F�#qE$�7$xz���e0�mx����,�RF�""�nE`ct��6.�6��V�\|��\jN��p�>]���k�;��r�& ��?�� `� �d|�d��c6�!��!M�d�]�l��\�����?{ѿ}F����WA����0�gq�$�Mv��fۘ�;;��F�,����M�3S�wK�X���1ks� 9���6�����6�G��^��	'��K$󏸯hI����&�FIS
%UN s���{�X��X���>ڈڭF�㍧�ӓ ;�f޽� �m� >� ��Tr5�G$�9$�;׵`-��ݶ`wl�P� 0�B��;�F�Z7n��l��tv�/�pm�Dgd����ӳ���+�͓�[����N��8��b;F�Z�m��%�LDb�U�T�q�@�n�����bt�l�n�����x'��{l�j��v ��z79�.����1����ZZ��q��ɡ�|Ag�����O4u���R�8s[�Ӷ�+�^�{�}�ﴝ��Υ���{h��n-�kR�3�N^�j��m��@pN y�{�ݽ�Q�Ӟ�H�uv�Y�����7f�[	�R�ت�k���&*�k�E�Gݷ����~`3[� ��V��V�����B�rp���x��� wv��{V��^{I�NE�p��S�x��0��\�����c��
Jby	Mɀw�j�>[k�>]��wl���&�i'"mp�, �l�>]���f�ݯ ���|�6&��὎z��m;����cƙf��g���:N�ao��w���7�
��������� ݶ`]��߹ϐ�z`�Dmy��q��	��z�����>A�Q�*%�� ���/�]��U{��0�mx[�)"Q8I$���x��6��������́��N��c��N'#��f }�f�mxWv�{g,�܁i��5��96��ݞj�9�V��w8��s�9]]��฀T��N��9ݞ^�^d���AVH\:g,ۯgd�z:�t��*�����X�ـvـ�:ȓ��$pMI#�;׵`�f }�f�����^'x��RF�o[�U}��|����|�o�DU��(U�PF)���y��9���K���RH��ԏ��0�����X�mx�^%(��q���r`[��]�������0��U�6Jស;r�sqvMV�7T�4�d��-�6n���Fh�D=pޱPTm5R�?ͷ���� �]� >� �ݯ ݰV4�'"$cr,�v��?s�uo��V���ڰ���TF��"��E�b��������]�MX�ڰ1�8^Y��$e�T��ڠ^f�$��?g*��w���` ����EP�
��ڷ���K���'��H��rI�n�5`gKj�ŭ̀os�vy������`0l^[Dǒ�n��ק���;dj/�^͓���*T�i��o�㘬���c�I�{�� >D��5Y'u�����1��Ⱦ$�wuߪ�$Os6`V��k�`Sh�q>8�i�4���ـ|�k�>�j�>[���jRD���$m�$��v��v��^ջ^�`��M�) ���#�OVf;$�  935�uBM�s�r��ATW��"���j��+� �+�"��������*���*�������

�(�0� �@"C� �(�,� ��*(H"���TW��ATW�Q_�"�� ���*�����
���*�����+�
�����
���U�U���d�Me  ��qf�A@��̟\��|\�       ��            ��	
QR��J�
HP��� ���HQB���	RH �P� �� 	
� ���PB)(�       R�_}(��A˻{e��n=Ζ��t�O].,���Ξ���vǼ>��s�m9win;��  !㞞n. �U�/M�s�.=�Vl�� s���yO&�ˑ�Y�+� 8 �   
� d ���O}���W.v��� 4w��e|�;��{:z�[�� ���f���/��r��nm{�>��}./��O&�v���{� ܧ��:rk��iz��/ z �   �
�� ����n�q9:����� 7	Y�������#��L��&�	�O��x��W���v��r�M<�5׷�{�� \�/  �   � y�gC���  QJ � }Jgt\��O��r�MJ�>��=ri����{���>����)Y� "  �` "  @ D ) ����� 0P� ـ�� � � � T@ T�@�@� � � �"  �`    	  @ Ru�>� �Y;��^N�m� �ϥ2��/&�c�����Ү�}��/���;�nyS��_g������*oi*��  "����o*�T�L��"��U*T�=@ɓF�"{RG�A���hb)�����R�  �M�)F� <S}D�_���m�}�C�m0���v�;ޏ{���TW�r�蠊��
�
��A����TW�QX(����}�������B��|ß���g��8_9I���<��<4�y�.�מxr�8K����O����O߈ޟ������Qf���M���\��4��|���p���� ���y��f�O����{1�`���'�� [�oa��������ϳA)�P�j����ö؜��؛k$�0�1}��}��s����/}���~���[�۰����M����$�|�'�?{�~0	ISC��`���I+��d�T�@�:� �(b��)l$⑹�	L�hjhV��L f"SA����
J�H霁c%$$R\�9�	W٥ׯ��!��~2{3ԉ ���O0��H�Hl�$������9�����I&HA���_O7/��"D�d�xF�C \ˮ	'	H�� II$�����'!w9�B���rFy�`B�!0��P���<��9���2�����r���\7�S���}�1Ӟq!p�,�l����$.o)��9���+�kɻ��s�$H�3�?~�����R����=�"�)fT.�����~$��IjJ'���I�YD�L�9��d�N>HJf��1}�Ɛ*0���=��OJ��B�@ A�
��?@���.Fe��i����������@�.F��={uO=7l{��$�O��&m%��{�q.��M����ki�9�LY	$S�D)�� �  �� !�$R�H�2 � ����0�A*����$Z�� �
1! "�L�)A	$	�bơ��&Hy
���6U�PH�B��1����M8`H �؅,u9�Ġ@������`i��'$�Be�928D�F��!c��H�d�HrC�$.X��:H�	%1&����Ym�28c��$.x�&� �c��9ZL�ĉq�I��B�o�H%�ɚ�-��d��,(R׏��d��$���(KV%�䐓p S @�I�"���2��O!k���BFBp4�&iō�d�#� ��T�T1H�N x�(�:�,��W�B͊����k9Z�<$d"4�</�?}�G���h@�8<A���R50"�0%�PԅLna.�	I��*��d@jhcP�!���JW�B!#rpb@"�5���c	(Ғ�A�d�)�C�A��P�_FՄ^Mp#\&k��04���d(������
2愸h�(��V	p��p��)H����,SG��"W9O�
��bP��B�`��q�"��J��\t!��Lt�bBQ�Q"Q����~��A�y�G��JxB翡����I�No����|���
�)0^y�^���0���_}�_��7�S9�ā
g0�]�)���J��`B��_#6�����(�����[��w�L���Ņ�-8�Аe1�H�#�1�>�i�bjj���zO8��ۻa!��ß��R6F3YL	F!b@�eIRW �P����ksx��w63�:g$ns@4�$��A��H�!$��"!�ࣷ{�#F�	dI��e� �r���Q5���b����1���
(���$�4�a�(�Ӑ��63��S9�"�`�
`i�Q��Ux�n]�=�c����FL?�CR<�y@ș���>BK��Ȅ�p�I.@�A=u1 �sbia�0�F_P���\�)	��0?z{&�13l6F�),l� A6��$q��v4��6Bi��<t󾛥������X�i�;+��	md�I�d޽���)o�9��6a23)푲bF��g9�8S�y������pi/6�kN��ԍ�}�ܧ����t�"��#6]��y�L�1�Ӛn��NS���R��������˙��$���9Y4w�����[�n����O�~�H$��oĒ�A�I�{�D7���x�HD��B��	 @�	I �
D� H�l��,H�� >@+
z�T�!�����"�QH�I@b�X�@��� �
�0
3$|@�0�BIZc��XA#�%�e�a	�2N@�;�S���Hf�ͩ# ir���RFprZ�t�BE���l�	#��%�!\$�pxJd��@��\f��������#����҄�hC� diBL1o#9(a,��l�B6ӓ���"�У	 FA#CdIXs���p�,�Zs
��GP����c��F	��!�<X�a5��ėω��<�	I\4�J���Cs#��P���g!!����)�N0�1ׇ��i��B<Hc`��NxK��p�"H$H�^��$0bBѤ��Ü<�IsN��
c�$�,Za�<�.oA�d��v0e�2\�I �k��40t�(���R�$�q2S1I���[ha��M	##i6�M��'8r��㮘H𴅰ic!	��v�-��K���43!����p$4� H�c��2o��x����a$	��%3�\�4"Ǟ%���p�.k�	�8H����$J#���<�`��5G�㰹#���ŀJf�'$��5�1a@%<7�J�*�!rD�C����H�HW<�2�7��!40�$�I�
��ޗ0a��CS���OB������`R RA��J�� I���L=��a����%�ja��7�o<֙�$$Ǉ�^o'��3y���.r��zzƙ�����������?Lז���Yl!�P���.p��cxO��	!13y<!0�s�.o<H���ȇ���B�B7P�8xp��I%0�O1��@�Č/7�����'²f�!L�nHj)��yOФhJi4�S�dy�<BD�o<?��<�H�+��W"o$'���"P�=�! �����7�w�?:�.V,~4��ԓ9��_�!��s�I\9r�����o𐡆��C�*"��¹��)$HSxx>�	c���i���$����I��S�����^��-���~�儑�C��`¤���ZBd6��(p瞄J��L�RK!���!+�� K�$��B��!P�?J��@ @b �b0`E�� ��`����{MF~����w���4� XR2�<9	l��~���xy��{��9�\��ܰ.�s<X$X�����)�<M\bVH���\5bL(ЏB51����,��`�HF����!��aM�ā\�|'&�a7$�O"D�%�Hl�4Y�VbP�b#P���YLBL�B$b��`������D��-��YId	!jR�bB�
�������"D�
���r!�Y�1B5��bhq��VRK��h:]�&��f�!VY	6�3Yr�*@�.i��p�I�jI�MȒ�SZ���bU�Ej&��#�0���8хHT����&����5׍$aHb�R�)ns�H]ap��k�ĸ�.iHD#T�V�o%m��p�1�Myo,Jd.;�D��
\�Ąt�&�R!h�\u�4�L#	&�����!p��	r�32"Iq$<�|�0�
����4<���9�����8�~L���C�l��'~}��~ӿG��      m�  ���V���aP�n�i�u���zW:�ԁ&�\�%�Ͷ��v[m�@���m�����#���\�Z��ԫ�.$\��Ilq�r ����F�l�ᵷdL�셠�&���U�Tu����Ʀ��<kF�=lR����pm��iMˇ4]S\�I��m [Am�)e����NX�m"��� �kl�]8f�r�ęsv��U^y�ԛ�CTc++mѡ��/�:z��U��H���� gE��'7(��..[i��\&�yz`�[����T]fN��l]�$�H�7��@�@T����pe�V�k���u�� �b*��;��g	:t7Z��Y�{�#� U�$%��3Pr��K��8��� H[y %��v�km�;m��$�ks��	V��*��
�Z�"�nm� l  @�U���imm&�I6��8���-�Ό �$�8�n�m� �I�Ā�hX��-U@vI8vu�mKkn�b�:M�v�ZM�H�:Kd�T��  8%�\��]�۶�h,��`�N�] I&ݛ��6�8 ��V3���nΒ�����l �L�Ԝ�`[:k%�#m� 6݁ղ�T�	�q���U��U�L l[+��84^���I6[m��ʭB� D�܆��T�Fm����m��i@e�V��L�� $ �t���?�zF�'m�l�v�Z�n�dh-��-ȵ9!��[:`   8�� ��-���`;mѮ8�u���o˷�	  $6Ϋ��ms���t�]�m��6�Xcm�  [%�k:@ �t댳-Of�� �:��v�
�5�  q)r��ŲQ���[M�7���m�Y�%��$�k'Kz��d:�x��!l�,ւ@l�m,���D�f��w�U~t9�L�f�` �e�]F�j��`��     }˵�Z����0 A�h���|�Ka�@]�t�]tC7k5$�4S�[m��Z�tU�[mԄ�j۔�Uvy�z�{BD�U:��[l�y�F��W �a��  ��q���l�t �6ۄQ��)�J��Z�(�+�S` (
�j�9,ˠ[m��9'i�Hl8p�U�X�R�u*ʴk�Em�� -�t���C������ջ[ך�f�     ����[@�� -�Ā"څ���bۭ�     BAm�`p��6�I!$�o<I��8�jC��h�m��l�  M�F�/Yim�  @ 8[M�I��dKd$4P� �3�  	��m�m�o^)Km(-�0� �a v� $�Xkh ��se��6p�ɹ8��4���U� ��]K"�����
�6���K��'X�k�b���� cR�UI�a��ljj��U�n]��𕃘�@��Z��` � ��  ��k=����Uf=�A5'���TsU$*��V -�[v�����X��a�T��L��m�m���d� �]�nm��&	5���m��֒[BA�͵�q�d�a���*�yf��ƋR�T�me�6  7m�ꀪ��c�AKT��@�e%�#T
i
VR�xe[h	�qJnJڥZI.��RV�֭�rJ[��@�*��-W[�n]�-����m�v�j� m�5[i kj���;f��荂�4uRk�t��a~�L��Ԯ�jyy�$ �U�
�;R���%�vj�Wմl��a�[KE� �[@5�     v��Ͱ^�e�m������Tm UG�P�C�=NZ-����5�u�Í��:[ɫRcuE��8kH�ǖ��sm��׭�[j�Ud���0�+�
lr� ]+f���`8����%�魢A� 	  l+m,� �kn�bn�jm��ًd�y��j�^�6��'d"۫l      ��k5l�V���`*J�UUTj`����e���W1��Σ�묢��i��W;g[pdi��W٦��tԬ�" ,��P ��� m�l l-�6�����޷m���Ku�  [V��Eqi��H M���l�]%T)c��R��4q������C�ld�e��Ȩ2�!A�*Ҷ��5b�[�mf��Y�6�Fڎ7b�2Zح���&Yr���D�j���+-� ���*5m�����   8  $ �m�H βJud�����zԄ�[V���p mt�E :�5jU]��-\�{۠l/< 	�!P*�$�W[��W�:����We��UP����~Mm��e�� 	 �K���o.���:�; ++��,��\� ��)�m�+6�IR�M�����R���� 6�٬�:�5�e͓Yȹg+)��e�kn�p㦃[Ml�q���jٛ������^uB�gv�Z���ݫW�u���2��e�"q�|�8Eis�SF���A���Ӡg�����iF�뮕j^;*`�+k����[\s��*�1Yا�2ᕧ29�	����<I5�@]� ���o��� 8�c�Ql�b�����<���V�]��UUT�l�sY�M��u֒l�F�R��iY�u�� �m�oU�:M�t��( �$��d�z�4�Ce��(moW��x��H�~��j[v�*4M�M�4icfCj��XI���K9Zk֢�Ω����ݶ ����� -�+m�mղtt�dmF��ń����l�ur�5/[b��i�^��k:K�n �4P�f��y���ڷL��@j���5ZC�mT���M�m�ս�m8h-�J�Аm��nuЛg ���l/el�j -�,�M��:ѱ�J�s��  �8 I�H֯A�8��"�B��6�f��h8Y-6�f	��� �J ��m�ְ ��6� �[wn�t�ի�ݶV� H� ֶ�M���� �X�iY��&�`9g*瑪���m& �ڶm�Hꈕ2�5WGR  �f��6lO�Hr5F�j��VRW��e��Wm[B�  6ؑj��R��U*Ԯ�#�[z�R �C�٦�HEr!0�j�h��S(� ���KC��@�r�K���[s[�7ֻ�vհ �  [@
Ѱ��>/C ���    7Z�  k�`�m��� a���lᠭ&m��!IP�J��Vݭ�l[Ă��m�[��4P���*Ԫ��!-�[�U�V;n1MTd%�gn:և   �oi<5�˦� ��   �6�"@$�`m��m� ���.[�Q*� 6mR�8 �moPcIv^f� *�=C@U@U*�U̩d�IeZ�R\���e�V�۩X���Ttf�J+�3�-)��<en�2��BG`m��kv����    m�   m[   [Cm� � f�   � ���l    ���H   �`�` H����m�   6�m� 8i�   [v @� [Amm���m�� m�m�,��M� ����$�d�[�i4�+q�EJ �	2�,T��J��vUj%'[@��E9�]Uf`�m6���m�   -�Ͷ  �`  �   	�s`@  v�@  ,�T��;����6�ְ��
��B�[T�*�R��Tkt0�� �v-�FE�\ۮ9�t����h ��Þ'l_>-�)j�fm�)Mn� U٪�@�\���2�(7m��m����V�  m�  � l[@�  [@�'@ �� �  ���`  p �B�F�ʹ��� I��I�m�V�p��ҽ��E��j��X2�%��]��s�s�l  ��� �n�� 6�   SP ! հ m �4쵷VʍJ�Q�aTv܁J�!J���U*�2���{YehYVUi�9xq�����j��M����l�m�<H� � m�-���l b�훶�Z��m��� 
F���1�5^��m���-�-� �i�m��N�>�2�D;+Q���V������\��[ �lu�����y��l;j�� ֤¨	]��ڎ�H��6vd%k"¨��=��ĉ@x�p���)�uK����o��XC&�o+MU��A[-���Г��,�.Ү�-H!WWU ���"ruH̺�a�Cj���!fmv���� E���/lGea�ͧk(Ԯ[\ku��R�%���6��ٶ� Բ��[Zޚ��C�T�{8E��+3wL�&I��m%��QQO�D������C��W�^��n(�D�ਡ�x�� ��� ?�OPS� (1<� �
�_��@1����T�W���x��@W��x�N��<@z<8���ptE�AG�*�P�t<@��@�	�!�p�MW�~P0����#�H
b@[���z�3S�T���@ �V��� � A�ň@!0�k΁����@ �≀E_ADc�? *�@*'���������!�`z������ <8��+���#V ����~��j �\N~���A��6$�K)-��
耾(/�D�����QQ�8��*����
��C�?�PEEx��!OE)�A�$@�O������UJ�C�=��9�Q�n�4�mt���:�F�����������H�`���{#��]�.����ISn�ZL�P�r���Q���9Uk��Is����+[��Ң[q�f]ی��=]#��.xLrF���;l�5���()pĜ��\��kd�r���Z�p�6�q,��ku&��I���l��֡�d1Zh8�.�S�v*���Am��q�]�Ɍm�;��l�t�Up^u��9� \�Wi�cY�'v�.��3+Uv��^u�RRWG��{�7R�۵�%V�Av	z�0mE�b�x6�d-խke'�]�mOkfr���Qm���{N���d݌F	��g[��G0Z��;v�t�UY5�#sC�Ѻ�5�܍��Ntz�UkX.4r��e��[zϝ#�\Nn|c�Z���;Fҩj�5UK�+Ҫ�M���z��2f*JX���=s��jјѻèaV6��2`1vY9���ˌ�F�H*ʬ�ت�H�\z:n	m:�m�KJ�nz�%�:d��J�Hb�]�Tt3:��sq���"���{oh.�$`;sG7S`2�  h�Ng���5iS��u�<�i��O����r2�5KC��n�`��I٘bj���4�/ s���@)*q���ؠ6��`����(
� �:�d6���yV��N����	���L�/E�Ӟ�
�(��"�үl��˵�㧇K��[7 ��2���"�HkXN�J�[ɶΣ���&���[��]&����  6ؓj�%m ���f'	�쐝�@*շG6[v� ��%��eV�ٶ �Vү���q�$����Y�m+�D���q���K$d$����L[$�	8n����̫ڥV�v%�f�R��8�L"�6�7l5HH;+/T,f�K�;U��P���+�K���fGO�g�)����X���&�#ųd�]7e6d�� �~��"�D1Π� �U5T�"�T�"�w��ܖM٥̥&�ݍ.�b��X�=y7��p5���Zs�Wl��x�9`՛�eGm�mb�ư[�ꤹ�jp%k��Z���1��k[3;=]l���|]㛧9�=s����d�ַn��y�#��{��'he�\�P�9�+��:���7&�pL��Ƚ/n̎@h�:�v������\НpA��ttIg�x�B��y����f��;�s��ca˻q���l����<C�cc1!���Y�K���}'0"���-J���X��2G&�Wu{�3���"���h.��޳@�˕��Ƥ���������� ���R]`}���1,y1�@��^�{�@����{l�.{�"X<pb�G��l������9��@��^��}O��v���z��n��F7d!:	��^8��Թ ����d�$f2]gn�s͕0<�[�
�.�Yy�}��Ƞ�A&n-��ng�%p�B�!fo�x��x���V�0W#Xؓ�$�*�^�{z���G�� ΢�0���D�A'�{z��>V��
���U�@-J�y|�O&H�rhu�@�{l�*�^�{m�/j��)0xF�Rۡ���$l#���+��V�t[���l /C�"0��I�����G[4
���=m��*`}�ܛx�ı,�jՕwx=[�X��x �]�&�4��,81I#�z٤�����M�EE��1IF�(J)(Jbodv� r۬��%\�$l`�	#�@/[4Q�����~K޻4Ԡ��G	0MH���� s�� }�� �u��!Dx��O����3c��8��k�/�=�o\�:�@d�R���([&-�޸��j�x"�$�����{�� ��h����E|aY�%#�zٿ��A��M�~�h{���\N�86�vw.��`_m���Ky�T�X��@��˒H�!0QŠz��hN���9$���w�h �x*!�:
g�vՠu���ǉ�ǌrM�e��o0/�x��%���e75r��nl(��;U1Hsv|<�fc\�Ζ�
��$��1flv���)��m���w�?���>�[��Q�:w���!d_!���$�M��Q���z� �����i#���$or`y�`U%��o0/�T���.(bT�ǋ#��I4>�_>�= ���@��M�wY��]��K�����}-���`y^`U#���@�"]l�j��.ɻE �V^�mU��S�n9�njT��p[:u8�A��Ɍ�V����f81�����z�V�q�da�PKS�ΰ�k��k��8ԽR�1�΃.�ƻ�3l���݌���p܅��K�V=�髲;�m�D�+ɻ[*�.���Aӭۙ��K�7w ����@�$�66�%��,T
@�[�1)��Cv��v�m�Jb��w�^��Dw?6Xښ��Q��5toB�A	�\�Y�nw����!�t�8X nl	�Q�=����=Gu�]���hq���1� M��=Gu�R]`Ky�}k��4�pd�nM����[4�]��wY�\���AcD��#�@?[y�}+�D��z]`}�!g*��c�$RM�����f�W�^�~�f��������s��'�Vꅭs�N������<\�#�/�^]��c;�,N<��Cq~�o�@�ޯ@?u�@���@�=.(`�,l�ɲN���9�<Q8��/�d���y$�}����� ΢���(��@>���[�"K�
���-Jcu"�2I4>�_>��r��U�^�~�f��h��L�d}�����.����/�����sk�]�-<��u��Yƭ��Н�Q�as���˺�U��&:un�������`U%�����������(%|���L�94�[7��<�H>ﾚ+~z{��?{�ESQ�;�wuw��� �w]a�IDEDE�f�~���J͑bq�LjI�E%�e��>�� ��`{�\\bT�$4F��@/[4�[4��@�wW�r�r�9���6�s#�&�r/I;$��c*�v��e��Հv#e`��i{<�)��D�D����女WZ�Wuz]���v7qE�Ɣ#�h����K�
�.������LU�1)0M94]�������h��}s,1aJ"n=�^V ~m��ֹ��Qi
"!�P�����$�{�e��wd�Mܺ�ͻ�=�[���������������30�ۆ��6P]�X�1�Pp��.v�q�\�Mc��n9����]�0"��/K��o0/��/6E�G�@X��@��^��g�$U�� >���?:�8�&��3CJ�+yi������ ����ʘIu�g\WH�#Jd���l�?W�h���9{���s,�m�7rM�}V��v��W_��~��$�bz"�]����s%�e�0�@���ݙ����Z�ځ����F+� �@��<.6:��۬������Ehz��s�[� ��cu��	:sa��ב�Ѳk�(�� ݂ r��cz�e�_C�+X0�ݷ-8!��q��ָ`���;�ٍ�+nfr-��t�G<��� QlK-�v�UH3N�y�"悭�"��ݟْNN^i6�-�2o����w�����0�F��'O�I��q/Li���mJK�99��v��zv@�k���&�q1��
�|�^�z��4��Z��9��x�B�=��^�}m��eL����Y�{s�蚴]�� ~m��ֹ�СB�r���W_���!dU51c�$RM벦R�`E�u�z����b��@x��@��@�<����� w��~���y%�p$���H��a���;�s�u�`���٤y�Im�l�m�(dn�Q�)��ޯ@=�f����ߤ�u`�w)%r��t�mY3���^fe�̟��������/uzjU��iB7&�����"������ ������o�j[��v0"���'���/0>��h�9��&$��{�h�!D%;ϯ�s�X��� �w�R)�Q����P�WH�W<u�9]"�p=i��֌��NC��z�sr-| �����Ku�OK�zYN6�8�NM�빿g�$U�|���h���/�j�"��dǉ]�g�� 7�w���/� �bE�1+���$X>
V �$H22 F
@��B@X(��B(� @"�F
H �H����B	H!�B! BHH$B DbdF+ ��`$P� �#`āA�0!"�2$ @�$�b2`I��C��K9�G�"F$j"B�a�	�>@O�{����DlIb� B��0`�B��R(�@"@� Db��2�		@�!I!�	$XD�!$A�$H� E$$0$#�H1$�Bb�R$#0a�I	!$$X�$Y$�!!	V@$HF!�Dq�dd��W�P� �OJ���|�Ub�(��DCIA
�D%����_v,�3�Tu���WSD����}��}׀~{l��S��� #��+�W4����]�ͻ�:7�~_�r�� 7����wx����xc�5�8��v5����jP�4���l�Q�������t����|w�1�&�d$�z��.��{l�����_���?��cIȓ��˺� �����`zΣ���ۜpG9�H���4�l�?W�h�נ{܅��H�1��rh���'��{y$���s�S�~�=QUz���C�y�7�O{���{�t���n��`z쩁r���=7��� ͭ������љ|f*�u]�u�vc�n���ٷnu��`Ǜ��muɗ�/K�
�n�����eL	�.(`� �' �z^����h�U�r�נ�[���A@s ԏ@�}~������9{k�*���R��&!ƔNI4��]k�*���m�@�4v+"�
F93����K�
�.�����Σ��w���[}z0۳/cL@Z�2�Vح..cZ6�=A�lk��om��:�%��Bn�si���)y&JƇtX��\�x|m	��cV,���@����]�8d��t���;���c�=�Tsu)kP�;���q��s�3]K���1����g�䵹�i���牂CbVy��P ����{�>L|�$+�Î] ����;��[��rkc�]�킕\�듙�1�1���y�trtD�)YI���kMG� x�ɒ8�W_��}m��uIu�����gvj7�V�k �����0"��/K��xBȬ�`c��Hܚ��s�*��U����@���\	�ٸ�v0"��/K��o0/�y�vz\P���bǊH7�W�^�}m��W������,�Ws�w6����Jrv��b���ý���0t1�m�s�<X9��dxHA��~���׌���
���-JmĻs���Iv�������"���K���hF��dYq�q��9w:���W$����������n䘱4��ۏ@��� �m�����uz��Y| ��9�7 ����^0"���.�?��f~�~���x}�ۤZǚ�^6��4�kpu�z��;@u�̐)��%;&1�ֻnl�+_�;{�`;��;���n���Z����Q���h�g�*��U�^�~���n���qC���9�r��$�����y��y :DD�(J!%S_7� �;��j�%4�xFA��~���n�˺�����s���&'n)$��w0P�BN���K�g�� �[�&�͡�=��PE�FD�v�fuŔA�����]PВ�=���3�GFs6|_��XIu�����P��n�IH��
���9{k�/��h����!de�,�ƛ������V]`U%�ނEdP1�I�n=�n�궽���<��ֽ�w$���Ҙ�7���m�R]`E-����H+v$��H��c��wR�k	L󰬧l��\�S�-!V�`�o>3ŻN#�Nw��?�����[��^0<���2a{��2<$ ӏ@��^�}�s@���@����R�������������m�R]`E%��%ج�Fd�!�3@���@���gu��Ok�� �
MMr���vWi�ݬ
�.�"���W���Y��w�����c,K�cC�c�Fi�$#=�����>�N�j	�l9�#���J]mt7"�q�#�[���c�����F��Z��^���P��a{
�[�ɚ��Rr���LRmX컞���m���Y�v�]v�M���v�D�^��p�ʵ������$���늴v���XQP���&�vn9��qmű��FZE�����^�۰Pg��w��a�yu�I�\�&�yz���ی�aX3ɘ�k�^�Vs�M�u�#�7"�������X�^,����G��}X�$�8�G�c��@����?+k�*���9wW�~ㄈ_��cƤ��m�^�XKu������b����݂9{Xz]`K�����mz�*�$;���"iǠ[���V�`E�u�.�V��,v���'jtYƭq��i�hm�^���q���Tkh4�hK(/\E���`����۬�.�	-����{�e7!7d�wNI?^���P?ER��IDM� �����ŀ~aKq��&9	$z/z� �h�]��mz��Pa����i��u��?6�`Kn�9DB���}Xu�|�<�E�$�@�m��=Vנr�@;����,���G1���_Uuu�lH�޺��բ�I�ۙ֞8���	�qHǓ#��}�����[���f�}�s@�=;0�Prdʛ�j� s��'�(��� ��� �[^�ge�bE�)�&�z�m��l¡B>�Q
L�n�?k� �+f

�1Ɯ�@��M�m�R]`[�	u%1^3�,�{�`y[u�T�XKu�}z��V�p��0�pX�B�d��c����vUQn]��l;;���2v����c��k9"�=���]k�/�S�����|�~�Pi�y���i��]k�/�S@�[^�Wu{�Gu�|�8yR�uWX�����u���]=ެ������"�x�ɏ$����\�����Հl�u�尡ZDBK�0�
%$�rJ!z>���`��uY6]݈�
�����>��o_��z��%T��sqCdm��I�A�(��m�m�Vm�qcX�qXX0�ֹ@�Im���<��{�j�������t��X��0��]�9[���K�dy�B�r=��s9(�6y�`:������#Ꙗ��W*�U�7k ;{����Շ�BQ�U���`~�,�R�4�Y2U�Wh����
z���:[������3�K���{�B�o��!Lsn=���$�{�/��׀9�u�R��)�N��A��T�H��@$�!	"B�Ad�bD D���E2$�� 
@� HH��08£�B�(��̑���@"�+��)�
B��JĠb$ƸJ�K�A� �1��x�F5�DO!�(T�$���H���W�)����HB#	!��d"��$$���*�$�"BF ���R`SŀW��!!L	ee\�"FT�I%0S,!�`Sd��BP�7T�&_AjČ`B��� �$X�I�����,d	�-���j�{Z;�n���գ���nΝXÓ<Nf��8d0�;	����g��r�3�m�����H�ie�ʛN���70�����k[[<�n���_6��eٍ�����v��}�٢�L���;��
���Zsŀ:놶����;4����Sz���)+�vѐvQV���t�渦Ĵ��F2%�f��@��$��[^���E�n{���Z�#³s�`
��] A���7 iܗT;,�Tk��l��ҚC�d�zSn�z����M�*�U���祙YV����te��ڌ�C/\l �vαcH��tC�`K��ƹܓ�����ۅ4=��,����;y�-u�p�Ц[gL��c�q�ʊԫ\8���g�6tU��$Y��Yx�vka��76�L�Y6�#]�D����;�n3��A>۴�eb�g�{r�U2�ͣ�lv�&\5UU�@ �gE����͹͎M�6�jR���G>�s\��f�n:����ۗ��Q�m�3�fܺ(
%�H�,pֻf� j�g`1��g�U�L�3quh�s��v]�A��;m���#��i7"�lŭ6V�j �����*��G�muhT�.`]�n��N��� MJ(�ݭkQ�	TGZ]��n`��n��ƪ��t�� q6����n@�Mm��mEƝ�Wn�B� 8���D�hmڮ\4+�rƑګ���k�b\�-�{�sR��j5��{f��W���c�%R�9-c�-�����A�YI	�3�A�ɷn��]2� �7k��]u�9�{k/g�EӀm�ӛl�Jۀ�VÆ؏�:��*��0:��l� �۱���i�h���[��i�PR˻>3)C�G���2P��\��4UA]6�� 8ڠ�󉝸�M�yU���R ����t.sq]=��9�.Í6�zZ��j*�T���mRG�{/i��t����;���C�q��<7<aZ�4wm��ywl���)i�[����S�DQ���9�TTy��l��iM�K�Uy��gtɡV�g�j&�+�v"iT����g�<!��7h�f��td垊U;8+�Z��j9���V����&��gԖ7]���vz��5��$�܎�RG���Z�p8m�d'*qrcg����[��[�BT�������^��k��p�J�N�͹h�k;R�&�rr�Ep�z�t��]��;c�d:*T|�������o���=�e�X#k��0u�h�������E�0�8����w%�u�)]ʕv����?��b��� ��u�~���Հ|�L�t]ڤ]M�eլ o]���
����Nw� ���X����3Ď�.,��D�ȰO�h&��;���(�(U^~�, ��� ��
Z��M+WSsWX��V�݋ �^���S��V wL��])V��mU�Wu�?�ŀtF�>��t�Հl�k�;�S��b��(�I�Jb�㏬s�1��4�Nn��-�Qi{;k���<��?>q�ݗFbs��r���
���9{k���;{�`�&��R��+UW$�]`w^s}X���2$H�`�`1���R@R@�$*�	(��� {���u���}�Pb�x��1���>W����w4U��
���?{�b�X�bǓ}��^0<����K��n�>�%Cj%�2b�s4U��
���9{k�/��huIx�QI�	#�¹o��}$������dJGIyDj�:tėiӤ������ L�@������޻���z��{�.9ƉD�`?7Xz�`K�X����(I$|�y�(,��m87#�>���=O]a�kQ�"D(̩�V �u���]���6���3@�^�@������q^����;�)�d��I�k/E�y}&�'�x���B�»�)	bJ���W"�qt��#V�=��}�ю�� �A�][!�9���x��R�`_Z��m�R]`{�,Y+�DC&8������
���9u�@��	���P�c�۬
����[��^0=�&(`�5	�`�z]���נ?�ŀB䐡%]�X �9�'+��R]�\�����ݽߗ�6{��
���{�x���!�b�$i��9�ՃS��Ҝ��+s��[d/;��k\ۂ�#�::�˷W%�Ɂ}k���XIu�#�hZK�XdS"O��3@�[^�T�Xm��}k��7&-��b��Z��XIu�&ڙ�_Z���א�6��0Oƛ�@���@����[�
�������w�s��;�qor`_Z����.�=3���x(�{{)K����ɶ[$!c�GH����u>��ȴ�.y�j���V-��a,L�I�u����|�� :ݨ'p"vsn�\�X��Z����V#������g�Eq�ie�@�e����z6���s<)�*q�)��
�q��#��[��$�)�����G&-�4�A�S
-��Җ��p��F�dn��;k�;l�̳&��3nC.�x :n|~;��;�cRv�Ok��z�����N�99%�N�e�m=;v1�]u��Wwc+���
�����S�׌����d�@l�@����v���s@�u�@<�{��E&9#l�ݬM�0/�x����.�
U�.((�IA���۹�z�נr�@�u�@��]��� ۘ��c�[�������׌��w���Wl8G�\���q�v���ql�Mv��5�l��M�zv�mi��k�+!vvn�wk�.�<�������-���Yw&�0�q��l�/��h���wW�{�Pv5���3w��}k���XIu�z[���
TL��$ԓ4WZ�
��`���yDB���� է)�UW�����f��;�����}����X��z���W��I$�q�HKY��X���\�k&|�q�4n��痲g��^����1��N=�v��n���^�WuzJ���K&8�Iȴ�).�*��鶦�����79\�U��`N�X��XJ�����U�_m��?p<�W#���b�XIu�鶦��)��k��"o��s"n=�>�@�۹�~]k�*�@�ަ&E��Iᑴ�I�+�$$�f�&�ӥ��ci]�4�`�C;����cq�1��br-�n��u�@����v��
T5&LcsjN���XIu�鶦����ߒ;8�1�}�R@L�@�[��=�j�/��h������j��by2aswX��:�p��Xӭ����̾f`>����������s��׌)n�*���mL����������L�⭍����]�R�\:�PT&M����8N���[�=�).�*��鶦��@yجPx��Ĥz]���ڴ�x��u�t(S'��sU� �쩫��>u�8��aВJge������?{�W c�br-����K�
����l���@]Q��;�Ě�f��u�@��z�������7��<<�{YY�
cX��9���D�n\ݴ�+v'�f+���έѝ����ty���#F�q��Wv�{8�ݵ�爰��ڝ��\ݶ���vQݎ��Ka9㇮�[�@�����b��Bu+,�u�Z�:�A�T�<���GQu��XFC�Զd+O��:�jP�6�ۦ��f66AW��[�P��;�!mlGE�A\��ȫ]W���޳����Ň|@la�Ynk�����Ǝ��m�"D�/U�d�fK�*��6.��<Q�k����v��?���鲦��`|���?L���)�$&H�yڴ��y��r�|������.D�c$b�9�z���ֽ?ľV���դ��$1����������>V���M�%=�ߖ�
MO+�T�]���]� �u�������ذ�u����{����i��֧�B��M�m�c�½�Ue�� �s�A�'��-�Zݸ��i�#�����-�s@�wW�����z�D(?��&�1��z�X�RQY�}����X��:�Ԡ��m�1�a1�&hﾚ]]a�U?Wzpw�� �|56�]ڵwP��I&�WZ�k���h|�ﾚ�ϯ�|)�$&H�k�-x�'��R�`}M��3x7yv���gX�8��ð����J���f���mbg�5>Y!�D�ȅ"r�����o�� s���%�7�~0�L�)����1&�h{�hwW�~�)�_m�߳1"���_@px)"lIɠt�Հ~{l�W߿D��h	8Q�C�F	T�
'��,`���""�@H�  � �$x����B"�F0�"�aՉ`����It@�7X*!֢AG�`�(���#������@?�<E3�<�~���O~��~�����
H�mǡ�������>���*�^�WZ��#ޢͨR�SV�f��9�b�=�ϫ���pzS@)�YS��15L�ߊ�1[s����u��bn�;�:�n�l�������c�cRL�m�h]�@�l��/D}A���`L�7�Wv�]��UAW|��mL��0%�� �^���bA�ϯ�}��GS�Z�}>4���н
���^ޯzp~c�j�.*���hm��*����h%�ݦ��4��a�L�q$���k�%�S��`Kk���w7��\���v{Vۨ�9D7VЇg��]��G���n��י�%�b�0dŒ8�@��Z����׌
�����,���1I�H�l��׮�U��_U�{�Pu��1�M8h���*����h�M����ӄ�Ȝ��UmzW�h�M޻��N�
G	�I@N=��h���8�wv, ��x�BB�!C�P��w=�����&\&K\�Z針h�Cذ��6٭�����m�~�l�z�g�x�x�9��t���h��/X'���n���wI�
5�#�y�<3v�/]b�լ��z�VP�Ų�q��j��h��61�r�ݭ�2q][;�vN�-��8w�b�ҵGL�-ٗ���w$�K	cMO�( &�������{Yݭ*q®�a�g���)]ݢ݂.ߍ�T��F�;�0�ٻ-�[n!�I�f��7b�;ۓۧ�mE0�ec���{�Xm���w�7M� /�rX�<��H�z��hwY�Z�Z�mz��W�E1Ʉ�m��*��ݵ0*���^0'�ˊ�o$j7$�@�ڴ
��@�n�U���!dƝɆ(��9"�*��[^0*��]�0=i^�չ�[��X6�27Q��g�Ġ�=@��.�\m��盭Üḁ��[�g����^0*��ݵ0*����[��a���nO}���=@D�"B�iD+'��p��[x��5M�q�x��rM��h���m���@<��W��FLqh{���Kk��M�=6D�3�LYrS�RI#�:۹��f��ڴ���ּx��Y@j$�%8��sҌڬ\u̓F6�[+��F$×@<�dxӉ73@;����h���z�h��Ⱈ@c�$�G�u�S�n�%���n�>�;E�)#rI�U��m��g���3<�ƪ����}�
��A!��7�m��VנZ�ZVנ^傦��'�LS	$� ��4]�@���@�������7�F�fY�����"och���L"�r@���n��l0��ݵW����T��m��m����?\���âpq��Z�v��w4��>����� �r���&��n��� m��ޗ�������ԕŷ3���*���X	(��������s�����%�� �)j�e�"��m7&�k�h��h۹�U�_�o�����0��Rčp��*�J��-��;sņ/<� d�[�n�t�畻��8�n-�e4m��*�����|�z�P�	�hCs�Z��hIu�nژ�j`Y
�n��̙0�L�*�@�ڴ�h۹�\���D�l`�H�G�Z�Z�j`Yk�R]`�I�n��i˱v-�����S�^0z^`Y����?x�[��^�ܲ�%˒�c0-��3h�-j�h{�*��VJa%�		b.��ۮ�]ͣn�,^�!�u��W!&J�Xs;�s4����.��9F2N�̶�۳�q��Yrڢ��n�	b3�����mn��6�¹��nN#p�1����A��\m�vB�bY����K��u���A��hz�v���C�U����1�����_>����n�6P��{X�˞�ci�!n���6���q���F�:㮳�ԅʁ����{��͵0>�ژ����<���s4
�נ^v��h���=�yqXH���q�5�fژm��e�Ku���Ln�L�'�@��Z�w4
���/;V����cMF�'1����ŀ9�� Ss�=�� �?C'G2m�����q'=��<F^���^�w[Z����۳%����tF���?��^v���Z��h=.(PN&�G�Z�[���DD(UC�np�o �[� ���:�&)�'�yڴm��]k�9u�@2��ˑ�S!R)"�=��`U%���X�j`K�+�x�H���6�hwW�r�@��V��۹�vfs�y�br$H���ˑ�A]nܰ�����<s���m,\�a��ɩ7NG�r�@��V��۹�U�^���&7aFL��8��0>��`U-�R�`{�B��NDa�̄�h�w4
�ק�g��T滫 �]Ӏ}�(�d�U��բ��`u��6u���s��"S��~����Y>Bq0hp�R=�Z�6������n�"$+�غ0 �+Y���Ƃ�skrx�|��*���#�]��'�x��D8LSN=�h޻�]k�9{k��\��F�r������0*��/[�6����U�G�<I��3@��z/mz�j�=�w4ރʋ"`ڎ.\�{Xz�`Y����\y�������$����i�݆��7f۽�6������n�"������9#�v�n�R�勧uld.N��v���ĻF�Y�9PUI�qX4c�7e.�I��+�R�`E�u�fژ�*�k� �L�*�^��$U�|����{z�h�.,�	����j]�����͵0=ex��[�˖��	1�i8��ՠ{z�hu�@��@3�\YrO'����LY^0*��/[�6����w��)J�hX{�H@(D���$a$	1 H�$�H=:Ÿ0��!$I�^�H2A� (D��zN =cQ��xB:�q��$XB$Y��H��h@� �H���*I@ ��T-#$�$
�,�$e?&F$0bI��	1@�1�#!I�	!$ �H�E @�
���bP��@�%T$�E @��5�� FF!=�����Ru�-��Gi9r$kf��@n�^�a+8�પ]뇲�:��3�D���v���t���2;,>t&��t�Ӝ.�y���AYndK*�וU��<N�PԵ �s����Q� X��UM���\��$;4
�ή��'k8*iӴ[.eF���d��v�9烰٪ez|�@��N����[�d�΍V��Ȍ��QlN�Ό.\v���v�UXړ���{c[����m�I@e���h�v5�����a#�2���2���s�!�VU��/k��Bp�ln�҂�Mŝ���CJ9i9�SA����ث�xza�=(֘&�m�ks���>�ƸTKn-u�����j��h(��=��`톳�{ 8�{ 3q�6�Op��M�"��8���[JDU���x�;�N�d7�.rm9P�v�z�oS�6ۡ�����UUK*�i@ݹ�f�芊�tE[d��gS�ە���X�6�����X9D�X�6�����Գ;6X6[F�F�80����[Gt���m��B̰2�mK�,�z@}Vh�.��6��n^ӈ��5���*���m��%��Y��l����:�2ǒ �!$��y�펈�2��������\F�v������mq��<Y:8%y�s����v�Vv�y�y�#
�4�����]�&vc�'�fnm]!vx�5�\ت�t�
�w ��+��
J��8���.�s�G(�U��	��Bcl�F�H��	9��n#Zʂ�D�ca��h��=r;��Z��+�YPe���m�M�3�,�ek��p�6�U���gd�2���� �UJ��U��˳�*�۴s�O[��7G=��I��h�[��!#�d��m��do�>]u ::�UL�p ���YI]7k{m�l�Cį4�D\/<��j�!.n^���� ���v�9 Ж�3����cq��2�I�9�3'�nl��6f#��:�� 8��烥 ��	���~��~I���#kۧWCa�8|��J�kC��ug`��Y
[��혱�@p5�{i���֤�s���DV�oT]��Jv�{*m���j���R��r�� 9s� �#[R70�E���=&�;(���;!�%�g�6N���D�wg�;���<Y��2̻Fm��ɸ�%]�Y3O9�h���i���ܥ=Jt�p�t �vɮ����w3gb0�m�CX���	���ܸq�� �(W.���L�:��(�4�d���pi��=W��9{.�,�S�+��ʋܴ�r��w�����j`}ex��[�{��cv%
dJG�^v��n�WZ�]k�=��(_"p�cs8�������n�"����mLx�R�&�X�SG&hu�@��u�=�� ��ŀr��)_h�ML��`����ϟ>o��ٻ���ݶ�*�x�3c������F{.�!O�m�?z����u���u�����)]ԫ�T�]`i��B�J ����
�נU�����Y�F&�Ӝ������.�*���mL	u%q܃�N4�i��]��wW�_]�@����?z.+"���6�s��W���ژJ�T�XH}�˭�n�t��0�ه�����յeq�q�,{u;+{Y1�m�㋤��6���W�
�����?���%��9a"�"�/[��y�bG�ߞ��|��h�r�q,lpyuv�;���n��Q��JR��9��A��Xh�J����Eժ�&n�tB�������� ��� s�� <�{�^$x�4�z�ڴm��]���נ\����XH����Q�U=��"Ͷs��6�mӵWs�	�;)O,�i0�HF�@�۹�Uz��Z�
�W�ui*ːQ	Ɠ���0*��)n�*���׌�yQdL18FӒ8�]k�*�kIJ�w�� ���X�J�4왛ɑ)�U����h^�Bf?1�DP|x���_�o�g$������&�&Ez�w4
�W�Uֽ����癋=�G�5X���O���u�{gv#^�n��4����k�����wl�ul�9&z�����u�@��z�w4靋%CpxG1�&n� s��y(Q���O�Շ�L�����������u�Ƞ��4�z������Тg��V��� f���Q�nH���h^�@��zg�/���_�K�?�Q	ƛ��1�U�XKu�U�XZ񁿿}�������K���Mzy��&�iK�]]L��s�i��b�^v97`�{qպ�ӣ[<��n��'6�q�;>=��v��M�N��P���3ˍQm��\T���.��kf���D��q�ml�v9y(:nk��g5ہx�-�<tvѝ�>�9څ[�NS���r��O-ש��m���z���(̜���;=���<uqm�ޫ����%îz;]��֨\�q�D�Nl^�mݝ��L�Ѣޗi����"i�~�����*�^ �o��J>����X���j�@*U36����/]g�$���݋ ��Հ9�u��DU��l�L�hEj��� ���`^��艗:��r���z�$�ǉ�6���f*�W�r���
�W�~��h=�%iD��cP���gu����}_����`^נu�U0��Y6H���#���%u�s�x�I�(�tbS�(������瞋\��~��V��� r���B��������Հ�:%zʪ�U3WUWwX��,�	)���X��� r��tDDL��%Y�Bq��s4���z���*�^�����;����2x�"i��D(Q;M�`<����,��X�y&4�&�%�dJG�Uz����}ߗ�:y�`N��cʢj��[��n�h�d��tm�����rp�nݵɌ�G��l�[�8Èֻrut���~}�� ��gu�D$�Ht���>M�=�kq��2#�4
�W�r�@���ozIz"*�&�~���Eբ�fn� ���`^���0������ϫ !��N�J�T�J�����Q=\����,�n���� &�����D�I��׮��y�?�����=�k�?u�'�G0DM���q�G8�'����\V� [yݞn[:�]���(ɐɉƛPi��*����^��\�~���b���O]ʵ%YwSWwwX���?yBP����Հ}ϱ`[u�
�(UC�U��YeT�Lڹ���=>�� ������ ��]`}��d�,�"��uuu�Т~��� ����'����$��
U<���9�(+�k����NL�*���QZ����Հ~z�`��*nM���j�5ˍ��ّ7E�:�7͙�,�l072 �����`�IǠr����� ����P��OwV G.讬G��,iH�
��@��V׀}?k��Q����R�����$�z_����k�=^�zVנui.e�(
Fۃnf���y����=�}X��`y$�~��� zR�=w6R]���� ��u�r��I(��ޯ��{ذ-����u�\�˹���W8nV������������dz�4��7Cy���:9��9���n�lց 3�n��;���̇V�b���I�gd@��s��,u�؋K��(�1�2/n�Nȵ�I�7X��Z��܆�]:�Ա�m�n���5�]n�h�`�I�6۷�L.H͛p��Y6�������&�N�rAt�g�������v��Э\s��6��=��L�盷`�:�]�u�9��e[�����Հ~m����Т#����!A|�pX�I����۹�Umz.��
��~�3ďiA}�k�Aa23�4��|�]��[^��۹�_L;���$�z.��-������=]�Xs��C�ؠ<iH�
��@�۹�Umz]��{ܱQ���1!G"�!����c��v-<����(��x��kk�\�~��qo�;��x�$������*���uzVנui.e�(	�ӃrW��P"������۽�9��� ��ŞP�G�.S�r�UUjcrI�Uo�@��Z�n�u�h���`��$�R`��@�mz�e0[w��	)t�V��*l���h�2&�@�m��m�.��
��@�3����0���o$i�R(%2�<3z�|�{m�O;S�+����=[cb��j�������}��*��UmoP~�S@��p�\l0�a&$��9w:ΈP�N����� n�{^I�844�zVנ~�SN�ŹC��JZXV��ۄ���zL@��B"�dBFE���CA8%Q���A�S`� ��""�$� ĀF$ b��5]N*��x�
�@ �jpz pb���}�I=����Z\A`�DO�z��h�����
��@�Ĺ�bj2���0�� �(t�W�:{����h��yΉɀ�#bja$m[�n�v�u˳�[��;��.���&9�^�犎.x���M�uzVנ~�S@-�h���bv@����U��>���-��Iu��D�p�j��#�@�]�@-�h���*���
��,&DcR- ������I;{��$�"-�����۲��z�J�h�9�L�@��� r۬�M� 7���
#��Oc��6$��tG<�m�s�v�f�A�[W
\g�7��vy�d)����Հ~t��z� ��u�	�bU�dd�<I���ڴ޳@��^�U���K�p�#��@-��Ku�U�X�*`}r�r�%R�
�����)u�Հt���=���z���,���"X��	K���8%���� ���?7Xy|Ϣ�b�\X�i�	�-m��ֻanme�T۵��ή�<Ҧ���{.���ݺ�ض�!HC؉�����%�.�c�<��v*���j��_Y�a02���؛j�&	�}y$L;���=���.tJǨ�=;p(����ݯ/+v94��6��WK�ݚU�A��.x�$
�T{p�S
4rQ%��O]m�ݮ�o��ۨ���̜���xT��b��Xa�u�m���;�	Tܽ���kmzt%�
F�O"qH���nh^�@��_�y�__��Ԡ��6E"@�3N����n�"����`\�;W&<"�JbRM����W�^��׬�;/x��I84j[���ˬ/Q�K/0*�� Χx��l��'�9�}��د�����=����\�t��y��EѥN���;i$�V�c��7g=�fS�����,PI�a&2"F���u�4
�]`/]t~���� ��.S�r�jT�i2���I���~��C����P��U����u�����\�Q�H�q��W�_l��[�hwW�~���cPI�P�=�e���.�*���LW}ˢ@��#��u�4
���9^�@�۹���x����jH��Q��f�|q@A�9c�=m�c���Φt�ۈ�Y�㍞�L�R<��+~zW��/��h�f�y�{�^H�I���#�*�[�׌�y�T�XZLA�7��$�$�z��� �٧���1*�W�UmzV%ȸE���q��hm� �u� �X����`0��z�UȊUh������9.���}�}��m�sⷄ��<#!���.����Wm����v4�9Gpnnݘ���n�d�!	�L��@�mz���u�h{���R�cP��U� �׋ 5�x����۬�ďiq}�l�D���93@/�}4
�.�"���W��	�u����	<IɠU�W�r�����?�ŝ8���o�o�o$���\�������5.�`Em������J��~����y?^z���Jxv��u��h�2�v�N;[��v�Yz]'g>[��J������`�� s���!~�s��=�Į/�D��	�D�� �l�*����۬�^9��G�e˦�j77V�W��R.}��[oh�BɕŒ#)�"����@��� ��`U�u��T�r�oo.㷵�_K�[y�W��V�`n�f癜��Y#�) �����L�ycB7m=��N�����9�z�:�U�h7�^v��1N,�}��cm8J9�mv�nƭ�.I���c]�E�ɜ��i�.{:u����K�Qլ���,v��=A��@V��ͮ8����(���O�����79�/��D�gd���X *ǈ�����:y�pW"��=�cį;��=o�܎\�pR<�pQ/��:�l��93n�b�p��rs��nI�c#Bxd���phi���l�*���9[^�_z���d�A��]�os�K����/��-��<�ƨH��i6��@�mz}�xtB�	L��� �����q48)Z��UUwX�?�U{�׀�z�?k����X�"�H��S$��4[w�9�]`-�����=ϿU+����=���h�(��]����n��p��t��wm8���{������.�3��-��z_z���a�DH�(�BQ=�� �`�`�`�{��o �`�`�`��ݲ�>ɳf�]ɥ���� � � � �>�����G¢�u@�G`��A�A�w�7��A�A�A�A�{���� � � � �������lll}��K��nf���ٛ��� � � � ߽���� � � � ������ ؃�r9������ � � � ������� � � � ��l��f�6��t�7x �������x ������� � � � �>�����ll#�A�{߷��A�A�A�A��N���v��3d̒�� �`�`�`��{߳��A�A�A�C�@���g�A�A�A�A�����>A������>A���Z�t���o6�Kt^u�h�ٻ{:Nͱ�944t왳IV����'G�.ɺ\��ne�����666?g���pA�6667�~�x �߾�x ����8 �w��r}&I���.n� �`�`�`�~�ﷂ�Dlllo~�����lll~������lll{�}�pA�666=�e���m�̹�n����A�6667��x ����8 �}Oʧ��B���q�QF"�Tx ���<�����A�A�A�A�����|�����ɿI~7M2\ɥ������lll~������lll~Ͼ�8 ���}�|�������>A����ݲ�>ͦ�0��Kws��A�A�A�A�>�����lllP�A �����?��`�`�`�������A�A�A�A�;߳��A�C��wx���w���]ܴ�����]r�a,-�� �n�%<��q�� �m�\����2i��.�pA�6667�~�x ���}�|��������PO �`�`�`��}���� � � � ��l��f��sffKww��A�A�A�A�}���� � � � ������ � � � ��}�pA�6667�~�x �O� ��A� � ��}'�7n̓sr�&n� �`�`�`���}��|������~�>A��A�A�{���� � � � ߾�����lllk��~�vL��ne���� � � ߳��I'����m��%�(\�B��}X �㢞}��1�#��@-�hwW�Umz{jǉ�ő�IF�#x'^b��q;r�f��D�ϕ��ã`�#ldq�0F�,Y$q�4�f�Wuz�ھ�������há�I2d�9$��S}_�ޮ���w���z"�{�Bɉ��&<Q�������f�{�����}�b�o#�1�����@=�f�Wuzy������{j�f�D��$�z٠U%��ژ����FL03R���m��2��Q.���A�@�D�*�)�x�|�W�|񠇀OX &/��HŁ�$���� �H���x	$#��ۻ��{��χ�UԫT�rv�<����h�����tD���Uak�j�:@�>87fݜڣ�wN�F8�Lyr�ed�[crez�{	$v�Õ8����\�M�]mʬ�r���8�v�k�ض��Qښ��n��1�%6�������.��xX����Fw[�uZ3WGj-xU�V|��m!X�ɺ�t�m���onԨ;;�s`�n�p����P�xT����w#�]��g�6��kg��Pr���rà7k���=�;��E�p
2�[��U��W��InX��ɲ�bAMq�V��.N��b��l�p�q>ŀ�(�i�w��t���T^\��]\U��<n(�U]-��=�J�@ye��٤ː�s=�8��&G����7n�R�7&�l@�0��nۍ�BI6ͶO�DF�@nî�	���lG:]��@�UU1��hY�g�*�UUR��VY]a^G�pH��IM6+6�@u�r�Hn�����`N�6�{r��pI�����@u)��ֳ]�de�'B�$�\lh�`H������ǝ�X�3g��]�k"�����V���s;���Wr�k�[��Rܪ�'I\�n����s�6�X6E5ӣ��9x�w��h�;�M���0nJ��M��� Fx����Q���g\�����G��j����գ!��q��$��j����ƜJY��6��Rqf1����X�����ݔ����:;aW�W�uU/;1Q��59�T���q�pYe����"fWTF��.��Nλ3�5�6N�%���:�H  5��l2�i&�	Вަ�̓k�8�eY�r�m�����34��U*Ӕڤj��y�m���ƪ x4ysC�j�V������*VVRg����JjiW�;T�@P6[������v�w �R�M��vñ���>	�n�Ľ��;i+tkx���C�m�b�î�ی7A8����h7j�e�3so��{��� Px�4}@tX�@���Az��Ν��IsL˻�ew<j5�vHX�,�=FY�*<�Y��Gv��p��{�Ar�u�s�wgv��V���k����.�Q�n.���+[Ok��Z�6Jp�NR�G�Unz��ڻk݄^jn+���Nո���%�n7�����a1Z������XiNS[�I���,Q!�b���,��[�)@k�g�����>7'��)3ôe�h�c�6�tb�y ���Brj�bd�uu�b�0h�g�U<�:YL�ށ�۬�� �K�呂ys�>�I�N4�JG�{�ՠ�w�n�������JdrqT�4�񹄎E�u�h��h{���ڴ�K�`���ɒ8ܚ�y�)�o� ��Հ~�np<�������7�A��d�s"rhwW�r�^�_z� ��h�]x'�mLcR��/n���ӟ�ڬ�B��u�vƂ�q����YM9�M�m��Kss�'o��9 k� ׮��_�:u�`oL���Uٳfl��ss�I����'�E�bQP"āVE"�	�@qC�͓��7�~�X��Y脡D��rO!e�r�����@/��U�^���z}�hx��$x�4���@���e� 7x�����׀�88�pȤ�z+���٠z���Т"'�)]T�]ئI��
p3ٸϱ�����+�k��'Ѷ��q�x7��w{�:<����x���#���M ��hw]y(K�}X�R5=b�f�V�q�4�Y�U�^���z}�7�3<�=���I��"�M�����ˬ���y�K/0=br�s��I8�W���Y�m�g�y����w|�(|�qBD�z}/0m�^�X[u�}awsś=���rЗ38�\��8%�pr�b��9y4��c����������E�5�a9? }��M�z��k��Y�u���I�8L$�@�ޯ@��������:S!wA�]E]%YSwXOwV ?���
&N���:z��:��4LC��r= ��� �w�9�]`B�	�/(����U%��1�d�nM �٠U�W�Umz}�4y�\V�Ʊ) ��Yضk���=�vwh�Wnٳl�G[b	�h�̓#1HLN'&�W�^�U�����m����'q�dq
'u�9m�z&C������;���Df$wT�C�8H�rǠw�M m�á$�z[��:{���j�e�*��wrM��r���
g������
��@/���\6)&L$�K����9%���������j� !��r���w-���0=gU���@��ƚc=&�l���p�ːm��$�;C:�ٸ˸I�X�[u�y�{su��3�8�ʉ���u���x�k��[��&����S:F�xO�Y����F-�m3�Jx9�O!�w%81`Ÿy�`�p=�C�϶N����=5�CS���B;��gXږ�&���l���GF��I.P�:z��9`kl`�㷞�:�����������]6�l$��jGc��K2)�DI�H��v�N*b�����ۚs���s�0jG@��= ��4�f�Wuz�r���S�r= ��4�f�WuzVנuƎ�a�� H�h�����
��@/�����I���(ۓ@����k��@-�h�!dn��A�ܓSWX��`�P���� ww^ 纽�ߛ�2G<M��`�S/-��f�b�1s�=q;,xE3�B#F8���ѵ4�"�	�������]��^�@��b�=QC"y#�'&�[�m��j�)M�ӏ� ��Հ�� צ$���	$�*�@����l��� ���284�Ĥ�V�`�� ��`U%������8�m9�W�� �l�*�@�mzy�:�9�H�`����7��U�""���V%���y��\�q�c�!��xI#��[f�WuzWj�*�נ~�t�21$�8㗀9�u���d}]Ӏt�u`�� �y#w��E�q�]�@��kV�q	BW�0�{׀9��`|�T�@���2H��@��^�u�hwW�uv�����E�O$pIǠ��
����mL
�n��
O�a��n:o����|�(�rv�g��ۣ���W%bŧ�n�[��7�Λ�qΚ�"��'K}X�np?7X�����J8cR�R=��mă�\ �l�}�?��<�H3�|o+�2A��z�}�������Vנuv+$7<Q��g�bWﾚ�ߞ�=��s�~W��Q(�D�P��}�٠w��2D�%�#rhwW�Umz}�h[f��m���$���wP�.\�u�ڊ��	���!�M��00��gj�Y1��}�N�%?�o�����l^�h[f�WZ�}�b�@���ԐN= �l�m�]k�*����Ď�����QB'�}��FR�`Um�R�`K.��d�y&L$�@��zVנUֽ�S=�׀�8��]L݅�3WX��`u��m� �[���
M�lC!sۧ�Kd(�V�s�ι�,U��C8�E�`.}&��{[���4���ˠ��⠳�;8�T���7I�\/9�tX^��&3������v�&�:-;i�An3\f�wK͕�[�s��Lf���7�m��!k)���cp�Ng�x�f�;��ݪV�bT���b���l[]����S�n�+c����m�W;�+��<F~Q3<�|�l��]��f���f� �H�Mһ�1۶�kb��ֶ{<���E���x(��m9�����z����u�D~�}]Ӏ>E.S�*�rG#������[^�WZ��WQ"hsrhu� r۬?�!%䒊���^ {�����dN� ����[^�yڴ�f�WZ�}�b�@��"q�R�����K�%^����z��f��,��x�kpX�"Iģ�Nf*��cr�D�������a��8����8�<=�[�Mݓd����%�bX�w��ND�,K��{�O"X�%�g{���Kı;�����Kİ{�'I͹�k7M0ۛ���bX�'s��8�C\U4Ā���'�b�~|��,K>����K�dL������<�bX�%�}��r'®TȖ%z}���pܗvM�nnq<�bX�%�}��r%�bX��{���%��C"dK>����Kı>���q<�bX�%췮a��r䛓%����Kϟ�B���������%�bX�n�"X�%�����'�,Kĳ���r%�bX���t�ْe�\�ۻ���Kı,�{���bX�'s��8�D�,K�����Kı;�����Kı?o�~S�NtY��]�гv�Ll���/���rŭx]�
nnC��������P�4˳swSȖ%�b}����yı,�{���bX�'}���<�bX�%����Ȗ%�by�l�.t�$.�ܗn�q<�bX���ND�,K��{x�D�,K�����Kı;�����'�	�2%���Jo�sٸe�&��"X�%��w�Ȗ%�bY�{���c�;�0�����Iʙ�dX��uT�yB���!$�(!V�eaYR$%%eB����D� �q�F[e�	%��$�$!ز�$�YHXHŉI`Y$�HXI����`D8	����u���0D*����(��z"�'��g�>臑?D����Ȗ%�`߻�jr%�bX������7)���i�f��yı,K=���Ȗ%�bw=�s��Kİo��59İ>�>�>��<�bX���KfK�5���m��ND�,K��{�O"X�%�{���Kı;�����Kı,��wS�,K��{�-;]?S�9�6t}u�$vݫ�N�ockn:���q�,e�u�{y���WiB�?����X�%�{߳S�,K����'�,Kĳ�{���<��,K���gȖ%�bS�>,��͙s&��n�jr%�bX��{���%�bX�~���Ȗ%�bw=����%�bX7��59ı,OzM=/vd&ᴙ�wv�<�bX�%����Ȗ%�bw=����%�ȫ��o~�59ı,O�߾�O"X�%��I�����R�4˳swS�,K?���>����yı,�����bX�'o{x�D�,}��|������r%�bX�{e9s��$6�Ɇ���yı,��ND�,K������Kı,��S�,K��{�s��Kı;��|/Wr�P6�⸛b��2O@!��!�5WN���'XP�4/C�l;���bX�'o{x�D�,K����r%�bY���~�'�%�`�����Kı<�z^�'��͓L�7oȖ%�bY���NC�@�D
�M�bg�gȖ%�bY��۩Ȗ%�bw?w���'��L�`����d��Y�nI�7u9ı,O���8�D�,K�}��r%�bX����q<�bX�%�����Kı+��^���7ffKws��K��`dL��۩Ȗ%�b}���q<�bX�%�����Kı;����yı,Jt�r�ݦ\ɦ廛���bX�'s�{�O"X�%�g��u9ı,N��8�D�,K�}��r%�bX��������U�vg5ڎ;L�7A���K���v\ck��4�:[�A�\=���=A�v���4s�ZCָ�u-��۩��]X;>k	��M㖓���r���iq�6��gcI��ׇ\�����hE��scla4�����۳J����L�\`� �5䝌�(vݼܡ&�W��^�S ����l�'�ғ�q���z�$��l0�3eɷ3�"�{�y��+�M�ꗱ�^'�� ƫ�k.�d3Y��u��*��]����%m����<�bX�%���u9ı,N��8�D�,K���t?��DȖ%��{����%�bX�I3�>3w2�srnl����Kı;����yı,K?{���Kı;����yı,K?{���Kı<�S��2a��rm��'�,Kĳ���ND�,K����'�,~ dL�g��u9ı,O���8�D�,K����\&���&f�"X�%�����'�,Kĳ���ND�,K���'�,Kĳ�{���bX�'��K�fy�۸i�	����Kı,���"X�%�����8��X�%�g{��r%�bX�����yı,K�������k3S�R��[I ���l�M�B�Pcjf�ݫ��+ar��7^��:��,K��{�s��Kı,���"X�%�����'�,Kĳ�{���bX�%};���sd��rd�w8�D�,K�{���=D~E+�6%��wϯȖ%�bY߾�ND�,K���'�,KħK�;�nf\�vd�����bX�'o{x�D�,K�{���K��Dȟg{�q<�bX�%�}��r%�bX���zY݅˻$�ݻ�x�D�,�Q dL�}��r%�bX�g{�q<�bX�%��wS�,K����oȖ%�b~�=���<�4L�^��oq���}��8�D�,K����Ȗ%�bw�����Kı,�{���bX�'��}�{���D�,e�l\��[/uƞ���ҁj��8X��mn�Rx��w�/�tq�:M���~�bX�%�}��r%�bX�����yı,K;��"X�%�����Ȗ%�b{=���˒l�0��nn�r%�bX����q<�bX�%��wS�,K��{�s��Kı,�{����S"X��:S�3͆˷ve2��Ȗ%�bY��n�"X�%�����Ȗ�+��RSblK;��"X�%�����Ȗ%�`���l�s��t����Ȗ%��02'����O"X�%�g�}���bX�'s���'�,Kĳ���r%�bX���^�l�rn���n�q<�bX�%��wS�,K��?o��8��X�%�g�}���bX�'s���'�,Kľ��^���m���\���8󂧑���f�b^zV����\��v��Y�U՜5^��oq���}�߯��%�bX�w��ND�,K����Ȗ%�bY��u9ı,OzM=�읩��������7���{����NC�DȖ'��~�'�,Kĳ��ND�,K����Ȗ%�b~�?s��y�"Z�w��7���{���{�O"X�%�g{���K�dL��{߳��Kı,��S�,K���Ngw)$6��.�nq<�bY���%�����u9ı,O����q<�bX�%��wS�,K�O�QA�P/"g7�gȖ%�b{=����f�p�7m����Kı;�����%�bXG'��u<�bX�'����O"X�%�g}��r%�bX������kg=(�=B\����մI��n��<s�m� ^6Fx2k��lq�-n���ɻ�O"X�%�g}��r%�bX��}�q<�bX�%����Ȗ%�bw?w���%�bX=;�l�y�Y�i�����Kı;����yı,K;�wS�,K��~�s��Kı,��ND�,K����a�in�L���Ȗ%�bY�{���bX�'s�{�O"X� C"dK>�۩Ȗ%�b}����yı,Jvι�3p�r�nf�"X�%�����'�,Kĳ��u9ı,N��8�D�,K��f�b<�y��:�3�bXE#����'�,Kĳ��u9ı,N��8�D�,K�����Kı;�{���%�bX�����$�y&�t�5�84����KR��7\ԩ�ʹ�+N�7K��@��^�� ��q�v�`)�s��`�����`�Dsl���u�%�][�)�)�=��n9��:�[2�	r�0ر��m���
[p��Wl\��p Ku4Y�ev��9����u�VR��]e� ��˃���q� s�&�X�������N���\�O!����(g����w�{���ǇU<&)�Eu�u8���$�O^���R�G.
)7rŨ�Nn��&��|��{��7���߳��Kı,��ND�,K����O"X�%�g}��r%�bX����v�7,&l�nf�Ȗ%�bY�{������,O�߾�O"X�%�g��u9ı,N��8�D�2�D���鎾�����U^��oq��N����<�bX�%����Ȗ%�bw=����%�bX�w��"X�%��ҝ.y��rf�I����Kı,��ND�,K���'�,Kĳ��u9İ?ɑ>��}x�D�,K�ﭳ%��f�swS�,K��{�s��Kı,��ND�,K����O"X�%�g}��r%�b]����v>�t� ��x�H�x��3�4���ݷb9�4��t=�o>9��Di�-��'�,Kĳ��u9ı,N����<�bX�%������&D�,O���8�D�,K�Y�}�Ks.���n�r%�bX�����y���r&D�{�y�Ȗ%�bw?{��yı,K;�wS�,K�����;��w7$���ݼO"X�%��{�ND�,K���'�,~�DȖ}߷S�,K�������%�bX��;�{�f�&ٗsq9ı,N��8�D�,K����Ȗ%�bw?w���%�bX���19ı,N��Jp�m0�n٦nf�Ȗ%�bY�{���bX�'s�{�O"X�%���y�Ȗ%�bw=����%�bX��y��LɰT�mw;U8���)�Ϊ}�ⴀ\��ncI(f���.M��2FkM^��ou�bw�����Kı;;�br%�bX��}�p<B�H=�q6	 �{=)��6sܔ��x$�H��}��;ı;����yı,K;�wS�,K����oȖ%�`��m�%��$�4ٹ��Ȗ%�bw=����%�bX�w��"X� �1^�"y=�;x�D�,K�}��r%�bX���nM͆�[��ws��Kı,��ND�,K����O"X�%�{}��r%�`�L����gȖ%�bS�>s�3p�2�nf�"X�%�����'�,KĽ��q9ı,N��8�D�,Kޮy�y���#�W�7��A�nF��:^r�:��Z�=Wfv��XF�VZ��T�3���<f�UT|�~oq����}��q9ı,N��8�D�,K���"X�%�����'�,K��Aѧr<��RG�i�#�G��2�����%�bX7��59ı,N����<�bX�%����ȟ	�2%������6����ə���O"X�%�~�٩Ȗ%�bw��oȖ%�b^�{���bX�'s��8�D�,K�����ɴ�4�n��"X�@ȟw�}x�D�,K�~�q9ı,N��q<�bX��	" � ������bX�'��J|fxl۸eҗ7oȖ%�b^�{���bX�'s��8�D�,K���"X�%��w��O"X�%�Ol��3�K�-�7wsBI�&h�Aqu�����'f*��.Ŏ��$�&pc.�Y&馓sw�,K��{��Ȗ%�`�����Kı;�����%�bX����'"X�%�_N����ne��2[��O"X�%�{�sS��9"X�g~�8�D�,K�{��r%�bX��{��yı,Jvν�3v�&�.f�"X�%�����'�,KĽ��q9ı,N��O"X�%�{�sS�,K���Ӷ����˛�����%�bX����'"X�%����É�Kİo}�h}<��,K���^'�,K��>�3�fɸn�ݗ7q9ı,N��O"X�%�{��"X�%��w��O"X�%�{}��r%�bX�Op�2L�T��ZF"DD�S=��v"��
�b 0��@�FD�`F�6�������1����D"�H�E"��H�, H#1�����AI�V6H�-f-�$x��/��V4"����BB@ F2B,�@ @"Ř	
�l�6�~��hH�J�����H�@���"H�H#"��dB,H�H��"�X�FX!)�B,���H�b� ���1AEXDDa??�MMX���� $$BBT��??*�V�A�"�\H��yџn�cx��٘Dة넶e�p�8��0!N��j$n\�[�u��Э��提)�[�٢.u�ݛc"�Qў6���R�z2+\��l=��[O'N�\�7��1���9�(a�.�m��آ��)�D��ۛH�%<��:��� ɍ�헷,.R�5��=9vk�7�z	��:[nυ��g^��G��닗�b���mn
]� *�����lv�d9ѻ[:�Q��>QeS��j�x���zUۨ@a�M@���eYp�q�n�2��b�>D�=���-�*����)�vIk�au�$��uV�/���t�ҫ��MғrT�`��n�����7;l>]6��Ğ����j��IUX8[@S��X5)7V�$I�e3b�7Lk�n'�V�``������������g�9�� �%[9N��k��ڗ��(k�CZ��8)�%Px��+2�Q�&Yx<˵���Y���sU��m��֩�܅Ƭ���f[�c WiS(�`��T�b[���0AD� �лZ]1�=�0�mgIwa�M��"ڍ�,�h��{�t��n��j5�n��g[<hm�S�3��d�()0����w��q��fP�4QM[[),�w\.�m��v�f��X9ܳ�b�C����v9�[r�l��[V��T jL�z���2a6yp]�jS%c8�	g���7ρ�;�1�pP9�v̫*�j�<�]:tG-[��)e��ޣ��l��ʜ�l�*kh�����/[u�V�l 6��g5�$ ����M��$��J��h(��9!U����dBa8��[UT�������P��]�)��k�+���v���'f���1 �i&oY�UuҼ`�-U*�˲�P`(cQ�T�-j:�kҰ6��J+�v�յ!'��^y��Pq��L�y%tc:�z���Ň�36)�s=���[�7f�s4�[���Z�*�F�� 8E\Q0?b*(�'��}�%̘fqͲ�2���3�n̸�h��n����=[���R%>�U3��\�v����[��k�E�����h璋g��j獷]Զzw/l[6Vh��WV��H�3�T���L]����Ξ�.HG��
dЍ|�\Wx��s�i�R��ѯ��=�o8�O��v
�Pb���Ǝ	y8ڶ�
S�2:��W���۬u�ݩN�}���������]�0�vsֆط�ܤW��('�n�`�guƫiT���t���ssO���,K�����Kı;�����Kı/o��ND�,K�{��Ȗ%�b{=��ܷe�fl�M����Kı;�����%�bX����'"X�%��=�s��Kİo}�jr%�bX�������n�J\ݼO"X�%�{}��r%�bX����8�D�,K���"X�%�����'�,K��ge�'2l�K�]&��'"X�%��=�s��Kİo}�jr%�bX��{��yİ?�fD���n�"X�%�N�u�ٴ�˙�d���'�,K�����Ȗ%�bw=�s��Kı/o��ND�,K�{���{��7�����>�j�-R�t]m��m���J�����w���Ԇ�Ä+�����Tf�3I���jr%�bX��{��yı,K��w�,K������%�bX7��59ı,OzM:Y�s.�wwsw8�D�,K�����!�|�W���O"X�ß����%�bX7�����Kı;�����%�bX��3���	Lܗv\���Kı;���q<�bX���ND�,K��{�O"X�%�{}��r%�bX����vn]���.i����%�g�2}߳S�,K��;����%�bX����'"X�%��=�s��Kı?Ol����fl���njr%�bX��{��yı,K��w�,K������%�bX7��59=���oq��>���v+4��a�L	�������rH(�]Uc���87'X�]weٗJ\ݼO"X�%�{}��r%�bX����8�D�,K�����&D�,O��}�O"X�%��g�ٓ�6i&f��wwq9ı,N��{�O!���,��f�"X�%��wﳉ�Kı/o{���bX�%=;�݅�����.�q<�bX��{���bX�'}���<�cSԀA�X��
A�b	+'D�$1��.2$�H�pU� 	���"�8�H�%��n'"X�%��=�s��Kı):u�ۛ�&�%����Kυ ��>�>��<�bX�%����r%�bX����8�D�,K���ND�,KޓN�/]���˻�����Kı/o{���bX�'�_�w�3��%�bX7��ND�,K��{�O"X�%��߿��/,�X,�f�Y��g����b�]cs�]I��*�Ssrذ7Y�z��n�r%�bX����8�D�,K���"X�%��w��O"X�%�g}��r%�bX�~��'vn��[��vnnq<�bX���ND�,K����O"X�%�g}��r%�bX���{�O"X�%����m�]�.l�M����Kı;�{���%�bX�{�wS�,KĽ����yı,���"X�%��ҝ3͆�2�K����Kρ`dL�����Kı/ӽ�8�D�,K��sS�,K
�ȝ����yı,{;|����-^��oq���w����yı,?�g�}��D�,K�w�Ȗ%�bY��ND�,K���=��^�UK���;n�pul����^9��rk�aZ&ى�kv�ۊ�bI�a���Kİo��59ı,N����<�bX�%�����Kı/g��8�D�,K��[ݹ�,�4�-��ND�,K����O!��șĳ��u9ı,K��~�'�,K������Kı=�4��܆nn�Lݻ����Kı,���ND�,K�{�s��Kİo��jr%�bX���vq<�bX�'a�v��$�n˻nn�r%�bX���{�O"X�%�}�sS�,K����oȖ%�bY�{���bX�'�����wvl-�4ݙ��O"X�} �~�59ı,?��w�����ı,K;�۩Ȗ%�b^�}�q<�bX�&(x�A>�~���vn�۳��2����pW��u&.n#F���sd:v�>ݭ�n��b��Y��vq����˫����֎��sX��t��J;�˥�W�p��iܝ�\m�����kE����F��]x��׶���GX�v�yb0�Vڹ@é 6��ܭpͶ���n���n��	�c�A�:��5nNn�wn֒Y���_gn��{u��>ws�����������K��
펶)�;w0�`���=����J&�
n�K�1ɭ��+��������D��oȖ%�bY��ND�,K�{�s��Kİo}�jr%�bX�{=)�3͛.�0�f��'�,Kĳ��u9�c�?ͩ�/�����yı,���jr%�bX����q<�c���ZQ#bn89�f�b<,K�{�s��Kİo}�jr%�bX����q<�bX�%����Ȗ%�bSӾ���.��73%��'�,K�����Ȗ%�bw�{���%�bX=�{u9İ?��3����O"X�%�O��>��ٓ0�乛���bX�'w�O"X�%��w�S�,KĽ����yı,�{����1b<��Տ?90� !A䑰J���z��������2ݴ4賌A���v�.�\�빶˻.�i��%�bX=�{u9ı,K���'�,K�����Ȗ%�bw�{���%�bX��,��a�3v]�wn�"X�%�{=����@]J�{��؜�`߾�59ı,O��>�O"X�%����S�,K����9;�sfY$�K�3s��Kİo��59ı,N��|8�D�,K���S�,KĽ����yı,Og�Sl:l�7v�ɻ����bY� ���}��yı,�~���bX�%����Ȗ%�`���jr%�bX�{=)��&�ra���8�D�,K���S�,K���};߳��%�bX7߾�ND�,K����'�,Kľ���2�7il�&dj�fU0N��h����"�KF�3pl�s:pu�g�X3�k�E������oq�}�q<�bX���sS�,K����Á��!?DȖ%��w�ȟ�TȖ%>?�m���]�ݛ�fnq<�bX���f�"X�%����Ȗ%�`��{u9ı,K���'�,KħK�v�f�i��-��ND�,K���'�,K������K�����"r%��;�O"X�%�{���Kı=�4�2�B�m��˹�q<�bY��! ����r%�bX�����O"X�%�{�sS�,K����É�Kı=�Y�3��%3v]�wn�"X�%�{=����%�bX7��59ı,N��|8�D�,K��n�"X�%���������ՠX���r����X.�n�L�{\\G�U�z�0| +�M6rL�͔�M.����Kİo~�59ı,N��|8�D�,K��n�"X�%�{=����%�bX��l��u�n�ۙ73sS�,K���{���%�bX>�{u9ı,K����Ȗ%�`�{���Kı<�zS��˳2�a��t�yı,�{���bX�%���s��K�THdL�{�٩Ȗ%�b}�~��yı,}��Û�r�\6�w59ĳ�T��3��~�'�,K������Kı;�}��yı>�E|G�
�J���x�>��ϼ�59ı,Jz{�\��-̗7,���yı,��59ı,N���O"X�%�{��"X�%�{?{��yı,O�	���a~�M�`�h�<�mYώ쭰�m���I�X�"��m�M���)�"�iM�9����i�˛���%�bX����É�Kİo{���Kı/g�{�O"X�%�{��"X�%��I��grsm�v]����Kİo{���Kı/g�{�O"X�%�{��"X�%����É�Kı?Ba�3��&ỗf����Kı/g�{�O"X�%�{��"X����>��8�D�,K��٩Ȗ%�by�N���wp�\4�378�D�,K���ND�,K���'�,K�����Ȗ%�b^�}�q<�bX�'����7ٷlۻ���bX�'w��O"X�%�{�sS�,KĽ����yı/�s��5<�D̩�0N> ��*�'��|��72[�n�3������ڸtX�u��:��.7��Le�n�ǰ��a1t�"��sևT�pv�Gmq�ݺ��N��Y+vI�b�康vN8`Ͳ�锤ێn.�a��U�g=�v�nb�guI��k�<k[����Pny7�y{nI���f�pYK��Kf�#( �Ulr��
c���ݞ#�Q)J{9��&�wve2Y$�n�d�}A���@_9���Wiᵳ���:[�s�_F���oY'�M�v�m3Rq�V��Ru�x�Ӭ�ٶŻ7�}2�Ḍ�}��yS"fTș����'�3*dL�9�{��?~��3*dK���oș�2&e�>���˹d7M4ۛ��yS"fTș����'�� V;�6&e��S�*dK�2&{�>���&eL��G;�槞T�jn�ȗ�z��>lۙ�m���'�3*dL�9��f��Tș�2&~�;���Lʙ2�w��O<��3*dK����'�3*dLʘt�{w.l2�i���jy�L�����7�w��'�3*dL�9��f��Tș�2%���7��Lʙ���w��O<��3*dO���\��)6�i�����=��)������2&eL��(�7�����2�Ḍ�}�jy�L��S"g��w8�Or��{��n�/�cþԙ�5��\��ېi�,��8��M`�e�4��%j�����)h��~oq�����]ND�,K�﹩Ȗ%�`�=�59��Ḍ�����2&eL���8rvm��i��s77��Lʙ2�w�槞S��}@�b~�S"g����'�^c<��c����d߳33��]�B�F?��$iLq8�~I%��ԒU�w�HD�����m߾I/Z��D�ٍ�rG�$��_��$#�ɩ$���ߒIz�RI[J$g��ǆIdR?ߒHGu�RI}�y�f}-���I.}����_��$���µ8bM(�$ڞ^�zٍ��im��nxv�H'S��[<o\�x�y<��H�I�$����^�bԒU�����B;���IgR�\MǍdɐI���I/]��I*����$�wY5$�~��}��g�6��F��% Ĝ�ܑjI/�_���$#�ɩt~i�g����,���z	�1!cΆ��T0 �$p��A�^~�]c��y⁈?�K$?K���H �� BBg�FVƑa A�>��!B5�
��@# :1?'���	� �A5Z/�)��P�H�~|� p=W��� ��y�z�o�����J���I.�2�"Ȱ�6�9��$#�ɩ$�����I/l�jI*����$���
E"�/LPnM����{�ym�
�g��۞[m�=���$#�ɩ$���x�X�	$`�i͓U���I�8�F�si�*�)��i�	tc�1�#�S�=��K�lz�J���~I!�MI%_�_�=�&5r�����^�X^`U�u�}m�"�¢�d�����Û�r�nl�e۬����w]`���~n����VDE��"$G&�Wuz��4���{��O�'���J�X�bHE�a`t x�O3g7���z��.m-4�e���$���I��������
���@��z^�L�A��)"M;uiҹέz�K�t�86��+.���H,64�bRI�nI4
�נr:٠Uֽ ��4�������&��]`&�y�BQ	)���� ��x^�zz<��HߋǓ�$�*���Ky�W���-��!g#6�Y2@����٠U�@�u�C�DB�=M�`ܒ�T������^�X�`U-��o0�	�U�#B"��9ٙ�n�M�9�B�oC��"8��=>�j�2HN9�X�y��/�]�d��מ��N�?�k������彬ǭ�[,���SJD��ٰ]�i&{9�lN �vLn�� N��W5���σ�`q��7:��Y�3n��R�w�l�E�����˅�m�K�[�X �ɴÜRV��eAۨc�R1��ƣc�+W�c۝�/V����z^]��]�.�vu����]��͋`:����ݣ��`�κ5/m*�\�gc�v�cN:�?�Ϧ�W�^�{m�^�zyq���2))��M�z��W�
"L��u�:���[� Z��x�<��z�h{����h^�@8�I��P�Ԓh^��6Mn�?k���ID��u��\_c��1�dR=�������٠Uֽ���p��0�����ϖK��f�P�/�'�![��7�S��dQF�XȌPrM�z� ���^�X��9U�.�\f���~���#��
(|��ٗ�}�#��h^�@��&:�FLx�����ˬ�[�
�.�Yy�}��Ƞ���1����٠Uu� |�� ���$��Mu��ͩ�K���t���<�%���ӯ� ��m��}�YW�X�$i��Nf��y�����H1�ُm�i��[K3e���&}=�px�d�� �M�z��=�h{��u��j#	�biɠU�Z�?I�w�9�]`�k�k�B�Tu�����FԊ<�Ǡz��M������yJ�/߇�u���8�R�N��c	�rh[^�~���*�^����㐲*�A��&8�z��w�r�������׀9m�������[@6'��â68ެ�2z<g]neNj����`�Uܐc�gZ�盶��`Um������۬�K�iAy�(<�#�M������*�� ~�w�9m�tDD��r�=d��b�����>_}������ՠ~G�f�gS�T�ŉ0��z�޳Bw��o$�Y���$����
��~T<?Y����q�0�����(ܚ^�X�!DB�(P���_�z{�X�[�6�=����0�F���u��k���[�����ޏS�+++чqJ�b�� ]����(�;�����s�.��������svb�x�x�ܚ^�z�����������
�ɲU�u���1�#�o�M������b\�~�����?w!d�a�x6#�Mحk��>�u� �u�DD$�g��xw����E���������:�u~ ��^ �[�R�ID%}��9n8.��vNV	�l�m=s��L肙��O;0�,:�Qc��m��<�K�I��t�]C�!w����t���kH�cqƍ�[�� .khK���:��wn�w;/+	���w;ks����d��xc�]��n!*u�Ͽ_y맵��Rt��mw��SC�=��Ѹ�ZB�;�+���M�919ܰ����]��l���;v]M���vfi��b ~���,����t�Oxl���u����9�vݜ]�GO�=A��D�+�6웷lt�+ȩZ������ ��� s���"DB���o� ��,�,I��$�z��������w�9��?�
d;�Z��EZ��MU��/����w��D�K� �ߦ����$	"dr=�;��*�� �K�
����ܛx�d�E�eU� ��� �BS���t���=Gu�q`��U&Ԏ<�H�-��v_n�N�=�;tk�+�[4�rJ���x^rFȼpy0rH��u�]k�?#��������b�☆��@�[��I.Y
9�����/����4Ԡ��Hԏ@��hu�ÒJd��^��� �|5u�ƛj$7&�WZ��[4
�נz��4:���"�$�DHN= �[�
����$���[�	�h�zvs�n�.�jfI՗���w5��V��n͆	]g%v�����8~m��n������`y^`U�u�}-��n\W��jGF��=G[7 ��^�{������� �<��wx�n��n�Ĳ/�BPB�IJ��(]�$��~�Հt���;�� ��@�= ���]k�>�[�D(�S��� ��k�UVa���I4�ՠz��hu�@=�f�~�Ԇ�C�1&E�$F)1= �v�iW�7)�:��2�������3�꧘�B!&��=G[4
����٠^}V���qC
�cMā�4
��X����eL�o0���^�Aj�I�� ��x��8rP�B�J����>]��@-J�t1�`������:"'k�V �o� �����
(@�_@�^&>^��o$���|_�ɑ�#�
8�Gu�^����h�U�Tux�2��$��6I͔g�W!ɇFⷴ���f�5��nr�[g���X$<��ɠU�@?^�@�����Y�\���`��Lb�G�Yy�fʘ��z�`zD,��8���H����h�m�^����h�Ay�(8�d��qh'�� s�u�����BS��N �b��׍�8 rM�mz��ȭ���/���O۷�%
"D���Q_�ATW�eTV�"��� ���Ȃ*+�Ђ*+�@
#��(�  �@�( �A`� � �!b� �*!b��P�"����"��� ��� ���TW�A��TW��Q_�EE�A��TW��Q_�����(+$�k0yy�{+�0
 ?��d��-_�                      � ��$"��"��BU
 J��!*�PJ�  T�J�R��� � D
*��B����T)E)I�   ��  � 
 �)J٠[QJD =�h A�R��N�vi�h" 
N� R )@ w�<�   �@��]�>��	{�O�Y{=y=.��T��WַzS���W��Tﳪ�y>�� }�  T� &�>���|�S���g����Ҭ ��q�{�^:ӓӽ�O{ks���Ҿ������ <��A�� ���˥�=;�.�<��� 4�r�{KŇ�'O[�/m� }�@(�P� ����)bޚ����yus��G�� <�=�w�Wu�����C�

n�S��ڜm{����o]��Q�E ���q��l��=>������ y���W_ݼڏ r  PE	   

 �  C�yW3���ν<�J�}�>�u����������0�}x ���z�m{k� �K�i��s対gN�|����94�}}94�q�G�  ��� ( � ����r��w>{����� u�n/w����FO��wy��ox>�G�(��h�: 4����%��h � �%%�D�@��4@ @�'����"R�M��R�� DT���T� �?Q=SoUJT   D��J�2`@��D�*��R*�!����T�Д{T�* �"B�JR��A��t�����k�����������$=���>׵��TW�ATV�� ��aTW�� ���(��� QO�>Hx�����i�������A�&�G�����ɽ~����2����]~g"D�@? E���+��ѣ��o��¢`X�@�8r�'n��5���pn��5�����f��\e��a
b�J`L�e�.t.$�e0 @ѷ�Lt;��lǉ
f�͵�*D�7��p��e8��
�3N˚J�57YM)�k`�A���h�h�3��ݝ�qe���nl�������(���ܝ!po���BlM�(BK������
a�n�?	s��-`�	d�0�b�os��;H���������D4b�*B����?B�	�������k	LYL%����%��S�rIp���)�\��u]�F&�cX`i(B�[�c�0b�HGL��;��o!�(�T D�.~�~4I�.0dH��VR%<A�!�H��D�2C��4C�FD I8�)�n�S��:�h�@�f��X�s}�;M��!~2q�	й�C��%�$�A��-@���&�-a%)BF!!C$�?��@f�g6z���1�/R$I��f���"H2P�ۏ�Oe�0H<�;5�a�wo���M���Ɩ���@,(z5��[�S.�@�˛���o5!7���p��; P�I ��!$�M���+�j��qmf�F�f�\�!\]���I��$	7�Km&���k\vxKCW��[=����8n� ~������8�0ѳK�5�OW�b1���ݒh���}2&�סp��P�oӬ)S�"����X��\A�  <$`\�Q��c#$� X�h�2$	G�sd�%0�;x��hE$�X����v���F��%��@m�\6qB�Z��,��d���B������p�����9B�)�rc�S�ZF�Ca�eqn�kQ�`WbI$h�����P���"XG	!q��$��@�H5�V��; @���p�6� B @ $z/l�$��*CGo�?~�g�94��vk]֝�aC���,{�$!9ן��2db�!\�]���F��n��)
'�6BHN�9����@��M<�}4^�:�]h+ LJ! I�0�Hk\
0$�B1%p<m��ڐ����D)!������d0u�����BId�hp���T�DN	�S���݌i������P��90�P��xE7�$�h@��l���\��HŁ��%�Helّ��G[�Yi��~;@1��&r7��l�Λ3�bсX���x�G\4�&�"@2���q�]6^!��F�JVYH�6B�a����!7nj��a$A��vl����t�?Z3{%B�l��l�+�,��d(A�I����E�@d
��p�2��F���0�U��06R��
`h0�$,��K��%��	L4oZ���~�$����3�D)�!L��fj��!���k��@�M��5;�dc
R�$�v~9o��#Y+����
�{tѸ^���_ߎ{�_�׭V�nOXS���������;���)�ڇM&&�Ė���!	�ѨĪ1`B�(�09��V�k��4nFA��to��SF�E prq�i�	WD@�(����\�;�60!!Ҏ����2�'�!Y`B��Z�RVɆ�|�,�i�rk0��e��I)
��R
nh��!�7�8����g����"Gl���HO�$?q;X��a �l�	��� ��A��d�Gj25�B���JL]������L�m�`H�p�"P�Xd8�s�Ht)�R�B��a���c��d`�VB�1��U�Q��e�X�a�h�!,Kd�e�Ʊ8��nh�,��d5���-��֒�!��No-�`���l���m���Y ��	8�s��6���s�a7������	)�alp"0b�4H������5�*^<v��6�2,���+$���st����w��l��ʤ
1��7��+�`r4#
< �[���k7�T"'���r��3��O  AcE���A��CD��"�DX�BHRa���%���/�<+�ݶILX�	Hi�<P����:vS��#�����C"CN��,y����I$�h�f�;�����hHG �ԛT0���8��D�L�jG"W�1�$�\�,�mu�CKa&�&I!���(U"� �)�o�0����Ƥ��NLX�i,��(a#�"B,�o��p4��RR����bC��v��0)���F�2�ԫ"�S��ò=����!�bB2&�@��Hp	RB�CP#�����w�{0�8�C%	��c$�6���	�"�doz���f�C �Ll%�L-r2�XD�+
�p1tC���j-�5����`C5iL�2���
=Ѕ1��7L�/'��~�8]j[-v���Y�F�F��5��8��$9��	q�i!R5%!�L����$(�V�a&�3&�'T����� �
��=��l�[��K!�;*IX��.����J�7���9_�	�H0\-�$�]-lR��jB,�X�Ըpc�X�������x��`�9ǟ��S�Y�ADd$$Cg��gh�HH�p07z�W��Y��ɷA#��\��N@+��m�	9$�r2R K,�B���:HE�$]�
��L��40�Brl��(qۙ$ٶn]]X$v��֎9�2�����Ԙ�Ȱ!!Z��j��P̚6�!�Cp�0��	c�!2edV[�L[5u�#.�g7���tF��f���e��$1�$'���##u.MZ��&P-�R
� ���E�1��XHH� � H2&:z*c��n�H�H�	 ���1I0���BP�f�H2Ʉ$H�tD��`�I˸C7!-�j�Khc�l�3T�K&�@�%̅�	7!D��l��$�,b��H1�A��2ۦĔl�ݦk$��I	�!���@$RY1�ik�kP*M��	!�G[�3v��!H�h��VLXSR1a$$1���A�������21 @,��Qq�-S�Q�� @"S���z�� �u�m*Snl�ԛ��LhmӰ6A�.��c2�[Y�����[C2�A��Z��a!��{�r�kd��)�(l:@�u�CD67ґ�(\[$a �(����Hh�f�k�O�AȐ �d���OР`MN�$�w{�k���!��aa�Yׁ��/�HƤ
������@��!�ez��q�;�w#�����	�DvV�����6s�������Z�a���F0,3d?B�t^n�'{>��9���\�QT�H�@��V���$�f��0a� E#0)�Tp"�1�łp�a�7���=		��� fKJn�
R� �2 Ѡh��\�� +��R�ں� ���;�������OH���!��0))��E���!�9&����P��k���ra�O�bD8g@�ġ �f�$Ѩv���\U�602�*Jf�~�@��#L�찍C@�Hl��401Ӳ�0��V��SA ��l,o���Ԅ�P�(h����~���ٷ %H:B4��M��)aG`RF��n����jXK,��?o���Mj�4��B�p&��J`a���I$�4?!5�@�3��}�?J�( ��      ��}�sm�  %�]�m��mF4�6ݭ� �N$mK\�uT82*��US��[]U[�	��\�I�A���5Hl��ڶ��l:sSa�Xi�kV�H8��`׫8i�kpq���V�mXI��[@ְ+n�m�*���u����j�n��V�F��S���R�;'mC��(f큶�k�.�� kXD�6 ����Cm���ۛV�$kխ���h���2�\�UJN�v�^�\:��AK�Y%RX*�j
�M�Ryz�Nk&��n�gm���R�5�)'e]#@=v�h��oX]�=mt  ��i�-�m��$l�m*}�E�ڕV��T��<�lr���H���4V�h sl۶�X׍��r��R�N4�UJ��Zv�lͱ�V�N&`4�(se(��P"�غ�A����~9�f� ` 	��   �v݉�e�`m��e�NҤ\�ʶ�B��e%�>�)jS 'l�G[հ� m�r�	 X H  �.�W(pM�m�l�}��f݃���zkiV�b���q۔*�ؔ�� ����j�׭���m��������mm� p�M�!5Vꚻ�Ȁ�vaV�F�8%^���oF�Z���+�g�y���[4��*E�ٶ *��ƶW���,*��U�e�x����U���R�V��v4��UW �����J4ïf��Z��kl��n�n���ղ��H[JP
���v� �.����UV�v�U�i(��n��6,�q�&ۛFXA�rF���%[�Z�I���u��[� 6�`�kfـX�`N�Ֆ5�m�
[V�-�!�܍���c%��L�*QKs��liL�]��| :�c���.�%�&��]t��mm��N���l�ۂ�km-��m�x�-�v*���eV�M`YW(�ʣ���	��ZtTt�ki�$l5��h  ��җ[yi�U��N۱��m��خ�y��5lt�5@l��n���.v�j�i�8���	���T֚ge���
dv�)�YVBh M��1�LM��lQ�:e��X5�G�� Ӎ��m�;-�Wh�@-���m��$����]��M�뇊Uv�-q��l6�ަ���֨`s�EU�Cv��6�n׭�' �ku��}���{) ���so�ī�C�� U�MUQ��wUp\�9)	$�٫�M�v�[���� 6�H��p6�7l��m�`   n�L�e��0�O���^��j��`ڢ�S[��E�m�!��VJ��I�`h׫lk��lN�:Y2@>�Tjj�m���PJd٠&ʯYyUz��8����� A�*��[l�ǝ�F�Ҭ�P*�^ 8ڃc@�խabiA�h�$E�mˈ��N�[�����yI�h·�e�v�����.�t��7` �]�UT�[,����-�m��^��֯eM�m��Í�`7jZ ��M�o���c��8'GdݫIjk:��0t� ڦ� �H�e��҅�U�##V�#٩P��a���Ӣ���
���T�c�UUJ	+U@]'PV�J�غ��kT�l��ʧ��s�������uUvSP�n9!��J655U&��ϯ����K�}�a= [z�2�;H����NpX3�S�܁sj�;�6�I� �@ ��!!#mzt�V��U�!    �-��m{)gk�Ԝ��D�] ��HZ�"۶�X�����U��q��ҼZl#�:7P�Z�eZ�@.\M&�m��~��m��cGo/S�u��m��s��:Ku�� og��Ӥ�̀  6CmҮ4����mm�)n���m���bI[l �lR�m[\m-��m9:�v�"rm���Q{�,:�#��F�T�d��h��mmT��R��V�	l�8�  $� � 6�ݵ�qλf[A�襷�t�J�,�܋ڮ-Oj� 6�6�;]�6��-�z�l [5�5� �]��m��طe�  <N�N�mh��6 jT��/2��K�0�am 7o�[I�-T�Ht�ɖ�5�0    q��Ç�lNqm-��>}o}��nj�m�� &ٗ�����W[%kX-�-��l��ݴ�m��H�m�m� 6�h[��4���4��S��7^�9�ͳl	 /In� j��� ���5��Kh�m��������f��W� 翍|W�]*���CU*�<cc2����UR�R��kҫWL�q�8/��m�d4�i/l�  ����e1U��V.©m��R8�`�a�ש�H�uyj;*?�_*��N��`����}�g���yN�-�޹��5�R�ŕ)�&�&���� kgD�%Y��m�L�ڰ  m&�m l�f� -�[S���a��۲i�b�t$8��̴�V�Q�C`tN����V[�ܣR�� pzGHu�.�5�d�l���UK��*�P �J�h���Jۂ�)Z��/��@�T�ɰ�>�nN�U�Ӥ�� ����a&�-6H�am6�����Hmm��l ��� mH���J�l�@m�  �J*��pU[@[=��@6�6��� ��۶������xR�\� �+T�gM�M�`�k���&�҂��8��z�6��   ��*`ݶ      H$�[��[rl sm�e�ݰ�[%$6�  ��v���H/��5 �g`
�+��T���v�R����U+��bUq���JL��S�+_�ϘĮ�7;/g�^�)ض N)VV��D�t�9h6�!��[d  e�-�  m��X$�4]�lt�m�
�*�UT  U�V��6�k��V��H2�lm�� S���� �Knn�Hmf��j���35�����M�r�5 ��j �Z� �hs{n�m�6�d���
V�0��l   i�l��k2��`A�h��͎p m�&���u[�i2� �ZKj�	��87 A� ����pN� �mm	 ����2@:�q�H��R��`s�T��I6KY4RBCm�  $Y�&�h����
%�<�PS�4�� �m�`m�8   �[tP�m�M�Z.� ����2�.ؐ*m�	��m���%�m1u�h��qm    �ֶ�nF�k�����kn�a��H)m�m����čۢ]��U�)��V��
�U*�D����p�U\�UI9�պE� ��έ���V�@[C� ������>   -�m�m-�!��͵�� m�   �� �[@q,��a4����e�ʬ1
d�aƪ����n�%���0�    �n��a�n�f���
PM+*�ɐum�)���Vm�?>���ru��k\��WN�l���g��[e�k  ��$S�p�� 	�6�m�    6�+@��e��TB����>u�Ui1j�P�#�r�u�i8�ֶ��|  �n�    f� KF��Ύ�b�톀��͆9ݮ����ə�䶶�L�U/� �2�͠
��jBjt�n�F�i� �   p89��qU��h��S��
�m�V2-�v%[lVW�lӀ�V1YݹV�BL��l�� �գ�Tq�{��|��csTJ�����)t����IrJ��+��*�M�pUUW*��ȝ.٫	w@��KZU�ps9�]9۶1r�PA5t�:S��qmM�2 �ܣJ���y��9�YZ���Yʨ� �5+U][���-�RsI[Q����;kZ�!cijڨ8UU���$m�Hm��   HZ���z��!Sm�o��m>k)�	B�q��UR�VԄ�ՠ  .��ړ]�ݪ� vĖ� �Oda:H u�\���5��u���N6`�\�T��¹%�5�9a��Ud�F�$    �8�+CKm������:-��4]���kn�d  UUJ�Dщr;&�᪪���eeZ����upVƂUm�@���yu�l;��vM��8"�p���Ӷ�m8�Ĵ^�3JT� ְn�  �ڜm��H�lH��Q��y�z�ڀ]��m� qV��F�ͻkdim ����(���B�q�.X\�#"m6ҽ������: ���t��H �sl[F۰��;n�M�� ��P�(�pU]l��ڶ$� �l���b۶�	e�t]d�Z�WUR�3\rD�R����$:�t�j��ZL ��lH�V�ͱV��+�@j��8���
j*�v����5 !f��l��Exݕt둖ꪀ�g����Q�8���UUW����������ʇ�H�"�����*���?�
#�
C�
����S�"S`�#�J��E�)�H�V$E�"- . A
)+������BH0!$��0"H  �bB0H��@"��FFBE �#@`��
��X�bH,$T�� D",a B��! Y �E�`C��Q6���&�?�|��Gʪ�M��8���Ѐ�Gc�4���z!��Ӣ�v(�[��)�B�D(�������A��.D�S�+�NT0P?^p���@*��^PV�"i��H�Hʉ�P_�uU1�<�M+���D"���P� �y�8��A�O��| �ʉ�v����Q?�@)� �t�������P����LH��:(� ���U��E<"��F�\�,�!��D�� �D4��~@ |b �� R�	�������q�Ev�o�C�H/�28ج&d�gĖ�8*:����Ƅ^UӶۨか��Kt�=n�$�ZEc����K���;^��a���&���'e��	q��� ��I���֋/���l�=$b��V3f�q�S��=+��W^6�m�YP�7ێ{u�x.���ۀ���ms���m��V���[����\���԰n�8k��8q����;���Z]���x�Ʀ�z-!geݕ{�m��ۧq�V H�7n�kl(9�Y���A�&�md����\M:	�G�>�����AN�I��e8-�x	&�:θ��ñ����.�a���ҩ���-��V�g�^�hs����U����ˊ6]=Tgv�y� �)�];/t��cYb���ucp���[t��OkE�GL,ev��)��d9��l9�/(e��.n^�i�G5�<r�����6�B��ݳ1�X�vN�J������Z��{GK\���5d"i�:��N5l��Y8��
+�I�7n��Y�W,��\�D�r�v��=�ku�G�0���Z�k�ݡt�& ��5��'@�D���-$q�'@�,i�i�C�u� PPFW[.�]|즩Yy����ڀwc�4���r9yc���n:;^�<�U��`�Wd)5�{g+�{-8��gf�̭ͽ]Z�j�b�
G�]���`4�F+������k�h`+i��E�b:%kL�	�hvMQ۩]����sӎ�52��q�j��34����j����M�ʆ5!�=�[$���u���i2��p�dre`�H�6�f��p�knNC��!�m�*�=��˃�����h�g��ƭ]Fvn^z���Fݐ�<K�j���/8�v�R��9��Vi�n-R���S:rP�F*7b,��v�.os5Y��hK��;:�Re:i��q��y�6ڎq=݇mGANۡ�\����g#NQ�7F359+ O�!��m�V�Y&���*�cJ[�ӛ����*n���z�?��z���B; 6*�8 ���v�٭Ir�F�VzlOn���N�`�c)	Ą���v��7���� �V��ѣU�!��G\i7"l��J�q���۰�A���5l�]-Ż1M(X�{N4���Zsڳ��h�y�펊6�4$�A���V7m��7k��
u���v�U+َ��Cg��[s��k[vb��fkD=X�Js�kg��p�׮�.r�<6��}�݇c�9^8\!�&���=�ݷls�on2��q�1�˹r�v��B����CPN�=�$A���j	 ��;�m=ı,Owٸ��c���~~��o�D��J>{�7��,K��]&����T��j%�s�}��"X�%������Kı;�w��������ow���tI��f�D�Kı/}�kiȖ%�b{����Kı;�{�iȖ%�b{;�;��{��7�������MP%����"X�%���7q,K���]�"X�%��ﵑ7İ: �"f{��ӑ,KĽ���kVjf�fhչ��D�Kı;�{�ӑ,K��w�ț�bX�%��m9ı,Owٸ��bX�'������I�˘\p\qp�7e�����m=��zAE�E��6�M���7B˝U���~Ou��=�x�w�ț�bX�%��m9ı,Owٸ��bX�'}�p�r%�bX�_����հ�<�;��{��7����{��r
gV����'���D�Kı=����Kı=���&�X�%��{g��fM]\�2̙��ӑ,K��}�"n%�bX����iȖ%�b{;�dMı,K������bX�'��n�$�kY�S32�Z"n%�bX����iȖ%�b{;�dMı,K������bX�'���q,��oq�����z���|�~oq�ı=���&�X�%�T9}�kiȖ%�b{�ޤMı,K���m9ı,OvI���jۚ��l�D�vU���i�2[b�V8�-��Y�6�bI�GW���]e՚5�2�&kYq,KĽ����"X�%���z�7ı,N����Kı=���&�X�%����jE5@��j�����7���{����m�q,K���ND�,K��k"n%�bX������NTȖ%���֥-�qr����oq���{���iȖ%�b{;�dMı�n
E@�QS� x�Ț�u�{[ND�,K���"n%�bX���y�=�q��������ow���&�X�%�{�{[ND�,K���"n%�bX����iȖ%�b{=��Ԁ,��;��{��7������kiȖ%�b{�ޤMı,K���m9ı,g}t��bX�'�}���p��5 nm`qէ�R+�;x�X�'�m�9��*�Ҝ�������˶�2��2fk\O�,K���oR&�X�%��{�6��bX����Mı,K������bX�'��n�$�kY�S32�5"n%�bX����iȖ%�`�;��Kı/{�kiȖ%�b{�ޤMı,K󾙖x֮�ɢ�ֳ5�iȖ%�`�;��Kı/{�kiȖ<THdL���z�7ı,N���m9ı,Oz��j�.�֦�˖ۚ�Mı,K������bX�'���D�Kı?{���K���+��҃eZދ.��E�.�u��LCh�Ě�\ֵ�m9ı,Ow�ԉ��%�b~���iȖ%�`�;��Kı/{�kiȖ%�b|N����I.�kY��QginvE΂:�$��u�E��n��<b�/;w�www.O���CE��=ߢ{�K�����Kİ}���n%�bX������T��dK���|��|��{��7�����^���ie�3Fӑ,K��w�I��%�b^���ӑ,K��}�H��bX�'�{�6��bX�%���j��e�2�	�֮�q,KĽ�}��"X�%���z�7ı,N{���Kİ}���n%�bX��{NL�4]2̗Z�ӑ,K8�@Ȟ﹩q,K������Kİ}���n%�bX��ﵴ�Kı?N�w#3Z��.L�u��7ı,N{���Kİ����IȖ%�b_{�kiȖ%�b{�ޤMı,K�m9h_��Y��C����SgٶS:ٍ�f��SYR&[�cX9��Μd�{9y����,�����X�Yݎڛm����ݱ�ے㱫�Nnݮ��#�2TU�R[/4^su�$�1xP�/d�rNDi�: ��tP��rꇀH��[��qal��Ņ�m�s�+�B�{�����Q�<d���F;��x�����n6��r�xݙyL����Dc�Heܗ/Iv8����ݧsM�#����vA�W;e�^]�a�.SF�u3%�u�fkGS�,K��}��n%�bX��ﵴ�Kı=�oR�'"dK���{�ӑ,K�����I�g�a���{��7�������bX�'���D�Kı9�{�ӑ,K��w�I��%�bw?{�2��:�5�������ow�߿-q,K���ND�,K��]&�X�%�{��[ND�,K��MȘ�B5M�����oq�ߟ~���"X�%��ﮓq,KĽ�}��"X�dOw�ԉ��%�b{��~�S����%���{��7���}t��bX�%�{�m9ı,Ow�ԉ��%�bs���"X�%��g�l^�����&����v[�3��W���T�սRs�i�*sl)s��������5�]'"X�%�}�}��"X�%���z�7ı,N{���g��E\}]it��]"���-������Z�ӑ,K��}�H���Ө8�&�X�����Kİ~�}t��bX�%�{�m9��2%��{ۙ��frf[�ԉ��%�b~���m9ı,g}t��bX�%�{�m9ı,Ow�ԉ��%�b_��̳Ƶu�&��֮f�ӑ,K��w�I��%�b^��ٴ�Kı=�oR&�X�%��{~�ND�,K޺��ˬˣZ�\��WI��%�b^��ٴ�Kİ��}�sR'"X�%������Kı;=�LMı,K���؛�����]<��錶��;v��i��]i]@cI���M�6�K�2�f�9ı,N��ԉ��%�bs���ӑ,K����17ı,K���>{�7���{���~�w�SN-�iq,K���]�!�$r&D�=>��q,Kľ��ٴ�Kĳ�u��i����:ί$�Y!#RkV�Z��r%�bX��צ&�X�%�{;�fӑ,~@R*���	�D�M}��"n%�bX�����ND��7���~�s]=�'٬��oq��K�w�ͧ"X�%��{z�7ı,N{^��r%�bX��צ&�X�%���g��̓Eђa�]k6��bX�'}��D�Kı9�{�iȖ%�bv{^���bX�%��}�ND��{���'Ӎ��i�C�V��@׃��3v�n��7e�)zٻIG8��OG}�wwϟ3��k3�fe�jD�Kı?~׽v��bX�'g�鉸�%�b^��ٴ�Kı;�oR&�X�%�t�fO��\��5�e�]�"X�%���zbn%�bX����m9ı,N��ԉ��%�bs���ӑ>ʙ��z�]e�ѭMYf˚���bX�%���ͧ"X�%��{z�7ı,N{^��r%�bX>��4��bX�'s���3,֍S5��fjfk6��bY�����}��H��bX�'k�ӑ,K�����K��mb@�"D^ #�wț����ND�,K��M�]1��j�Uv�|��{��7�������Ȗ%�`����n%�bX����m9ı,O{ٲ&�X�%���|~3�^�ɓ59�V���-��
R�m��=��j<7��Nucp��#`�/�9ı,{^�Mı,K�w�ͧ"X�%��{6D�Kı9�{�o~oq����~���ѭ�k�Q�n%�bX����m9�? )]D�K�͑7ı,N���]�"X�%��kڱ7ı,Nw�=�&d�.����Y��Kı=�fț�bX�'=�z�9ı,N�^Չ��%�b^��ٴ�Kı==��!3Z��)��u�7ı,N{^��r%�bX����q,KĽ��iȖ%��&D｜"n%�bX��;���Qe.z�c��{��7���߷��7ı,K���6��bX�'}��q,K���]�"X�%��@?����>��ޕ�v�u�'f�7gJu%�츥�O&�S��.����2����g��ԖV��ƭ�,W/1�B���xk@���kKҲ \l2�E�=u��.z�bMմtn�q<Y�X���s�����L�+v�av����k&V���N^a� q;d��e��ݭ�[/On��]�=Nvgb���T��9h-Es����̐�KU�r��;�w��Vό�'�#v���d��Rk���Ƅ��4'M�lC���*	�z�����KĿ���ٴ�Kı;�fț�bX�'=�z�9ı,N�^Չ��{��7���}�M]�Ke�����,K��l���%�bs���ӑ,K���X��bX�%��}�NG�=���'���{���_�R�P��ڭh���%�b~��z�9ı,N�^Չ��?�(C"dK��}�ND�,K�}�"n%�bX����kY)�Է5��u�j�9ı,N�^Չ��%�b^���m9ı,N�ٲ&�X�%��k��ND�,K���2�k)s.kNkZ�7ı,K���ͧ"X�%��G�}�"r%�bX��׾�ND�,K�׵bn%�bX���9�����f���'c\��)�X㛈�"jN^���ԉ��w��ww8z�����g��Y��Kı;�fț�bX�'=�z�9ı,N�^Չ��%�b^��ٴ�Kı=����f�s�.dִD�Kı9�{�iȧ��#���bw���Mı,K�{�ͧ"X�%��{6D�Kı/����Z�˓Fֲ�ӑ,K���X��bX�%��}�ND��0ș��l���%�b~���m9ı,OOk�"QG2B!
D~�?b?b1.;��5YP�[�k�p|�fe��v��y���=�ݵ�K������"�G"��=]I��K�	�̢������́��	n����$�46�q5g��s�\+$$n<�I�I� ��Ɓ�ڴ���g�߳Pu�s@���$�L�i��fb�=Ϲl����"�:I��Z�Z�u�B m�?9"�*��ܓ���nu��|�Pi�P�b5	�I"b�%�!H�`�!B2���1 E�F,B$ �H�	  B+�ӛC}�C�"�H@ �aF0b@��1E�A�|2��:�����"td�0�Ieb�bcE�#0p���21� E @dHA�`B��bH;ģ0 I�CX���$@$"�E��	a	1 ��D"����#HI"@ B�� �#���I��	$dd�D�$�$1aT�		�$�X��"Ab0�@��D�)�VFB,H$b�#"`$��E�$� B 	��	14�ā��4	 �ă�+H����
B0ciBP��E#��A�R21 1I�U@M�3@�
D�(�P��+��C�x���6�? hC�@JxUy9�?v����'�{_M�m����he6VSI����Wwv��?V�$�>P^Y?{�}78� gٓ����(y��j�r�����$��wWI�2~���J(H�wM�wu_�}u~��"����Q��k+[iN����c	�S��ћ���n!vW7��]uP����ު�H����Tp�~��kIV��!����OM��,X�X�5��E	ʪ�H�t���]URRL����!*��u]]��46��0x�cOš�����?]U�ԓa��%�U]�$Z��j�X�^'�	�-P�{��'�}���F���k�'S��}��E<���@6�_UUu�Z��}[�UUU$}�f&'�<��kV�5��'_��NI<�}��_�N �~���?~�l� ��pJ8F�!�E��.�76��Kq��u�&�����Z�����Kؒ"pfI���Hm�ى|}��?]�{�~��H�ZJ����d4�p�2�h�2L>P�Mn�I�{훟"ե#�h�2�� �-�wUT��b���&�i�feh9˻��H��E�U�%�uWWQ�"�wd6UUU�A����)��cf4�h����d��BE����K���E.��� ��"��,O)fb��WWt���@�섪����G"��Uut��tZ�� D����ԥ̗8M3R,/���.����{[;cC��2���.�p����Ye�7Yg�g�%�y�N$��D���'QAȇ��e킸�]tț��;gT�1p��-c���(Skƶ��y��ATF�����mp=��ۮ�|]ڹr;j���J0�g��cO`���qmv�Y��z� [�O\�s���V�zL���d�s<�k��U���w~�����v5��M�cOi^9�㦫;6t4I�͛v�q+����,�;=ؒ5v���f���U]]������#�K������>���#����xH�wCLX�^'�	љ��Uui9��E*��� �-�WUk����:�lM�<�o0Y��e�]RG�}�$R����d4?]])2E�.���R��x��e]]$E	��섫���G"�˻��WO�oE�{�*e2�FSI��ЗT�ݰ�$r)u��}�$S�]���Y�bǙO���ߋ�QRI�݅э� �����`�P���c�ݧt�6�x~�����@����%>�h���=�m�$JL���s��]�E�� �P"�"@X�D�����';�}7$���[3?bE�ʲ%NA��hN-�K�@����%ZR9��E�ys�D�H�J1�E�w�)�Z�Z��ZT�h�SH���N4&Iqn���[�o�� �Ѻ]����8�v����n�D7,��y����.�u�;���c����ꞥ�����;���5�h� �oR �� :��2HLX�ra$�@�����M�j�<���<�e�l�)�^Y���z�ŸNUQU[ˮ9^bP](����{�ܓ��޻�w�=f#�x�6��߳����v�����Z���4�s�e�nF%��<Z�~�J����"�{��ՠ\�؇[o"�1FD,�yv+��vf{i������Jn�Y�Cp]d�c��9SМZT�h�Jh�M�������6a�D�m�h��M�W9Uv8� 9��E����Q�ND6G�j�<���*��@�zS@��W�6&�<�(���� ��n �-�7�ʁ���W*�U�ܙ"������)SM��Š6�p�9UU�؟ ��9��߿�{�	�b%8��ܬd����`WkG6��ݽO[a�Ǟn���1]n]/^Y���z�Ÿ�kp�n�;f#�x�4Ƥ��Z�Z��ZT�h�]� ����rE������n���[�y�Ur���ʀ_]�@�u��QIS�	ŠUE��YPŸ�kp�W;�Em�h�]��j�<���*��@���:�RI�K�Ɉ}�⬎Ջ��6n�O���W2�p�<L���Nv"��=^���͡�v׊^Wn�W7��ǝ��I%ӊ�$�H�KWq�#�Bdf�n.nY�$z89�8��Ј0<nqY�s�jv�Zm�^9M�۝\�����*���ts^�cR����Mې�jꎙ���Y�9`h�Ķⱓ��h������F�!u`a�%�3Z�J\�e��rp�ߞ�nݢq[s:����J��q;�YbTIk��N�4���yí�U��}�>�ܓ����I���_�4�'�/_�4��F��ǒH�NH������}���� ��0�!1cM�IzT�h���-v����+U�l�F0X�Z�* �� ��n�UW*��n�;f#"bx��f�k�hW�hRՠw�w4<�M��I�d�X����nj�'���<;un:��yyH�ӱ{&7��L�)#�ԑ���YM�Z�{��k�hμ�)#jc�M\�ܓ��޻��τ;����f~�Z��Z�vq������w�O��Q�BE�{�w4]�@󬦁U-Z��4�8����iI$����z��n�Us���_�f����#bR<�Lm'$Z�e4�n��Tqn x�ze]8\k]6�gE
e�38+�z4y�n4[q�їwV��-���w��|��m�Qm���m��-�=�ʀ.-�>ש ����x���J�CŠ{ݵ���$r-����*��@��l�aI��X�;ڀ.-�>ש�\��W*���m:ށ�u��}�m�$JF�NI�B~�s���� o��۬���w+����&�!�#��U:����k�:�h��ߒ�dx�
H,x�����'����n�9�.��٧N�PH62�W�'�9�iqh�]���hu��*�U�y�SH�X7M.��� ����+����z��kpo]��|�#bN27�rE�y�R �kpn���� ��+�t6��G�uZ�Қ���Ǡ�6ɍ���� ~�����{���~�q"bi,M-��M�?~̣�:�hS��<V�@��}sv��/cf�零�b��nݓv�b31sn�j랉��I��8�Ƙ�p�-�Mβ�T�{�4�s�e�rHE���4���e�]$E�@�vC@��4�^U$j"`5�8hS�h��q�������n>�h�2�����ō�K#H��@��S@��4:�hS��=�����A��RGޔ�<�)�UN�@��Sd�<��A4��H�A�IB2	��$��.��4��BVP��cϷ1885�Cd	BFA!I��Eq Os����?���SmO����u_�|_�<q�,�A#"�"�H����"2$H� N �$�u�;M�RA�H�bF5�&�ZI!�B"Đ5��"�n4���#�E�@) �u"��t�� ��K"k���K�#�h��4@��_g8�,��;���f�ֵ�[%��MYT�r�NI�<��
�N��4s�3���F�>7O�~:C�p�2��֮%F7l��Lڥ{1���qf٠��'5���p۞mR=��4�%��6���e����퍀�3�ḯ�\9:z�3Q 2�Ү���nUV��g[�K�8�av���¨��p��bŒ��d�k/3�l;-��:[�:�&�r�ݫC91�(V8:�{*��gݼ�\n*��J��v��3GfJ�6�Y��/<�9���T�Ү)��Սe��Hu��[l��/ �Vݻ+�v��ъ��D��G|y����њ�5p�K5V�}|��v>o��󭵅��n��N1��ݺ�>^��=�9��`��l�V(}Q���4Z�t�cJFtr]�]���]��1�/�ѭlC�<�NT@��X\+T���g9v��H:�g����uq�%�l�P��ȷ:kmI��H$�V�`�k��d��Ӆ�ix	��nE��V�!��:B�}��t�����@l9�k�c�{+惰�;p���kh�RlJϬUъN�#vͺfE��4�r�$����R�,�n��[Z7e��v���^i�U�ڇ,�}�(2GV(���m;�+Ź[��tW�v��n��Ƽ���!^�V2��h���k�3'��U@hTѴ���E,h̶�b��v	��v4����	S�b�gf� ������ԛdk�rī<;�Y�6�.%YYIj�ٚ:UU�ڎ8����f#RK�9�m\�Ȗ�{vZܼ2���U�k	l�U �lո԰�82�fw���r=�c��]�v�b�ܶ�8��ݨɸ�����^��	�lOAJm<��� �!��$�W	����G�U�ٲ�MSF*l uQ�;F�6z!�������\�ҫ\��Z nb�FƗ2P[m6��S�Q=[�ݢ���Ō�p�n�+Y�,��#�6z��X+��Bm�j%�t���X"r��*0 �D;0Т6:T���O �?�s��k�z�7W	ۛШ��A�x���A�+�[];3�ӷv�sܜ'�#u����tl�;�	�ki�{L�V��չ��ݚ�Wz�]�����|�Z�:ⓛll6��MYI���	�`43��v4�Y�k�WqstQ=v�ɘ��Fݙ�j@<q�x�����2d�V�@��}��s��4t���%��F�N��nݺ�"�ӿ:��.>H��n��Վ�6
�6�݅�]���=p�u.Gk���[�ng*���9�I$��E@��ύ�Z�{�4l��u]Fdn�ӓ�� �-��r�˳۽H� �^�@�Z�2Ă3����=��;�8��K�L��$Z�>�Q�&�i�G�)�yl��U-Zw]� ����rD��Ip�<�R���W�n����H�޹���:�"�ٹ^!13������o�vR�d�ksۙ@��=�*x��L@E��� 
� /R o��`�ŎA,�AŠwt���߷����! ��F��I ��T(��|!�?~��}�ܓ��_T�o߿~H�ߌ�F2	Ȅ5#xh9���8��wWT�&w-��q�{ϕ$lRD��)$Z��h��Z���BU)&�@:.�+31$4��D�UKV��Қ�S@��M˖��)�AĔ��Ț�l�ƹ+�z�%�N*_@�8ny{Wc��m�Y S�X�ZwJh�M�e;3?g�T�V��;f#��'�1�� W� �^��[�{w�?Us�9�a�>m��"nE0�H�4��V{�s���|�B�� ����~�����@��g1�Y�fQ�bxhJ�ReH�wd4�ܴ=R���� ;��Rb�&	L�Z�� �g��r���~�|h��h�\X\Y��F8+g�]bn�x	n�Zä�'%&.�v�3��&6�2B1�ND!���m��<�)�Z�ՠ{�)�{ϕ$li�$Q�&�4:�hRՠ{�)�Z�Zj�Cib�r`I�Z���Cj�U˷1n��Hַ�Pn$��&���t��k�huצ����F׷��]�;���XMa�ؘ�p�-���e4
�j�=��/Q#��3#s,������J�]5��ۑ��͍��q<���=��\ާ�uԛ�0�H�<����*��@��S�f~��vS@�W�QI"&Oɑ8@E��z�Ÿ�� �Zl����AŠ{�)�Z�ZWj�*��@;�222E�����:@�/R �-�7w� ��T���0�G ��h[)�vg��,[�n�* �� +�ʯ�*��U��{�����9=:C��qT�aA0����vWk����y9�+�Imt�8��>��Ǯ�msΫ���v!�N���8��g���)6���k��p�8�.l�,�8�Y�v^셻fʘ8��٥m�8����/�\c���8kTv�vΜ�ku�a-��9�ۮ7DH5������l�m�l�ٓԖ�=8�
��]�[dG������x"� �+k�2[\�ul�Kq��J6���{7��%�d����8r�h����?��{8�;�r�� ��!�)�A8 �ı48���-v��e4
�j�<�l�aM�lLJ8@�/R��]���wz��s�e�rFE$iŠyl��U-ZwJh�V������ĦOɇs��[�n�R �� �z�6�ߦ��ۓ&��W/].4�e�3;l#��(˹���A�ۑ��=,���1��h�)�Z���e;?g��L���d�c2'�r'3@��Z�#�e4
�j�;�S~Ď���s	r	����O��uZ.��_U�Z��A�b�C@m5����n�� q��5,�M��3WrN��ٹ'ʪ�B�~�L��ˏr�<��Вh��^9[��_9�����i�+�x��m۵�J=�m��	�-����1�n�bbc��E�yl��U-Z.���xm$M�$�5"�<�S�>_�Uo�@��Z{�f&��ĦOɄp�*�U�N��ٹ���T� �&����'}�|h�jM�H�ȒɄ$Z.���ܴ��Ƅ��$Z��
�#1��$c�8�]�@��M�Z�]�����7?6�Ą�r�;M�ٳq�v뎎t'+VQ`�)n5\���:����B98��<�S@����uz�ՠuy�fF�,m�LMH@E��U]�{�@b���@<�����S�X�Z.��]�@��M�Z�9�1FF�6,i,ǡ*���I�-�L��ˎ��@�������nI=��g�k3k	$�8�-��;�V�V�˺��j�/.�cm�������Q�"b�n���n{�P��-n���4�A5�E2̏�@����uz�ՠyl��w���5#"K&�h���.-�>^��[�o�R̾�X	�O<zs�Z�vq������h����T��I�7 )Z��� o��׺�qn�V�271cn'9�Z�Wuzs�Z�vq�m]U��%+�O|�t�#k�f�؍К��v6�dݴ��Q㈄�p�-�zy#��kl�k���3'�dh͵�!���v����mnM�m��=�EѫmM��tt2����t��e]�ǷE�s��N�d<�ڮ���0�]`����  �t�<[�'jc�ӈ�*��{��GtXm�� ��FڛW������� յ����5�Jg����;�~TO��Ӗ�;s2k&k5�2h֬3Ɂ�Ԉ�Wkj��y��tluʶ�=<;t �tbpXFcX�^˻���V�岚T�hs�b0���m!��z���U��� �[�m� =�M�䍼��F�Z��hRՠr�@�ڴ���ME$	�`�� m�~� �p�^�7�أ���%�H�^�z�ՠ�ݚ.;������"���b����E���d\�!3��&�v�kZ�=*2sY�2�˫f�j1�'�8���>���^�@�����^���Ks#�`&� ���ܺ��wUT�$Z���@�ڴ�:���@ۉ�I�� �-�6��@�ν�|�Y���S�X�Z/z��j�<���*��@����<M��/�����5�h� ��� �������]j5�+��6.�sM�6�eu�1�� %݈�����W��R�-�?r�9qܴ/�s�u�H�Z���ME$I�x0N-�Z�^�z�ՠy_U�w�أ���l��ӽ�ߵ���2��<�r�*'�z��"FB`Lbtb���
�sC�g6��",l5���4���aH�#E`�# E		X�! -%�E"H�"�X�"��02��A�E ��D	X R,!��%�A`�#��RD����
�AP�mGh�� j��T� �A��Ch��T�)��#������~��z�{�@�}Rƣ�q�q��V��}V�k�h���^�Thm̏$q�qŠy_U�Z�Z/z��j�OpK��M(���1������⭅��V]��-�9ضp��-0��C�X챧�@�ڴ^�z�ՠy_U�y],�bpX)�b�@��W�Z�Z��Z�ՠ{�혰�Ƞ�X�R=�j�<���-v���^�{�&�rF�H�I#N-���qn��r�r��s�pVv�;}�'�Bqh�V��ޯ@�ڴ+�{�CZ���q���"ǐ�D�X�ޝۓ�[P�]4�:b�e��j��NTQ2)��ޯ@�ڴ+�]�@�}Rƣ�q�q��V��}V�k�h���^�ThRD�H��@�@�ڴ^�z�ՠu|T̍ōc�Dܑh�n��r �� ��n���/:]���h_��J�2E���-$��޻�mS����׽��3-�5k��7eJ8g65��z1;N-����9#���:�	;:ې���y��эa���Zq�;m ���m㐫�;C�8�u�f�sٱDDq�[su��ŵ�H�w:V;&��:��ەhŷ.�ug;�HF .�-��{=mj��s��x�����m�X�.�c�St�JkqsRʚ���9��7�]���qƹ���l�����wwmo���=Z!�v/sh��W�5�=u���=Q>;u�#6��\nĥsۗE��ґ�:���<���-v���^�{�$ҹ#o$y�'��}V�k�h���]�@�z�C"�6�6����-v���^�k�hW�h�(ƤcD��dR-��\qn��qn���e�)'�i�&�k�h����j�=�h���\{kHdC���9��]�fnÚ��Nݎ'�;���Ņ,뎠(�U5"�@N8�}}V�k�h��4]�@/��fF�ƜM��h��?��
H�@�b�T`," ��!���ﵹ'�g���~��Z����NS��7�y�@\[�{٭����tVa��&�0�Mq[) ���hψ�wM ��m$m�#�$��=��Z�� �������p+ǹWz��c2]��&*A!�M�eW��!Pfcm�:�M��Se���	�u��c��������/z��j�<���;�lQ�H�B~��@��W�Z�Z��Z���;�T�����F8�@��Z���G{*ꮩU�U�n��)��/U�4FH�M�	���}V�k�h���]�@:��pn)��n �� ��� \��9��=��߼�x.+1�0���+d��.&Hk��Ս'u`{&e:ͮs�쮯X`�xpfv��^�5����qn�c�&�#���ґ��V��}V�k�^�z；E�x�Ȝ��� ��n ���6��@5��{��f,Ǎ��I�x�%�R�:- �߾���{�r~TJ��[��ܓ����H��ɑH��m��ՠ{��]�@�ՉaV�"9�C�-ٮ�{2ݢ�`x �T������<�
&��"X�m~�#qǠZ�Z��Z�ՠr���9z�Q�H��� )���=� \[�z�� \[�yՌ��p�4]�@�{k�-v��l���t���
c�<��=~\�.-�=� \[�yc�&�#��c�@�ڴ}��s�Z���@uW*���֕bHK{S�譧f�l`-&R{u�!f�� HMVB����m��9��Vy�$u�[[
���r8;5���E5տ�}.������tH�TlI�q��N^�7ER��e�r�"8��z|�����ax 0u�F�N�*�J`��q�]������rnν1�L����y;	˄��#���zzzv�#��窒��)�L[�������KΝ���C��c㑚K����8P΢ {4&�ۍv�;+��(TL�7�L��'���4]�@<���j�=�QH�2C����-���&h9��{��>���4��H��l�-v����k�h��,j6�$��4�.-�7u� \[�+��6أD�F܂rE�wu��-v� ��٠w>�J������U��VVr�a�[Sڶf%��@�ml���֍�E�m�³`K x�31⧏�cy_��ȴ�{ \[�n�*���/;v_y��L�]�'=�kx����`&��j�/_�4]�@����d�6�0�� �p�� \[�m� =��h�#i�pR18�-���ՠr�@�ڴ���2)�$TXw����ou����eM��~�7럸\1���q��vNe�3;l%�f��jxx�3b�h.t0֜��`����n���qn��p��K���8�c�8�]�@�۹�Z�Z.��y�F�&)$nA9"�<��h�V�f~K�J�]�@:��#��ә�Z�Z���@�}�B]U���~��8L��
~M��@=�٠Z�Z�۹�Z�Z缄��cQ(�&Dg�֧�eD�F�M�]�vI;m؏\�y+�Ӷ��Y��ˤi���9<��-�m��-v� ��f�{�&�rDۊA����=�ݨ�� ���Ÿ�;f{ۊH�&L�-v� ��f�k�h�n�޾��jF<����{�ܓ��z�I����rmD� l�6�y�ݺ�k�5_�q���rh�pye@�{�@>�Ծ����:�KI.�v�i�f�fo/ ���Mh��d�v܎���%j����Q��ʀ.-�6�\�.-�u��$qcR"L�9��ՠr�@�ڴ-������N$)�7�N-ou����e@����f,M6Y�C�Rd�@��mh]�@��^�{�&�dM��"���p�� �ps��q C�&�D$A2FBD?@��Y��3$@H�@4��œ�ݼ���������6N�v���7�P6�$��!4���	��1��BYm*@��їX	Y4$,��$I	H�`�Yh"YH̀}
dB:HHBa�I!0N8�m#B!��K�E�H��)BA��D�
āD�!	@`I!�$X1��"H�a2,H������B�Q
M��"�`Ұ)VEY@�}�9[�kFݰ�t�Z�2Qe�n��ٴ��L�\���N��n�ۡN�s��N%���q��s�:�N�TPNV�ݚI"�!rD��vգ��H祌�Y弯WT�!�5�ոT������v����t;om��h۩e�:�ڳ v�#���2'^�Υ�K�VW�}Tp�M����C�3����85�*��<	��=Ρ�V6.��6��8��Z��;Ӭ�������}dD�n��l��,	Wm�z�vS�vټ�.�T�*��p[p-��J##��s��m�A�RYE�M�����3A"����n$��9K�.�P!j��(�x6(����jtٸ���[��x:Nd��s��Ѵg�yc����m��E�ۤ[�&�gFX�{.Q,qF!yTR���;V��Bn�7OS��ŃCQ�̫\QŐ�F�y^��*�:������uG�����������8�f���-�@��������Z�4�݈�V.�R��["�g =��i��c��^���N
볳�kp��P���gNu�n4�%�6�m"�΋nAL�g��f6�L+��Ѻ)Z����a{g�cV��(��J��[j]�)ܾj�Ug�-����]iͮPeZ]���)h88�@Ve���[�<W75�ڊv&�\��[qǮ��������t4�mb�S!���$zn5g;�n��GT��LEr��;�誣u�U[n��`�*������2�!KU��fU��cn8(퍢��+��)�q������YGY̖���ڸ�v�q-��:"1�bX�����+Jq���#�n�)]��5��p��(<!=&��M��c��f�<�cn�0���:�].ݶ��ixk+����f*m\2�e�d6^8f]-Wmٶ�:��� ��7�;��t`:�˹�)d�ʎ�zQ�C6��X9�j�*r)�[��ܖ����C4k���I��t�e��	N�ZmJ����']�C`���-Q8�Ԧ��V趑 8�-r��jɺ�]�[�k��E�МY�8P:3�&��{pk\�f��М7���E�G;`��.Myܲ��ͺv�!%�ⴒ�i�]�\����^��,���`XT�V�[���N�ݱr����.i!㧣 � Xm������ƕ�͛;ce_Mۡ�"�����m�^v�ϲ�����;x^ٍ�g��}tW&J{�ֺ��J�:�1ѝ�m�g$�V�����nI�GO0���4gj��8v���o�f����Ÿ�ʀo��N��#FL�ԋ@��^�k�h[w4]�@�_T�����Q`8�@�-�>VTqn���ۛoo�d�$�� ��h[w4]�@��^�k�h^�c$q4��!"s4Ÿ��Ÿ�ʀ~�UU;W}��V&i�]Frƌ��+�����c�����/*zm���"ٷX`��9�v����Ÿ�ʀ.-�7�]��l�&���G�Z�[߳�����EhC`���w{7$����䝽�z�riDԙ25"�@�۹�Z�Z.��]�@�z�C	"���с����p�� �p���;ޖEDHcĤZ.��Ÿ�ʀ.-���_z.,�E�ޗJ��΂:�rB[gm,�Uc�i��)�PrJpn53?6�~�~�6�[w4]��Uo�@��(�#�$�H)$Z����j�9wW�Z�Z׬XƤ)1HH���j�N��ٹ�CI��~7��ϻw$����?wev^	�K)�tŘ�%��]�k� �c��+* ���7�q�t�(�l�z���<��h��@��^��9,��bxE"YLCm�vy�]�7�nSι�����N��9���"�Rd�〜Z�����h���-}V���؆E$��L$��Z���uz���<��oؑzϡ �,u�*t�Šr�@�~��V���s@��~Zz���F�!9c�8��n�� ���9ʫ�W9�������v��@�u?�H�̒I$�-��@5����n���������u���M3&j�^-�ڃ�et�!r��;Y�s�����/i�5�1
��?���˺���h[)�yl���<�m��-���_�m�|��h��?��j�;�� O"����1�Ϲh���%�%#�h���{�H�&�I�)�Z��h��@��^�ٟ��K��/_�!��9#o�Z�Z.��]�@��^��U�z� �=y~�F����,K�$u7����۰�'M��#DL�I���^�0�gr��tv�V�n���<�/\���`��F�k=w)�\푸g���Nسh����23HV�f�F,;�s�H�{��t�%�v�tq��xٻ�V��ձ�
-�� b师z�.�X����G;��=�XPEl�ِ��n2v�{[5�h�W��#��<-�U������w?��=�ߏnp�늺����Xx�-�����m�%�h�g���:�9"z#Y�Y�����w>�~��>��꿘}���Ns䩬mRkL�x��Ϲo�T��&C@�ȴ/{��uwI�&�#�$RH)߾��է��%˪�[e4��b�!����>�r�kո����z��� �{]��x%�����h^�=]��I6���!�w>�~_����N�tu�y��׎Y4ju���������tn#>H�x���	�Cbx1H�l��岚��}_]�]0�O��t��}��c��l�� �z��\�]��p�� e7�߳3/_�!��9"o�8h|��h���-����h�K	�c�X�%��%������$�h[)�Z�Zz���X��G�7=��k@�ww_�l?#�h^�?�o����}�=�tn��7,u��bٛ�4���Ѷ#�8�Ӝ<[tl�:�IB�E1��!�yl��k�h���3�g�I2ӡ�x�k`<Y�������z���?��r���W9�o�e}��x,ci���"��wvq����
�������ܓ��޻�w�ϕe�b��t1f=��ꔓa�{���@�ڴ]���ɤYlpĳ�-�vq�J���$_����k�hzvL_�u�Hq��N%1�����&벪nܐ�:�m��i|�>9om4gj�8�ư��ՠr�@�ھ��������/Y�$�<���H�^�=���"G"�?��hϹl����"��LX�Cy���o3�����M�j�9wW�{���F�do�1hK��_�l4	�@����pU1 	W�P�*����k�Z~��q4�R�C@�ڴ���t��ȴ��Ɓ�����=���vk��]��n*{y�]k�ٮ���OQ����l�^q\)�2�ͷ���zs�Z���U�_�9���œo"��b���V�岚��h^�=���뺫l:D�/�7��〜ZO�@�ڴ]����@���L���<x��1�.��I�-�tzs�ZZ��a�w�n,����3��Y�@�����������߾_�{��@�}�@����QwuU^�&�C�{I��#Ʋ�i3���p�x���Wn�Au�ڂ,]ku�è)�a��h�eu/O=WO-�i��0��n���v�Ӊ����v-�!n�t�y��]%��3�vܢ�ۦ"��	�ӭ9�E 3=�$�rFt�넦�Q����l�=Y�6���k� ��u������A�	e�����$ؽ��ٷ���;:N���[t�7^�,wu��Wbؖ���d@Z���`1�U�ӱ�a�qo0��1�G"�?wgs�/��<AU�=�b�&�G"I�E$�h/R �� ��r ��?r�v��5�86�R�C@��~Z.��
�W�yl���,�&(�x�K�m� \��/R�W/� ���d�Ȉ��b����@��M��h���<�*�	M��w�|�]���%�XMm��,���m��,f��p�.��su5Ks<3+1�x����gƁ���@�����uu�S��;�4�a����\�Rk57$��޻�	�*�I�����9=u��rN߽�nI�{^����~ؤ�d�%�H�
�����ԗ��G"�<���1bM<ȱ���k�hu��-v���ٗ���>z��6�o1�x��1�Z���@��L�~�tzs�Z��W/�8��k��k��ݙ�n6�k[;Jݢ�냡b�eݿ��|�rP�U�hx�?�Z.��]�@󬦁岻/�X�n�*Š/{��wUwi?�Z���Z�Z�����Q4�0�� �p��C�q�Uo9EW
��E� � RD��mB�B�E�hLEL�1��
&�8����	 ��B �J�(� �A��rXbD�� FF�VI�iЕA�D�# �y� �1Ah�
8�6�O�A�!�j�m��.��y�g�w!�^�{�&�dC�&7$�8�?��톁#�h���w>�{�ݦS��Y�T���;��hUU_>��#�-�e4
�����E��챲u-ڙ���`�C�v�k���-�t�֐j(�PX��@��^�k�h^�>��$}���b�16c0�fgr ���>^�qn�����]��h�8⑲)�@��Ɓk�h���-v� �ԍcR&ӒcO30Д�΋@������@����BA�0 <��]wUTt�����쩗�̬lm:T7�@��r �� �z�Ÿ��9\?~�o�M�'�w����"����n������8�7\�P��;�/������[�]�R>����-�e4]�@��^�{ܚE�92L��	Šyl����#��-�~zVנw�t��I���ǆ�������s�U�������;޻�QI2&��)����]����H���Ƈ�vH�^��!��e`ř��^�z�_�l?9ȴ/{��*��':(�$����:��j��xvyf�=`8��=��9�ȼ�.A�I�n�N�����΄�����nZ�_cȕ�8������v���vqq`�zڲ��wi��F��דDN���fӢ�y�d�l �m��ق�յ���:(wh8��0g�k&s�XN����E���in8D�X�f�/���2 �t��FwC��y�-�3��zd�rk�35�JO���͵t�vڲOSnܝ1h��wn�Wj���*i�����߿w� w�j��\�[o�cR$ӎ��^v����ws�=ݜl�����|^2����P�\��?�̀7��^��[�.m��!�o��;$ZI��/;V�������,�8����Š{�8�%N��9I��}�@��C�9��6�8.�(��rVi�	��6eދ�jv㔅�狶�k������� �-�6���� ��@=�]�A���6�I)�����ٟ��߮��]UK��s�Z��h�ܴ/�sLQO2QH��ՠu��}wiNr-�����.��(ǀ�$�@�e4�ՠr����b�߾z�|�R$7"m8�7#��yڴVנUֽ���=�rO,rAL���5�4bnX��]�v�t򎧧m�)��Z�Yz��WK�x��m�}�����������U����@���"&6�ǠUֽ���/;V�����H�Z�G�$���&&��/�w� w�j��\�{u�k��x�n�xhE;$Z)#�9{��}uWk��h�d�0k�Xڥ��m\�7��^��[�~�W������8Ɋ��v�.y.���s�v��i�v�nX���P�n�L�t�������>W��h��@�mz�sV&��E�@�e7�#���@�$z/w=���� �c�፷��p�>����
�נwYM�Χ�)#M&ذn-�m{$�｛�w�צ���V�AX���߿~ɟ�!{n��ʨ`6DLm�w ��u�@Ÿ�\�z��w}SBb��\
���պ�7��z��S�˷����a�e���xY���z�qn�W?r��X~���j���H�m<��@��Z���
�נwYM����οF�m�`�2��z/y@=��z���bb��M�b�G�Uֽ��h�rЖ��@=����0Y�<��Y� �z�qn�W ��r�^?�@�9~�;Z��+i������:����m��ۇasY��M�k��wf�O���L�Z�ܺ�2��A�B�1��\l[��'7k�$$�FӜ����fX�\�.� �D�,���M��m�#i���k�q���͓�|l�Zva�xo��.8U(�<��[�H��p���ɧkm��3�<;
��nƇ7�N�p�t�ғ%I�~����|��~+˛ө�6"�浗fn����ٍ��%�l.��x�r�C={��r�>%�U�~�_������
�נwYM�Χ�) �M�X��@�[^�WZ��)�^}�e�$N|����:Cx��G�{ݜi�]RS��@����y4��I��ǙI�z]]R�M��9ȴU��
�נy�t��I���;� �-�=n� oW � �v}���3��๫����܏Ma�=Y�;U��m=[�s��T���{���>Ed��^�_{��Ҡ��|� �� �}�M&�H�Nf�WZ���߳�����f^ŠNr-����?���D� �!�@����i��.�mht�@?wsXbX�i<��'�B]��t����@�O��^�z����y�W�) ؛Ʊ7�׮��w]��>��>s�w�r�?��y.Mt�3��L^x����W�Îlsg�vgl>�^�5��"ݲ茏ak�m���~����ՠu빠{Z�4�"CM�y��z���˪���E�t鹠Uֽ���H��1��8�w=�'}�l�?�X7`��"� ��0�M�5�V T�
UR*��E�*���n���O�=�?�Z���qfbǘ�t`_{pu� oW � w�{�bȣi5�E�cs4
�נ~����϶|���?�Z�ݵ�~�u���	�v���I�z�]�7d�������`g�4O��&�PQIH���_U�w�r�=��U�E�= ���1,pQ��m���/;V�׮�WZ�s�-�#���f`�����-�M�����]�R]E�Nr-��<v	�`�M�V��U�\}#�A�lll}���؃� � � � ��}�؃� � �(uD�H��  �BA����6 �666>�����lֵ)�35�jfk6 �666>�^��A�lll~����A�lll}����A�A�A�A�=�ٱ�A�A�A�A�g���3�2�M]\�ff��G���J	�Ƹ�wo9�B"6�rj�OnF��k��ֵ�h��.j�A�lll~����A�lll}����A�A�A�A�=�ٴP�lll}���؃� � � � ������˫�֭�&���؃� � � � ��}�b �`�`�`��{�b �`�`�`����A����k��EP�A�A�A�}�M[�������34lA�lll~�}�lA�lll}���؃� � � � ��}�؃� � � � ��}�b �`�`�`�~��~�V�ԙ�����f�A���b��A��]�<���������y}�lA�llQK��}�y߾�������C;���������6?{_}v �666>��p؃� � � � ����؃� � � � ��{��A�A�A�A��:�t0�dC��0 ���;��� �A��A}�� * A�R�!*���)a�I:1��a�!�Б�+�a�c$T� "Q1d��hHȱ5����
�^Z�]$�%�
]��rFf�Dn�8�g���W��� �z��:�x��3i���GkR�\L:N��RR����N�-0jT�F��M�Nk�ʤn���<�&���//cu� -N�sW5��K�G� ԛ	@�K���s��f�#P^�Al*nvB��aP�"���v�d��,����+]�-�u(�cx�4��=�hܣ��ۜoi�GgT�h���lj[xIӱӥ��[��GJ���n�L��*K�t�()�R��d,i�mN���1R��sf%��TX�LN�n4�krm�l�=:	c)�f���;a�i�2tv��6�P:`mT�6ٻ;��E�G��r\��ꒌw.\p�f.���d�:��0�+iN3�˥�딶`x�K�)���]�[m2���	�W)�ݺ\����:�{e��"��\ӵ��ڴv5��=��v1r�����[�*�.ԔKg�nۜ.:7��-$Н�^Uqn�55l[�rԢ�;���Wd��zz�s�νrF5[�1)�9�\WU\ڗ�m���X�)78L���70Y6��UG8��۩W�t�T�&Vꌋ*�r3���m\�λq��*ʼڀ��<;�)��6ͫ����z���j�v�)l�YYjP6`��^�Yvp����r>ZuK<�M��z��ɗ�v�ݞW��v�2����ۑwiխ-�\���X5�om��&�R'Cn�j��)i{�UKkTc�"U���I2�U�.��� h�و��-�#mؕ#=�N�S&��bC�͉kMZr�e�Ss,)�5Z�]�]q%�T�^�<c�UE���/^B��Y�R%3�cGF��O����wc���F��e��9��*ݦ�Pgst\���&����o'.��밲M�ٵt�J���sbU��ץ��݀�l�m�v���kmf�r��Nxs��W]���X˵ ѱ�l�6��"5�|��]�=�X5e�ѩ�5�-՞F�	�8�� 	��Uq@6��Q�O�k��H� Dð�I�06�(l�=%;%�jXB�m����Ŕ6ŧL'"�!�.{���fV��vbpc���sקN�=i�l]�<�����:K��
Վ��ČM'lLg���W\�@�Y݋\6M;��z�2�!�;�tY���v��h��Av�9n��xtKv�D��m��nLX��'[v�'Lúb
Yfo�:��(ɇC��8�v�s;u�vx�;�����}�v����^��i�#s���mb"[�=;N�+���!��f��cW��tyŭL�sK���"��666=��p؃� � � � ����؃� � � � ��{�@�lll~����A�lll~Ͼ��.M]Y.Ks5�b �`�`�`��{�b �`�`�`����A����k��A����{�y����j���f��L���kS3Y��A�A�A�A����b �`�`�`�����b �`�`�`����<������͈<����}�4d�֮�S4fa�5v �666?{_}v �666>��p؃� � � � ����؃� � ؀�>�^��A�lll{�}�]je��֮fR]j�A�lll}����A�A�A�A�=�b �`�`�`����A�������A����~��Ⓞ՚�\՗55�5k�v��v��d��JX�ob�ٵ���k���;z��M[��kN�V34lA�lll~�{�؃� � � � ��{��A�A�A�A�����H!�9���ᶪ� >�5�f`7�e,O���[Ȁ,@	�6�V,B!	��*A�R1I��UH�`D"Eb@$@�D`��h�qN��Lr-�N��9{��ꪤ�ӣ0Ĥ�x�R5�@���-�]�������/���RF��Ɠqh�����@�?rЕV��E�E!0	&�nL�*�^���Z�ܴ��q�}U} �R�bW�R����M���N.��k`^Sڽhx����`.�'<�C����"H,i�$�q�����Z�j�/�)�Uֽ��La$��m�Yۀ;�p�Ԁ7��٭��vo_��	D��7�`�Z�ύ�i3����wV�k�=�udj8�YF19��j�:�V�yڴ?�ߕ�~� ���V'�'�e#3��}� w��* �-�^9�yy��FR�F{F��7bb[��{N�A����AE�w\0C��٩ւ�D1�m������* �-�5�n y�o�_s�5�bn-�]��h_U�^v��J���HbMɚ�j�=�ܴ�uV��"�:t��?�˵	 ���n'���Z�j�:��rqL j(9��w$�{��2MkSZ����8��ՠu빠^v���F�;+�dM�cs�Әk�@�Tݩ���ݐ3%��n�1s�.����lA2�0�@�n�z�h]�@��Z��:�5X�n3����[:>�@��Z�ݵ���� ����8��&"Hh�~Z�j���K�M�t�Z���x�'�6�f,O����S�E�t鵠w�8�=��h�u~��44�4��@��s@�Wu:l?��Zy�-U���?Z:8ݳt��eی�/c&�۴Nuj	vB�3�%G�;Bl�[��;q�q�q��ɳn]:��iu9�W��ȴr������ש��fL�;RQ�9ꍉ3�"��Ƀ듰Q�q���,��ZNSl�6�4�GL`���u=3�Qh �-�8�Wj�'���'=��u�=�O)�#�������E����ä�=�i�0p']�����6�5Z,pZ�o��6�'N*�]v8�-�]���`G���c��ŏXP6��I7�_��2W�h��@��s@��!��&�M�����Z�j�:���/YM���I�Q4��yڴ�w4�S@���ΰ��G �D�hz�h�����Z�j���ő)"�q���h����UUUWL�9ȴw�k@����{%�js]�8�2�sfںl\h�S��2�U�X���P��.`�a�Z�5�`�5��� �YP^� �gH)�W��c���������������w����nh_�4������$hi�Ɠqhz�h�����Z�j�*���@I���4�S@����hz�h�R�0�M��p�:��@��Z^���)�_X�1�q�ƒ�LCN(�k	�7!3���q���=�S����٫	�U\�DrF�cN-�hz�h�����Z��� (���,p�@��ke�]$N�����Z_��b�D�mLb��^��W�i�3��P: '�>�}�ܓ������Qn!L��9���ՠu빠^�����H���)��o;pqn��������o���.�+�,��r,��ܱB��L�
xsmp��8�]ed�{'��@�]e�go���PVT\�����J���H$�I�3@�n��$U�@/;V�������?${yJ��H�i���}�-�hz�h���;�����m��Z��}g�]�=��ٹ'��lܝ����f~VJ�o]r@Q(�#�ĜZ�ʀ:��� w��W����1:��cH3�OGn�sVnn7[yt���ۆM,����\Y���|���Ӊ�e��?;� � w��* .�R��n1����W�h��@��s@�e7��߱ ���H���)"�Š}_�-�]����:��@/s�����,i7�׮�^��������;$ZRa@�f	$�ܙ���W�h��@��M�?
�~��=�]j٢K�u��̶zi�]���,��kq����cE���NI$xYx�>yՇr�����y[�7l�!�em�
[<��d-�Ju�-���Xᶒ���IS�����X��z�˥�q�(����}�^��XYm��/�@s����;��u�[� S�1�69"�v��m��X4�*kp�ɩ+�v�k9�F�^70���ԷZ%c�Ѫe��T~PfM�|:x$�mu����V�,�Ŝ�skZ�r�3ǷD�k�A�������}��}�@�{������&h�"x�H����i8��ՠu빠��W�h޺�8(�slx7���mh����.��n|��@�}>z�u��%$N&�f!9�W��9wW�Uz��n�_xu(���cU��Y�@��s�>������|��������yؗb��'���JC6�F�Ηn��9ztGWmmX�G��蘜􃖭���j@N=���[w4
�W�r�@/s��q�O4ԏ@�۹��6��LAt?9����f����˽�~���H�uE�a��m�m�E:=�����uiE:=�wۚuR�@�$4�m�ǡ������>__���빠Uz��ʞ �&�QD��zW��<�w4
�W�r���<��۪d`�9&D�	���U���D�p�d׌�J/H��T���{�5���J2dm��q��_�4
�W�r���*�^�w�f,�I��3���\�m�\�6��eO��U�~�(��ؔőa�@���@��zi 9<�H{�7.JB�����
�a+),�@��h��)��1�RVX�
P�@��`B�� E�m�!IIB��B���6�v�u�s���	�S8��'8�D18�Np<X�R��"�:i ���
+nb��0CL
���A&����A���X0"J�&j�XE��\$�F%����U�;�|�x�A�!���'�C�&�_� �N��vnI��{7$����Ս)#i����zW��<�w4
���J��\����qV0m��_{���@u�ߵ�n� �?޻�Q{R�7AИ��k�gI\i[a�����`���,mK�ˈ�w9t[���+��"�����z.�?��� ����-�?�@�$4�m�Ǡr���*�^���M���l��	"N'"M1�������IUiE:=��=�zY�
%$i��q�g����~��}~�ٹ'o��7'��8"�7�>���o}1AD�c��9���]���G��G�~�g��:��V#��2-h��-���.�P ������ZZ��9�Elrf$:v��F�~m�O��zW��<�)�Uz����#b���ly��=��sߪ�꫶�}3�@�_}��^�zyu2
8����s�܀|�R ���k��� o��X'FbM�6���G��˯�@��^���M��D0����f<z����U���?�d4^��rO*x�F� �,�%�2K�i�[���q;���V݆%X;��3������e�A�r��ew�ƺ�m�Inc��F�.�*6F��jN6'�ٹdN���Ch���23N.�l��~|�6�M�޹x <Ì�;s=e0Q���%0ޮ��-�k(M �X7^P@UjQӳ��;%W�]ugqz�Ǎ���,�qsk���l�+H��9�n��v�^�*:.�-�&f�,��E֌��
<C�K�Cp��0�%�Si�q�h�a���^A$HrGC����=�Қ]����� ���@�߶LpQ$�A�;���@u�ߵ�~\��$N&8�c��*�@��W��J)��Ӳ�{�f6�t�(U�@��W�Uz��ҚW��=�.E��M�@N=���~�����S��<���@?wu$#+1,a��^��Ԛ��D���ۧ�g�	.�����L��&(&���z��4
�W�r���*�^�U����Lm�h^�V~��g��͜�W�Uz��Қ��"I,m��z��������*������"����[�D�'"NG�Uz��ҚW��9{�����RD�cI�r�n� ��� m� S��o���Ԝ�6�훮ͰF�[�V�'Y6Й���݈�UM��j9nΩ`�S��j ۮ@6��@u��X{��T���$mA�Q��^�zW��<�w4
�W�{z\�4)#hm)$��nI���7$�}�M�8(,"?)*EH1B#P����=�~��S��Rb�o#����H~\�7���\�6�7]�Ơ&�54
���u�@�����Ɓ$�*�E�6��X/���|A���k`:V���j�3�4tJ �9�OB�D�m&ؤ~�����z]�����W��ޕ��,�ȓ��� u�@���\�.���RaMǠ^��^��
�נU�^����PD�1H��n]�ҏ�=.����z��wU@�c"�*���ߦ䝾����e$bXL�ǠUֽ����S@��^�_o�4���M~R% ���K3�e\�&s�M�й�4�\�Im�/W�	�	������
���/YM�mz]k�*�S �DM��R=���7��z� ou�n�u�*򚀛x�p�*�נUֽ>����_+~z���z�����%�cM1H��r ���e@��u땖�"X'"NG�U�^��빠U��y{���]���$�b��y����$6���j��[@�qQ��D+�f�a��ۢ2zF^ca�m��m�9^0Ob���u��^�����������ϵmv���N�d��)�Hgc�t��6��v[Lpu�rܤ]�S�v=s1�|�r:u�4��4��oN������ݲf�y���O$ixD���c���,j8��У�#'gf^snP�4u�ՇM{�������>�{��� ��g6S6�·�Wd:��L��8�,�Β1�4��n�ͨ;-F�d4������ۚ^��^�zWj�;޻��!�H���r���k��\�|��۩�{�h�"7�q����*�@�۹�U�@���Pdr&��s��-� �YP�r����5+��dI��#�G�ym��*�^�˺����g��<�BFG���|�_(*\�Vtq�:�M'n�Cm�k��d��8�k��1<jm�rL��}��9wW�U�^��s@�[���,���#�@��r}_�Ur�}�W*BZ���YP��4:�1�I�H�r=��^��s@��^�˺���f8�jd4��@����*�נr���*�@���PD�88�RL�*�נr���*�@����=�|*�dJbk����ל΍�WY�9������a��Y�V��0�ԡ�	tf�����~�~Wuz��.x��� ����mF�bs��}� ��q�U�@��W��AN�|)�E��#�=�ύ�={ٹ���M�yN��u�^�U����� �54�ۆ����@���=���C꫿����4_g�P	"YlR=��^�WZ�/Jhu�@��Q����hJf���qVf�nBJJT;w>�槷=�] k%�aɍ"H�G2F���[^���M�k�9{����b�A��A�Jf=�{8ؑ���������k�LD�8��(�Umz/z��k�<�)�z��d��Qēj!�cЗK��=)#�?w�kAUU_�wWQ]�V,�=��icƝ6��3;��r�n� ��� �������%�u�Ӗta�YFn����=SHg`[��VWhV�۬Z��ˍǠyz�h[^��ޯ�3<A�����w>y O$x�LmɚW��9{��[^��빠x�ej$K"bm�1�_��r�示���M�/����,ȑ$D�F�r=�k�<�w4
��@��W�[�d��7!��jH�/]��k�9{��{���8q ���(�XA$"I	���0��\ ��B�֤Y����
zQ:!�h$�� H@�F0(���B!��$�B�
Ċp��4�H�!y�$?~�#��D$�H��
�ő*@�D�a,lFH@��RK +@����*Y��B��~C�4(Q�5t,b�Sr! � L��i�*Ĉ��q ������D�@�	b��BD�USdE��h!��� ��b���K�SN�X�% �WCJ�,� ��
A\����9�R� d`@�E IH�H� B Eb�U��#��h1 �ňA
lA D����b�
̅n��ĉ�+$ ���
�wo��x�=���㿀T�W+9zW�B��RL`7Q�R	LU�jt)��ne�T�T^��l�: �c��㥲�5�Y�4۠-���Z5�v{@;��E��u��g�T46�����ݮ^�H]!�q�d @U�uq3���(�6�U��5-��rt�vI�kX͘[0��T�L
���	�h6$��l���ֶ�ʖEm�
.��]n����mڂ��v�X����wj����	�RXWn���l��|��nf�us�՜�f�3����^�TF�]��0��-,�j5	5m��S x1��ڭ��=���M�m�u �űr��N����E�=[5X���j��P�!��mΉ䪣���c�z}v݉�mktpvUt^`FF�&t���$���c��u�������Ko���
,�m�.�k�m�u�e���b���۷k2nke��8���[�����
����m����D�$Dmeh
�s2�V�� tjWjEh��B�y����4GnWM����<l�<d����vB�v��U�V1ш�u�ꕞ$���"7vV+i8�
I��g\�;�V����Tl,�YP�ۤ�I9�mjJ�5��P:�
��6%U��i���jV�;��� �ѤL�mR��'R��Y�n.us�\��͆Ķ�Ѷ��ʻ]q�Gvմ��3 ⇶z�{(�L�:km��k�p�2�*�v�e�q ٸ��Z���72��R�mtv��r��@UA��P*��v�Mny�X5�);1�gF˧�Z[�m��}�Jm:n��N��mBڶ];l�J��+�q\ؔ�1��*�5�.��1���-ۥ	����7_>�Ol���y1r�W
�ף��M�xȸ�଺%X��q��N� (�U��K�nWW��k�n�nf� w-l)�d�Z(�-��.̫��V�Q�۴Q&tu�:�/;{	&�$L���:0m4���e�G(p=�!r�ư�	.�Ľf�7[��8�֧�>j�#[A�$TN)�( ����
s����>�& ��^��l��1ڎڷ0ZJd��v��n�8��/j������볪��^wVX8�sY����3YŮwq��$A�������>6��j�jU��av��:7GdӸ[��K{Y�v��{�wC����1����my��JԂ�87k!��p;K<�sN�n�mwM���Vg�m&z=�Ɨ�,<��=�S����7nK�I+��30ה<5�N2�4p����:z;t뚳sq�w<�;����Bj;Q�E������a��~m�����r���*�^���M�m#iN���Cy�@���=�*��".��Ӳ.�{�U$zvCcK$�I<��zRG�~�g}IE$z/tzT�d&A7�cq��/Jhws�<���C�Q��#ꎲ�N�&�o ���4�럺?�.���Jh��ʚD�@&LM�����[�3v�Jݲ�sƳ��e�'It\��&��$��94]��+k�<�S@��z��2$I�L����@��{+n���WUU}_�~�Ɓ���=���U�I�3)bX�o+M,�z���k�9wW�Umz���LD�1<x�1��B]]�_��Ͼ��I��9wW�_l��궵�F"cɑ��$z{�@��� oW |����~������I�n����R'��۷<] ��um�\s����U��&@n�?0r�s�;��k@���? ��=(t2
 �8cq8�-��]k�9u�@��z��W ��G���ܙ�O^�ٹ'o}����B8�6!��0
�j����LimV	8p�W9�}Uۗ}\�y�T�Zs�A�ī��c����s'�=�>���������,ȑ$E!J8�^�z�uU�'��]#�<��������S�x���<����h�-���u�-��Tsv�˗Z�Ħ���?>WKT���~�}��WZ�]k�*�^�{��LD�1H�9&hu��"���@�[��=��h��U��&G�=�Z�
����1.��4�#�?����4��7I%�1�}uv_���7$��}�rO_��nJ���1�/ʧQ���[��>�N�5��R\���,Ǡ~]���?H�˺=���������}G�.�"Y;N���vt��6�h��Ʋ��<�*{s�f�;�z��6�TD�q�{k�9wW�U�^�ⶽ�nW�,Q���@��^�Wuz���
���ߒ;��"D�Y�JH���=�mz^��]����b�Fԑbx�n=�mz^��]��wW�y�]�1�F�H�G�U�@�+�����=�{�ܓJ@?����������>�v\�ٹ�����-*�u��t�-��X@��y�;mv͸����܀��w&��]���\N�lhM��pzT�v��v����;\!��6�uc���l��^zlu1��.���R&����y�(D�l..�snۍ�F{>�nu�W��,k&�o*�f�̛�0n����;]�+�����O]�'n��G]��N+�׻��kn;�&gu�ҍ�"��]��ݴ`۱k��uH��v�`5p�Ή�g��0��6߇���U�^�ⶽ�mz��F�S��������{�RG�=/H�]��^u1�&$�YN=�W ��ou�z� �Oy�8G����q�u�@��^�WZ�?����>��y}�|��fbT���w {�@��֮@���ށ�~��[��e㞇��Ma�0�y-i�fq�la����<��iV;�H��z� ���z� ��r ��kEպ�3V˚�nI��{7��U������O����>_}��9{�����Bc$��q�$�@��z.��
�נx��@/pʣ1LpQ$�BU�R���H�˻�����@���Q��4�Bq�u�@�[^�WZ�^�z�θ�Y2d�&i��nq7L���K�H��>-��͗�]v�^�Ύ�	��C�Ǡx�W�U��@���˫���.����e��鶚LN=������*�^�ⶽ�nW�,��m�G�r�נr�s�������]]�����z������ͪ��*��3ǏCꫫQ�@����u�@�z�ޖLQ(�rx�r=���
�נr�^�WZ���!V���n"8��Ƀl����İc�=����)N���]����/��u#$�E$��>W��z]k�9^�@/pʣ1HLMƄ�@�u�{�@6�r ߗ w���
c�r&�D��wW�r�^�~����^���G�r��V�<<Y܀m���r����U_Us�Y@�(����f��t��K���M�'�U���W�Umz+�����EI%[(���2��k�k��8T�gEv\�8�K�ňm�
�)����{����lxĲ7��)������[^���zVנ{��o.F,�s#q)�r����ۮ@z�b�F��ld���W�Umz}��ݥ�tzRG�{��ff<Ǌ�9#�*�����
��C���_��}F|�1G�l�=�����ۮ@W mUU�ʮQ�`������3z5,���]�ɡ���4�γRv֤wKێ��u�kHzc�عͫy8���un��se \e�5p�:�f�EU/0������Zw�^�����e�듷�s�n5���ɗ �d7*1����ή�l�K�j��6p�.�0M!*f�E�8�^vâ�q���[`�n͂�Q�g�����̰��&jkXYff� ��P������������n��_\v�$���݅�n;]v������l��,;M�M��U�t���#�?����@�z��k�9^�@��L�����q��W��U�$E$z)������wt�����<�M��LO���_��@�mz��z��+q,��m�G��]R�:=)#�<���%ҎH�T�mԬb�O)��=�w=뺺��"�=����]�G���rͱ�F��Wd9����&�<n6�LcXf��;]�V�j�	j�.5O��}�������� ���@��q&�"#%ֵ�LֳrO_{پ(�D�L����rO�����7ı,O���6����7���\��:�t2�3;��{��ı=����r%�bX��{Yq,K����iȖ%�b{=�dMı�~�~�om$l��2FF��g��BX�'���D�Kı?g���r%�bX��{Yq,K��~��iȖ{��7���?u��[r��g{�oq�ı?g���r%�bX|(��}��'"X�%����fӑ,K��{�ț�bX�%�Ӷ���f���kF��p��.g+�ob�Yr�ݘ���^hmc��+]^���E3���oq���������ı,K���6��bX�'���D�Kı;��iȖ%�`�t��k5i�e˒�Yq,K��{�ͧ"X�%�����7ı,N���r%�bX��{Yq?�Dʙ��;[u+�ǔ�ĳ�~.�t��]G>�D�Kı;��iȖ4*P�ᵲ(oΰզ�C��8���#����'��U�K��Xw�}OxL�'{��;�.���gH��V$��<�T��8	� �"f���#�����8W{��v+k6 �6��c��ډ�)�E(��". �:�� A�hv�x⃏D�M���"n%�bX���ٴ�Kı=��\A-R�Ʃ���oq���~��iȖ%�b{=�dMı,K���6��bX�'���D�Kı;�߿���H�4��~oq�����=�dMı,K�T#�}�i�%�bX�g�k"n%�bX��wٴ�K7�����}��V�S�ے�|��.t��q;;TŚ�n��<�Ah��Tu�Xs�N����Y���D�Kı;��iȖ%�b{;�dMı,K���6��bX�'���DߪdLʙ���kY��֌�Z��5�fm92�D̩�w�Ȝ�L��S"\�}��r&eL��S�ﵑ9ʙ2�D���e�r'��� oz�|��=���g���ӹ�g{�?vD̩�.}���r&eL��S�ﵑ9ʙ2�D���e�r&eL��S�ﵑ9ʙ2�Dﷳ�u35�fe��%�f����S"fT���dNr�D̩�=���v���S"fT���dNr�D̡�<	#,҂�YZP*ʲ��?��D������"b{��S����8��TqN�~~쉙S"{]߲�92�Ḑ�	�ﵑ?~��3*dK�{��ӑ3*dLʞ�}���Tș�2%��Od�}&t\��� ���v��sM� J�۬� ��`��r���a�eW��v�m9~{�7�ʙ2���k"s�2&eL�s�}��r&eL��S�ﵑ9ʙ2�D���/�w��)�w�Owߧϵ��.\lֲ'9S"fTȗ=�f����� �w����S�_k"s�2&eL�����ͧ"fTș�=�粧9S"fTȇ߿8�"�UY������=��9S�ﵑ9ʙ2�D���k[ND̩�3*{]�eNr�D̩�.~�[NDS��r�����:��X�jw��2&eL����ֶ���S"fT���ʜ�L��S"\��f����S  �� ���s��dNr�D̩�>Ͽ�R��s$�SW�w��)�w�Ow��=�9ʙ2�D����m92�D̩�w�Ȝ�L��S"fw�ֶ���S"fT� 6�#07�I��d�ɛ���6�����&�G��p|�~;*�xn%�l��i#qm�n|�͵g/`�\:����k�]�����j�t���\��Ȯ���mIF���9�L��Y�p3�}�N�@�p��"8+p�U��V�&������.V�I�`�axt�3�sF+����#b�;�	6z��p6��g��t[��v�7�m��ͅl��]���-ǰ�{���{����~ �I��������vg������˞ò��.40�f��l�L�'����;ܧ������[iș�2&eOk��D�*dLʙ��}���Lʙ2����T�*dLʙ�߿~|﷬�<�#�o����S��veOk��D�)�  1�Mj�D�Z�ٛND̩�3*}�g�S���3*dK��[ND̩�3(�d��3WXS3.K�dNr�D̩�=�wٛND̩�3*{]�eNr�D̩�.{��m92�D̩�w�Ȝ�L��S"t��3��5�\պ�fӑ3*dLʞ�s�S���3*dK��[ND̩�3*{]��'9S"fP�P�����6���Q��=����q#8ˌ�{�?s�2�D���5��Lʙ2���k"s�2&eL��k���r&eL��S��{*s�2&eL���p�-֤�.[s&�qWk==�c-����A�7<k�Ɩw��ˡ��c
��U6i�{�7�Os��{�߾�D�*dLʙ��}���Lʙ2����T�*dLʙ���ӑ3*d�)�~���N���S�ߟ���3*dOk]�fӐ�G�b���<�MD�9�ϲ��X�%�y�}��"X�%��ﵑ7ı,O�����]s��VcT|�~oq�������;ݸ�%�b^���ӑ,K��w�ț�bX�'}���9ı,Og�zjZ.�S5�f�5�7ı,K�w��r%�bX���Yq,K���]�"X�%��ﵑ7ı,O���i��֩��ܹ35��"X�%��ﵑ7ı,>A>�~��?D�,K���ț�bX�%��m9ı,N����]��!�i�rp:#�3v�G,�0v<�t�ŵał�y���α�'�TqYq,K���]�"X�%��ﵑ7ı,K�w��r%�bX���N�|��{��7���>�o�A�7]�"X�%��ﵑ7ı,K�w��r%�bX���Yq,K���]�"|��TȖ'�]}�V�浬̙��ֲ&�X�%�}���ӑ,K��w�ț�c�܈H���F ��q7�k]�"X�%��}��{�oq����?�~�WT����[ND�,K��k"n%�bX�����Kı=���&�X�%�{��_=ߛ�oq���ϿmjS��Qjț�bX�'}���9ı,?�T����dND�,K��}��"X�%�����7ı,O$�f�2�Vɚ��q7�؛�懟m�e�j]0���:��{pZM:������{��7������7ı,K�w��r%�bX��{Yq,K���]�"X�%������Bs&a�������D��}��"X�%�����7ı,N�]��r%�bX��{Yq>UW�.�u�6�^�&�ci��m���	bX�g�k"n%�bX�����Kı=���&�X�%�{��[ND�,K��OK35u�32��D�Kı;�w�iȖ%�b{=�dMı,K������bXQ4:pVD���dMı,K����g�jɭh����Z�ND�,K��k"n%�bX  ?ª���kiؖ%�bg���&�X�%��k��ND�,K;���=��y㭧7au\��M��XLn��v�-ʦ������0�x1U��*6�kYq,KĽ�}��"X�%�����7ı,N�]��r%�bX�v�~�?b?b?b?b��P�d���]jf���"X�%�����7ı,N�]��r%�bX>�z�7ı,K�w��r'�����5ľ����ֳ)�a��\˙�k"n%�bX�k���Kİ}���n%�bX��ﵴ�Kı=���&�X�%��;�ֲk&��s5���Z��r%�bX>�z�7ı,K�w��r%�bX��{Yq,K�P��o�ӑ,K��>��[����j/w��7���{�߾����bX�� �_}��Ȗ%�b{�{��Kİ}���n%�bX�:@_zs�nS.GZ�2����t��&���S�[��q��Hp�q�ù,�����z��+:�
p`�al<�W�����^E�7�X9�C�ر���*x�z�{�3�Wϫh�geHΤ-o9ڻ�r��t��Ue�q�.b(M�Z�뭠2���`Ν��r�;��I?�>c�ύ۰gC���l����ƺ�ۓ�M�7���I�Giq���vȗ�������w{�ٻ��s��x�����];:F�4�������X8�,Fۗkx;�W��V�32��ֺ��bX�'s�k"n%�bX�����Kİ}���� ��L�bX��{�m9ı,��'���k0�f\�Zț�bX�'}���9ı,g�t��bX�%��m9ı,Og������(9S"X����%f ǀ�Ɩbۯ��.�t����I��%�b^���ӑ,�dL��}��&�X�%���ӑ,K�����A+:p�(��7���{��;��[ND�,K��k"n%�bX�����Kİ}���n%�bX�����
���l��������ow���D�Kİ�Q>�~��?D�,K����Kı/}�kiȖ%��w�~��}�凚��p%�:cW��-��@��
L��k�K4ҺL����je��ֲ&�X�%��k��ND�,K��]&�X�%�{��[��&D��QɌ���H�Eןt��f0�e�jf�ֵv��bX��޺MÊ@֕��T�#�D�K��m9ı,Og�����%�bw��ӓ�oq���}~��U��Q{�d�,K������bX�'���D�K�Ta�2'�׾�ND�,K���K�]"�_��]��f,Bm�����"X�%��ﵑ7ı,O��}v��bX����Mı,K���|�~oq�������i{9W��Kı?{]��r%�bX>���7ı,K�w��r%�bX���Yq,K��}��\���3W�+�z^*Pz��3�+x�3��n�[�s�܍������|T�:�[$PQ���oq������}t��bX�%��m9ı,Og}����%�bw��ӑ,K����$,i�L1{�oq����~���ӑ,K��w�ț�bX�'}���9ı,g}t��bX�%�����
Z��W�w���oq��^�Yq,K���w�iȖ;]�B)� A#Ea�bF	0�c$ �����LRđ0H�,B0a�H�%V� ���B������7ı,K��ﵴ���oq���߶�)�]7@�;ݸ�%�bw��ӑ,K��w�I��%�b^���ӑ,K�BdI�1�Z]"�H���efc1����f]kZ�ND�,K��]&�X�%�{��[ND�,K��k"n%�bX�����Kı,�g�n��&��SE87Rk��Ff%���:��Fc�ZmӲ�2�������|����Fb�~oq��%�}߾�ӑ,K��w�ț�bX�'�k��ND�,K��]&�X�%�����:��kS.L�%�kiȖ%�b{;�dM���DȖ'~׾�ND�,K���I��%�b^�����K��w�~þ�M/'*������,O��}v��bX����Mı�D�Dȗ�{�m9ı,O��k"|��{��7���>�o�D�j����D�,�Q d�ﮓq,Kľ��kiȖ%�b{;�dMı,
�� "'�5���{��Kİ}��y$��s�^��oq����{�m9ı,Owٸ��bX�'}���9ı,g}t��bX�%=�����'j[�◎n�z��gErN�2[֣�:X�I�ɦnW��u٘5@����Z�r%�bX��q7ı,N�]��r%�bX>���?�Ișı/����r%�bX��}�SZ��kF�F��fj&�X�%����ӑ,K��w�I��%�b^�����Kı/W����#�#�#�[-���)��R�Y���Kİ}���n%�bX��ﵴ�Kı=�f�n%�bX�����Kı=���k4j�r�乭j�7ĳ�FD�}ﵴ�Kı>�ٸ��bX�'}���9İ?�A��{��Kı;��>ө�5us0�2fk[ND�,K��n&�X�%��k��ĐI�}��$�O���lI�?��TW��TW��D���*+TAQ_�QE�D��D����H# D�0E b,B �A	P0A�P"U��(�� ���AQ_�QE~QEj�*+�D��TW��AQ_�QE�D��TW�(����AQ_��PVI��e�� @.r�` �����Y?�          6G�S�     ]�@��   % �@��"��BJ�AD*�@"@) @�  �H� H
U( ���    (�@����������]����κ��}�z�|����_y�v{>��>�;Żlۛt���sץ����    �à b  �tѤM &� ���  ��M4H h�@3� �  ;�� )AEB) �5@0 :(�b �(C���@� Q#� �Ҁ0:6 ����wo}�*��Ԯ� ԦN�W�;����m��N� ����s����nm�f緽�| }@ (��B1 �R�r{�N^��ܯg������R�>츷^�u<������}Zs��|��ݳ�����{�}ϓ޶�� �[nMDͻs5^ۓӧ�}{�+��\{����eק��{�|����  $@M i����x  q   c��n �q{�t�k�s��﻾��� ӥ��À���:w��[χ�� z���9��л�v���r�����{�O&�9�N�:N緞��} @P(@�(cb�5����ž�r�mv��7+����. ;�w��w���9wo�<�{����p ��7����|x�{�ӎ;9W Nu{]��q����������� >�{�O���t����\}����=F�ةJ� h�P�ԥ* �O���<$FF@=��#�*��db41O�BSmT�* �"$�JRD@G�z	�>��?������o���'m;���{���Ezo�� ���� ��� ����AQ_�E`�"
�}������IIp�[�y��@�>��&����%1�S���GvG�ⰲJbk��HԞ�t�H5Q+���"@��4��aL8���+�i�9���=asRz�Ohfz<i�!�n��N���� P���0�l�nixK�k�p5&d���@�g��~�y�b�(�Å��+
E�)w�OX�4��y2k��q���!H�ȍ��B��� HH2R{���@Ć!�E�M�(�I��z{�d��2��<L�`�B�~1?B�Ü��`�0���@*�Nq�乁q�Sǆ��������5�)>��F�MxBHEi�H�\a�
H��!		�`P�HT�`y��聴����/�8y�;?/9\ux���"`o<a��y��k�2�d���!��A<b!4�i��O���'��\˃����թ�Cv~�ĉ�sOe�H�)�"HF,�a�c�F�����2aS e8�%ap�[��C�FJfO�'���o��2p�<)|�2´N,c���&KE�MBXʜbfp�$��0 r��t��8�A�p���N>pJE������)C'9��qݦI��qt�p8$��k����$i���O&��$��@�'���0�
T��<��jDˡ�8A�(br���ZD���ǩ �A�0�,�6CHp��f@}�"1X�zq4�?J�L�x� ���=�'��p�ɨ�C-/���Q��)�z�B�xE`�B*.
F�dF��xZI��fM'��11!Da���@��X���hl��F2�򄩈D�c�!�ٹv�9��� �`��$�S��0H8����� �% ��� ��Č�X�h�R�BH	׉(��������H԰�@��ơ��)!F@��ЋH(0�Ò$Y�,1"BiCHG�p#S9#�
�IM��Hюk��fJ<i��b$�Nl��W��P0�1��#I#�ׇ Wf�2���$8�J�2�����g�%1J>����Cx�{$k�*s-Έt<¤)��ƪbBH� c���Zk�
`؄�@*�:� Pq�NZ���#[&$�`�H�2�МI���2���*L���	�i!�@���ӌHČ HF���6��(�7xXg,1��¥�K� B2��dyV�2Jk��@��H��%S�A�o$�d!!�p2�E���� �9Ν1�"T��B�I`г�Z:0�<�аR'������^�g�`�D��H�$i3a��H�p#rHIS�p� T�<�b��.i4���hI��i��!RĐ�=MXS!w��ȏ�x��X��c���K��֞�ag�%4�,#䙉���%�6ټ+�m���K���w����s'���#Xg4��d����~T��o��do���B{$���G�z�1"�"��"N,�b�0��cC�ňċ4�NT�B2J�		@H2�C�!�&3l�� q�dB@�Ò�a�# FB0�I�r�l�
��!q��F�M���$��$�A���K��0�%�-dd�$�1�##�4���4��!ŰI�-���ZVW"m�Z6I`x��
�1�BH��5�Ӟ$��Ğ\5b������-�bF}�|�gngeB�(�M��Q�L�DB_B"�P��q�u����>.p[��$g�ޭS���d��r�� �ȅr]U��M�؛W�L#ot���5��9�ܥ�S�*jI�%YE���D��}
��9��V�PE���[/����؛�K�7c���"������ݚ��b�[9:Ub������ffL(F*#k.4��Q�4ҥUa�q[�=�A���%dg|DV�]�]�yd�U�����D*��I&L����n�MT�Y5spQ%�������&E(�N"���+�O+�[�x�}�X��!B�P *q`�%����,j¡-��	����$L�%T��W��"��s�g�� �	!K�hB�c�&�X�c
!"t�\&ְ��ڱ"8�h0�@�F�A*a̅��"A����1��KP�-L�,-���k���r�@� �u��H�HB{���Ǵ2kx�x�$8�II͵�����<L?SI$�����q<V�^$.[u�����~@�0hF
DH�P� F�
�h�"E�� �b$$c#��b� ��0)�"�*�2C @���BM+�"����8E�h��䎐*:�"E��ŀ�R�U ��H�T*
@�bXRX�"?�������A�d�1k�Sf��8����i���p������H�0�g0��<�VV\�]�n��	s����p�\�sn2��+
�D�i*@�PR V%`�W ��4X!H Q`�V"EX�U� �D�"��R)�:!.s�<��g�!� �	|MX�7i���
�W�b��|Պiگ?G����'�\93��~	IR�Oܧ(D���F64 @ F�\"D�"D!�% W�S0��QŁ4����h�+0,\H  �aLhF�bX�	I�@�BC�p P�`P�(hD ������C����+ h ~R���H,�A`�P"�"�!ĠD��*Ą�~�Ǿ�,����?y���Ca��)�x��r3�|&�l
9b��< fH�d�xq�B\�9�ԅ8jK��$.i���`F�0�i��8�F�1	�W4L5�N��#��� p�14`��b ����"Q���u��bW9���	f�?	I3�2=���r�`E��.��O�	�j��R���7�_��#Z����y�da��%�Ic���XK���5%6:�5%2H�\�C6����"K�B�+������(i�D!�J`��97�����ѕ��5!] 4�BR�@B�N+�5wiN�MZ&ڱ�F5�����(k
�H, ���i�K� ��!F	�Q �VH!E�H1! ��0R
F)D180j���k�������)CN#L4 �H�04x�`�#_���t8���iǉ� Qp3(cNs��c�p��� B6D<	���� ���#���EJ8:D(��@�KK E�~��Sz��;��������       ,0  ��H  �        ��\�sH��T[6����Ϧ'2���C��T�UJ�t���%�)�X*說�
U�6�AoP�m{m��&K�������    ��4V�   -�-���hM�z���`�l [vZ6�i-�   M�    ��m1��l��#�LY�� m.� m�-��Ŵl�   �	�   �    -�Ͷ �,�;mm��lv����hE��מλl==UiV���� �Z�r@  8��  ]�݀�\]n��  �` � l-� @� m�� �� ���   H;e���/Z������HH� ඛl      m�M,���eIղ@  � ��` �[@h t�� l[@ ��^��m��6������:Ҷ �l���[R �[%�o`�g�بN�<�Y:�|m�>[m�f2-�"��ȅ5Mmx�`�����v�f��suյeN6�b����F��V}4�3��qtQ���r��Rnc���#t<íscr�˃m7b���G�5@<���*�ڜ��
e�.{T�k+�4��KUQ�-!f$�CC�&eh��W��������om�H�{ �N���rV��m��(�p����ir�[7�t����m�v�޺B� ,��J�Z �k���xYYU@V�)�y��D�/Uj9e�vT�# ��m:c6�p��:!6�� p�29'-���  -��n�h�z� Y���' -���AÜ�n��h����P,�t�K=m���U���[+j��P8$ �Ͷj��MU�����f������@Um)l����6-�$-��hII����  -�ܴ  l�I�8[d i	!&�3��T��U���6�8��c���)��}m[F�[m�� HH�mڪ�6�m��Ld��JImm���� ٴ�$KM���5]���4[h	 %�e��E�@��hܛl ѥ�5��n7k�,�PUV��P��Ɛ�UUl�� ��  �u��v�8�8ɮ` ��m���|�r�p@J�*�rD��X��Cn5Uԫ*�6�MT:�`:�cj�AmmMU�˦� � 'YD����  �v��ewmɪz�!��AĪ6���6U�� -� Eu��� R��m��`�����}��   d� 	6�����y�BT�eA.�u�m��ʹ���m��E9�m����&@�`�m8I�@�� <
��݁�kn+j�5vԨR�T�C�ʰ@U��B���-��vm�ڶ�` ۶m����K�.�`,4���
�S�*�;*��F�6e��Ԓ�6�`  ۭe����6���ﵲ0 [%�  M�m�h�m���
��P�VQ��^j�Tѳ -V�U=���88 T�UU�*�ʀ�
i�U�v^D��FE��u�8n�kȡÀ ��-��]��:iX [&���|-�E�nv�aӣfUv[�ٗ��X -���e�lh�e��m���    mm��m�Y��M��+kz���(r� ��		7ju�i6RJ��mH@�0����v�^���P ݮW6��I��� -��β��� �fT6 B��^�k�\�Pq۵R��neV�T˴A�#']���.�bR�iV�U��4�^�YM���i�4ڭ�(B�~�����4�Zhj�#a���,�����oҶ�U��[z��i�b^e�A�N2	����V̪e�2�@Uj�1^��� �J��1:NIY$ګ`���N�TK	(pʵ]We�yx
�(r�'�1+UW]]R�hŤ�:�n	���\�[�bO,Sv]�Z��[�U��C�9��wQ�U��<9�
��@�#"�m R�G�� *����v��
8�������� �ؖQ"Aa��fU\��� �l�[�� �<J�� �����X+��7ª�0
ps����V���o�i7|$ �K.8�`   ���(�����M� �km��   m  $:�V�nצ��m�l&ݤ��m��  m��%�h���j�m��ݒ<�t�O5U�J�R�5t��lmlvZ�hI�� e,��m3v��	N�-R� :�*����.��Q/�;T�9^|��W�L��.�k�l[Kl�D�����$ m*�[[l�5u�v�v���EJ�zBWc\���N8V�Ԯ���vM�Eyj펩��V��ŝ�ѭ�m�����>�� :K��h-�n�`6�� �5�{kd���m��ml� �     ��   6�6�@�a��Hphl$�����I9Yyj�T�PT m��8  3�
��Y���kj� ѶŴp[xl� �` 8v��  l    � q�o8qm*��e봋@�Ů
2�m�m��l	�  $m�`p�> 	B@v�lm�� ��.�\[E�HImͶ ��k,3m�m�m���WB�:U��jCk�r��-@ ��`  h��"e�p�M��� r�[dm��m�һq�D��ہ���$lpo�2ϥ��oP��jU�X%]���uU�UUUΉv%�PB�^k��H�k6ѺR0��l�l�h�Ã�߾�� �` �H-�H   �` 6�m�   �|   �$ 8       � 8� 8�m  �   �`[@-��� ��    �@	�   h          H [@       -�t��m-���p��J)[m� �`��6�j��U��%��]�n	 ��bC��	-��i$���H m�@ k�o���	�m��[@�/ZHkm& -��ZlH ��v 6� $ :k�ZXa��[M�� ��� �� � [x9m$m��`� $ ���l ���H/[���(�nYu��D�U��@wD��UUV�	��( x� ��6�  �� �� m�m�ObG  �͖)mm����� $�p $     �a�     H� *j�m6:Z�U�����W%��Gmjܶ�Kh $p    �l  8  ����       6�    H   [g�n
�����c �̮2m�m� $� ���     �UU+
^1���!ض��m��ʴ�oc�m7+J�BD�P.��-�   �� ��6����m�l�@ |-��m��            �l    ��    �         ��           6� m�	    � � p[@� � -�� �gm������b۠6�mcQ;�΂�U�N�h��2-<�Ѷ�y�뫚�6��� �@p[@��/6l  [D� �  6�m � -�	 2�   [E�M����mkn��  ����N3P ʵ@��麪  H p  �۰  �3!�$����vԴ �VΈ �`;m�&� 8p��rD�*�W�_/�n�h�5�0�`5��m7k&��-�m���Be3�����PP#ӵ��d�  6�[k̀;M�ku�p8�%� $$����`�ޝ�	��� 6�m�`m�Zq��p$   4j�i�a   	'$kF� m�@��a��[K9̶ͮ  ;YT�oH�`��U��AěY��ڴ�lHH���-�H5U]@�� ���P$�k#YN��B�Y�]j�t���<�e�M=7�$KX�8���CLj��,睝�Z�
�	Z��3c(�;���j��j���)X ��\�@F���� h�gN�n���1Q��` ^tUMA����V�p�I�ƣ��S�U|K��XćM*偠 �ء{jR��љ7d����EQT��� >C��_ ��
!��#��z*(b���MV���z�C��Ӂ�x�"�]S�b�`�H�@#~R�.
0 � "�J���� �H���H�0X2# I $�1"�� � @H�|���] 0C��EAD}D�5f� �z'��<�5���N���FEP���(���A��)���=:��~U�,B ����*�F������p�!��*���Z�z��O����C�ʀ��@S�"��*���������I"�X��V+��]P��A�<DD�t�P��AA=�ECJ)
 ?��?z�'���/���
�����t� �Q@<���t��P�4PL�j�ǂ��Q

'�P��P�/UN�����tA���EtG��F��
w{n�wn��{���~�����
� 7K4�ĳI;Y}4�Ieݶ�l��)CZ�k�,�]9F!c]�"J�I-[��m�[m�$��-�؟k[��d�p�EL�ʁ/[]�],@gUt��஬����8�&��ѷ�wTv�'�y^̮��Y��yV��s&@T����v<q��8���t0X�ԥ˨n�i�����v�n�#��'*s��V�0*,P:ц�r�ԛ�4�9D�9�<ոEx��9
�-��@���J	0\�	n���k�Wmg(��4�-�9��m�:���E�!˂V�,�m�%�M3"��ɔ��/�9rQւ��*�5Zl�<��3���+��Ǌb��ݤ�ǂXw4��ѹ��N�hkX㦞�����P�Q�sU0l�5��n����
��5�r�홢��Y��^�r�Jڪ[z̾'"�	��4���K�C�[e{y�l�u��skq�m�:U�����VR�7m+1<W���n�V�S��]J�ڡ&�a����u+�B���a3ܚ��g�sZ���.훳m��rX9��j��ճ��n�va��Lu$!.Ke��v��=��wc6nB��!$�@=�=���i6����[v�D�`YR�',\�Ggr�ا(�� ʫčKQ�UU*ք�s�"@�vP�UT���T�[vz��M�(�#�h9�j�mu��펉SVq+�5�n0�nw'fP9\Ck��趐t�p!�ru9��9���9ۃ�z^P�K��!t�������v�6rG�e�X�B޼
ƶ�i,��m��R�� Xv�n�H@���m��[�À��=���@s���`.5�V
vW����z�)�1�eT٪�]٬�l��v�ݸ2��]��%�	4]�(��%��Y�Ĝ���n�-�['�;�=l��s�tqVB�S�"m���v[��ػ��ٮL�ƛ�ː�'�b�pA=D�
EP����pGUG�^�S�h�"��|乲�/3�Z���hR�$�X�=ٺ��W:�:�MGn.�q���v��3���v+��<���ݎ���vѹݮ��^x��ۧ�:3v{b^zVǥ�윬��L�����c���-+�:.�8��K���nT�э�cfԯU�:��H����hδf9�D7O�c���Ij���G;c%�	<�3is7sKf��ir�������۝�9A����>�x���|���������r���cm���'�-�s@=�p������s@3�NX�'�8�m�3@=����t	$�$�%A�]����V�빠}��A���r4�jI�}��(�� 3y�@�� >�qE�'�&�qhu���빠�f���B���Vl��r���-�t�S.n������7��@cmB_ӣ�}lx�<��R����H��(L��sb��9�5�T&�slr�M:J�5w���7��@c��ڄv����eӡ�T�v��f�D%
�*b��@O;����{��O}���{���ԊH��dN-�n��s@;����Z�UW�2)#u4�i�ٯK�Jd3w���]�`}��h{(g+��7$h���}�}F��(�� 3y�@7�.��K=8��<՚���S.z7�r�$v��l�U����c�iJ��s�sj��@�� c9Y�#J9�&�qhu��޷s@=�����6o�"b!$���SΜ�i�t�S.[V��Հ{3]�	B�Q1
aB�W� � j ��w��h��Q*�ԑ��$�4����ܠ3�P��mB;�L��J8�9$�=�j�>��h��������*dWēT�MSHM;s�h�lֻv6Xn���,�&.���F���{�'	�ԊH��dN/���߷4{��wu��v���Z��)#�7uWp��� ws�ms�6� �P�W��	4G ��4s�6tD$������j���Ł�b������i�9&��v��n���I�(��8��~�T�_������"��E#I�Z���l@���M�7�GU��f�{q�Ŏ�u����3v�`��8(dg�3�B�'��������6vbkT�7�� v��7>������7�&~MF�QF�RL��Y�}��h^���빫�#��fM�H�����P�P��� ws�~�i.r�ٻ�wv�nm�
!U_�}��������P����N���6���j��S����[גO;�xrI�QP �'���.�l՝��nv�m֨�����{\O��Z^��x����ۑd��gD�hb/:k"�`uޅג�����:����k�mvLn���#�me����2;Y�̏������%���5��wp�e�ID��`nr��j���{D�s�؍,dη.�i<YY.5��mt��D����A�6��h�,���@[-�U�K��:t����YnzE=����t��ŋ�\��6�R����Cv*��K�����6�Q�	4G�-����v��n��g�،���n9�$�@ަ����l@�� lob�n9�&�qh^����h{��=�ՠ�Z��8�Y���� v��7H���|� ;�U5�EN7&h{��>���6Ձ��mX�(Q9�u3R�M&+�jT��
�{vֱ�ȭ#2�/ION�ז7g�`�يH!(�$xܓ�=��Z׮����h{��>�Z�[p�E&۷6�I�}�|x@�D `�A��w��`������_D�$�<n��l�H�M����߷4��hVנ}z�hvx3����	4Ԑ�;y�e�H|� ;�P��&�"*�6US)�`zwv��IB(�o|���V��vn�i6ܪ66���\�.3���l�t�K5N��������׆�}IҤؙ��Hg�������@o6� os�ms���:��j��iE&h{��{�f���U�}�w4{�Ԋ(�i7 ���$�����|�����TC!DA�	+-��`f����0�,rE��BG��4s�hz���e4{���:���$�I�Šf�����j�ܠ;h����F$�lJ]�<)��'k��3�{VB�2�A]v��5qƢ��{���̛���E���@f�P����\��ڄ���h���jL�=�}�`}��V�͵|�DB�<�F��ʚ������j��OҀ�mB7����s@>���
AI�&�qh~����I(��w|���V��j��,P��D(�TDJ�ͧs`�k]T��鲦nn���B�}�s�F�OҀͷs@�,*�bCJbD�ȢO�,L��v3���=��z�V\W��m��[Uv{��HI(�ꦮ���� 2w� 3[P��繠}�V����7 �I��}V��	B������j���Ł�fڰ=����MH��ȔN-�[��{���{�f��v� ������8�q�p��v�����ܠ>�#菣7�� �Q,���	4G ����#5�O�{;�X�zX�"�If��w�Ɛ��h�u���h�+�������*�ә^FuE�8��#�hS>۱�k��SJ�zj��ޝ��N�kz���3e{��Ь]�n���ɅOD�7nI,��9��z�UusBy�`��(g���݁��k����y����a�9d���WE�����d��s���%^Bi�uA��kg��ϕ�f�r�Q:�'�)xVɃ�~�_G���_��9�GKىh�,n��\&�'[�#i�8�<�s��y:i�K�m������-�[��{���{�f�{<�Ǒ�'�$ێ-5��l@�����"#菢 �9����r(����h����DD)�����j���I�;U.��mp����9u�@���h\^�w4���آ`ېq�rM��j��	%���|gu� �f���g��/�,ឝ>Ԕ\�Nnx��	X��6���\�nIW�˻��{�ح�vh�]w6U] 3�P��mB ��hv�>���PqIi�ܙ�wu��Ǚ�D`	P�`x�=�o$�����u���RYkDnH$�Rf�n�ηH�#����mBu�R#6DU:l���M�LI��ڸ_D�,K�{�S�,K������yı,K�݉Ȗ%�b_v��M�sn�ۙwws��Kİw�59ı,>������%�bX���v'"X�%��?w���%�bX�	߼�7 ��b�%\����PY��j��oC]�㡷����*@q�%3���wMO"X�%��}���%�bX����ND�,K���x �D�,K��ND�,K�Y=�훗v��˗st�yı,K��v'"X�%�|�{�O"X�%�����"X��ȝ�~�q<�bX�'�K�frm�.fn��77v'"X�%�|�{�O"X�%��{�S�,j�m2D�E�d )���D �i��c"A�!# ��21$bf��Cw�SF���!�1!	��"�H�E+A�!(P�� !4���,�`�!��@�@H$�! B1c�%X�д�A�0	0�K$I�őH�A FH�D��@�����c�(�"�X���c"G"U�$RF!�+D�� � E�0"�c�$X0��I �@�d�H Ad_�3��Le�e�,�<���E1J A$	"�" B�JF�����Ȫ�����O���> ��xfIRV��̶a)H@�@���/8
�5��DT��� >�⁁����SJ=W�����tL@N�3��3�*����O����	�&D�,K����<ʙ���~�.�M˻�7inn�<�bY�VA��xjr%�bX��~��|(���D�,K�~݉Ȗx(�Uh�$U�?}����%�bX7�;�ԙ7wwr�|*���O"X�%����'��U�DȖ�G;�۱<�c� C"dK���'�,K���p��V>DȖ%��*{�����Y��.��he�K��2���:�Gn�UVsғ���]���~��.�/'2ܓs7v\���T!�2%���݉Ȗ%�a����o�Kİ~��4?���&� dL���xq<�bX��D鰟�?��T�sSC)�B����$)�w;��?�5؛������"X���ș����yı,K�~݇ʢ�ȑZ.bdK�'m�g�6\ۻ��n�n�<�bY�DA��xjr%�bXx �G��ߎ'�?�"_���ND��@BDȞ�}�O"X�%�{��av��3sve�QD�g8jyĳ���=��O!�P�DȖ%��br%�bY�?}����İ*��'F"�E�W�ϟ��=�jr'���S"X�z�����]�˷.]��'�,K���,ϻ��O"X�%�UC����8(��$�}ߴ�$C�,�=���|��۽ߣ�}~ؐ25�W�\�aD{x:s���+p�f��YK[��2|��ffm۴���>���ș��wﳉ�Kİ�,�����,K�����?Dɉ"dK�~݉Ȗ%�b{��r�3͛�wnnߑ���x��X�%��~��}�Aʙ߾��'�,KĿw�� �șı;����yı���9��d/�����3s7MND�,K�w�����?�9"X����؜�cP_)bd�����g�Kİ~��59�Qʙľ���$��ݗ2���yı,�3���Ȗ%�bw;����%���C"d��ND�,&D�����
��L�bX��	�ϭ���ݙrl�݉Ȗ%�(2'w�}�O"X�%��~��TȖ%���}�Ȗ%���=��؜�bX�'��������gd�O$��sf]n�U��7�r�R۵�#��rtdӷkr�7;��h4������{X�5��a�ݗVv�]�g�`�n��s��l�wY�vKDm`չ�\�l�<ՠ����B��m��<v�:{Y���ñ��6Fk���)6�Z��dH79�����jm�SVS�����>?%`�x갤P��<�.J�%�g����.c�w�}?6;����:�67X�ѡ��(J`�r�-�V�[@U����sn�9�a��J������{���������Kı?{��O��L�bX�߾݁�I"X��Ȟ��8�D�,K����v��3sve���S�,K���{���%�bX��{��*dK��=����%�bX=��59ı,O�����n��ܻr���C"dK��۱9ı,Os���O��S"X�{�ND�,f���W����$.\���說r��3wbr?*ș��=����%�bX=��5>�D�,K�߾�'�,K��-�����ND�,K���g��IP�e�����7���{w;���ND�,K��﷉�dKľ���ND�,K���gȖ%�ow���cy�b��Jc���g�$�x�)@S�۴�T��#y�m9L_knji���S�,Kľ~�w��Kı/��v'"X�%��?{��yı,#3m8VB������5��ET�ɪ33w��Kı/��v'!� ��TO�\P^DȖ's�~�'�,K��p��Kı/�����'�`�Ȗ'�B}3�i377ff���9ı,N��8�D�,K���Ȗ<B"_��w��Kı/��v'"X�%��;&tٙ�wm�����yı,}�ND�,K��{�O"X�%�{�؜�bX�%���x�D�,K��i�wfٛ��-ۺjr%�bX��{��yı,K�{��,K����É�Kİ}�xjr%�bX���0���[0��9�]s���nR:�B=�f[v�s[�Bh777��x�0T����������b_{�؜�bX�%����Ȗ%�`�����Kı/����yı)���˝|ۢ�USn\�M��)!X�%����O"X�%��{�S�,Kľ~�w��Kı/{�؜�b]�7�������夨h�k��{��"X=�xjr%�bX�����<�cPu} �?'��2%�����Kı/��w��Kı,��q�����ܹ���jr%�d�|���Ȗ%�b^���9ı,K����'�,K��{�S�,K���'{s˻&fn칆fn�<�bX�%�{��,K��{�~�'�%�`���59ı,K���x�D�,K�w��ff�Jri݄j��rnj�ϱ���m��Z�v��gm��t�[zl��r�}ı,K����'�,K��{�S�,Kľ~�w��Kı/{�؜�bX�%���:l�ۻ��nn��<�bX�{���#bX�%���x�D�,K��wjr%�bX��{��yı,����7d�77f[�t��Kı/�����%�bX���ݩȖ%�b_}�w��Kİ{���bX�'��IgN�ܻ�n�\�7x�D�,K��;�9ı,K���<�bX��{�S�,K�A�R 0AC�&r'7��'�,K�w����_�\*����������D����Ȗ%�a�{�S�,KĿ���Ȗ%�b_��v�"X�%����Nv̦��f�م�.f���gNwge���u�e�W$�dL޺�ṣ̘�7wnn�s7x�D�,K���Ȗ%�b_?w���%�bX���r'"X�%��?{��yı,K=�ْ�Cwv������S�,Kľ~�w��Kı;���ND�,K�~����%�bX=�xjr$�,K��{���&e��nm���'�,K��w��9ı,Os��8�D�����{�S�,KĿ���Ȗ%�bw݌�;m&f����ww"r%�bX���q<�bX�{���bX�%���x�D�,K���D�Kı<��m�gM��wv�˻��O"X�%�����"X�%�w��'�,K��w��9ı,Os��8�D�,K���˙������q�fCusu�����2v&�Zg/B۞;3��,��m�8"L�{(���E�s�fCnn6�F�ϋ�`r��We�q��&ˋ�q�xH�#��7gV���ւ�u@��0��y�����1mmV66x�&�N���{$Z�\j��>l����rE�n7I6� pHPm�˦��[8���J�.����눙�KM�9P�&���K	aR�%��wY�	m�fDqn&����:hࡑ����&چȥ�,�&���2ݻ��"X�%�|�﷉�Kı;���ND�,K�����@o�%�`���59Ĥ)!eb	�9�����uM�/�RB��'s�܉Ȗ%�b~���8�D�,K��ND�,K����'�,K=��}��G�p��GSG����d�?g�{�O"X�%����Ȗ%�b_?w���%�bX���r'"X�*H_/n�2W�u-���N��)!I�2�}�Ȗ%�b_~���yı,N�{��,K"��=�{���{��7���~���}۪�E��ND�,K��{�O"X�%���w"r%�bX���q<�bX�{���bX�%���Iݲ�wvn��6�i�� �������,�<��#q��-��E�;�[n�2��6�f�Ȗ%�bw;�Ȝ�bX�%��{�O"X�%�����"X�%�}���Ȗ%�b~��e��i377ff���,K��=����
��tǑ9��y�S�,K��=���yı,K��v'"E�,K��v�^�ٙ�wm̻����%�bX=�xjr%�bX����x�D��"_��v'"X�%��{����%�bX7���3.�L�ݙn��S�,KĿ�w���%�bX����ND�,K�~�s��K�r��ww�²���$/V �����ɻ���n�<�bX�%�{��,K������yı,��59ı,K��{�O"X�%�}���d��*uq���ɹ:rsp����ᶍ�r�v⽻U���=;��{��9;,��݂{�ı,�{���q?D�,K���19ı,K��{�O"X�%�{���7���{����}�c���h l�yı,��59��DȖ'��ﳉ�Kı/�}��,K�����q<�bX�%���R�Cwv������S�,Kľ~�w��Kı/{�؜�c�:�Qpț��<�'�,K���xbr%�bX����nywI�wv\̙��O"X�P�"^���9ı,O����Ȗ%�`���Ȗ%�by����yı,K�[3(�t�ULm����$)!~���8�D�,K��ND�,K��{�O"X�%�{����Kı<���4Q瓔;cs㮇��n*s+����0�⡚�<u�\�	�'2r�N��.An�ww8�D�,K���Ȗ%�b_��w��Kı/{�؜�bX�'��{�O"X�%�{헳2�t��ٖ��59ı,K����<�P#"X�%�{��,K��=�s��Kİ{����Kı/����w&��.�73w��Kı/{�؜�bX�'���s��Kı;;���bX�%����'�,K���ə�3f[��n᛻�9ı,O����'�,K��{�S�,KĿ�w���%�`| ���؛�}��,K���~����wv��nnq<�bX�{���bX�8�g����?D�,K��۱9ı,O����'�,K��������L��Lnƛ�Lq�k��	G<�u�e����U�j�E�[uQH�f�Ȗ%�b_߻��yı,K��v'"X�%��?w���I�&D�$Q�֜+!I
HRB��U��*��\˙�q<�bX�%�{����DȖ'���gȖ%�`���59ı,O߻�'�,KĿ�;&ge��t�ULm����$)!z��W��bX=�xjr%���$L��߾��yı,K��n��Kı;�d;mΛ.l��s.��q<�bX�{���bX�'���'�,KĽ�wbr%�bX���{�O"X�%�{헳2�3sve�wMND�,K���Ȗ%�a�
!��byı,K��x�D�,K��ND�,K	��� �!#P��$T��#_�� 8p>�XA7��Fi� ���s��# H1BzEL�D�"�#"�)�� "d��L�8����ĀFA�ŅNi�j�X,2 Ȑ�"BD""	�"�*H��?!����T�E�H�@$#-*�ς,D�AS`�+,��V(�=!@�����	�|�
���������6�m� .��ʝ���$�i�Uٹ�T%.,;M4���n)D��M�;tƺeӤ�n-ju �ċ^z�y�C�5n�y����QTIv���.Ka�m���]*�0HF��Ʃ1�gl��m�뎶����Ҏ낲�rg����Y�Ǉ�Db�����<4�r<������ȩ�͍�1���s�@�69�]����O��-�M���,\���m�%U�`6e�c'�;>��V�&[!e��-C� 0��a�m�W,a�0���='�[�E��Թ�]�L�j��*�b�eD���л0ԭ�4a� t��Xͣ���]�:a0v3�p�Bm�:i�T��;�����L���v��t
�L�\�Y[SW:��zl,�eks��a�ʥ�[,���e�^�T�MH	N�T��$4c>��;��˼���i���c��g��L]��ug���p�Z7\mм��Q�CA�����'f܃&�[4��U��#���'i��K��:�hpF��ɣX��V��	5�Û*=v]�-4��8Ӭ�Z�j�7�_��t�lz�x���V�a�G�]"ʲ���9�3Ȑ]��ǂ��+���v۰��Ŷ/T�vLV���Y�̮���
�J9��uu�[v��(d� cMj,$�Ŷ@�rl$q�m$������F��;e؍M�Y@7WI� ���B�-'F�֓����Z��]�;^+�P�4�[j�4cPMJ�Ç.�m:t���G[5�%�*k,�l����m�j� �im���]pIs�A-mRd���9��,�S��p$@��l�0�z���Tn���f����A֋�%f����j�ƅ۶cL�g��J�Z����p��+p��n���<��p�*8�=[��]@Dd*;[���#�mʖn�krNq*�mƍ�89myݤ�gq�/&����h��;.��6��e7	%�@��� L(	��(銼Ӈ� E�W�~� \�M!oh�{D�F0ut��b�_�m�����d�D�v���9�3Wg�ps�n��g)u'n�m1^���q�h:U����,�=,�c�mѰ�]1�[���]���sH7T�;MS j#��]��v��\��E�s�F4Pm�?4�ݭ�i�u�G�����Y�ʛ:Y'��K��Xg���8�FX��v4qŶF����嗃��ɩ�E�N��"u��8u�����:+e���ی�m��[Uv{���:ٺf�m�=O�,KĽ�۱9ı,K����'�,K��{�C��DȖ%�{����%�bX���ۙ�.nMܳ77br%�bX���{�O!�)�dL�`���59ı,O����Ȗ%�b^���9ı,O���7m˻�7i���O"X�%�����"X�%�w��'�,KĽ�wbr%�bX��{��yı,K=��2�ɻ�wr�nf�Ȗ%�b_��w��Kı/{�؜�bX�%���x�D�,K��ND�,K����ٺL˻�ܖ��Ȗ%�b^���9ı,*F{�{�O"X�%�����"X�%�w��'�,K���w�Qkp��s͐D�a�t�]\5ew@5U���Vӫ����#*�Y����r%�bX��{��yı,��59ı,K����>'�ı/w6B����$,���I�L�cnf�sww��Kİ{����>E��n�Q�P^
c�KĽ��oȖ%�b_��v'"X�%�}���'�>r�D�oݲ�e�6��ݙn��S�,Kľ�����%�bX����ND��$K��{�O"X�%���Ӆd)!I
H^���1���f�kw��Kı/{�؜�bX�%���x�D�,K��ND�,�fEVws�_��$)!r�u[�����ܹɛ��9ı,K���<�bX�{���bX�%���x�D�,K��݉Ȗ%�b~��g!
�fJYr^:ɀ�hљc����N�3rv&�n#���9��P�hk��{��7����ND�,K��{�O"X�%�{����Kı/�����%�bX����zd�ݻ�sm�59ı,K����<�bX�%�{��,Kľ���Ȗ%�`���Ȗ%�b~=���=Yl
�{�7���{��>���9ı,K���<�cP�+��C"l����"X�%�}���Ȗ%�b~��3�s	���30�͉Ȗ%�b_}�w��Kİ{����Kı/����yİ"��{�	B�tڙ���lm̕M�ݨ@$���lE����w�ؖ%�bw��D�Kı/���x�D�,K��_C�u�b�3��.�j���*P�L�@�e��m�5=�7������3Y
�bX�%��{�O"X�%���9�,KĿ�{��yı,��59ı,O2�.w&��.�˹���%�bX��s�9ı,O߻�'�,K���xbr%�bX�����<�bX�'N����\����r�͉Ȗ%�b~��|8�D�,K���Ȗ%�b_?w���%�bX��s�9ı,N�t�|ͳ.��ݴٛ�Ȗ%��ȟO����Kı/�~�x�D�,K��r'"X��z�?�"w��Ӊ�Kı,���S�6���˓ni�Ȗ%�b_?w���%�bX}��byı,O}��O"X�%������Kı/���˙�k��ל�5zoh�r��δ�Ӧ��*�V�<��f�nu?)�ȳ`r����oq��%�~��؜�bX�'���É�Kı;;�$�bX�%��{�O"]�7������~�x�������,K��{���%�bX���ND�,K����'�,KĽ�wbr'�TȖ'��}�����ݶfffi��%�bX�O��Ȗ%�b_?w���%��2&D�}��ND�,K�{��Ȗ%�`��e;�4�3sveܻ�'"X�%�|���Ȗ%�b^���9ı,O߽�Ȗ%��2'��2���$)!z��ms(m��*i�7i�Kı/{�؜�bX�O���É�%�bX�O��Ȗ%�b_?w���%�bX�ʿ �Fz,�T��� �y�g�6GI���e�:�Gks�W["6��=$�*Mv�\IڳOA�۞]�ڌ��5�]M�qI4�Y�'�4j�O�;����$�6˼XJ�Ƌ��p��^:�}���Y�a��{]��'N�r[b%-'i�7E�$�:�kt�mՅ�;BfCrv{i��!mʠ\��V�@�Ig�hPzśv�q��"(�sB�.Rҗ8�z�����ǽ��c��(��@.��6�n�x��\���x�R:m����jLR��qٓ�"ff�ݹ�sr'�,K��?���É�Kı;;���bX�%��{��O��'"X�'�nD�Kı?���y�f]ݹ�i�7N'�,K���xbr� G"dK��﷉�Kı>Ͼ܉Ȗ%�b~��|8�D���,K;K�d�ͻ�sr�ۚbr%�bX���}�O"X�%���w"r%���4�2'���'�,K��}�Noq������޾���p�9Z���%�g�2'��ۑ9ı,O}��O"X�%������K��Fa
������$)!I
r8�je�4鲳�܉Ȗ%�b{�{���%�bX/�	_������ı,K�����yı,N�{��,K���igɅ��3���Nky5L�����fm�\��l7��m�Ք��{��@�εZ�ʫ'�%�b}>��'"X�%�w��'�,K��w��>|T,��,K���'�,K���m>˚M3sveܻ�'"X�%�w��'��>+�6%��}��ND�,K���Ȗ%�bvw�19���M�bw���.n-���'�,KĿ}��S�,K����É�K�!�2'��br%�bX����'�,K7��}�?t�+Q
L�w��7�������~���yı,O�����,K���{���%�`|"g{�mND�,K��%>�vܻ�sv�fn�O"X�%��w�19ı,?�+�߾���ı,K���S�,K�����q<�bX�'C���ZfI7%�YEC$�x"o<���"�vY�����o=)�G���yc����֨dt7>���7���'�~�É�Kı;���ND�,K��{���I�&D�,O��p��Kı/�e�3>�n[�se�n���%�bX���r'!���؛��~���yı,O�����,K�����O�*dK��e�KK���30��"r%�bX���xq<�bX�'g{��,�#��@_�(a"y����8�D�,K����'"X�%����e�wf��.f\Ӊ�Kϕ��>�}�Ȗ%�b{���q<�bX�'{���,K�?��￿�8�D7���w��`��3Y4�ϻ��,K�{��'�,K����g�O"X�%�{߾�'�,K��;���bX�'�gl-��	�t³2�l�#ǫ��b�J�;2�Q�l�Y��&�V<�A8n�wt��l�6q<�bX�'��8D�Kı/�����%�bX��{���DȖ%���s���%�bX��WUUESn\�h�d)!I
HS���'��C�&D�=�}��,K�����yı,O}�p�ȟ( �L�b~��S�7m���wm&���yı,Og�p��Kı?w���y��HdL����"r%�bX�����yı,K;K�d雹���rm�19ĳ�O� hlO{�����%�bX�}��"r%�bX���{�O"X��pX
u=�Ty�'��Θ��bX�%��/s3��nnf��n���%�bX��{��,K����'�,K��;���bX�'���'�,K���;ff��<�מ����r���8���Y���n��]�dW��ʁx�]�iw77ff���<�bX�%����O"X�%��w�19ı,O?w��	�&D�,K����d)!I
H^���&:cnd�ow��Kı?N��'!�ș����xq<�bX�%�~݉Ȗ%�b���w�(��D)n��(����fY���'"X�%��߾��yı,K�݉Ȗ?�4؛��oȖ%�bvp��Kı;��ne��m��weٙ�Ȗ%�02&w�n��Kı/����yı,Oӽ�Ȗ%�by����yı,O�:K�s30��ͻM�݉Ȗ%�b_߽��<�bX�1�}��'�,K����xq<�bX�%�����Kı4�o{�����������@&ԋ\˴�f���S�X�a.�a���u݃�ױ�Y��9IFt��h㓠�J�5.ǝ���Nض��N��-��mp�ӽ�GS���c��X�]es֐�o��~m9���`���q�r<)�[H�),��2/F
��lt7"�Ύ���u��Kh�b�ک!�B��ɎВ�g��-ƚnm��Y32�)r� �Uns��Yz�3����Vn!�����,4I��쵪q�f�Ͷ�����>����(�����Kı=���Ȗ%�by����yı,K�݁�șı/����yı,K>�|S>3s7s7.M��'"X�%����g�|+��,K�����D�,K������%�bX�Ͼ�Ȗ%�b_����ݛ�.m͙�n��yı,K�݉Ȗ%�b{�{���%��+��=�}��,K�����yı,K�����nn��7w7br%�g��@ȝ��~8�D�,K���19ı,O��;8�D�,��;߷br%�����S�\�鍹�h��j�|B�,K��xbr%�bX|�$}��O�,KĽ�۱9ı,O}�|8�D�,K����9�\ c���幃�i�l[��^�x(dg�70ɶ��r�I�M3sve���br%�bX����q<�bX�%�����Kı/�����Q	�&D�,Og�p��Kı?��L�e�7Mݖ�Ȗ%�b_}��NC����,K��x�D�,K���19ı,O?w�O"X�%�ӽ����.fݻM�݉Ȗ%�b_߽��<�bX�'�����Kı/����yı,K�݉Ȗ%�by�{-���7v��nn�<�bX�'�����Kı/����yı,K�݉Ȗ%�b_߽��<�bX�%��t�t͹�sr�ۚbr%�bX�g��8�D�,K��wbr%������w���ݵ`o�K�hsR%>��뇦�܃r�G�6jj���+�V�n�cW��o��;�1�VT*��o����@��w����@�'�L�ێA�G�.���]� ��h����%
d��I�ɕLmʙ��m��֬ۺ�B^H��D! I,H-H��aU"9�HI�8ŀD!"#�0� �$Y � �#�1"E��@�H��D�I$b��E!�D"`0J0�
A`��N���Y�Zd̙����x@�*1 �(E@"
�X�V��MUL8��@�W���*�W�N @�Oʀ���"�Ґ���Q� h����"�o���u�f9��4��:l�.���� n�h��h�� >���n�IɎD�Iɠ��@;3G`{۶��3���f��4�C~����s�J۬��ဴv�$��Y:���]�?�Xؓ�oqEI$���=��V��_%
�@��vn�ԕt��I"���n�}�f�{�� ��&�g�W;�7#q�D�h��v�n�:!%2fw���`XT�TXӊA���4�[4޴���j�E%���`Ѥ�*]:�*h���@����� f�h=l�--x�$X�cihY1�yd��Psv���L��#vC�v��2t�z���������@n�P�3[��ݠ���>�E�W0Y#�h�ɚ����ݠ��@n�P��ږ��j�9NǠ}�w4/Z=�빠|�k�.{�+�Sor5�L�<�iH�j�� f�h��WW@�H�JA��]� ��h޶hfh�3ud�T�!I-L�e�����iz��}���T��0;�	�6xxv�n՘��1rgڮ��6�CN�6��lLK���s��mȱA!q�<vLx�q��f]�t
���·\Z�=�q=�mӡړ���� Z�{k���سlv��D��:�x����{P$t�2S,	�܅غ����V��9��[�B*�@�faR����h�߾�w{���>>^����ܜY����5��&��Q�1��&[��mMgq�l]/'.9�����.j�@��z�kv�7[-��s@=�T�TXӊA��I4�[4u���� ;[P�#>d�L��[�i��&�{Գ@���h�w4�[4*��XA�I$�$�=��� �� n��\�������4F���n�}�f�{Գ@���h�",lM��&I#�)�&�0��4S�)��/�j���-��7g�vn���"H��z٠�,�=������\z�xېq�M ���~��(�)�BP����y�j��μ��l�/Z�=�0rE�Mw���55�@�� GlK���8�"s4..�r {�� �9�>��s@;)��,i� �mɚ�ݠlv��mB{����x)������x�o�ºΩ١3f.���F�!.y��W,h��)��f&ٕw������� 7��@��'��Y�$X�$L�@����;��h�l�z�hwe�L��4J�Ձ�ݵ`���I*P��!%)B��BD��d$�$���zBWf�9��֬=��
�IM������ n�h�7[P��繠{�M3[Xېq�rM ���u��l@����>���w�@c#kK��¬r=c��ve�u���n@���=W����i0��6�䓹��l@�� �c�b\NX29�2'3@�[����@=�k菤3;�X�&����r�US.�@�� �c��j�� ǿ���r9$�@>��@����=���6>�I��������&��$�$�=�w4w]� ������w��LrLX,D�om:'l�%
d�ԍ�[���17q-�7�جKr�3@�u��=�w4�K4z��؏a��c�$17�ݵ}�J&C3�vgu�=�j��ë��6�jL�z�h���z��޷s@��q���'"AT]�7[P��mBu�u����Ę�F�Qɠw���=붬��]�{ۮ��J#�	B�!-���w㦨<=�	��26
+u�B7\��֮�E7Y�9��g�:5�[�ɞ�vӓ@�<�X!���|���-���A�(Cmu�yr;�8{m=�	v��u�����T�f[��ۭ�� ����;m�=g%CQl�����-�\�;+b1�.�.55�vJ�y�X�aª�����-���N��[1m a������u���޻���v�_��G8��l�VN��t�6�:��6�r�Z\�y5�5�dN)�9����ۚ�R� ������S��+F�G����j�>�5��
"d3;����j�����>\+cX�RE�2D�4�n��� 7[P�1��;��	w�r�@�u��=�w4��z�[4��ؑ$�"X�Nf��mB%�� �n��� =�{��.�� �'Y펈�H�,�7�5���mhnuR`����u!���v����ݠ����Hw{��Ҧm�TԶ曙EP��=��}�Q
؈I!DD]�>�`n�Z�=>�j�/�P�I�H�i��޶h��:B���:�3��h�*��s�8�iI4�n���W��Y��f�V{�
�,Q� �M9���� n��s�kjG�k� ���m���gj��j�{�FQ���O-�a�j����VS�Xixb���:~ n������@d�:@c��1Y�c�A�#rhwY�}�w4�R� ��� ���$�� �Hܤkj-��3�����������nc�,�L�>V���]�ә�a�}��+��L�����4���Qt�������ڄKc�qh�Y��f1�Ș�f<J&��iJ�`+�e�h"�k���vy����6��%�\ 6{� 3[P��lt��� u1sMR,�� �mǠ}�w4��j���mX�ͫ�2t����*T�t쪩���ϼz��� 6{� 3y�h,�:�<N)"Ę�dz�빠zs6�{6Ն�bJ�d��\B؅
 �Po�˫=�AN�2��eIT�4���t�������ڄ> �s��]���ka루�㧖Ŭ�#�ve�c���X8˪�8��n�ЋGe6R7��Kc�o5��H�:��!��D�I3@�ZW�}�3j���m_(S'oJ�}5@�tۙ������(@l�:@n�P��v�/�qW$r4�nMًٟ���y�B%�� ��h��5,�ȜR��z�빠|�+���i'���I<]7���ЩX�����S�`��BHF%�#ju�"?F1
B� �!	#S �1�:�k�@�B��� �P���X��A�a"���-0 I�� ���P2h�f� D��`=N�����a��7�̷�����Ke���P���BN;d$R�(Ub�8��P�1V A��E0b�~��#�D@@��G� ��4����� s���4�/km�MW^v�u&L(�tp9�-u5�m�T���nl�OZ�	��(N���6`'�^6
6<�0U�Q@�2��r��\D<ʰT �Z�UF.�j������n�v���t��x��nڱ�\��'1De�'b�+��s��Ճ��{rl�ln4�v�l�P]����˭R���+b�0<�݉�%�T�%qۑ���P�	����qu�\�v�.�z�j�j�d ���rӛ�.�B�<�l!ù�c8�w<۶��7.���v:$\.�[ZZ�˰�S֠�rc э�:9�P���yM8T�M� �n[���'%����h�{v��څʜ��v^^¨[�k�rn���R�Ҽsݦ�]*��j�ɜK�n4Lظ����b���3�-W��v���,�lON�NrA�8\c9R���G]7'�li�a:�.�x�m8.�C�ix��Eѩ���-��9�m�V[�Y�t�y1<�-F�3�U���^t�Xz�h�GK�j`�iHi[8���c����#z9�uϝ��J#k-�]]g�� �Tڗ�3��Ʊ�8e%����1M�Tʚ��y8�E�Z�H/J�p,��*8�Wm���c�z1�%&�cA\s�`�N���-��@�la�׮
�/ 	f�,q&�m[BX�8*�Ҡ4���Pnð��W\���KP���T��[�n�YNc��X�NY��`m�`���:�sg�]����*���*8��v����<�#줡;@*Ԑ]7`�Hm�m[U���������Y+I`��I6$:�ŷ���l�	 M��	 q[R�*���@mu]R�*�m��r��&j��6Ɛ�S�M]q��)T�+Z�VX&�u��Q��]�B\�p����vv䗭��:��e��{ 5n\Z͜Wm�΍�t��x㋞��k���;�)8�;�t���kcFq���I��K�vIwwj���At�`{�pO�D8�u=DO�!����D������s3&�M���+�%�f�bBڹ	�W�v�ᖆ�dh��\�jvz�3�x��>y�1��Pl�0l��S�Y����8��`��R�y��	���ɺ1qv�qv�RW�[EtLvzN9M�M^���l��{n�9�̃���@�[W��*����7\nl8v��8;J녎%`�x�$�n (^�:A�\��
U�ug���Gfz�ܩr���8��v8��{�V��	�u��x�Sh�g�U\�ۯAY8���MM\ �e �v������B��2���$X�RH= ��f���t�������L���O\8��@��ߞ����hW�z������%$� �H�z����� 2w� 2u�@o@�ER�J�����j���t��Y�_����>�]� ��X��!B8�"m��]tvۍ[7on9a�L7ge�Rv-	&o]	��4�*�rG"Q)�|���/Z���s@�����.
ƣ�H�NF��߻���"�6���A��Ps�(@t�2�;Η���3�g�Y�A���@�_ۚ�uO@�{��z٠rV�b�9��s4��R'y� �n��� 2xd;�<nE�9�h/uz�u��빠wU4�����6/�X$C�OQE{,�\k�n'�mxxi1Bt�u��'\Z�U�a9�ԑ���4��s@>�T�K�NoU��Q�9��m����H�j>sh��H��H�-y�bs�d�f�}z��|����
 IBJC7����VٛH�ʩn�t��Sr�9D��z�7��{.�{�T���ě�H�NF������B ��6���t�p���aعe�uָ�J ��ز�q�0�������U�[�����u���-VT+�y�B ��V���t�7�����X��A���3@=�h/uv��v�͵�(Jd�Yҹ�4��ە3M�r�NoU���6��IL�oZ�~���>�b�N)�ԑ�O�j���mX�6���&#T+J!"�1]+��}��'�'�'{6���b���{��}z��|�k�>^��ׁQ0s��N1���nn���t���V�خq���v盶Y�D�$� ��S@�zנ|����]��ŊX��7�r)�|�k�P�d���Y�Q3��j����Հo��Jģ�H�NF��u�@���h^ꞁ���@=R�[t�"qH6җh�j;�i��� �n�@rV�b�9��s4��Ǡ~]����os�37mX#ab��	JII��X2[��V�j��=�'����F�e�[v؎��P���+����:K�&�<<=ck"��pnUث�g�O;nS9�j<������m��la�r�͢�@U���n×7d�@bVv��i��.�X��#s��z���3�4���X�v���m�m�
���Y���N V�#�#$ݧ@�ni�܅�34��Vټ�9�G{
=���w`��m�L�r�ƩL���P���s�,ܙ:^k�wl���`�I'>v�7��sjo:�OtI���H�nM �[4�w4��ɠ���`v)&9M'&��ڄN�G}���Ձ��������<lm��r��&�{����^��s@�qdt�E$�D��$��n�;ΐͨ@9�whꎩ&
>�4÷7�:�ͷr��O	n8���e�x�fn&��2����R,���W|�~����Ǻ���u�@�[���1�,�� �mǠ{�����0*�Y4u��>�f�򈈙�$��*]:l����O?]�7������ڄL;^9	��H�&I$���h/uz����u�@����f�RTՈ��(�� �;�� >������/q[��6�a6�#c�34�)
�Y�f�5cbos7 sɇj�5�����ڄ��v��v�N�Z�,=�I1ț�L�*�Y4uzXz�f��nھ�Q2v����-�ۙU2�v�zՁ��6��D5)(T�E�BT�؅
�k�VOf�`�Wn9#�7�4����u��*�Y4��s@=B�:E�8�m��@n�P�s�����@f�9@v�/�ٻ��&(Lc�7�����)�v�� mڹ��c�*F�z�r�v���d�f�-U\`�~�@f���\���B�j�rp�,I���z�Ϳ���V��� ���/�D}2k�^N)��s4�M�u��/�X���s@���arc�	���>�m�}Y����jÒ���LĨ�!B��z݁��R��2�T��m�6�� 3y�@��7��������\���6��g2rs�p��]�����g��s�{f��^	�������� ����B6�� ߮;"�9#�7�4�l�>�]��Vk��fھI%!�T��)�9l��*����k��=��������|ث��Q� �M����t�������y�!��z����E�8�$��빠|���w]�I;{��I>�����n>�	�c����f"Xx�A+�Ӹ�cA�����t��u��:ElC�WCN"�>܊t�C"��9���N�P�q۫v�[��I�[�S͔3���=��b�h
��'��f�4�V7I%��Ԑ)��B�]v�tga�s�F4Pm�Xun� �\my���v�G!�6�q�zH�6Z�rH�e�&msŮX��\i�]�����ۤ2�)�n]�廌��Sp���l��J��Z%
l���lW��2�cn%�<f�d�NGC�#��U���{��W�ɠ}�<�+�Lr!L�� 3��@yՠ2{� 2w� ;���=�92H)$� ������h{���u��>�e͎3"�I"MwV������Bw��ȉ�s�Z ���:mө�eS��fڰ=�w4���˭z*�yDC#�j�]�N�["c�v�h���6����L�f�G�ǤY�A$ܙ�o�� ��m�����2Cy�B ��>�T����.e�ӒI�}��*�$T?��6_�Ho��� 2_9������*f�tܻ��ڰ>�m�:!D�n��{������uf'#���RG�f�P��� c�6��DDL�{ր�Y:Nd��7$�M5`f�ڰ?D)�oK�{��{6Ձ�nR�s-:��xȦ/b�W3�&3L�7�>���hnuR`����!+�mMR��D�M����ݽ.�9�h�j�P���p��m�3S2ܻ ��w�?(��U��Ձ����s@>�T��G�ƛĜ��y�������9=[�!	*0+@<�G-ꓑ3�p�&�9��G�` �
����D�j��uG�� 5!C�"�\aL�dHڔ��.o<a>��<�?0�L�XZ"��@bET=|���T%�r[l B)��qB"���?h�'��~���C��-�C�~��
��r��[4��t��I7"���DB��{���n�>�m� �eĺ�b�9�M���U4IBJw���{7�X���jV}����8��kf�\���	�ۊ �[��5v�Z�c2i�e�I�s���m�7��6�{菢2@�?M�5\��cr8��4��s@�n�}���7u�(��=+%j�s%6�ܓpM\ ��9�ͻ@f�`b��UJj�M6�cmXrQ3�ޗ`����ٶ�-BJ��
Q�7����� z��!�sϸrI�ֆ�1�9$�&��M �l�>�]�����ꦁijZf8ю��-���+��5�ٛ��$�j
ъ���2���3t[$M�i3r|����:۹�^�h[f�^¦:E�q�)���@smB�D�o�����h�i_�%
d�"w�e�6T�t�V�~�@۴~�gy�B��P��|�H�H�'29����u��3wmXtDϻz]���L���t椤]U�7��6� |��6���<U��'�6e��&arl�m��
��ӭ��Qʴ�vK4�Ӈ�(�q�y�)���{lxz�	]a�L�԰D�ɍf�F�ݪx1��eή�p��)@�cRm�AewS�>t�U��Z� �]�2��Pe͒��c�&�۪��\��uW)4�pm:�۝`��N�GC�p�Ud��i,���ml�F�Ɇ,4�n��¶���㢶�Ώ�{��x� �<A���/�n���PM+֞�P�iٗ���h�:�H6������N��3\ѧb�0������ �ݠ3y�@w��q	̒$�4��M ��`{5�`n�ڿпU���n�4�m��2�Հ~���=����̥���������΢rFܑƓrh��{�������� ۴�P�K�M���5`n�ڰ?(�WoM|߿~��빠\�V��ڐX$��m��H�ΰn��e�ε��xsv��vx5rV��"j#q�4����z���4��s@��� ���98I$�m�X��G�K�QY�j���`|�T���.+�hxF��>�[V��9(Jd�oK���`}>'[�)�M��&������{������
!)�o|�ӹAWS� �I3@>�T�m���h۹����TM��Bc�"Iv�9���r�E����hv-@޺sG1p��-�s*�e�v���f�,��]	,��)��e?'m�i`ܚ� mB ��6�n׾�>���隞nT�t�-̶X�֬�͗e�$���&��3smX�j�*v)Ӧʚr�jâ�
gٽN�;�����h�Z�98I&�ۧ`����	(�����wwZ���N��P���d4GʥHH剹�J[Jp�<\b��3�ʬqRi����擣DF�����X�`��C�7'������[n�_us@-�hy�IW91Ȉ�SV���Jd;7��ws�>�m�ݖ��=��O$�4�������>��Vwu��l	�y$K�@-�h�w4��hw��Nd�u�6��9$�ܔ�n�횦�:�ESv�6Ձ�%�������@-�h��c*k�'�s�"m��`��x�3ˉN3�X�3��M�_>���lI�π��~���@:�4��;/�9��I�}��6� ���6�.�鐍p�*A��Ęۀm�{�@=�ۚ��4�	ubrܚ�]�3vՀo�]����`{��ꪦSiȈ�9�[w4����������X���DQ�cmᒑ�ݧ++�(��xA枞���F����N��!��sѝ�[�
��rn�wYv�C�W��Y�%��p�q��NyE�s�5�gHf�rl*9z��e���Nb27<ce��`um"���Q@%F6s<��ck�:��t�c��Ğ��Kfw8A���U���q
��Lv���9]\S[�%�ۛ��2�d��?	|���	���=]�W\v=�����������j����M���Oo縺��O�J醊� �~���@=��ڄ�v	��D��I4�٠_u��;7mX�5�(S'��Ӑ�s4�n�QUv��?(@w6� =�h[v�1fL��r�ӦɗM�V��
��~��ߝ�{w]��͵`�#Q�N�njj��� c�h[v����ڄ��{�)��D5B�@��.��Z�zyZ7)q�zY�+Y�g\��b�~����I$�r9'�/����޷s@�s@=�@��$gX!� �A�@��m\��(�7{�Xf�n�>��	�n�I�w[��{��[f�}�@��U�o�RdqG#V�$�s7��gw; �ۮ�Q&[��}�[�	`ۙ$K�4+k�?(J?(J+7���;�~�`�k��~���7יf��\l��6v=���J�q�S-g�[5B5.�wUrOG�iF�Ce� f�h�� �v��m� �s[���8��nM���������n�2{����v�ȜSKb�:l�����ٚ�N�՟�J1DB!DE
1�
��"�s3��֬�߭XJ�ֵN��r�i�۰6[t��mB��{��3jfH�d�麙��:�>�zX�DD%�DBK���/ ow�`zwv���S�T�hK�h�,8��qķ�n+i�5.͸Zدnz�Ąbpć��2,NC@�[����`zsv�!/�37�X܎�*���ӧ2�j�>���&L��3z�@�[��^3�ŉ`ۙ$KI4�n��� 7�P�3[�t�%IrIXǠ{�w4u�����I���9��ϳ�I��o{�0Q� �r9���� ���˭z��s@�ۇ�����,�Ӑ��YL�����έinW�e�����sWi���n^��9�rg��ߦ��ֽ�빠{���*�u��$�q�&������Հw{�ͨ@��YS0�㑤�F��=��� ��� �[4דu�I��"�h{舉��d �z�<� 7y�@kxU�<{�rcq)$� ����Z��m�ٻj���K�">��S0�a0��b<H��c�����8�5��< �*!@�I"$��b����(4�b�ӆs�)�s*j�Xm0� f�Rm��b�"D`DY� �`�8"C���O�B� ���ww6l��� �v�t�2��ݭvU��{$]�4Q�ٌ�ӌ;j�U��v��]uk}�D��$Hڕm�۰�@U+��gEJ�jz��T.eYvvv�j؞z���9�dÜ�kvRK,$�I�B�d�I˻n��艴�-�B5��������A�Ԟ�D
�5,��n�u\ܹ��=3һ[;ܪ�HRE�/Z@�Ų�����x�V{la���H��%(��55*vn���
qt��eƑ��mT�T�R�n��p��r�f�a��%�U�8����8���#�5�ɬ������i�:��զ����S5O]�K+�v�H�HVQyu�gD��iچ�q��AU�C��ei{��1eg�742�ƃ��ډJ0�z�^Lgg��V�Fj�>+h�&1��x4�uV��'iq��%v�`gB�[��L�ζ�����v�űml�\���U`7P;�gd�Q9[�s�b��7X�E`�s>�,,�Prc=Ėz�\���)j(�'9{S]*�N���)��u�S���4nP1B݌�+�T	����%���>-OA 4����Cvfm@T�K̨z����������U��]����u�Ѷ���y˺���4���q��j��{�e8 �������t�LE��l��s�Uy'��x /.�Gh	$[VЖ4�8���@iWWI�tC�戶����ٵ�Fp:�^-��)͸�ܻ�	=��VP'�[�pN�
�S�3���x��i�[UUUC���F3�V�T9�i!��i�k�.ʘ�ڤ�Ws���$�zD�o8m�$sm�� p���A!��W�Zj��]�X�g����l7����E�u��U�H(>ؠ"͍J���瞝���uQ�#��z�lb����hᎷF;r�#
��jJ�Cq���s����AB�A��hr��5� 㶺���p���n���W�ݛ���P)�*�_O@O�D�
�|����P8�D�pP�1��D ��~@S��@��CP_�\ /B�|��D��ی=��s�L�.���s�u��l9�`��"*u�r�wo&vu���<쵐S��f�.K8o=��*�9:X�3��xj71�6��{=��S9Q�Gb�5��]���rc�S;p�4�@����\�M�6�j�Km���՘v�)WW<^���BP���n��E��T��F�"r�m�6d���%ڴ�vi+�n�C���yp�s&�bv^�,[v�@�=c��R�����g��CQ�,�$#�bX6�I�rM��@�u��=m���Y�}�Ë�cm�i|U]�;y�@>mB ����� }�K�M�9����/[��^�@/[4�e4#/by�q�4�SmXr���v����m�
P�sw��*�x��$X���4��@�u��/[��^�@��*�p_�E�u��9��I9q��
m����49̸�XۉaLč!�q��o#rh�� �s_(Q������_
�$� � ߿��,���\ӂ�A�A�A�A��}��ȏ���K�d�lQ$B�!�@x�	����|��������x �}��|�������J\��ۚ\ۙ�� �`�`�`�}߷��A�A�A�A�wﷂ�A�A�A�A����pA�666?w�8 �����Ͷ�34��f]����lllo������lll~��xpA�666?}��|��������|�������77wsw7-ff� �`�`�`����Â�A�A�A�A��}��� � � � ߻߷��A�A�A�A�wﷂ�A�A�A�A�M���w��2H-u=��l�՗k+Y���5Zj�����Wf�l�۬e�f����A�666?w�8 ����x ��~�x ����|������fO���ݙrl��8 ����x ���}�|�������>A�����Â�A�A�A�A�=��p��nl��[�swx ���}�|�������� �b*� ��b����Â�A�A�A�A�{߷��A�A�A�A��߬��̙����l���|����
E ������ �`�`�`�������� � � � ߻߷��A�A�P���s����x �������]�3a�K�pA�666?}��|��������|�������>A����{�� �`�`�`��C���H��y1�ױj���Ɇ��d�\�w6⍦��7Y�0H��Y�����W|� �`�`�`�~�~�>A������o �`�`�`���}��� � � � ���xpA�666?w��d�JL��wm����� � � � ߾�����G�X�dr6?�������lll����8 ��{��A�666?�}~&y������k37x ����>A�����Â�A�A�A�A�{߷��A�A�A�A�}���� � � � ���Ϸ3����&�ӂ�A�A�A�A������lllo������P-���y'���	���=�{#(c�9�Y$���� �٠_[��[n�s��p+��S�nd���	��p܃up��uuA�c��ګq3s��x���-٫��}�ݠ��͵�;@f�OIC��t�L�eSv�v��P�S&�u� �o�m�{�hv!I�O�`��7vՀnf�:!)�{���֬ܪ��pI̎I3@/u��٠_[��w[��z�f���2H����� ��m�@��}�{�����Ս���텁��]�M�A�v�q6�+�+��8�
����mA�!��ɘ�lݕ�í v����}��Ǔ��]V�d�j����<@v��v�;S[������f�:`n^�(ks��'��9v���U�Ql�9K[Hݮ���a�̘�/��T�#�v�!�.�y�Z���CӣuV�R���WCF��[u�,�����q�\��Qۤ z�n��-{x��l��e�S���1^��X�ƦI$�GX��=߿nh��h�@� Ϗ,-cx��H���w[��������m_�'l�
�:l���mXn�@l�� ��ͨ@��\M�]BH�'�hu�@��s@�n�^�4��:�c�F�9����v����0���y�@gu���:䓍r��&�m�dfLu����ؗ��
6����&۫��8y�+��l7|�}��j�v�s���jØqQRp�曛37t�w�{��r`�"��N����j��ݵ`{pFѠ�m̒$8��*�^�}n�z�� ��h{q=rH܎4��@zڄ�� ����� ͙�m��8䉵��^�s@/u�]k�/���*�+j�$c�I��-��:�\�&J2��l�mSX�a&d)�v�dq� ���3@/u�.����h�w4�/*���RE�8ܑ�����m�@���>�ꉎI��F��;��h��h��,�tC��On}�rI>��o$�A�v$��'�@����� ��4]k�;��h�+x�5��1�*��@�����kj�P�>���_�u0ٸ-�T1��λn9a�u���4[Y�j��]N�����l�l*����[�P�;y�t:���q�i`7���M�/Y���h{� ߒ��bb�9"n)V ;y�@�� >n��؀ߚ���T�[d�&�V�L�o; ���I<���? =R(5@]��~� ���H�'�h�f����ͨ@����'*Ț<lh�R�n�n�#lۙ��2ڽD��Xݜu;���ۄ�G-0ᬵ���>�����h{�����ܒIؒs�NC@�n�w�� �l�>�)�wU[���'2H7$� �u� ��@c�b�j���W30UT�"D�M �l�>�)�^�s@;�f��\z�R7#�/�4�Jh���=��su��D(=���ጀ�ղEn��ؠ5#\O=iт�+GG=���v�v���wGc��7nQ�k�dnZ��.w<�O8�%ٺ�ɭ��mrn�.ugn��Z��^2���F�i��Z]����Ұs�'cp�6��<��8ܜ�+�dWN�`.����qƲ���J�K����뉎P�v:�9��;uok�������|�*�q՜+������w{�|�-���:)�7�\�����M��і�+�c#1�����K�7�8䉸�����ۚ��v����$�}!��Ł��S��8ԐI�$���@-�h^��-�s@=���	1H��	��[v����m�@�� h�f�ܱ�"brɠ}zS@��� �u�m�@�X�s�����@{�_?^ {���1�� v��\�g3���4':�G��Q�N�Y�CnuYM\f���xp��H�{�nhj�����h���ڄm�@f���)������7sw�I����
`�@�?GE� y;�yÒO;���~�� �VF����`ܚz���w4׬�m���¨lQ�$M����w4׬�m�z����;#(c�I�RI���h���n�m���T�ȱ��C�
[����ezyZ��䭹sm&Y�s�#�T�x9D��F��RM�k�;��h۹��f�{��H�nG��@�[��[n�z��Vנ���$��ɆA9���h��w���!�jAcB$�`�� ꚰa�j�#8euHRs8���$$d�2Hvʐ$!��I {���RA!���3�z���`˂��� Ŋ�B�)�����(@�� 5T�"0���F	� �C��@�qA�qPʪ����H�T�@�| � �C�(�|z#������&{6��7{�Tʩ����s4�`��@9m����P��pʚRL��D��Vנw���-�s@=���脡B�'���9̶��S�E;KKs�1�.��aL���l�Ի�U�CSn)�Ȑ7�^��s@��M ��h+k���h�أRH�\ ;�؀s�Kn�[P��2�ceq� �mHh�@�[^�}n��қ�=�y_�c�91��>�	D������Vf=,%%b��'}���'{���w737sn[�]���j�l@��%�H���o�[g����k=��f��NV%l�[�c�*n��mg��U�5s�!��M\ ;�؀s�Kn�[P��ݩS4M�M4ۙeS,s5�B�2z{����Vf=,��vJ-JSND��������wJhwY�^k�d$rG"@�z���wJh�@�[^�|e�Cm9m2'3@��M ��h+k�>��rI��	�R�g�}.lۆf�m�H�7�Y�1-$�,ђH��:,�3t0�4�:����<�����:��h9J���U�(H�FT���'Iewd��FW��uƧ��َ���f{s����4�X�ۤucr/t���Wgu�e�WEn�r����h�3p=j���ݞ�j����e(]nٹm�� X�;T��j�0���ݟ���сy��j�"]=�:�٩l���(����=�-P�d�)UKT-I�G;�ssZ��b粀�H�\��^#�������5$m� ��|��@��k����|X����mSn�)U1��-�@cmB������:c�+�F�q�dn=�n��Қ��h+k�/�<HN�G�90Ȝ�w[w;@d������T�qSM6�sT� ��v(^��wZ�77mXN�[��dmU6	�q���������LW'N���K�V!��s62c�72H��@��z����Қ��hqʱE�H�H�`}����+P�R�%�������|�נ�t�6����I��7�؀;��'��6� Q�R��8�i�ؕ���<���@�۹�^�s@�<9;����prD�n��P���b ��h��*��r���t�N-����6�&��p���q5��?��N~|KR�)�'T��=�֬�zXfk�D}!���?s�	7�2<�ɆD�h�����=;�Vۻj��(�;�~�EQ7T�ne:�Xw~vӛ�g舕	y%��Q	5
���V�=,{�U6�����N����ouX��V����h�9\q��rG"@�zֵ�}�� ~�Kn��ﾈu�����1��*�)�v�v���;YZ�FC�i��k�K���=rݑb�m(Ш�Wn� �v��m�j&^cT1��Lm�hwY������?�~�?~�j��ǥ���4�m�uUUݠ2[t��ڄ~������@o�r��H��G@�F���g�/ow����ŀ{3]�(�J�R�BR��?�N[����	7cJ(��dNf�����o׀l�ޤsj$o��}��s�x�b��̜iX��5:����K�i�.u�����?�����r���4]UY��Z%�Hm�@wu���¡���E�I4���[w4���@/�#QH�D������#��L�߭��z��4P��#m�s4{�4��h/Z������̱��r4L�e�{3]��G�;��=�֬~�{9$� y,�A�� H��F�~���[,�۴��2�$���K���r�%0�#��tqpogd;y4gd��G�6|�,�S�6�=o1�h������n�Fmfl�uG>�=�w"&��v+��`-����.�@`�T��W%FӜj��V'<��E��rj�	�,ms���P[��@'[�v�S���X#��`��Z#YNź��f�Y���\���&��S�qɬ��F��K,�b��؉�s�	�Յn��6�S�	d��$��%�vN��`l�~�����|f�9%�����y6A��q�F��>�w�艓�߄���:�/�6�"j���"ra�9��Қ��4��z�n�67�"s�(������9�=���ׄt8=����E�I4��z�n��t��{���QZѤ5�#Bcƣv�ţ�{x��[��8�&
c��61�r΍D㑹��>�w4{�4��~��yw��@<Z�����#M�s�l[��()�Zg��@g6���yP��	�I�h���>^����}�֬�|XHx�m7N��ST�Kn��%>����j��c��=�f�oLU���q�9#�@����=�)��@�u�@��B����4�.��|Z�n�;s�a�%�N�=4pS�V�6֓u_�����m�S�������wY�|�k��[2��X6�܍I�D�p�{�W����[��{�i|�L�i����nSm�ӽ�`}����
3�BP�BP�+w�;,7l�;�7��8(�nD��������M �u��ֽ ϻ�UarG3SW3w� ?}-�^���@cws@���U5B2'��l&G���X�gؓi����9nښ�V.�L���S�2R	17!��f���^���s@�t���
��G����h.�����j���ŀff��	B�2t�.�ȓ���hrG��߿nh���@�u�@���&ݐX㑋"�4?Nn�����7j��BP�I|DLB��Q�]�����
�j�t7S.�`�����j�l@7�v�p�M��1�+m��(��nyz4f�6Z��Z6��7g'��f���;�}!���j�l��d�����U�8(�nD����������?m�4��z�y�F��$Ӊ6�{�����
ϧ;���wZ�=���,q� �Ĝ��wu��ֽ�n���M�(W�r4�!�˭z����Қ��rI����3U�x��bDb��w<H��dRMV���C�R�<����?V$+��G�i�"�h$�+?$� 8��,	c4�E%J4�JJ$�����ӂ6�����l��v�2_Nc�HO&��X[�M�;m3ZL��)�-���ᴻs==�f���0"Ь� 0�F Db����X@�;���wwKm�� ���l����}n����k<H�e�V��K2��K��!d�.��V�i-[��B@�4�[�7P7F�5��`�I怊:��`�U�����"�á��y��uҨ6T-�vU1�F;b&؛zN�k�uu�i"���m�Fݮ�ͷb;A�7�ۜ����l6�*�u���N�U�uq��6/VgN�� �[`�F�j�5���VH��zS�55�[�C��Um�Vy�g�Id�T�$M��Y:m+�o��| �,ɦ�l[�g�뮧8���5�5�x�JӸ1�MU[g�5!M۝���5�yR6���	ҵ��s�sn�����A����0�R��qqn�w���o��+�!8�g%;���خ))��:�e����۬��.��JD�=�U�0�K`�����vM^�{�`��5���9Y� ��ps`�GvL��,a�ml�t�rE�B����<�n��!��4ܼ�WoS���8&�Cs� 6��tcq3�M!2�v���p��M��0õ\�/�>|m�s��q�5�.ـ�F��K�����j�Н����E�9l<R�UJ�gc3�d6�܄�l�/�G-Pm��9�γ�vպ�-��r�:Ѭ��\r�n9xR�r��Am�ջ 6�� ^],���m'i�e8���@U*��hȔ�(��f���@T
÷�u"������OG ;�+��k�P5�p�������;r��r�n��Ȳ��UT�U�:7KpU<�t�@HHm�Zgl۶B훒8�[T�It^����m~�72�p��v��۳� t�,;Y@� MT�R�3e�6���@��3�B��F(n"�Z�X)�W[��M�B�OlPLiV]�AKv�b5$�%dt)1c�l$d��x��K��v��vU��*;t�k�iu���b��X3���k�[&�2'%��rp�in'smwn�tew#K�3\��A*�!�SV<A��C�)~�����DN/���y��!I��3dۮ����)|rG4�ۅH2W�������v���-�!���gۓQj�X{a�i�Aq��o�6���] �YVq%��q��ewb#V�m�[���|a�pu��5#�%Μh��S���ʷ6�a�{kw$[K�ZWn`-���4����:�rm�iۍ��%^U��uh2�(�띛�,��s�H/	�Y���	6@~EP�s�<��6+e��wsf͹�q��^f���GM��.��S��,^�I�w��f��GCp�:w����{�S@;���ֽ��%òr1E$ 7�ؿ���G� ���6_�Hm�_�DB�3vz�����N���T� ��h�n�ͨ@ou��t2f�����M�ֽ�n���M�������g�m�4��s!T���ڄ^0��@d�t��sqX]��͆�M�ێI���K�#:��-�F[��7U@��q����7?6�K2�Q�sw� ws��ݠ1���#�6Y*�Kl��j�,35��"�QM]�d���o$��p��t���1#�8�����l�rh�z��P���b ��h���Y%7MӪ���nÒ��J����V�?ŀg�]��3��v�ӧ6�T�%QuW� �v�3��>jx�X@I��LX�?����ٸd�f�zƫrո�o�\��8yK��M]U�����������d�s�Ɓ�.��ő7#�����>j�l@���t��vL���s0U7`}���{�b��
" ��4�[4>���(�q�Ӊ]�߾���o��@~�h5�@c�@�"�*���	1'!��@>�#5�@c����6L�eT�����8:��0X�.��V�$Hn\�MyĹ�g;u:�~��w_�>�Hɱ�v�G䁽�Z5� �v�q:��A�$��G$�>�w7������ƀ^���}�� ��qd���I���� �v��D}2k���~P��:�����5��@;�f�}��I<���?�ET8�P>T.����s���(�.j�Ҫm�sv�����# ��� ��h\���-�Y�թ�٘��g�	X�ZxYN�v�Xa��u�9$�S..-���|� 7�؀;y� �n�7ESRF�j7&h��9{���٠}z�o��~��Px�A�&�y��sv���B{���':�87#����@>�f��빠{�S@��@��u��$����ݠ1�P���b�y� �n���}��~���&tK����{T���)eu�#u�R�n��k��Z6�;�] =a=�2e/�!�n��.z�&7Z�����8��s���G���?�2��96��n6gOmi���`[7<I=m�˓��M��\�ݹ�]�:U��h�Xkm�U��흞���Mp��r�P�2��[[ف����Fu�U��zr�!W���c�0�F;7e�-�3�+��I���lqb��$�J{f��z�l�5٢�6��lW�6X1Ӷ���!�-�6�����H9�@c���j��X��6�dn/uz�[4�]�ُK�(��=�$�Sj\�:�M�`��@cmB{�����7�%��q9�/�4�]��Қ��4�hֱ�RF�j7&h�l@�� g7h|� 9u�(��N�/u����ռ3��:��צ�%�wV�<��֡�r�<�3Y-ó���������[GLs���M�u5T��v�n���B��(K�	OwZ�3u�`����l�tԕN�n�IN�vۻj��c�Έ�Q(�M ���hxY[�A�A��w޶ �v�;y�5�i��q�I�D��4��h��h^��޲�����<&9ɍڃ��;'=�\3v���s�m��uG`��\!4�ɉ��$x�@=�@�۹�}�zX{5�$�d�:FO0sM�73��ݠ7���؀;�� ��h��t�E����ɚ޲����'A�y��(Ow��;��hsX��x��A�����v�7y�5�l@�rcr9mĤ��u�׮�����w���I܈�"DLl�H`J�-����3k��p�X{�q-�����A7$�6�XG&��빠}�)��@=�@�ʻd8�n73@�v�N������@f�%���rH�dn/uz�u�׮�������
��n&ۈ��H���vۻj����a��$	'�� ���"x"'~߳�O>�]�w��ȗ�RM��s@������^�{����F��ȓ��L�GpKv�p��k]�,�Xl�\�磩���]^ɨ��D�Rf��v���� ��4�]��gex�f(�i�8���H���1�P��M��L���{�܎F�dR= ���׮��v������g�MI$��K��1�P��v�N�������m�qc�A��s4z�h����uwM���ڰ<�D(X��5@�5%
k�.�g�"=X(���v�62�]���KD����vCpT�Zz��{�
��.�=����5c5d���d]`ܳhP\f���
�/P�4z�,��m�k::��v��5���2�Na�.����Y�����Xp����%��7��k3��l�:�d�(\F�f�d��$(6�gb��gd��N+�7&�M45�˯��w��-��(�,3!��v�7%,�.ff�9Cl��7��y�#��Gj�ۆ�)��M�äA�"���<�_�@���@����f|����h��6�q6�D��G�n�r���Bu�;Η�d����QG�dJE�{����{�S@��@���@>-�g��H�N%&h�؀��t�ݦ����D��F�1G�MŠr�W�w>�@����>�ՠ,��G!XLq���XB�v.�<�Vn\�l���׶N2t�u�L3�ؗ�L�cr9m�H�������>����s�;�]�?�jI$m���������FE�7&�=�@=�f��}V�[ͱ�\X�j��뜠�v��r���B�Q
����Ei��w�������s@��V��p�mc�n!ʊ��@wW9@{|���o�ޔ��ѷ�ߧS��Wv/O\���%�78^���G6K��:�He����1:S��ZZ��@c���������� x�\��9)���9�Ձ�k��3ٮ���vl�6��P�M�J��b��M�5U-����z�f��JD��L
 ����^pL9���$kB��T�X��#'	���	�S�N.�H�9\p�$d���7�)��;���y;�.��û.�@��!��O9�W֜ �p�-c@b�⟨� P��"B@ �!bEہ!q�s��.���0�0����"@��D_��D�Q�Pt] h��/��"�|0�(��P	�� |E�s���?�,�{��`�gIԦi�u5T2[v��9��lv���ץ�(Jgsy��른uR�m�JS��͵`~P�g_ ^����;V��������4�6���e㮸ݡ��Rf��y�cGM�[F�a�mFl��cq��� �q���e4��h�h^��ױ
���rH�n9,@���M�5�l^���֤�#�n!ǍI4����>�w4z�h{��R����'"r)s-́��ڰ>��,=��?DBS��Z��U�g���8���r��j����`rJ"w7��fWt�nm���G}0:�I�M��N��5�x6�F�`�hYxo�mM`�c3VP��sI��dT�0���7i�@c��!�������)N���T�[v�۵��
d�oZ�39�`��`g���j�Tے6�QǠ}z�h����Y�yzנ}�a��x�i���޲���v�۵a�!%�D(���������14�NLr
&��@���@�smX��,�>�]E:&�t���=�(dK<�Vճ��t1V����yΝ�gsL1����s����zi���~ip�|�Q��c�ju�ӣ���x+q�-Ӏ�wmq�y��<�:��*:��l�m1#.��8�tu���H�r�k���l�s�5̓��H��۵�+*��]P�r�n���2m&�!�L !4���b٬a��,P@m�Ӳ-���	v��w�G�B�����2̦��Mݺf̶��v��N��X\6Ѵ�4v����F,�n;69S��q�RO����@����=�)��@<URLw$ND�Q����ھJ!B�39�`�����v��W,�m�rH�q)3@����w��?∙���=�֬�v���S�M�5U7b ��h�n���A�������� ��1��r4�8��@���@��B7(���1��.����,: ���OK65��L���H��W���ȃ����Y��~~���}��v� �u�.����J�Ԙ�7f\��ӒO;��⟓稡SwĦ���J�'�$����|�^v�Kq��� ����]�g�$�'�=I%������r�RI}�*�7�	7���|�\�V�$��߳�K��-I$��ϾI/�,���c�$ND�Pr7�V��}���[o�+��ϥ��m�{����sߣ� �~���o�X�b�f�;\-O!�#:��/Nі�FK�#\ν`����'ۏ.Y��D�nL��K�9�Z�Iwu�|�\�T�$��߳�Ig��a[X�A���$���>�$����I/��g�$��zM�Q�%	�39�)ESm�U*��ym���ٜ���{�<��ĂD�) �P��<߹��'-��~�?����{���KUJ�S/����}�IwY�jI.}���Iy�[Ԓ_^�I�&8�n73�K���RS>��ݙ��z�L��6�3&fNw0}v��.;	ǌgV�m�\V褛��6����:�b�Ol(��5�b��\�����v��$����|�]�n�K��V1��I��#��K��ޥ38��̙��v�S33���3�EUIq�&-��9��I/~������pԒK޶}�I%m�RIy��T��H�j7&}�I[f�$��l��J�'-�G�H@���	�w�{��-��0?��8�i���RI/z���%�����M����L�����/�����h���̓~�����L�0:K�:y[�ƭ��j��:��<��m���]zlmأ�I+l��K޷��䒶����i%����� ~���7��4�Ե| ?_��;�K�����^���I.�o��"����F���M��ho�� ����[4z�����A���"Pnf����`d��X����D�;�V��By�$�c�"rh^���gw���o{��v�#�ᎆE�UZИ�ph�0"�O\�Z���]�Z���s˛���]V]�9�P�rk
.$8m�5n�y�vc���v��N��.��cN�/N	�vj�9�ڋ��z��Cn$�Svm��،��UP�Y"�{r����P�Bۈ���;8�U�1ª��S�6p�cn��]�+���*�?�|#�\Cg��"{A�*��S��2ܻfi��i���We��sK�/f�axYN�q��5.�'5�&�L�r)"Q'����nhz�V�n��QHd��X+6��MK�#�7�4�n�{���}V��nڿ�L�Š��K�M�5U-� ��v�ٵg舄�s;�X��V�d��ŃrH�nI�y{��=޷s@=�f�Wv;!��H�i�$��ڄ﷽� �������F����b��z�m���5ne�z�c�q�^17�$̓������B+���@��gy�u�}sF�Ni�M�Ӗڰ��z�8�@�1�M @?
��'o~�rI�~�s@���hw�O7����Mgy�j��g{�P�rߩ���=MB9�(��@�۹�}�w4]��^���^�?�dRGn7&hݱ������j�炙������ǮxSN����v�W*��p�Z��`�[V��sWb�#�q�[w��/U���� �����<� 1����{�b�q`ܒ6ۑ�4]k�>�w4[)��@>��f20�9ni�6ٻj������B���"&BT~P�R�J�]�����V���VZ�E&H�QI�����@�v��DB�ww����.h�e6���rۄ�����P�P���ﶽ����v�ج\Y��v�fum����n�-�m��u\�u�{��Ӹ��&���u�Ҁ�ڄo5���>��I�jH��dN-�n�����""d�~P�~�ms�L>�L��N���6���j�33]��(S��=�֬yh,�UJ]:l���mXt(_�J*���3k�M��nڰ� 1��V�
"/�/D�7��{����ؖ&㑦܍ɠ{��@����=�S@;�����p�`=:N*� �ƇG����٤'-´�ր�q-���ӡ�AY��oϿ~��=���fk�Q	}!�]�`b�ٞn�s$r(���e4��h�j�>�w4wb��d��I��h���7��@g6���B;��D��ӡ�M��9DB��=�=�֬��j��L��;��*f��cm�ne9��sj��� o�`,��@#�E�E�AQ_��AQZ"
��Ј*+�" ���B ���* �?����A@����������"
��"
��TW�D��TW��AQ_�E�D��TW��AQ_� ����(+$�k8�d`5�0
 ?��d��-;�                       �*��( 	HP(P(		*
�
�B���
T%R%	(( ��� )DX  4� @ U(SO��W6����e�e�����7�7���)�y�y���t��}��=n}O>�f}t���{� �w������� ���.T�}��w+�{�E�� ��ӓ��������۞ܩ�  �  � 
 AX��}�=w��T�ӓ�Nϼ
O�>���w�9wnqe�@n}>��v�     �P�}�� H tw` �   � �(;�� D @ 6`  �   %�� 0   �  �  m�   � � @��w6  �{ 3W'ӽ���w ��*ݞ�K�ܽ���Ez�Z���
}�rjLL���ەzr�7��(    ��,� }�}3�%Y��3+�r  E �  �};��������Ͼ�R����JW�=�/�g< j��>�u>�x w�W�w�,w.m����� ��qn��νzy=���� ��P��%@ R�� �VgvS���q�8�n�K�
{����;��]ŝU�����N�t�����>�M|Z�s{���>��}..s[���דӫ��U��Gz�Ynv�e��^.���}��m� ��=��*��db41T��45J�4��Ǫ�T�&�� Ob�Rm�L�O�BT��*U  ""I��)�@G�z��}�����������ܝ��������AEEz���
*+� (*�
*+��`TW�QQX���������4B�&�l��b˖��X�����i�������4�����X�R0Г�m 1V$X��[&&��䗎�E�d�] ���@�#\te�!CN0+�qXsN1䜼4���1�#$����d$,m!%��N.���I
`k)�.B����͟�Ց:��aC$(D����$M�<����ܞ�<auГ}}=�A��0HՉ H��I$	"Ԙ�J���=!BB4�d��!.��Y�2��&2��`E�%VHQ�X@�֌�b�(�H4ÇN��hq*h&�1�">��i�pN�,b��� W8�H�$
�[����u!	D��$� �A*!0���k�/:0
$i�����8� z�E�z����0,���j@��K��! 8F$�d�H�@�%H-m�4���!0����
D�n���p�х��H�Dp�� X���H&���4"��� �H��S�C��;���E�@���`�#�lS?BZ�Ȓ+R0�4�p#VB,��V�JU��H���H��$	%6g�Bx�Lp�!1�N�#H����@�XЁH�p�$$��
F+$,@7'8K k�!!p5��4��A�"A!LC0�HG��
��F�H1`@�R0���čXSXЀG@ A?,="	�g?~`�} �	�D�CbB0���4�@�c�!
`B��V�V$��!-��̧�DH��$�"'�����%pa	X% ������x���o��q!s&����0�́�S�y�E9 'H�q�'<�[�.3�ą`���_|�2��?z�bJ£�0�s�4}�O�`���~O����	pՙ��.x;q%��5�n��Ӂ��B�8��V!L�P(p�����)����,V	�'�� T�Ny�)�R��%.�ǌ0��ᤕ�L�Ӂȑ#\�r��]4�B�D��xB���� ͎S(�2X�i����ȴ�N�&�#m	&���8P��^0�'����ӏ8>n�<7@�$ܰ���)2�S)LX\	�d0�pa9�R�K�nB$.�+��������C�+�B�0��v�!! �'"D������X$%�-�a�%�1�)*0��8f��ˑ$����P4BB7t�$'s���w���L�+.���9�׌&���Je5�H+-��f�Д�J淌���`�W�����1�^x5�&�$#d1�)V V�-%�k
`�cW�ZNq�s�/)���n��L�$qH1�GЍfm��sf^��xB?aH��o<��M������I���0�+�CT�H`�*I�!�,���#��F��4���C0�m!㧃�z@�B���"��p�0�������9�%���)����[�3�(ybL�����ߘU�S\L�VR!4�B�b��0�5�sN0�i���$n�3�*�&��$� �(Ɗ`Sk,)����Js�Lח�z���
`B�i
���#8�����W�'�eHG����CsR%���HJf�Z���Ă���S4����^>��۞��<R2f��3�	�盻6���9������&�&y�'k���~=�4�H�<=?Ji��,��d�K���<�
��ha��H��+�+�Bi���ic/3Ɏ��~��9�Iip��)
Ğ����B&��F0 �b@hb��c�`H�&_�J�s�~�$2��F1<!se����<�����~4�P�����I��! ���]�<��%!�:�a���X�#Ja��=����)�L�a��/���#���rE,)IZ:�\�U!f�$�w�b�v�bxA�"T����"F��ɧ&�$,� zB��8�)�����)��)��ƤH�(ጦVF��ɺ2)�
�ʒ����@�
� F��#�8H��0�y���Y1$l�<)�p���B��<C��r;�^ʧ�8$�B�.Z�
Z9!�B�k3��0�y�c��0Hk���7.��ܲ~5�X�y���焘����vynK�<=|��at�@����)�w����VL��~���@���LĞ��?y�C�y���"A�����\�%ɛ�&m����1b��e1#X�t�M(_5�9Ą����uY�
�Ja�.��bF��`]�-��x�?@����S!x�x~_� �g=1�_!��!.9�&M�z����&�����)�|b�`��"b�CǄx[��r#���F�+�1!!		"�!"�T��8Ġb�d�p�q"�G��PɄ�����8,ht#W7�s��K&n��<8��<�M1���|�kI���Ò$�J� B!�8���%�B%�y�7�)�}�ՈE!Hf�(2��4	L7 p���B^I�)� �f�a
Sx�Ą�	p�4�r��p���e3�'W����,�Bй}��$b��۟���?��g�{���f0�<���������, �
f��|��M�YHR�`J�~�.���"�B%X���¸+��p�?y��e�d�(���I��7X��IL�4�zn�y<�����9�H���*�k��1%�癙�|4G*�hŠ�#�)�sx#�@� �L�T04#\5O\t�VFE�O%p�
2����Ns��HҠb�M��~��a����x���I8,���@"�$���vs���C�J²���xp� @�c<	d�����,dR!d Pb?'�,
a뇤+��J�
���X��
B�$�cJa��H"0�@�*E"`�j`)��!
`Ġŋ�ƄB!i��A�O3�^v�D�xF��20��B$ՂG��X��@b��!p�Bŉ`p��
@�2D���^~�f�������#X#R%2�7L#=��O0�+(Jo�y�< �d�6������E��y��R����K;����5�0 DbPbT�%HS�,	M�?���B�!\|H�a�RYr2a�L�y�_58�`x�0
0)�! �B䫉
c�F�k�#�!���.eq ��x��	5"_P �H�� �@��[F$7��a+��%#\�@�B�(B��%��9Ȑ�Is�!I4#P�YD�B7!	�d�+�B��d��y�%:��fVFA�$HB$I	$0d�6CX@�0#`�)��J�Ţ��*1�X�0
��;��=������ 6�   /���8     �$    � � �V6�� $�i�7m�l�	p �` �c� �I��h$       H    -�l� �Z/  -�� �m��!�        
�*�� إ��\�$    m�6�6��`�[%��(@�	� ��@6��m��m��Y�:.��e� �Fݷ��m�"�-�޶�jE��V�U���ۧSǶb:۽R[p6�4��9m%Z�)kk����m��T(	�����l�km&��  8�Ͳ��m��*���T��eB^\� �m��� ��/�	���F[m�	 -�H6�  [@�����#�g�}�v�u��Ž��n� �}'�|H�j@ 6�hIJ �-��zM� �kn�/Qr�'U;5UU �'�� [A���c�     ��� �l�mGP��9Ʞݬa]�E�7-��m��z��5�6�8  .�I ��$i�T����[J�(� I���$I 9�'Xt�m��k��I�v��[n^V�$�@� -�  ��햰p�m��x8m�m$�f�뀷U�����ٮ��}��UT�6ٶ�n� ��l$Ă@�m���k��`N�;a �k$1�l[�a� 6ۀ[B@:@�S�		�m��$ r���L��amImm�� �� ��q�4�$�m��g�o��  pH6�[nu�ܼ:�瓄�՟�;��=[<���
�ץ햪�j��f��6��   � �\pH� � �m-�K�Aŷm� �K}z�m�m�m�,6k5Ŵ    r@m�nۭ�N��%.h -�MZ��-����	�N���Nۛi0[���l 6���Uٺ�6��G:�a�j�	�4v�s�\��ܧ_V��Ӥ���$�b�V��a.P8�0>&�ڲ�\ �+/3��UI%�m���6�5�!�m 6�ZR�\��h�&����-6�h��H��Cn�)���t�   h H����v[E�@ )K);l�*�qخڪ��h��6�I& ��6ͰHH�D�����ݶK$�Uӫm���m����l�p� '(�m�Y�yg����5TM�Z�U��h � [@l  �N�l�6۶�jV[[[ @@T�,�` ���� 	ea���E�;��6�o6�A�S�p�  ��c�� m�f�c��6�m�-� m�--�@VV��u[R��@�%�L}I-�ѭ` L�4BK� jG ��j�6��@�I�J��,��j� p\�;AT] �ʸ@$r跀 �Bڶ�� �.n��8 ��}~��I�#�/[*�ζ���k5��L �n��֒$�;m��9m�U��xHI�f�;h�Eqe@8�7f��D�-�C��=Fש���� n[�V��I�#Nڀ4k�����mf�`[@� ж�R�4�dp8���i% ����ڶۛ2K�x���ͮ�$8��t�+@Y���8��e�UT�A�<��$ 6�٧\m��}��!1ph�����M�����66�`��dsm�h�L��m�_6�Ti�-��_�:^��I-�V` �Y����`헤�����H۰6�M�h;m�E�� Z��m�l��p��   �	 .�ك��P'pp3ҍ�E[��������
.;M*si@zBB�5�v�޳9ÁoP� -�Y�9Fa�]��^Z��Ku��� -�X�Gs���d�r���VT0��).�y]�mL���(�Rc��\��N�e�֠�\�ur�BkT�HMU���Ѷ�j탐I�m�	$���F�gO9Wo��}T�D��^�L�6��ګJ�­U�U.�U6y]�l,s9��h i��� �6�$"K���  ��0$N��`			�.�&��H  $ݪM&p;m��u�v���  �-��+[v�?6����r��m�l ��^��m�J�m3[��$    Ft�n�m���ޫh �-����a%� 9���P�1����UT8�n���É�9��m�`  -�k�l�Ku��K:���M�i5�X�6�H�kGZ[%���a���
� k�ձ��`��2�
�T�r�UUO$�������l�e�*�綈RΑ�xe��+7R9��(q�7 JҐp�����R͍vޫ�zܪ���
��]��e��@�� յªU�ƙY]U�F�M&Z�Î�`��l���f�M��8����a� 6���A�4�    |o}�|�U���2l�VT�Z����"�mt9i��      86�m� p�Kn���kXH��x6��*�!5J�4�� � m[kp'@�����u�m�#��h��kr�%�  6�m���-�    jL��e��K�ǭ��� n�t�5�,�Z 6������#m�
Bۇ#֫���۵�.�+�P��.�m� ⪄�j�VBxv�A�5r��j�,J+UR뎗*��	�Z��J�z�h�^f�t5�/B��4u�i��7-��ᴝ� H��������6��v���eF:6bj����[@ -��@m��j��@h
����  j`.����b��j���UoV�[i&�  �5�À6S`��0`[x��'5�S�	 ����h  )�Ut�mN���H5�n[R	�h�@ �ȧej��\�� �U[*��  �o0�[��u[�  �J��UUN��x��˶܀�   �����n��II�i  A����_��6�a�mƵ�m�a[l�K�$�����Vn�S$ � � H ;m�f���h���`����Ytk�<  $ֹ��v�[�5�K4ت��{[�D�q(��[I	���8-���˚z��@��nع^jv�q�
K�L���]UM���p*�`��t-�����|]jiZ�Bv��p���3m5�l��Cm�����:���k�*1r@�4�J�S�����}�p�`-���5�7n�����d#h�GZmu� �$��!�!:��J[o[��8 
������[o/�JKJP��l�*�WA�a���ۜ�mP �W�Ãm�����h�|Ѳ��u�  ziq�UV��lZ(
�DOZm��  8mb[y�Kh>� 	M�ղAl:�l8 �&ʹ�[l�veT�g�U����kd&����J��K�±�m���� �.lݶ$  M��`'�Z�u��
��UA�m��1��[$��U$�ɦ�0� �h�$[�H/S[qm�j	2 I"� �    I�!m�M�6ء[@UUR9
�	[���8 � �� �  6ե�Y�e�ٚ@�    tt�w` �$�^ݯY"�^�=��Ӂ $ �@�qm �  �` hKB@ �a�f�ڶ�V�8�NnY�(��kr��n]ҤZ��@ Z�p $   m��m�` ��   @   � � �� Im���)���m�m��`*�k��iV�Y�j�p ��   �>�}�	   H ku�ĉ$K5&mm�       �7�.�mE��c��w�5V�QHV�e�4d�n�Y�f�ISS�H| m-mZ�6��k�Tض���$ m�ݚ�
ږ
�y��ضU�gkh��I�-���n-��Jo]��a�e�hڶ8q�[.�����cm��K�[@�S`    &�{l�e��    -��A��zݶ��� [�66�[G�@H� [@   m����r$   l-�yX�` m$���XZUUꪪ��@� |o�� �Y� m -���۶˦���  �A���h   @��۶�  m�  ��ݭY�����A�7m���P��m� 	  �@    ml�@1*�T�x�h
�W 0Hl�( �6�,�)z�� �
v�nZڀ�R:}���жN6��-�h  �Z�m� 6ؐ�nm��m��۷a�K`ⶕj�xT�ڊ)Y@j���m��P��YY[�F����>�Uj�U��쵐�!�k��{������1O�H�A >�1���P�x!����P�@4 ��~Tj?�ߖ�AA��0�TL<�P�TC���Ax��?�8��E@*��z��� ?���"��*�H=x."��~�B'8
����� �U<C��q���"~���"�Uز#�Ƞ��9�?"��u`DBW������uO߁�Q}�/US�q@ ������(STP�FF2$B+c2:�&��<� �H>*x��S�* �T��h�PB��h����` ��"�*���D�j	�G���z�X*1����tD|��b��@�����S��~C����}���!�P��G�� ��������y����" =�:�#W��N��q_T��8�B	���tTWT��+�"����������F�t���@��-��e�UR�4�˰T���;����/I$������H���5v�ۦ�-�F�ٛۮ�j�.n�gs]�s"�<�a�gpl�N�99vf��S���*�a¬�ۖ�v�hA���6�nۦK�{$B���^q�I�����z4��[��*@�vz��6E�l����
nI̱�T�/
���v���O4$f\	�yۧ�ݹ�{].�m���ŹaM�Ļ���ZD����[/P�� ��õ�'�ܸ�9�gDKK+;3�U���! �vv��u3v�EE�#>��
3�NWz��J�(�ɂz�� mMuˡ.м��`g<\�Wn�7C�k;<t��z�ɮQ�KN6�����ʠr��8��6�m�a���rn�V�nZZ�c�9FeP`�z�F�I��^��Pns�Ӷ�pM�Ss۩�(p�U�e�Avg�H��e�c�򸢰�q�Ǎ�.:�;-8�Cҽi㞯$:�c�K�hr,Gm�Sj�;��*�M�
g�z��.u��Y���.N�M{<]�!m�Z����e�X��^��n&Mp����7bCi��ŀ�Qe����Sd/2v�i6�NQ�;s�ۯ-ţZ��:B;{��\�4
��#l�殺���&��[��j�rN��V�W�¨�cp>�í  \�&�SO^#M���Y8��ۑ��ð'�6�䝂��I�儎t���a+�Յct
Òݵ����L��qZ�&Ɗ�m	���ӛ�s��T@��g��ZMrΎh��.��/ot�e��d��V�$UX&�Y�� 	;kn�D)$����N�A5!;T�J���G���,��z,��T��;X��:X�#�k&SY��	l.ۘ��rKx$�#v���6jJq{8�s�K̭�*jn����U��&Qꔕ]����z�+jĶ췁#�l�s�#��b��j�z�ɻ�@��tmyn�#�t�t����P=Tz���� $X���ES� ����'�>!��T����I/2����[-GQ���f����d�&�nM�p��9;0�K�;Y����l��L�U^:��e�a�nК�m2p���ml��,���$���p�ź������<�.z웶-�
�цuû<�n�qۦ�a�nV���נ�똽w]�&Wgs�Z����]����*�)��âx�c���v�Fѵ���L�76�\�m�����@H�}���G����d�p�C��.�D�W�8��y�\��	�����RC!��ՠ~� ���_��IB�!�]Ӏn��=�w77Ew$���m�:"!D)�y�,�]Ӏl�נv*����$�q��z���3jD��Sw��
�U��+�UЮ��ͩ��L޸06t��U��^%�0d�8�^���p`l�6�LQ)=B��c��U�07��v���)���;����و�Z5щ�IƠ�E�ɋ�n=��MgG�mH��J`j�T���r���I?w���<< �����bH@"-�")$%j"!,��/k�w]`��0=�W�by&h��Zyڴ�.�>4����w�J�I��& �WwV��"`n������6�Z���Z(�k�N=��MgG�mH��J`}�}#���X�J���.�& ܨFx��:��K<]�\���"k&8�,cI��I����s@ͩ��L޸02TD*�w�^�*�Uc6�L[%07z����M�X��)�$qh�kП�{���4 ��B ,����҈��;�{i��?=ySeVE�ɋ�n=��M׮���ՠr��@<z�8�LLXF��8hz�`�78ϛ��v��!:ޯ�n��Y�;g%�I������t9l��+�@;vj�յn�ˊM��)��ng�د�u}�`r�)��.�����)2E$��#�@��^��YM׮��YM��x�q�R!U��;f��L���=���.*����@ԐN�Jh󽼒{�;��1Q>U`	~�� X������D��ID,��r2�]��M���j�v�Lڑ07e������}��Hs�-׋s8�ϙ�=�����&�$�����h�	Ykh\���m,xu�Ӏ{�l�<���H{k�p}~֠�E�ɋ����t����s@��j�;�ՠ=]j7���*�����6�Lڑ07z��3Ǒ����D�I��;V��v���M׮��i+R�$RLA*n�p�7XB�y��7�b�=�n�I�ES�� @�P�
B�+q ,xU�We�UU�4���kFG��kHOR�l�c���ưٜ�-�'b��/l�s��R\�3�K�n\�i睹ლ�6Ӛ��v��*�m2r�nؓ1/	9�GSۣu�.�"�ݭ�Y���ĞVx����<��Qi��eӽ�qa@t�Md
�F^3ӎq�d/�m �5FOb8�'6\=Ȱ�����[b9%�F�m^�2E��^�^x6��5���"t�g�9#-��0��[-��V��[12����ߝ/ၳ�ڑ09l���(��č0hiH��z�����ՠw��@��S@�]E�2,�q��@�˃��L�p`l�)*�+�ı@jH)��Z�e4^��=�)�~�u�7�a2b�$�@��� �׋ ��� ��u�}�_��{9q���ג�ݲf�ۉ�[6.��)=u�l����&cv�,,��Î�g���O������Sv�L�l���5sd�7k ���*"?�R�Qj8����3�� ��np=x��B��2E$�����v�޲��]������<V��(�E�%V��p`l���͗mH���免0i�H��z���>�Ģ����=���=�`�-�L��ꮮx�&Ϟlq�4QK�ܵ=�\r�u�\.mat�ra��L�0bp�?z�h�j�=��h�w4
�c��qJ�
�����7���B���7i�����������֠�&LX��8�z���I-P�"�Em]� �;V�x��D�LPXAǂqh���"`vԉ��] ����Z��!Ǒ Rf���ՠw��@��S@�빠w�y (��N6����;,��uc���ңָ;[e��ћu<�)& �IZyڴ{�4^���;V��<V��m"F��@��ٜ�(S&��X��� ��u�����Qb�5�b��4����~�hz٠{�)�~����
`8ɻX�$��m�N =���f�C�D�<=O'y��$���ɝ��vLp�"����@��S@�빠~���;�W1��4�d1�k���bk4�ٸ���L���b�Xd�b5��L����1b�#rh�Jh�w4�v� �[4ǭrd��x7׮��IL��� {�x��� ^���bs��I��;V�w���Қ�]���+b��bԑŠ�[w����"`n���\"���I�94{�4^��?y�8�n�!$B��"n�U]�ԉ,���������=�֠9ǌ�c�@ج�X-qv�YI:��`�<�2�����&��-��w��W\���M)���s���{I�����c�ط���C�1l�
:�v87j���p6�vv�yh�:�2ok-���/;��!"žM���y���F���R��)�yǤvy�p�Z[��c������S!���u�[^
�/���ߔU�8"'6rK�l˦�4�lʹ��\(ҏZ"�f�����z4+vG��of��H�M�F'}gƁ��ՠ�f��t�����7�dX)��J�`fԉ�n�l޸07e����<�(I�8�޶h�Jh���?yڴ��q�q!L��I���w��p`fԉ�n�lOU\Ĳb��<���YM���@7d��\t�ЄU�*�3�o(N��Nb�ٷ�[���9����[�X���'Na�q�N�;V�{����Mץ4�ĭ�HAɀF��s���1(��BJ2.�f�0��f���ՠ{���E!Hpiɠn�����ڑ0�-��Qp�bLi6��4^��?yڴ�l�=��?WQF�L�0bp�?z���	K����0=�`߾��Ö^�x<��R[��<&w�[[!�������f��C]�]Sqαf�k '}��7z����mH��u�ƅ2`��#rh�Jo�ى��s@�?�Z޶h�U\Ĳb���V`z�`�M�[p���H ��I%�1��B<D�+��@t"��
� u�5�2�-V���bD���]T��F$T�	p�"� �=����*���L%�a�S##QA� B%��H$1� �HU�| WX�FV0U��8';D�����0  �"���!,��8!� Q �qE��?<	� ���� H4QC�T=C�`�+��H9'?~���u�M �y�#�cp@)3@��b`�[w��p`vג��ݐr`�#�@;����Mץ4ަ� ��s�3v������J����w/!Ypb�G&���*�aX͹���;N����u�q�m!��'�;���=zS@��)��f�ت�YbLi1�N�\���;d��\��|����"0bp�=�w���Қ�Jh�:��1I�8�|����0=�`R�Q�H�G���
(~���䓽�r�.]�M%����]�7z���l�03jD�7y�߿���P)պB�]�Ζ��nˮ\��l8�>�z�g��kOg��ɤ���,qe]x����#�6�L�K`n��@3�B���
L�?yڴ�l�=��=z�h�Ց̃��.��զ�%�7z��������Z��H����Қ�]��v� �[4���&�T��X������R&�%�7f�rI��"�ߗ�l�3<�ɻ�������}]�3��9�aኤ�i��˸�v;R�ͷJb�36ùfQ�NrJAR�Q�98�u�szm���u���8�BҘ3$�LA��N�%�]�d�kv5�3��f��A�b�X��pb�փ�.�\wi����t�ԅ�o<y�"{F`[>������+8�[`�c>3	���)�v�P%��V4��~��߫����|���	簺�=<�k��+kW����nv���g&��6��^�rh&蚳��?}�N =�_�7z���;Ͽ, �鮥J�\J�Swe��t�=�w���m��N��NϮ���6���uWy�2n��o;��=�j���@<{��K&(, �UX����H�l��ݗ�<���a��Y�{�ՠ�f��YMץ4
����SĜ'����G�rt�ڷs�gO7��b�V�D[���ds�7 NG�w���e0=�%�Cv�� �
	�E�\�*�V\���;f	*���H��m��S�@;��⫁e��i6��4=�`�78t%�L�{� ��� �]�Sy&D
`(��{�ՠ�f��YMץ4ڝx�L��cRYui�v�l�p`l�v�L��~_������c��gG6�e4�rrGbۛ:�Z�$u�Y\�����RK�~����06u���R&�%�yqdɊ�'�@��M�v� �[4z�h{gXG0�n,�!5f�Ss����/��HzK��%舿���0�l�7�$�9��i�����@�����Қ��Z�5���������$���?�]Ӏ�� ��~}��Ͱ��͛���"F(]�	FV���:/Y3�I�q]�\ű�/ ��*� ���ڑ0�-��.�.�L�"0bp�=�j���@�����ҚmN�d�r%v0�-��.�p`n˃.��<P$�dnM޲��Jh�78�DD*�wn�ޝ*���M�"q��4^��=�)��f��YM����"9�@�$I�XS����=�kP�l�C��z�E���7���`����׭ Uf�_|�l��ݗޔ�;��������#�@;���06u���R&�P)<Uґ�X��@�����Қ��Z޶h\,V6��i�18h�)�{�ՠ�f��YM����$ȁ_�]
�`nԉ�v�l�p`l�{9$�������#D4�����XZER�t�bv jq�{f�79��jA���#'�6��#�N�=�&�7I�v����n��0ln׷0ܼ��Ӡ����X�c]�r5�7��y����v��v�&������ ITs�n��rsqnK��.g<͵�6)�ѹ�qa��0l��]��c[�i�n8-ӛ�VD�շB�؎�d�p�/U�����[�~���Da�����D�{fn\���|�.vf�z�=�]���R'�<��cNET��@�����Қ��Z]]Px�I�,$��� ���?�S&�0�� �7x�.�Y1AdN<���Қ��Z޶h����ydNa��YV07jD�;d��06u���x�Y��ɈNG�w���e4^��=�j�=κ��m24%y��q)��.��%���s�z�h�WF�����8ԏ����e4^��=�j���@���b����ڑ����}��
(��@!}`+���PCb�L ���*� � s&����I<��� {�S@����L���b�N�ۜ �7xtDBS;�|`���ܲ<���D4�QŠz�޲�=�`rP�v�� �}]6R��)EڵWl�p`}>�� L�K`~����^h�mw���Y4�6}dB�k����9�l�n��X�\X�g������0�-��.�{9�'0�N,�p�=�)�fbA~�M���u�M��.�'?��6����z� ���
�Z�E�7x`�e4x+AĤi!��&��YM�Jh����f�qU��co�ld�N^��=�)�z�޲��,�J(��cǉ��D'��:- �/F��kK7n��̓>��E��[N݂�������4z�h^�@����ץ4ڲǒ<s ��Hh^�@����ץ4z�huuA�&�"rh���:����YM ��h��n�d����hzS@��� 5�Q�%��
`�)���bb@
����Y��4?�Ўa��Y�{�S@�|������m��ZЮf���<Y�(n�<��ڧ�k6����.:�g�z�(B�ֆ�Q��\��I??�����`��ߤ7z��7B�{��I�pmɠ{�S@�Қ�e4�Y�\Up�X��6�bp�:����;f2>}x�_ڝ���F�F(��{�S@:���e4:%��0��uһ�v+SSWs7f k�x(IDn�q����=�l�%Zz�`�""b�����I`Vx�HF&`H�R����Y���<�� F$D�6$�P�!S!%Č��8���J��HF7VňH�F$P%��`��)��B HA#$`A�Hĉ��x��h��R���
�	д�d��H�����$!�;��4��RH%F%�%!B	B���ǀ� 2F3=���!��W��P�!B@�	���)�$$��c#��|< �����q�i��1p��L�&��BF���	w�1$�3�����-�O���$�$# E����FBI! �HD��
����ȜK��t�?)�ǪA���␜� z�N< D�S�
$ A�>'��F��ۓ�L�P!V �"ȋ���$&?���
�0�d�Ę�JJ���X�H�	b#
",bD"�g�����M��n-��H𷝶�mK@`�Uٜ�5R�
�[q5�[���9���nz�5�ӹ�u�]���r��۫v�J�q��f�8����^2񆶻[�=<a�� ���'!�uµ�};m[�%3�uJD���Bx���M��٠�VN����zw5竌N�lt66Ɂ:M�э*N,�;vC��.�-��.bQ�`@6�.F��x�l���X�"6�4nh�<r�ځ��t�v��d}�@l	��V�[6'�h"8.�fuѻK^�Li�u9�����)���5�2R�:�]9��,H�z���D�8��]x[P��X�N�'q�ֺ;e1#sܺ%�C�k������Սth͓WA[�〮,�u��v�<Hyۧy��V�@�1e��{B����q�p9���͸��ݦ��ź�Y ���t6˳oS��m�u������2/Q��զ��=9=�S,�۵�Eѫ�֑�v��{;�v�z)٤��W�v���qÄ���d�&a�"�{`~>����f{m��e�vK�����n7+lV��s-�Q�m��WR�RМ�ϚY�H$''Xl��Wp�Z�����^��}Ӊ�6�����v�mm�<n5,�&�s�֩��l�ޑ[F�l	��m3���ۋC�z�[h[S��O]��W۾ه�j�:�{mUz�  ��\C8���Ȇ5���8'5la���I6����m1Ҽ��X��:c�v8�	�*�FY��;D��m�M#+Å��j^���	Xagl5a	8���]��閴��6,�K�Ts���×Q+0 ۣBdUVVu��nE�ꪪ�dy��2�
F�;L�J���S���8&�mՠڶ������{�M����\%X�`\�ҭ���;i�`�!5=��H=�#I��@R��e��*k��+Di�r<lCR�N�ջ],���`� )��9�`әnM��[�ٷFe.(A����9���M����3L��˦�h5>O���u<EO��<C}�+�*	��$���wn�K72�I�2���h՗p�͘ݳ�L�)�;6��ˇtth
%�Ȝ�}��W:튼M��T�m�Y���n��7l�v���q3��gûk�^�rn.�����]V�ݲ�k�����Z���r��'[��\�LnGq���F���۵p.�  VS�	�\��.�z��y�ᘢ���0��m��7@m�V�qOS�-�b���m���6F��y���՞�ut����i�Ya�I�Bcq���@������|hzS@����u�4�\6\Y2l�&��Uf�m��%qF�_ ��4z�hq��0�a��Y�{�ـ��
gw���0�)V���RO獧��u�4z�hzS@�����hH��i86�`n˃=�\���:t��l_���Y��36��W*:�[��W[40����e�+D�6�KP�:�1�k�f�;f k�}��_2������nE7D՘��(���C_T0@d�����}��@׶��!���Һ�v+��Wsus����7e���K�07e��:]Jc�L&D��=�)�u�M�v�I(�|��vYTr�jl�SWh���Ӯ�p`:[v\����h���4E�\Eo�.��՘�㫻w]����� 4�q��y�\�Cv��A���=�l�z� ����"��]�U�/�m�����N) ��h���5� ���:Jd�
	����������w��^�0��DZ��o'�@:���W,��&�H���%/�q�n�����>v��,��6��Q����t���M���^��=���LqF�o���y��n�3�,��=mNl��1ƌ�Zz��*��ď$��biȔ��u�4z�hzS@����z�[(`��"r�������0�-�i���Y1B<M�n^��=�)��?�:ݚ�e48�u��'D�j��v� ׮�y�0)B�K`!
 B K�P"� �}8��?����i�!�z�޲�W�h���?V�JL�2'X���ܼ�	���ܚg���(��qg�d�;��gml6Ԣ��86��=�)�u}V��;W���� :ݚ�W	6��c$bp�9ֹ�P�dݮ��ϯ ��� {R����6�F(���=�j��f��YM��ڬy&8E�NEL�K`n˃�tL?��u��`}>�ꢔ�]�@�W5w�{�ـ|�_D.�;����N k�x�B��MVU+�Vh�c$�ё�	���}t�j�
Ƚ���k<2�H��.�f�u�n���z	Sbٶ4
ڑH�[�gkveezm��(C�F��q�M�X/3��봰rQkv�kgOn�[�c�uցݸ�nXõs��M:ɥ�M� ���f^�R�m�$Cjź7*g��E��N1՝u�vY &����=�`��;�\m��#m�@�an�|�� ���n�˷�h�uZ��vY��FL��n�r[zƪ�q4	Qrɐ���bY1B<NL������z�� ׮��Hn��	��Z.��ő n-�v����h�O���^�Z�s�9?�&��- �������]v�LРR��C�nM޲�Wj�=�j���⫁e������4���ݩ �%�7e����ڪ��(����[�gk�M���h��fU��������IZѮn�Tu7)�H�Nh�m����> �l�=�)�uv� �U�$��.\ݻ�y$����~���ٿ�������=�ns�IBS'o]uQJl.ы	2'&�����:�V��;V�u�h�r�bY1B<NL���ڴz�� ���t%��� 3S�W7a�q⍃�h�h[f��YM��huu��1�p��`Lx�N�]���my+r�6'z�'a�������=R<m9Z�٠{�S@��Z��Z�h8���86��=�)�uv��v� �l�.*�X��M��Bp�:�V��;V�����3��@��M�Y��i��1F9��Ss�ۼ�v�_��g�N }�O�j�U�*�����\��� �7{8�����=�j�?z�1���y�&��7�����e4�rrF(��FN	7j9��ؒS��	0ń��@�����ڴz����?H�� 4�=V�U�Wt���5f����	(��v�� w^�;ft(J"d�����RUқ�
��v�� 5�:""��_�}8ς[������J�j�p>J>J*�������]k��Q�J�%�%�~�h|�Q��rh���5ֹ�=�np^��>��Co:�Um��왳qX��p$b��xf�s�
�5=u��}6\�JG{��_lwҾsF��wӀ{����wпHn��t�M���j#cqh�o���4�Ɓ��[�A��}&I�d�ӑGs��^�;fBJ"&_S��7k�t�:��@�XI�94z�h_U�{�ՠz� �{�sɋ$x��'���t����~��e��/ � ���';�������	�Q�af�f�z� �fH��߼o��s��JUm�����r�6�uM�:�b��ա8��n��	ۭ���msƗqXu�Z�C���t�.�C��ƶ�sB�n��i�k ��nť%�A�Y�ûz�Q��7O+"�ml�ݠg=��<t��y�+�=��r�k��S\ӌr�-9y n�J��s����6<Q��;[A��y��?����Y���&�fl��e�.R�n��R�cθ�$���sd���T�r��(�7����@:���[4���9x��?��6��- ���l���]v�&w��jG#Hpmɠ�l�:��@��U�z�⫁e���َF7&��>�Ӏn���z��%3����i��hq��@��U�z� ��� �Z� �I$����\L��T���b�ŭ����I�X�~7�3gbh{-��k��bvr�ush�h��6����o����f���Z������oa�&�7y$��w��>=�tH�ey%�*�?y�Z׬�����b�@NW�h����E��4w��@8�dN!Ǌ6Š{Ϫ��f���S@�����+cn%R����� ׮���q���p�R%�ﻝ�9ı,O����˷.���2W�ew��Ss��J=��힅�r��:����|#9�6K͙wsw%3ffn���X�%���~���bX�'��{x�D�,K�w;h��*_�6%�b_����'�,K��3��IM��nd36[�19ı,O{���<�bX�'��v��Kı/�����%�bX��w��>Eʙ��;N���r���36�<�bX�'{���Ȗ%�b~�{��y�D�}X0�X�0�JRE�$) 1d��4%HAHPa$c$#BH��T�*��N1�t��R����q!����p� @�*x�4hKV4#�*1!�mb����M�E� @�spe%���0��
�	
AXD,3QCX2 �13�I!�1��°��?� x���58(�LE"��QD�S�P4P4M�	�}�<ꪆ"�? �U>�6'���br%�bX�����yı,K=��l�3f�lɛ�smND�,�D�{����%�bX�Ϸ�Ȗ%�b~�{���%�bX����S�,K���w�l��[&�M��'�,K��;����bX�{Ͼ�O�,K��n�*r%�bX����8�D�,K����ۮ��Xl�&�ͶS�=	�x�Fƪ��Gg�+n�E,k�=��]���kM)��]�36b~�bX�'~�����%�bX��w��"X�%��=�s��?DȖ%���~���bX�%�|w�6��Y����36�<�bX�'���Ȗ%�b~�{��yı,OӻىȖ%�b~�{���%�bX����w35�f�3.mݕ9ı,O��{�O"X�%���٩Ȗ?"+��=����yı,N��ҧ"X�%����/ve��ܔ�ۻ���%�bX?�����bX�'�w��O"X�%��{*r%�`p�?o��q<�bX�'�;{%7s1����nl��Kı?{���yı,O}��S�,K�������%�bX?�����bX�{���������U-4\��ˈϵ��7a��3��Ů]���6ٲL]<��v�&�'\Y36���X�%����T�Kı?g��q<�bX���f�"X�%����oȖ%�`����͙�iw%��n�Ȗ%�b~�{��yı,���ND�,K����'�,K���l�XB������:UH��	����s��Kİw{59ı,O��{x�D�,K�n�T�Kı?g��q<�bX�%'�s����6�.�36jr%�g�"{�}��yı,N��ҧ"X�%��=�s��Kİ|�RB����Z�\݄��uRfm�yı,O}��S�,K�叻߾�'�%�`���59ı,O��{x�D�,KqX
 UD�
�����۽���{���Vl5U�u�TRI�-QPr�nF���Q��u.��+��A�˺,��=vǷL������[j�8�֕��^�$x�e,C˶���Ӳr�Le��
���{g�;^ݛ�H���&NC����J"�Z��cI�=��}3���B �3���5s�u[5��t�n��N�4�n ћbd�s�!�Ĩ��u�jͅ��f�����4�͛�|��.����Xm'D]���'@���w]8�t�,�k�#բ�9���Ix-g�k�*yı,Os���O"X�%���٩Ȗ%�b~�{���%�bX��w��"X�%���R^�M���Lݻ��O"X�%���٩Ȗ%�b~�{���%�bX��w��"X�%��=�s��Kı:giқ����fm�6jr%�bX�����<�bX�'���Ȗ%�b~�{��yı,���ND�,K��Nܝ�6�[4�ɛ���Kı=��eND�,K���x�D�,K�w�S�,K���s�Ȗ%�`���͛�iw%��n�Ȗ%�b_{��Ȗ%�a�~��SȖ%�bw�����%�bX��w��"X�%�����L�7n���@��X	�o5��ugc����q�����5�ծR�L�i7d�M�nn�<�bX���f�"X�%��w��O"X�%��{(}<��,K���'�,KĤ��ni����-�%͚��bX�'����<��>�[!0��"~�b{w�S�,KĿ������Kİw{59ı,Os��tۦ��M̓sx�D�,K�n�T�Kı/��w��K� ���59ı,N���q<�bX�'p����]m�nnmݕ9Ĳ���� �)��٢H$���}��@��Bns���)!I
HOY���-]��͙����%�bX?�����bX�'��|�yı,O}��S�,Kľ���'�,K�ﳲ^m�.�w.�I},à�ҫI�b����:J��uv����O�i��n\nd36ۛ5<�bX�'~��8�D�,K�n�T�Kı/��w����2%�`���59ı,O�����I�2٦nM��yı,O}��S�,Kľ���'�,K������Kı=�{�ȟ�2%�߮��tݛK�,��weND�,K���'�,K������K�E`�!��`%C�U���X�~߾�O"X�%���~�9ı,N��3�fI��ɺm��'�,K������Kı=�����%�bX��w��"X��"g~����%�bX�����r]ۆ]�\٩Ȗ%�b{�����Kİ��{y���Kı/~����%�bX?�����bX�%�~��f�[V�Ex��]n���]9��u�>�����C�չyu�hn�j{K�������o'���Ȗ%�b_{�w��Kİw{4?�����,K�����<��oq��׿�_���S�(�c��Kı/�����r&D�}�~���bX�'~��x�D�,K�n�T�Kı=��Z[��ww7-3ffn�<�bX���f�"X�%��w��'�,~Aa�2'{w�S�,KĽ��oȖ%�bt�ӥ7s1����nl��K���B����Ͽ�Ȗ%�b}���S�,Kľ���Ȗ%��� � *C���A�<���Kı;��ے�����3rfm�yı,O}��S�,K��P#���o�Kİ}�~���bX�'��{x�D�,K�=��Ɇݹ���Z��lc�r��0q�XĨ��mZܽ�K6iQ>T�����7f��K3v��SȖ%�b^�߷��Kı?N�f'"X�%��w��'�,K��۽�9ı,N��gp�6�M-�tۛ�O"X�%��w{19�A���ؖ'�����yı,O���*r%�bX�����y�r�D�)=�ۦ�4����\ىȖ%�bw��׉�Kı=��eND�,K��{�O"X�%��w{19ı,K��{��t��w	��fm�yĳ�U`dN���S�,KĽ��oȖ%�b~���ND�,���s�^'�,K��	�3��2K���6�ʜ�bX�%���x�D�,K䏳�}1<�bX�'~��x�D�,K�n�T�KİC��O����ݛ�,˹�rc���ht�����Q������=iƩ���1��pD�J�+mn��Ey��]�XκY�-��nM�˞.9���S`$��5v,���n�`$&��V�z�1u�l�p��õƴ�hgMJL�3U���:�p�u.+�[n�vw�63�-�ֵv���^	��qc1E��u�_e>�y�c�y������������u�?q�8��sעܱNf���unM3��Fr�x�g�{;N������w�>�n���]�3w��%�bX�O��br%�bX��}��yı,O}��S�,Kľ���Ȗ%�bt�ӶM��n36[�19ı,O{���<���'�"WblK��J��bX�%�����yı,Oӻىȟ
TȖ'��v�s2Y�nLͼO"X�%����T�Kı/�����%�bX��w��,K����oȆ��n����]Z8�f����{��|�"g~����%�bX�Ϸ�Ȗ%�b{�����K���R�O��J��bX�'�����3��Kd�6��Ȗ%�b~���ND�,K�ｼO"X�%��{*r%�bX�׮�����$-ۚ�e�eX+�
��4)+vk7mI�m�-�]��ih"b��M��w��|�w\P�V�g����{��2w��׉�Kı=��eND�,K��{����dK��}�LND�,K�zw>�t���.�I����Kı=��eNA����KĻ��x�D�,K���br%�bX��}��y�ʙ��	�3���K2n.mݕ9ı,K߻��<�bX�'�����Kı=�����%�bX��w��"X�%����[�廻���6\��'�,K��;����bX�'��{x�D�,K�n�T�K��dL���x�D�,K�>�ԛ�1̙36[�19ı,O{���<�bX�'���Ȗ%�b_{�w��Kı?N�f'"X�%�����na6f]7B�9���A�Ի&�d���nd-���T�Z�����Ͼ��v�ƹ������oq���n�*r%�bX�����yı,OӻىȖ%�b{�����Kİ}����7f��K3v��S�,Kľ���Ȗ%�b~���ND�,K�ｼO"X�%��{*r%�bX����w0�L4�M�nn�<�bX�'�����Kı=�����%� �� bDdU�!��6'{w��"X�%�|��'�,KĤ��sf�4��fM�.l��KϠdN���x�D�,K����Ȗ%�b_{�w��K�����>���bX�%���}6魙�nfIsoȖ%�b{��ʜ�bX�%���x�D�,K���br%�bX��}��y=���oq������Ey�m�.y����6���!�%o-Ƈ�3\�yctВ÷���=?L�\��2���SȖ%�b^�߷��Kı?N�f'"X�%��w��'�,K��۽�9ı,Oߤ�/{����[&l���O"X�%��w{19��L�bw��׉�Kı;ۿJ��bX�%���x�D�,K�v��ݹ��&f�sf'"X�%��w��'�,K��۽�9ı,K�}��<�bX�'�����Kı;����zM��v�ܙ�x�D�,����T�Kı/~����%�bX��w��,K p"3����	�u~���{x�D�,K�f�sp�6�rY���ʜ�bX�%���x�D�,K�U��y�1?D�,K�����<�bX�'���Ȗ%�b~����iq�ҡ�L��u���B#��[�5��uآі�Nʗ;be�Ok����'�,K��;����bX�'��{x�D�,K�n�P�'�2%�b^�߷��Kı)=�ٳr]�3&�6br%�bX��}��y��
�M�b}���S�,KĿ}��O"X�%��w{19�r�D�/g�s�M,3p�̒��'�,K��n�*r%�bX�����y��R"{>ߦ'"X�%�߷�^'�,K��I闻�d�f�.\ۻ*r%�g�*@ș߻��<�bX�'���br%�bX��}��yİ?�FdN���S�,K���6K��w7v�$͗3w��Kı?N�f'"X�%��w��'�,K��۽�9ı,K�}��<�bX�%����$W �U���D�����F�B�E,�	��� @O@�\R��z�@B� ]��H��EB�U!4�A:B����෺P)��&�#��9(�� �)�Sԑ\\�=<M"��]�A�"�p��1��P<!��`���(g�y��ݓ0���&�ݖ��I�m���-U]U@�\ lNQV�U26�J�������%�T���d1AƓ��p��uj���	Q���b�d3��r���{l�q�"�:s@g{"lg�N�V���ݞܗ�:8%���{I��F�Ckx���K�%�Q��s{WY�9&5��.��d�u��[ɻ��p7�� -!pN1Vt�&M�:���#n�����K][\�4#�Uz4�/a�P��G�N˲VӋ��pT��>�Iٝ�f-�, �T�ۺ�l�6�S(�x�|=�x[;Um[x�.���]�Y��.IM�����70u�[]�\�]Fڶ|q�.����*��T��S̓��^E�哎�U�vm�� d�cd��� (SW�Nm�.�6�UC�z����m��z��.�5�qN͂��x�۟6�;W1�g�Wcdf-��Ջ�qp���!�:��;=%�(ஃ�g�-�s�l�'�z�ey6\���I���Y�V���k��ִӯV֐�'5�Ժ]2nƽ�:ˑ���8�e�᪨d�������ɷ�Ls=���B�pĵ�Y����c�n6��Җ�f,�.��Vܣ��`���v�6:����oj��j����^���NS1؉v�=6(��lP�/E���}KKR�t�m76� � �yRį5���;l�p�]�%�mDD����k&�s��q !F�d�=�'�e�%'M�\�c/ӺI4;q���/Q�]��q`ݒm�eçtJ�s�����z6sWB�Typs�f�� %�c�*�Z�ز��vej��+�N�VI��V��PK+�GTu�Z֐6�B@6�C��&р���C���d�k�2�:�.��͒��1� aݓ� �Ի�uR<��#��;i6',u�Gk-���s\�R�]PL�Hpv7���,��9]4��U٘��a����R���kO85���g��MK�j����E/'��O@�_q���=�~{�n����]R�;��;U�#CP��<�k�w6�ѵnq��n��Z3�4���b��]9�;$7l;��dܰpI�;�gY�6����YWwd��;u�zM�S��g3;ɕ<�q�h-ڹ�]SI�[u75G'Q�<�jOkA��64њ%�13�'���[����hg��h�w.���0v�c��]��\����Ѭ6���j؊�]����7��vL�v�v,n���rf.�W�Kii	4t��4�r���O�ἧ)9�1�d��nl��%�bX�}���<�bX�'���Ȗ%�b_{�w���L�bX>��MND�,K��;�/��̗K3rfm�yı,O}��S�,Kľ���Ȗ%�`���jr%�bX��}��y�Aʙ���s��3v�rY���ʜ�bX�%���x�D�,K�w�S�,K����oȖ%�b{��ʜ�bX�'}�2��7I��ɺm��'�,K>��}��MND�,K�o~�O"X�%��{*r%�`|�ș߻��<�bX�%'��6nCK�p��%͚��bX�'��{x�D�,K�n�T�Kı/�����%�bX?�����bX�'���{�q"j"L��\k�K3���T�XĵҒX�#wc���t����y�]��E��Ի'�,K���ҧ"X�%�}��'�,K������Kı=�����%�bX���rwsL��ۅ˛weND�,K��{�O!���T*�Ï"dK�o�S�,K�������%�bX��w��"X�%����%�r�n�,͗3w��Kİw{59ı,O{���<�c�C"dN��ҧ"X�%�{�~�'�,K�靧i3nV�3m��S�,K?���;�;��yı,N��ҧ"X�%�}��'�,K�d~��S�,K���N�K�73%�ܙ�x�D�,K�n�T�Kİ��w���O�,K����jr%�bX��}��yı��߽ߏׂ��D�\�S�V��
�j$RRC�6*[n��6�]:#n�<���f��"X�%�}��'�,K������Kı=�����ES��bX�'�]��9ı,O￹���n�-�tۛ�O"X�%���٩Ȗ%�b{�����Kı=��eND�,K��{�O"X�%�I�����iwnwIsf�"X�%��w��'�,K��۽�9��P��P�� �� �bdK�{��yı,}��ND�,K�?�I�i�&ộ%ͼO"X� 46'�_?�ND�,K�����<�bX���f�"X�%��w��'�,K��OK���d�f�.\ۻ*r%�bX�����yı,>����jyı,N����<�bX�'���Ȗ%���~����ʏA���˻�ю�%{��=>�6׳�Q�΋�[��ۜI���:�%���yı,���ND�,K�ｼO"X�%��{(}<��,K����O"X�%��S�Lە�d��nl��Kı=�����%�bX��w��"X�%�}��'�,K������O�*dK��;�/��̗K3rfm�yı,N��ҧ"X�%�}��'�,~�`����"X�%�����x�D�,K��������K3v��S�,Kľ���Ȗ%�`���jr%�bX��}��yİ4��+�!�	���ȟ}y�*r%�bX����K��t�il�����yı,���ND�,K�ｼO"X�%��g����bX�%���x�D�,K�O��y�n�77r�f�=&k;�A�ܚm�[,����&��e����ә�f��ivn����S�Kı>�߿�Ȗ%�b~��n'"X�%�}��'�,K����jr%�bX����;&�e7��36�<�bX�'���r���]��,K������%�bX=���"X�%��w��'�,K��OK���d�f�.]��q9ı,K�}��<�bX��w�S�,~HdL�߷�^'�,K��g~���bX�'���oon��0�wK����%�bX?���ND�,K�ｼO"X�%��g����bX!2&w���O"X�%��>�ԙ�+pə��٩Ȗ%�b{�����Kı?L���,Kľ���Ȗ%�`��{59ı,H/�u=�`�yO��H�U.��N����n�Q� �<1�%1ɲ5I��g�]�gâ͓֝t)tq���^Ŵ�w�K�Vq�K�<q)u�-��
�'6���ָR�y�=�6��Uu�b�Gcx� ,z��	�� n K��-��<�Z�<�q�VI�'��܋��e�N����0��Gu�U�Z܅���bܴ`�Q$f�K{7E�Ԧ[.i�͈
~��'$�y$������]��vv�kݛ�Z�7ejqi@ש���]���+]�nC���˛��X�{�{�oq���v}��ND�,K��{�O"X�%������_�[�&ı,O������%�bX?M���3v��)�M���Kı/������ G"dK���S�,K���߯Ȗ%�b~��������L�b}߹��0�&�JM�nn�<�bX��ߦ�"X�%��}�gȖ4X�'��jlD'����$A��s%��\�\��$���w����yı,Og~�'"X�%�}��'�,K����jr%�bX����;&�e7��.l�yı,O����,K��c���o�Kİ}��59ı,O{�;8�D�.�������~�d(��6J�)]�y��ú�$ź���Eգ�ݎ�5ũ���:n����Kı/�����%�bX?���ND�,K��������*�&ı,NϿ��Ȗ%�bw��o���ww&[7K����%�bX?���NB(4Dk"X�'����O"X�%��g����bX�%���x�D�@*dK�}O�3nS��6ۛ59ı,N����<�bX�'���r%�bX�����yı,��f�"X�%��v�ᗤ�̙���36�<�bY������q9ı,K߻��<�bX��w�S�,K����oȖ%�`��w��f�72ٺLݸ��bX�%���x�D�,K�Q��y���%�bX��{��yı,O�=���Kı=���L��wp�ӧ����!	�o-�Ӻ�<qS���\����d���.,�v��v����~����{�?���ND�,K�ｼO"X�%��g�� )<��,K����O"X�%�I��f��n�6�����S�,K����o�r&D�=�߮'"X�%�{�~�'�,K����jr'ʋ����,K���M�ir��nd��x�D�,K�>����bX�%���x�D���H�U=�%��7�Ȗ%�b~����<�bX�'rz\����L��˳7n'"X������oȖ%�`���jr%�bX��}��yİ?�D�o~���bX�'���~�f�l�.�s7x�D�,K��٩Ȗ%�a��G�s�^'�%�b{3�\ND�,K��{�O"X�%�ﳲ^m�7%ڬ�����\<n��4��:Eg�`n�M�Ā�����:;7�)F^ﷸ��%��w��'�,K��3��ND�,K��{��~��,K���S�,K���N��f�L��ܙ�x�D�,K��{q9�#�2%�{�~�'�,K������Kı=�����'Ȫ".�lK��w�7Lݥܖn�7n'"X�%�~���x�D�,K��٩Ȗ%�b{�����Kı?L���,K���Kن�4�Rn�sw��KϔRA���jr%�bX��{��yı,O�=���K�� dL����yı,JO��nܦ��i��K�59ı,O{���<�bX�(�}�߮'�,KĽ��oȖ%�`��{59ı,K��=�Ͱ��h\ͻ��ti�;,k�u�WNH����z�|q�:�Pլ�5�h�n��fm�yı,O�=���Kı/�����%�bX?����@�DȖ%�߷�^'�,K��;eɟf�Z��mٛ��,Kľ���Ȗ%�`��{59ı,O{���<�bX�'���r'� ���n&�q�ߟ������1\-}��oq��K�o���Kı=�����%�bX��{ۉȖ%�b_{�w��Kı=3��&m�a�2��sf�"X�|�$�߹߯Ȗ%�b{3�\ND�,K��{�O"X���:󋅄)!I
H\�S�'�7TU�*�fm�yı,O�=���Kİ��@R�������%�bX=���"X�%��w��'�,K��?YDb�$�O�ۄ�dݛdܓ5�"J-rm6�R�Hޒ�v�k��N�0�f�pu��;K�1V�rf�u�u����H��'Y�ֻ^{��G1�9.K�^:�O��MF�x��^�,�a���x���nm�MĞ���^�p3\וK���]m�b�la�a�;�S�[��u�Z�`�q�\&��IN��ky]�6�N�����n޸ K,�7���m�͛��s�<����/'jq��k�rs���{;@u�0@چ�-a̓�IYe�%1��ia�'�,KĿ~����%�bX?���ND�,K�ｼ���dK��g~���bX�'���o��i��n�sw��Kİ{������"dK�o~�O"X�%����q9ı,K�}��<���9S"X����nܹ4�iwt��59ı,N����<�bX�'���r%�bX�����yı,��f�"X�%��=����tۛ���fm�yı,O�=���Kı/�����%�bX?���ND�,�I�;�;��yı,O��S2}����%�3v�r%�bX�����yı,��f�"X�%��w��'�,K��3��ND�,K���V�V�M<�n-���\=[�L�s��� ]`,\�v��÷���F��|�f۶�n���%�bX>�~���bX�'��{x�D�,K��{q9ı,K�}��<�bX�'�v��ݗ.s.�6jr%�bX��}��y
-@��H�1(�b�@R��(|�"X�����,KĿ�����%�bX?���ND�@L��,O���a~%�ɚY��3oȖ%�b{3�\ND�,K��{�O"X�"C"d{�MND�,K�o~�O"X�%��gr�p��]�f�3v�r%�bX�����yı,��f�"X�%��w��'�,K�O���\ND�,K���e���i���6��Ȗ%�`��{59ı,?�߹߯�Kı=�߮'"X�%�}��'�,K��s;�v�l���3tښ�I��r�yu[���:�j�\-L\]������o3v�ɦK���٩�Kı;�����%�bX��{ۉȖ%�b_{�w��Kİ{����bX�'��zf٦��0�ܓ3oȖ%�b~+\�,AB�&_>���� �Z� ��,��/�"��f���{9=^��`�x��Pq���p# �"@�A F0b�#CB�� b<�ӫ'�=�~SЃ �c�1���؈p�<V�at�!]L�#N�#`B@gUS� ���J��ێ��c���J��n�%���b����~D�D"y��1�8��E���F ���@��P��Q	d$�W��Ӏyֹ�=�u.�M�� �����>J��UϿ|`���~����f��Vr��8��wD՘��8�DB_-�;��}�M�Қ��bx�&HA��C�&��k�{
��;��������l۱������=1��vQ�������ߖ�u�4�J�� �;��>�5��y(�I��hN�����tL��?�y#���_'�ɉ��@�gƁ��Z��� ��hw�n&�1�X��7�}o� �S��z��%j IBK!P�P4@{��g$����wf�r<x�`�Z��� ��h��9ֹ�?�B��o��n�J���M� \�vٌ68��1-���6�5��m�4lf�}���l�K����x����w�S@����}V����'	!$�@�m�9L�����}8�]����YVA8�J%#��~w�~�����~�M��\���p��LE]W8D(��Ӏ�^����K�}8wS�J�\��$�E]� k�x�	%�������78$ ��{�!.�ن�Y�e�n�d�6&ݪۉ���X����i�>n��wF�����sX-�H	��slh�qmI�9.�έ��fټ;s���ga�\;���cW�ֹ��'>�9�9+�s�u��^�\F�sV^�3v��H= ����ձO��Jq�j������r4"U�\���:斢'�x-��Xrp;��9�s�+�Έ�38LtF��ǽ��w��}\�KWU�-uƋ �<�5��͓Z8�v(����������6�\q��������'��:��@�]�@:����[#h��,RLi�@����v� ��h�lϡGЪ�<r�_Yj殕*�����7����z� ��f��������MT]U��t(�|����u}V���V�{�U��)�wwx��0J�}?��Wt��s@����?��x�R	Ⴢ14�=6��#��V�4k�f�e-�v���e��N�@��'���ڴ�Y�����-��@�U��_ab���Z���E ������;��I޳�@����Q�YE�4�L� 5�}��:D)���pu>���V�(DLX�L�ɠwt����������|����Z��T�Bn�5ֹ�>Q��� ����)�yU�N"RLP��7+�\ع���O
=�N��4�*mڦ�\�<x�`�Z��Z׬�;�S�������p����u����
,����w�n� �s�~t��B��L�rK��s�p�I�[gƁ������D	��s���Ow��K���b����U]V`rQ��[��=��8�n�>�Q
[y��ҝR_`�c���7���V�w��wJ`u�p�]���q3wEU�]Q3sw�:��窃�Q"���}�BkQ1�t{#�[�O����EQ�eʺW*n�U�*�t����we4W�h��h�j��B"bŗj��ݶgB��S&�>��]Ӏ��?�(���=��W7!j��Swu5f�O� ����P�������r��Ț��#�-�v� �7x��0=P�_$(HB����qE(�Bϳ��N��g�}�*�YRQe]� o��舄�y��7�~Š~�ՠ{���l�R7ywv���=��$��V�kdz�W2c]Zz�@a�S $�rM��4Wh��ڿ�
!/�$��}x��t����թ�N��@�_U��f���L�G(������JQS5Jj��=��p���ޜhWh�֬{G�b�D�9�w��{�4Wh�>���^�_����5�N<���d��@�u� ���?:�8�n�P�������n���~�o�o�:�H��(��u�YS��qtN�;\��͵��\
��v6.��1�\�4[[L:��f1*�݀�4��8��9uҎ�L%�h%��ђ�����I��Iщ/h���(�m)y��
Sx��t�R]�3M�A��\wnz���yS[�O�G��3�e'p<���h�V�^H��q��";tq�:����ZNUG]�J�}��m�ag!��j�L�O6�\\cU@0�>�/	�O+3���������Bms�T��`}�=�`d� ���p`r�y`�&����̋@�]�@;��wJh��[�GsB>���&��]� 7�x��0�B����Ӏ{�~�J�\��I�ffbm��r��?:npu��=.V�,18����'�ܫ@�]�@;��wJh�
�$Q�S�:;u�m�b����T���iKɮ��˛i���p����qd_���w[4��=]ʴmX�,�"��Ȱu��(���Q0��R[l�<馴�ڴ��<�"&$dnMwm��4��g�]Ӏ�^ o�;W5!j��Swu5f(J�_.��]���f��Қ.9��yY8�9�h��hu�@��M�ܫ������B�e�T��ۖ�$�Q��Mv���V7#>9��J���1����(9�w[4��=]ʴ�ڴ��EuLN)���nI�wt���%2oW.��]Ӏ���r�P�SW7V�U�5f�M9�?:np�
#�@��(�A��(b0F)Q�C� �'���?��O����9!UY��(���qdZ�^�}��~�h�)�z��hڱ�YFQVw8����/���������t�ڴ]�cljI�L��I1	��r�a.����8�����&a5��zF��)r�H��Dŋ$�ܚwJh��Z��_B��}׀z���HZ�jT��MY�y�Ns��]Ӏ�^����	%	"�V<�#������̋@��n�x|��m��r��=�\���Ȑ���hu�@��M�ܫH��J��~F��~��I=����)��87$�;�S@�w*�?Wj��f��P�$9�HHH�m�D�'k�����1�en�!5���М�;vN�	N(�,q��@�w*�?Wj���G���t��T��M�]�j�W�L�"`�[���=�(�;��eخ���(�
�� o����=]ʴ�ڴ
�YbyDZ��uWxB��q�oW.����	(�o���WZ��*�XJ����*z&J�0�-�����
z�Qq��H#C�@z c���t�B@0R	T�B1�"�hu�\A���f������z`�	��9��R�<�"qj�VH,m8�8x�I��H�P�X!=珍�.-��n�y *N~x��<W�&H�$1�d�b>@
��ǆ� �(��ƣ/�BX��	�=�;{�����w~@ �l9 �h
6��^���U[UR�&�.��U26��j�`.��7T�c;l@9#X�-Ӓ]�m��q8�
A
���;1Yًai��n5��Yy���vѲ��QS���*��s'qY�H�j1Z�sֳ����e��S���ڹcD�a���og���<���q�^:�L�Su.�ݶ���*iԚ�tU;l�S��.a�A�΍�a6{9*��!���vy���	<�O+r;v����5T<�=;w!2�m�f��U��iݕ��L���C�:�`���Yɪ�J��m�(��kq�M�2p���ut7Ӟqd�n���_&6�g6t�����<ݎ��\�mϥq7 ���Qɑ�C&긷a�[gq�t܆�ٹrq�C��<Nժ�ڪ��bݶtX5�aVC���ݲ�r�'P�ɐ:�0qq�v����s��]GC�D��2����B�ƘQ��[m
8Bc�6�u��+�d7i�ѱ�n�U��ѝaַf:C93n�!h����`|m���7��e�t^��N�e����]V�N��s�j4']�\������b���a����N_�h۷m�ו�7�,�����&����S�DV;H6�6�6�u��8�����:�&D�֋����F��-�lkR@��\�n��p�HN;'4:��M��`�`˯\����BX�5�z��̥�'۬��9]*l7@��]�a�څN��k=��մʙ�t��kY�0A�vbq���q���Lsɓ�L�`��Z<�b৶z V@.�V��>l.�a�U���@m��oP�S�Rj٥Z���	bT`�zؽ�!�n��K; �<�ѻK�*�V�t���k��m�D�M9ڞ�ۑ[tTn��������:�iv��V��;�н�20s8�ZY��ͦA6���r�Z�j�r���;dmm�q"���$p�m.�V�ײ�3���(~;��b� .�P �EĊ ����.M?)�$�*��p�������I�j�S�<�^Yu��M��r��:��Z��pl= �3�B��E(�x.�@.˶�4���n=�bI{��g6��v퍛��9�0�U����z�z��ۇ�nӝ��:���*��ں%�;�p���; �+�vm�.��C�L��(�Y�Ӷ�T�*�u��y[�)/B���2M�ڃ[�����Gw��׻��cpwx%�����Mv&�Y�to'��G��yn���{#L�#k#�2-�;V�w7x��>Q�(I/P?����ԓ����6�4(��Z�l�;�S@�w��79�%�M���:�nK���hWwl	%�06T�L�"`�[��I�ت�n�J��j��!N����=��8���}	$�����:�=��r�C����V�w[4��=]ʴ��bc����Œ&�Ln��\����{kո�M��fn����Ŵ�.�w����wVl�G���~ �女�Қ��V���V�W�,O&)�	�]��l�P����$�!BX<�����s���r�	L�ޮ�sJU���܉�h��>Z��Z�l�;�S@��1���6����̋@�]�@7[�wm�	%;�˧ ݥ3�W^�yAȴ�٠wt����Y�?:np�DF��t�\M���S)������v^�ɦ|9�δֵ`;%�i�\;}����Iꈑ��6�rx����ܫ@�]�@;���\$XcqG1c�N��V���V�w[4�ΈIL�=)�)�uWb��*���Ͼ��O}�w�(��$��Jh��Z���?�����8����l�<�8B��߳�@�+�g�'�İ�"rh�)�uw*�?Wj������c�s%�uSU������<�a�/K��˝��SZ,�..���Q��Yj攫Ua*����Ӏ~u�p[w��A�0�:�9](�x���̋@�_U�m�{�4��[���H��/���bm�xE$����7�l��	)��˧ �S��<��EuDH� �MI4�Jh�:v��[�o~�|����؊`�h.��AϹ���� � � � ��^�f|�m��Lܷ6pA�666=�~>�|����﷿^>A������>A������N>A����{��p�i�����4�l��˻"�4�0INۂ�,G_����sþ���\�c���l��\�3M�?��`�`�`�����x �߾�x ���}8 ���^>A�������f��)7-3d���� � � � �����ȏ� �� �l~��N>A������?� �`�`�`�������
"�A� �l���?��viv�fmۛ�|�����}���� � � � �����A�6 �#r9����A�6667�������lllo}�>�n�6Jfn�f�>A���"��A��������lll}�߿� �`�`�`�{��o �`�`��(\������� � � � ߧ~�?��s.̓7rL�o �`�`�`����ׂ�A�A�A�C��������A���?� �`�`�`�߷���� � � � ��	(;��;w����o����.�)dz����먞S6ġ=���SVȭ,�N���5��ڡt0��,�%���zt�R�-g \^�\p��e�v�ٝ�2಻,������Ev�;g��;	�<��-֝	�K�'��:VI����w-R�����r�s[>�2X��$k����%B"�vL��ZN��l���V��K���|��A�<[v��!��W[��T7x�{��7��x��F6��n�9�^u���+nq&.'mt�{;a��ͪ�vu����#��Y��A�6667�����A�666=���pA�666=�~>�|����﷿^>A������g���7sd%̹ww��A�A�A�A��ӂ�A�A�A�A�������lll}���A�6667�}��A�666>�ײٟ.�͔��sg �`�`�`�߷���� � � � ��{����lDllo~�����lll{�y����lll~�ӹ���f���ٚm���lll}���A�6667�}��A�666=���pA�66�=�~>�|���������wvRnZfɛ���A�A�A�A��ﷂ�A�A�A�A��ӂ�A�A�A�A�������lll}���A�666?�������������T��z箼Q��'���:9�k��BG����rj��P�k�q�mۛ�?��`�`�`��~�����lll{��}x ��o~�D �`�`�`�{��o �`�`�`�{����a�l����͜|����o�ל@����	$���� ��h��=�Ȳ70n49�h����O���gƁ~g�@�<J�ن&�F�z��`v���ҧ�`:[V��*+D�	�ԓ@�t���e�}�/���4��@��ĦO�@���i3v��)tuV�;����[�K�h��;S\K�*[$QG�4�4��Z����٠w�S@��sx��$��s"�ͻϗТ�;ﾼ�_���s�~��'�$��4���٠w�Sg8F.D@���lή�Z��4
�Ybx�17N��R����Ӏ�w�ۼ �WX&�cɋ�7��V�~�� �l�;�S@�8���'&@-��.�O-�ٌ�'�W���Us�N�#:�U����ך�Y��7ȿ {ﾚm�@��M�r���U��14���E$�m���e������h��?ٙ��ؑ�䒪�#��mI�_�J���d���[TGL˲j���UtMY��%�_}�/� 7���y$��{��OE{!$P=Ds����{}����u�bqdZ��4�f���M�r��λ?����x�A�G'�7=Rh�7T�����b�]P�&Br���#I�}�}I��.�]L����� }��^��f �5V�~�f�W�,O'�cqɠo�ـ7M9��]�m�rP��=�� �	�&,nF�4�g�@?^�@-�h��
{�WȜl�8�V�p��x �w�n��%
{���h�I}��&�(��m�@��M�r� �m�r��[d���9�;U�-P�����á^ٍ �n\�\��t]�2I+���	�N\�lul���e,����6̜����m�a�:A����\��9����۳��O�%4�v3\k����Vz�Srm�%�AS�:�a6Ef��r7�:-/;v�r�ҏ���ǳ��8-ۧ�f&J�dQ� W #���f�v�P��n�@�z�v����5?*��&�7�$�s&�6�ܼܞ�6���:���.3�W��OS���=r@(�q�9�6���O��r� �ۿ��!$���}��uL�3��Su8��Z�U���@-�h�)�r��+���"��ȴ��`m�%
�"IUwu�`}_/� �z��I�id�RM �٠wt��k�V�~���WVG�'�Ƀw%������(P�u����� �٠^:\q��6���J,�I�5l�����	%��am�4n���fs�bj��s�'#n��Z��4��@�빠�y\K#q��c��~��� ~<W���E0'��Qr�׀{��k����(Q&�	/��1b��E$���M��0���}\�p��x��3.]��WvUSSwx$�B��q�>�]8��4��@���+�7pX���OD�2Il�����i��_���+<��-�u�����ݕ��psGYey5Е�s�N��w{������K�s"���h[f��ҚWr���'�$��1I4��@�m� �M9��]�BJ�:y�R�B��Z*�n�� z�]4�M(��$PE�!jB~S�xB��\�I���C�E�4��)B	��c$KJ�3�_���H����!eI@�	RcFIP�I@%`U�,�H P�I%acT��������$�x'" ���X�h$(��0���	�,�|��y�hA`T�B5b��"�daP�B[k
��(>)�8�D1�4� �����D�J�(�*��
�����B���*�(`��
��Az舄@R�/� ��p�v�PH	��U1y����y$�z� �Wdh��b��M�@��Y��]���������0��ɍƁ8��E��Y�m��m��i��Q�e�B���d�NqLQ�̸ѩ)�,������6�e�BT��IR��V�x�/E_����?��m��0tӞ_D(��@o���\�����1�0����h��:��h��h[f�y��W#n%"X�����s��w�D(����u��ŀ9�[T��*��J��*���DDL��� w^���*�P���|��~�Qwd��e]�7w�ۼ�Q
!.����w���p�n���j��]]�w�m�])$#N�<�����uWM��]��n�-�
d$q�xd����7&���s@��U���@:�4�]sh�Jԩ�����k����/�B��Po�}x�����w]� �.t����x�8�V�p�n�[w��Je�ذ�˧ ����˵JJ���ɹ���%�JO�����ʞ��d���%-���Wv�UT������Do_.������� �QQ	$Dz����1��I��w3wv��ĥR�j��0�Cy��s�8�lp�
�P+'3ڲ��4FZ��K�5��e[f�w��/Z.��n�`6���5�N�ֆ�[X.1ն�%ύ�����uѲc�Xn��:��]���s���S��fC��mMM�T0��'���6�e�C�4���i���B�EQ�獛\]Ӷ�[i�c'��zѯ���|�G�;����{��1��7$�e�ی�.���+�^��ۅ	��I��М�;8ѷ�,q�L�=��>Z��4����J/��ŀt��U'+&��J��*�i�d��t����eOD��z�j��aX�JI������	D%;�˧ =�׀9{N���]��]�BP��ߖ�\�p�nhu�@;��16LX��ɚ�4� �Q>��� �u���`����1��ܔ�,�$,�&]���w)�	����bS7P��{pBړ����s�9�u��� �m�~�ޮ]8._}ǌc�!����ٯ?�?��)Q���W'[�0ur���]`^I+Hؤ�X6ӎM��4Zi�B���}X �u��2�F���f�e]�5f%�����/� ��}8�l�/�S@����\�xF`���[Ҙt����ʞ���?���b�֥OS��z����m���k�X+u΋gn����Ŵ닿���>�����C����� �u��m��4��_�7�@�}_�#�0�7nM�t����(S&�r��7׀��}
&C��bl&<��9p�;��|��u�o�f~��͙��hzS@=�Β5��'ȴ�u��l�?wJh��Z�����x�8�	�&�w[xB^ל~z�t��k��[�=�7�g\��������:{.��&x��4V��d���8����K��vTf�@oK�`l��oK`�[JK����d�N��V��� �_��[��@���*�9�W �F`�*�i�f���%�3z���S�0?6�&���E�ʫ�����"�2�u��|`tӜ��^D$��ZP���3K�vh^u�x2, ��@��p`l��oK`�[u%!E�N4S������՗5�g��&�<�ܹ�QpY-Yբ����,\.�=q�B���*z&���t���� �]P�k&'�72- ��@;���t����U�r�n�`�8��9$��� ��x��
}T���Ӏ���<��V��I�m���u��=]ʴ��� �h������e]�7k ��(�k�� �u��{��j�}�*����b ������v�v�w���f����V����ƨk#�d��!u�	E�M/���6T��c�۫=�nXzԌ���R�ܥnb΋<��Gs�N�Y9t�Y[-Y���h.n���r�CQ���8�O6��-����pwGS�jK�d���Q�6}d�q�4���n�����%� n!��p3���IS�"���^�RTt�m���Th�n�`h���w���m=�_}E�G3�Q͛�Ļc.x����Q+.���:�����\��!�r7k�:^.��;��?���� 7[������!�\�pwtb��aX�RI������h��Z��f�U�^G�"� �Q�4ޏ��= ��l�K`:���	�&,ND���ܫ@?{���f���)���Iɉŏ�nz� ��l�K`f������`���7���OXy[��n/Z�=z�m�,�؍הb�vX�Qs�&�`T��3����%�3z���S�0ޖ��䒴���`�N94�빷>���y�*�.� ��� �n��e9��)��4Wr� ��@;���u��*���r�f
!̋@3z[ ����*z&I?5_��aX�RI������h��, ��w�tD%w�W뉚���Wu4Tɞ���f9�d᭎��Mv��%L��ѹ�5�.<�E�`7nO�{�ۚ��@?{������ ~��bx�cɋ�Uߘ������	�[7�|��C&FA��M��@?{����� ��F2)"+�%���4��Šr������q�rK��w�~��0:֧�B��ϵ��<�$�����`�N94��M��Š��hz٠_uؓ�(�utn�����n���Lu����B��ve����eǒD�b�MAH2F'��Š��hz٠~�JhU��+�o"�tU_� ͒�l����euŠ~��j��aX�Qɠ�f��t������޶hZ���dYcqF��=��@?z١��`�E+ ��
g}���}�����Ǔ'"rf�����޶hz٠{�)�r��8�B(������M<�f�c��Y,\c�����ut͜�SQ��I�H�LL�q6�- ��f�U��wJh���,=�\Na�'�W��=�)�Z����l�?/$���#�o�����jp��B�<�� ��Հ7S+T�&��#JL�-}qh�h^�@�u��9r�o�7����Š�[)Ҙ��WO&�~��<B
� z0Q= !��¤B@��--H�cp(CX$`��$�h0f��ňā)�B0q�A��ʺDC�a�FL�����`���RS����HJ�
j�)⿉)�+SX�Ax��b�D�RbBB�Q��c$����<�_���PHA"1 �wI�������~��6���m�Am��]6 ��]��UL�*T��d����ɦ��l���2v�q<��Q��8�]]��F�]:��iĦ���4M	�:��E��o�{����u[;u��=�%;1ǰnUhq��� s�-ʵ�e	�m��vɐxq	
K�A�mm�ɑ�)nK�����pAq�9s	3N֦�v�nω;��'��l��.Zڶ�W���Ga��ʹ^��n1�&�UY3��D7d(��O=E��d�7TBUU���ː�t����_��1���K#�+�;bY.�n9ܺ�Y}�u��M�;)�s$��.��2X��]ZL��;�yL�/6�I�]� v�=��nbz���t"혳̫�b'V��ax��m$&��r��:iAZ�zC��B�mY�s���*�+v��;��*��pn�  ��vmDZ�S���S�N3��ev�ch�hݣO:P�j�� �
��N�gEm��9�X6u�Zڠ���n�fب"�hۣ�J��M:�zKzD�L뜒$��i�N�P��G�W]7�*�!3^�`�j�&�6��$�6�J�Mո�f���be��g��ֺWw<۵˟�c��4�m�k�bVs�CǤ���ڧ��ز
;�OQG(�4�sF�8������.Ӟd��IL�\�e��m�Wl�#�����1.�q�+n�s�r� ���`p@ˤ���.�I�<��˰�R*ޝB��ZL����B��2��VtUJ�O���Ѳ�Հ:�5rF�S6��1luJW8�)�����*tF� ��ݫ$��Z�9�FF��l �Zd`Ci�		����U����������n�� 	7k,N0��6�t��Un�;1�:6`0X,�;u��tTX��+�0/�����/��[l�S���p����T� ��7V.u+F�{����)V���Z^C���A�֮L��H��H1��.�I���l�v�7g���  �A�M����EZz��5U��"z�z�y	g��7m�3m�˺i�z�����۶:K��3�/f�ի�͓�Uz�q�S�.mc6��[Rm'.�{Ev��n1�z1����V7���`�8�i!ѮۄٳQ�.��qk�nxW��ے�MD��NfN�o!e�&���ۄ�p���4�,6�t4���Z�J9�g��}���Y��E�n�G��m�W��l�b���0m@tӎ�;�Ѻ���H3i��fZ�m)���7�篷����G'#ͫ:S,�;{������q�&�gﾬ�׋ n����n�-��<Dsq��]����~�w�9z�?��!B��W�Dҥj��SWsWk �����7x}	L���w_�4�s�"Y124	�ۘ������X���DOu�S�T���di�N94
�W���7_~_���p����V�������ǭ/�5Ì��\3sn���gs^���FLj$���#�o���]����~��@��z�bL�q��ܗt䓽�z^|��6��+�
"!T����O��`��Y�29r�y�27�LX������@��z��s@��Š~��j��a�ģ�興����V���֧ ?y��*�ב�Ȳ ��(��=��-}V�~��@��z�����<�c��S����z:��1�Kq�ú��Z)Y�������Ǔ'"n����n�/]rI%��0�]qwR�&F�8�qh�[7�������>4_U�rgY��'&'�o}�rI����Ƀ�b
�D1>#@�i4Eu �U��~Z���@���V�L�F���u��G�I*o�|`}]�����W�~�Ǌ�8�D��'��`BJ!O�����V��f�5L��h��X���n�!�\UЩp�X���A�k�+.�v��w{؎���u=�V�~�[)Ҙ�p`I]���S���N%�W����Gu��;��޶hZ���q,Sn��]`��0�\��ID�����V y�;���j��SWsUfВ��Ӏ����u��$�(�Q
+v���:8�LL�91��~��@�(�����|`ֹ�5iM��&���&�Ѹ��\�L���4�ύwZ9���y:�B�AdA1���' A8��*�^�����0ޖ�ũ%!w~���
��UwX�m�>��d�Ӏ�נUz��bG}�,��"F'��N ~����Jg��V�w������d�"���7�~��@��z�Қ���?[��#��3�G/ r���ל~��N ~�w�R�w������O�o��gE:bkl�"�a%4�w�QyV�+����kU�.��ɭ�̊�l���r�K/n6��w:4t�bs/�~��w�^-��`�ݑ�4����t�cl��nG���3���ӛr��R8��9����{m��nmv���q����r�"�$��mù��VF�P3&;��&�Qۇ���c*c�����{���u���]نw7��줶�d�tu�S��!W#�]�m��v!��jg��n[��'��	+�`�[)ҘΩ��cɋ�7��o�31 �}��>__���t��S���Y12<X�ʪ��3d�S�07z����&#��"�1D��$�@��z�Ҙu�p?�Q(��}x˙�����8�CM�r=��M��h�[4
�W�r��9��b&H�ǈ17��lr�@.���r�k��y��ttl��Yj6;	�H��Z�� ��f�U��{�4\��5�y#8����]�(JT�GBK09�^ ���uZ�nhْAdMbq(����@��ه�;��p��x��ҺE\�S8�rh�1w]��;�~Z��� �[4�:���cɋ�7Һ&�%��-���.RZ���F�uB�.��.�2�Kd2�ϴnn�ፋ�.*9�il���9�V>�o�������=�rQ�Cz�N ��\R(��D�rhz٠{�)�z��@?z٠~^I+I&G#���@��ـyֹ�bD%䄈KE(�>d(�f����� ��J&�&�칒���0:"'z�N y�� �7x�t��UY���<��cqh�u��%�3z���]��)UX��C\u���]���싱�����֍�Ol�r�8�뛵��w����컪�B����N��`f�����&���IR�o�0c�7&���)�z��@?{����@/��4�ɏ&,NF�4:�8���IB��^�w� x�:8�LLPX���Z��f�w���m��J�
%�]<�8�ɶE d��rM �[4��Mε� ~���>�
=�=�uq7B�Av����s�	��v[�s��]I�!�����B�������u$��L�G�I�'��������� �[4�
\��W�UcetL'K`�[��7��/�7��$b��Z��@7��DL��� ާӀ~m�*�wb�14�޶h��=_U��Y�UkT��1�q���;��y� ?6� 7���jP�~����������+�N)�3��v����l����i�l�XӋ,��=A�p�avl�������%�a�l��ZFܽm�Щ^�rr�/�u�s�v��k(mn��W�Ξ�.��O�{�l�	��L0:��vq<XjG�m6Ľ��e�ٺ�k��YX��v���Q�F�r�`��vZz�d�kq����8`Ӭ��sӻ �6���U�a�[O�w>�{���ԇ߬�8�N�VZ��#GM��t�ƝjM&���s*.��fkl,��\�������}��x�n�ݶ`�m2��Z�Sd��U5f ~m�B��A�u���z����?�>\��H�7*��`����p`l� �%�?/$���#���qɡ������V�� �w� ~m�BP�^�^ ������p�cN�Jh�^����}4��wu�Ǒc�"�8��Ivۅ��I�źҲ��=\H����s��|Yk����eE��dyHq����� {�t�=���zq�~�}���pX'�q�$��w���� ���u�}2t��_��X�q���=l��=zS@?wY��f�_WZi�Ly1br*����3�[ �%�3���4�:8�Lo9�4�[4��}�}?�ύ�Jh����8��#�a��6��̽�}g�7��n3���'=������tcI��E 1�<"M�4�٠{�S@�Қ������I29 m*��`ou��;�:K`d����#����$�I�@�����w��QJ$�~ Ơ�@����� d����BR$BH�X�b'�( ���M:�!�CH5��H��SD�=i	F�ĉXB)��R	`������XD��H�%?[�˪@#$@�ҵ$X� @�FB#����$+��*��#	 p����嘀Y��?h���&�T�\�'R{���5=��	R�:B��xQ�C�?)���A�E����.+��X����`�X$l$��v��*)J@a!}��Y4N H� E� �x���<A1H���+�~P?"�P`(zB��N����"#Т�ͽ��v�˝%M:Yus%Z��0?�g���ou��m��B����=��bԱ��x�rM ��������sw� ~�� ��:ˀ�Hr�t�׵�{M��٭�Nl��Q�&K�^�c-m*Z{0qvs2��on�0�l�������xϫ�4�&<��9p�/t��~�f�_7x�m�ДD|�*�c��n�V��ر������4�٠{�S@�Қy�]dN`�8��6���f���f�Ss��D"��"��|H��A����Q��ƌ �I0L����'�*k"da0$@^�w�sy$���_|I29 m'���4�fs�����x�7x��w�&��\ȁ�����ٷO5�N��`�KU��۳p�sW<$�1䁏��a �N���|�:K`�[{���yT��WW2U�U]`�n�舙���5�� �^��=��bԱ��x�nM ������T�L:K`E%(]xq,S8�rh��<�W��١�/{� 9�qTT��Jԩ���� ��u�����w�{�l�2D#�"	�A �D	��m����.�)dy����h�0�hj3pc�T�XV@FK<N�bwj��봎[���!}��	t�S���[q�RR�u���\��l�㋟�mr�}��\�/lmpގh�m�C��������՚�6navZ}-���ai�,�d�ٛk��\0*b0`��Θ��ݰ��n�w7b�	R�mm�����&�WR�~�w�G���^n�������K�fB��ƲAv�kp���t��+q31�O	*�qb�5���m��������@��S@�^��<K�����su5Uw���?�Dɺ�g�V�~��@���V�L�G�I�&����Ҙl��;d����	ƉN!8hW��޶hz١�����}��E���4�C���f�l�K`n����d���;�HSj��d�:�vM�Bvh��s�����]��j�',�;Xx����x̋_�ﾶ�\�J`�[.���72��E]]U��m�?l(��DjJ/�!~���z�[��y��?K�V��2b��m�@���@?z٠��@��S@<z�YX���ɉ8�l��7d��\�"`nג�"sc�6ۓ@=�f��w]���wN {���	��"�)Z�7I��A���baM��k�g����b6N���}�U���uʉ%!$��x���r~���{�ՠ��@?z٠w�.)A8�!��*���] ݒ�l��ݗb����1��i��޶h�[��TaN1J���w{9$�ܵh�\Z�9 �'��mɠ�l�=�)�y{��z٠Uլ��1Z(�����=�l�:IF־����@?z٠{��F��?����Y�B^g���M�l�E��M�X馊���e�\�"dŉ�ۆ���@=�f�~��@����x�'�ŋ91'�n��l�03e���zSv��K���$cn=�����YM��^���@��$�$��6�R�;f����=>�X�,P�R�ߡ8����������R�q�C�N��� �����޾0�v�|4��hz��sɎ�=���g�*�z�Z������:H���x�6�K3�ȎeZ���03e���.��:yjX�Ğ�����S@�����>�@���jI*���<#F)�"�3K��	��ݾ�1}�ߪ�]��m$������$���ƈ��)#NRIn�E��B�*�I,�ᘒ�����i$�[�b��2<������If�Ēޫ�i$�o��I'������~�
���[���۞�k�M¥��ya9�I�p�avm��z-��b�4جz��q;:ݔ��j����@;�ˆ��+���c��:�en�Y捛���3̵��m6@���9��օ�bi6���Q�q�:]�m:� u�[T��f���1v��v;d�^�N���q���M��3���$r@WH&��۷D!��Vn�%l��%7&Sn�f��S�M�No�V�.���N׳\Cacm ˓g���Y��5����t�ks�g��n�������K�}��I-�&�K%�_ǿ{��$���5$��I/�$��6��ߒKz�	���}bId�i$�zg�J�����I8-I%�Ϋ��[����߽��ꪝ>�f$�J���Io��U��f4�i��~I%�v�K��=��]�pM$�K�KeD1z��^J�t�]��K��{1$����I,����I/YbԒ^~�0cdj8%��8�e�i�;;��t� q<'@�O7N��k�����J9��$�s�Z�K��bI-�-}�߽�IN�g�K��Z�QvM4��ܹ���o����x�RW�"J�r�����[m�[o���> �������:x~�@��i$�zg�K��	�����$y�]dNa��Yi�!�$��g��%�W�Id�Ē[#����䒐��]]אU"�ى%�W�Id�Ē^�a�$��g��%��T���b&I#�=���O�+.8.��Ꝺz*�2����6����&���)NRI~����$�˖�I.ޙ�Ēi$����x�E�J��J��I%�妒K��{1$����I,�ᘒ[*!���K�_��-���m����ym����yo]CPG��{���!��Ē[.Zi$�IG�W��<�)U�u~�I.�&�K'803e��!K�ߖ��ʹ�Jl-Z�7vU]02u���.ޏ�[%0:R?��W�u��]`s30�[��x�:ۗ���+:m.���壎v�{cvG�oG����:��7e��v摹�ۙr{����ʪ�����=�)�~\�V�L�F�*���X��������޾0��`�)��Ԗ���&��:!)�<� ��� �kŁq
b��A
���&g{��t���'w.L�幸�X�ݗoG��H�:�������[�]��y��ۮxQ<j瞍�;ɲ�j2�9%�b&��gGFX�vE�]&RUc���v�L�p���b��@�}�1��(�(BG3@���~��R{��n��o���P�OwvU���dŊHӋ@��|h�w4�]���Z����x�1a��z�~`v����d�N�0n�t�UhRUҹ����o�ـ_B�P�{��=��6I翽��'�
*+��
*+�Ȃ���삊��TW��QQ_�AEE�EE�EE�� RDP0ATB1E `�A�U�����TW�tTW�PQQ_�QQZ��� ���������
*+�(�������􂊊��TW�
*+���
�2���K~��:�����9�>�D�   �   C�             �|�TP P 	B(
*�(��B�*��  @J@(��A@�I@�(� ��� %,   �     � i�@�������,��:�yu��� �y���t�\v鳓�}����i^� ���/6���;��u��wy��\ jL۫k��i�%Y�^pAN�s{���۽*�w)����ټ   �   ( d ��J�o���[�nm.��� z0�9��*�ܸ\���=�Ӏ �J}۔�{��5�׶��]�� �{�+wy��u�}|�qΓ� Ӷ��t�:����7��*� }�	  U�P  G{�7Gm�n��<���}ξW�K�W���j���yc�r�0 �O���=�� W�5Ebj�,�Ҫ��T��t�SҔ�Su@uB��:��\���B��J� =�$( �     'B��Ezv�iW-B�e�UF j�X�      {        \� �  
bҩX �J���b ��x���m�� ;�U�޼�ŹK�����}� }ϾSɠ�}y�;)����^�% 
  *�d =�7��w���y5'K� �˗v�����x��\�J�x �yqp�M�  ;/-����_w���� n^ӓק�wr��\qe]� >�ޭ9r�qk��i-���Ҧ�*R� 4 ����ʛ�T�@ 4 �~=T�$�� ��'�T�i"Pd24d���j���� �$�R�� ��=�O�������e�y�����.@��j��z3��u��EEz����Q؀

��(����Q��DTVPAS��� I�BG����;����	1���0����l�)R �p4�B����v�fCѭљkh�!� ���0�e��]	#*I�!�D� AN;	1tPc.,8�L!�Ɍ������XƱ�	r��Z��#0�1�-�1g�0e���[1˖�7Ř�	JB��#�$4,�Nf����|v��H�C���% �p`�F�sz�X�F����#3[��z��Q��qѭ�{�^<�%�ٷG���:��h6gķ��H�bY�4����f�oF��:9�$b�5�6�kf��	��K���pфfi�K1���F�V����5��YQ����a��!s:I�Uf����0�3z6r?p׎���'l��h�c&8�� �}��9�:��Az�l��|�_��JU~���n+��^RhSK���6��i��'�i���Lca�c#)�%�`Xh��8����a���M�1M�H��dd���SpXp!����L9�� ��hٰ���F���"q�n�'Fԗ�7��0�l!�vI�M��RN<-<Y$�� ���N!
P8�2ɍ���օ�ƛˠ��dፎNca�,2�sI9�h��FLӷ�014,8��0	�!!�hVq�m$�ѷ	� ��'Bb&��#�B��\$�cc ��׈H`M�'35��h�͜�o��$f��.:-�if��x���'�<�3L`�k|��7�G�5��=�H�<	a �����֎o��%��I��	\F��9�Xh��!g����04n�L����r�觭&��];N+:��ғ��`S �GJF&��!�4� ôa�4�"���Hpt��� �F�<9�аѴ�l��dqӳ�  �F���Ĝt������'JÁ��)9L��p���r#[9�9�^{煚�������p1ѷ������?$��h6��hv������Á£Ӂ��I���q�p6N.�l �`�N�0\�Fh��Y�M�Y���'��Fw����<��?�~T�Y�s��{�=��^�O�r����؏�A.��&�"���i�j��<&`X��L�0d�FN�8�	8o�����\x���#<� ��Kd�0c4���c!	�ł��=s��M������h�y�צo�?o5�~c<��n��߉��_�7�[0���� jSH�Q����q�f�j�C8RY�	4�����3h�##4%��4�:.kZq]�f� �����^����RXO�u�����K4�is_�4~:	�IO���M��X 0�vhH6� ��[�l��I���D�&:4�����2Á�[��Zi�5�H���N��m	15�Vx3�8�A@F�/�3[NI	a3-ԡ�0�5ÄY�7��|�ޛZ4���X�|�.@a��ℰBBF	Y$ &qt�&��a���܁k[�$�h�Yb�b]�I�!	�
$$�:x1�6D��H�x~b_K^V&��N,�=9�у���*|���'���4��O# �o�,P�!�DqI0ӷ�Eh�0lt�c��qB=���b%�B�,[/ӬP��G��cc��G�h6Nknk�xl��,��~X:!8S�S��	����#0�J�2L]��0���a���3A��,2P��n+&�oW7Xe��x�T8A��͐bI�8Q�{4�a�0ԙ�e�f9�A�%"L4i�։�sͱ8Yc\�<���lSiJl<Gd�l�� $���Ő!�1�le��m0�H�*���IƤ�����#'# ��a���1	b0,I"��IP�$��a� ��,c�2&���%�	8���ւ��<lu�ִF:4Y��Úo,,��#`�!��G4`Ή���,�Vl(	cyf �畦�k6�<q��!���5a���<xN@Ӂa�r%c4��ፔ����4�8�'#9�i����vHDD2�v�����,2��1`�4�91f���� �"3[��5��p�c0ű� ���!�*1��1?��j���4߃`z��'HA`�lԙ���z���^Fq�6�lܖ��f�"7.�0_Ǭ��@3dG�v'�FW�&.�i�d�o��s���k���k5��Z&��0fM0V%��4KH`L߷�As�2(���xX��F�m6h#1��@�4��7�.�����5��<�y�p#5��8oA�Q��05��p�nu��g30���7�K�Å����Mj��|�,"���#	I��Bp$�pă��#;	� 
S��	 ��	1#�1h%L8[�J�nxx����Iu��B0d!,��l��5��c?a��K|<㋮S
K�� D9bY���X##������3��< 1�A�f�04�a��~4x���Tsif�xkkqH�BBBsctl�I��u3��RL�
�$�p��0Ƭ3|��6��6�Y�21�,�M�� ��p4��ǜc|4�V���C�L,��#�q�C��K�`���I~P#Ӡ�N�h#|�5�"0u��s��&a���g9����������LJ�x��8�w�.����Nݡdч��8�t�����]$c�qa�f����H�C����x��hI���V8`���ȑ1�g�B��]�3`Y�j4�#y��i�La8FAĒK���ʌtae�j�� ��$�3�U��e�L��¦5xq�[H��i�d�X꤭��W�"4gi�̐A��H��I�<x�ya��Y�rr3L�f�I�a��`j��韔`��p	q�� �`��a�pf��H��6�c �l�c�����itl�vh�	�[�41���ӣ���h�స���dt��AF],a��BK&:4l�sF��[w�#{����9��w`�Zvi�wF`�k-�ښh"Gp�"�<!�x[Œ�,�0��N����OT�t~���I�N�f�6h!�0ѭ��Y����١0�sٰ���h04h������Éf��vh��ps#~h�x��pMr�5�cT�e�aB HL�:@��B�� ��HŜ	����\0�lZ�5��$`��c�����$ᤰ*�0d�`�tC�{��1���������t����?W��   �  �p�� ���     ��  H     	�l��9x��,��8�V����]7\U A:E��[�ѵ-+��pm�v�8�f�4�.j�BB@  ��-$8�okl�m�h���l    ��5��JU���q�� q!m l-�  � �� �m�� m�� ۶�l$-�m ekh
�h��8*��lH$pm�oյO,�P��5T�� ��{Ͷd�U�!]UA�*���t�+�=/��^v�5Id:GZkx��#4��@$Zi�f�	��fͰ�m�*�S�z�pU���@F��i69m�����	 �  8�n�խ�I�А�o$���l%��� ���-�-��ؓ�� � 6Ѯ�E�K.�e-�5���-� �)ٳ���[{  �-m*���  m�^�H�;l��<m� [@-�m�lN�(  �۳Z�J�Ux�W)-�k��u�[TD�kU���n��  [G/[�ǃ�  ���̀ 	�� ��Z�B@[@-� �["tl��   6Ƞ� ڶ6� �  �[�6[���ѶͶ��    ��    *�m��l��n� [D�u:�l	2NΎ��֎d㫶��� Y:�m   v���r�V�   kRsl���`n�k��Ԣ�D�L�T�j�Y痕jU���Vѱ�8�[%8ÒTUJ��5P]=����.�x\]� �@@��8�#���]���D~H��,p@O*���T��WUX��m[-�m��i0�p��ޫ��kIn�s�� $d�� �` $$�UM��^'H�1˶�s�H�h�`m���� �v�m�A ��� p�    ��gN��Z�r�4҉�X�i�l� �@� m�d���    �8H  � �m.������NCK�v��5��0	o  $  ���  ����۳d
�v٪�8w(�C� �m&�m��88z���ܦ�q�&f�3��n[צ�A&,�ki	�ɀo%ĳ���V�nH��m���5�栣��\p[}�*�Z[���k"5��z� 4���` 86�ܐ[G[K���[@^�l�U;�b�=0u*���; �����n�H��m��n �T�L  d-ɱ���6�@ �m-�j��@(��^l3��m��  �m��i��I�-���` �� ���@H $����T�::�U]���l�� �`  l����t�i0��H����W`���U��B^Uy`%Z�����6h[Cm�6�t�P�$h��d��oIm���7m�LĀpHA9u�YF������iIt� �`����k��z�� H�H�  m��m Ă�KW:.��5l��V���RZ�V�� 
�  $ ��M�$�kee0a��RE$��cq��6��m�6� -�{�y��jY�m���[7M���ݶ�Hl�
���d�
nz
�g���� � ��pu[*�V�j7j��M[l�/-�xv����zڪ��l��$h�	�ζJ�K	,kD�e�n�r�� H^�)@�� ��m� m����(��-*��;O9k���}�� �v$�ե�2��]mu'd��-�`m�	��9r]�6� tZ �mF�n񽷳������`�mPR�;ih�gj�t��m 6�!��$s�5�������@��\�z�h�� �  ���@�"�T���Ͷ[[f� m��p�A��8m&ֲڶ�H$Āl�  ֛l�qi�CUknݳ�Zl :Fݲ@[_l�ilp�����   d��p h�i��He��6�͂Nr@R�K@    ��l�l  $k�Ă���A�m&�L�$�W5�i�d�֤^���ׯ4��	l 8�l l  ���`l׭   m��|[@��Ҥ��m�Ͷ6���g2p���t�� �-�l  .�l��@  [@��V�րl& 8���ml����i3�l�6�m]Ap����Ӧm�`l m�m��hm���h ��m��n�H:�7m���qNh[)ۂ� �`l%��,��h�[��l $4U�0N�m^� ���H�ɹj�V�Z^P *�������:m�`�Iv�t�ݰ�M��m�H����V���'��m�{l�u[��֫���:%���m����{x�V���F�bBF@ɶ۶�O���i0��E�M���a��D�S`�[-� �`�h6	Yp ��h��a�(�I�r��L$�m 6�m���#�i��8@ "B�jڪ������A��yض�n�A$rmH�i�\�J�N�mq��l�>�5�@	  ��tؚ[�6A:�.���� ֶ�$� 6�m�D��zk.�]T�J��8�sN����suQE�������7*-�5UG�*�/;�R����.�����Y�`s�-;kw'u�Np5\�@U�@B�ۧ�� ���v�ػ4ksK�K*@wl���ӹ���9Z�5콕�/-��(��^Ɛ-�����,Z���\�)[jџ�R�U]�vy�"A�i��g����H��T��NI����T���m�Hm�)�ֶ�kn��9��J�t�U@*շ�,��  ����6WK6�V������@Hl�^�¶��i�O*ձg�ӭ�W��g.��@�UJ�@Z$8��[qm �v�s[p   �X6�@���}t�� �`�uV�m��8Yڛ r�����UFl�=����Ү�PÉ  �f�� �6��)@NY8�I�� m���	  ���Hл�8�[�[�6�5��m�L-�|����֐�)�z�*Uö�䆎6��#�� 6��J���%�$ m�m�bI@7�`	8H7m�-��l �j&��-�� -���%�m魓�� ��U��$��=�%�T�3P�; �*�7j���l  ۳��k�Ͷp�� �R���mUH.�`RUZ-��  �m�f�F� p��aS`mjڶ�ӥ���]�%��[K\�-��mٶ�kzɀn���z�H�H��i<y���IÀ:�HV�M��jĶ�aV�Z��j��+G%���m���`H� �i[�-� � H�a�!�� ����5�'�í��h ��m� -� [E�t��� ��f
\��cY:�5��:H$����v�I��i�ۧl� nӴ�����V�CZ ���� 6��� �     �� l �z�qn�ڽX	 [m�h�@�x 6�k6�-�s�ΐ  �Z��;n8I5��UY8�����`  l��3����|[@ �۶��À�Tڶ���-66�D��  ��   r�	m& �86֭�  �      ��6�jP/[#Rk� o��C�88*ڪ3�jh�2�@+*p[*�[ ��Z��
�l@   sn�-���Zɵ�"@    � A�ŷ�����l��M���o`$�:t��  "��m�6�a�i1����ŲP������hS[��am�Q�UR�;Q�@t��� m��� �m$���hӔm�l [B�Z"�5��I˱5UnʻW\�@��X�$��E1e�>�[:V��eWmm�5�nfL9#�r�����<ڶU� �`.�n�Hk�эY�kU1\�[ح��hh $e�#���.����V��ڀ Hm�`�m�I�� Zv��ڴ���Z�4r�!�UR��uӵ�mݳ[vn��  � H���%���� hHm�$Ku���z䀶ɶm��ߑ� ��   t���6��m���ړ���m -�H�M���'I6    6�AؒJj� �$  ��i$��m�H�8�BhZ��,��2ɭ4���m�KV� *TU
���T�Tm�Q���G.l�G���� -�ٶ�ͫkhm�'�o{x$ 㭺����\��j��-��M�֥`��͕d`y-��� �my�
�P�	��/7f�`������*�"�� ���AҎ(��������~ g� b�;|<�C��/��D�>�
!�v�����a��m�j��"�b.(��'�1P�����"l �P?����D=EW��P8�4�x���Q�2��T��T}TG���= C�)��"��b)T=D|�0z��z�&���PG�%Q_@6(���R	A���X U�	�IYh�d��$$HbFQ�ZB�	e �	��v���{P|0Uz�qN**z�ht�D�)�_� &��a�M�)����"~POM�hW�T>��/�z��PU����V������D���� pU���@WU}<��
����P���E���=M�p�*��m�<�H��"��Q�t_Ѝ"	���w����-�����9as[�skc�bM�<\��&��3�]T��q�7E�У�Z�/K��s�;g��3�D�Mn��n�6��ظ�wiν#v���M�)]��+�0����t5�(�`H+�Y*ˎ��{-msCi؞[�{X�uۭ�|�K+R�i&FEn�A�Q�-�Rm&X�3��;L;qтU�v;��K۝�a1�7a�x�����U�E��s�M�'�<��[]Pr�]jf�UB�m�-����!5]l&ݳ�^vc��X��T���Ca��e��6��9��F#c`㍫TP�s�q�]�'.���0pv�\sܻl�A�Ӄ�2���>A�[���n�1��j�m�e��@�R��]ϙ�lڛ�w���ˣT��v8ڳ��%�Ӻ8nت��ȝ<�hd7��#çf�`v�ZPr�A\�iʲ�Wk�H(M�r ���*�Y;	:ն��L����Kr4��zhӥ��V�d��,��b�%�m�Nм���F�Be��v.h�.��u��gqm�[bݰl$�8�g������s�]�=]lz��E2��mnW��m�6n��'��nS�H�s���5Ϋ<�A�O��:�����Ur=F蕵���m�aj����P��pڇ�s�f��C�7+Ek�i�id�';8eʠwTgq���ΰ�`M��j��Q��p�;9�֑�O2d���/5����%E;K���DGo���]"J�m��P�]OK��[o,1{���i�6�1��9s������������tF�U��L�:�vˇ�m�q�<����^��i�t퓱�l��V]t�u��[s�,�,�A��4b���5U�:6�F0��clěNn]����-,j��v��Fٷ:��n��q�P0���`�R�w=͛��b�@pHRN�З X���eے-q�m2��C��_;;E�Ӱ�A�^��	�rtŻM���و���W��w���0 C23,, � L$#1�0��)�� C���v?
�������w�?��գ���u�tƳ��Í��6�C���뗎����m���-i�'���\�H�0�N[<�8[�XN۝&@^��XzwE�A7�஺�20k��`��cn�5�lܣ�i�R$�I���4��ۥ�C�C���x]E�v��e�+`��:(�#�
���ŏm�ó��os�����}x�a�fb���TV�������p`p<��9���Q{���G�l��n<4�&��X�~,k����G�w&������������"!~������L��V�4����.J��˙��۷����D(���/�ԒJ�ߧ����v�I}xvbp���<i�=�$���RI.�g����v�K�v��$+k$�G�j)��MI$�����K��jI/�ۇ����RjI.��[sȦ,�<m��$������q{�Ie&��]��C?��~e���K�ל7@]�F�xN��.r˸`��3�=md�-�Tl���vzF�-\�`v���eT`Z�m����7T48m�_�nݩ��>,I#~ ����Z p=U,����׬�=��Z�u��Ģ�*��`���3w]�S?uw)�7��z�d���b��ܚ�٠{]���S@;����fLd��7���$������Q�I*`�4k��c!#s'��!����9e�6v$���ےӞ.T:�x�%ۋ���NR�6�-����@:���ۋ@�z�1HD���(��f�u�4k��ץ4���s�(T��n�75���T�)E	$� �8(�(4�*�� �2�4�%��J?~���`l��X�3]9�#NL"�I4���ץ4]k��f���kq�DAG��f����,�ݫ ��v�[�lDD|���m�8����d�'�lr��m��H]a$H��b�l��-ݚ��ű�qrU�@]����o-�`Km��<px�Ǎ���Y�}]���)�r�^�y�'�4�""�M��6n=,�P�vw��{���9يd��cJxۘ��S@�־U{��|�G�Q�LDa	 $� q3����*���q�$"YSp�9u�@;���ۋ@��M�E�&L�Ese��:�9�;������Z]�x���܎�E����,j8)��n= �hZ�S`}����6w���g:r4R�90�6��>��Z��h�נZ����Z�Q���4�~{��l��KS����*�1f��F�&7$4]k�����Šu����fO �51�r= ��D%����{�Ձ���`lD([�"
�!�	�0�y�W�:han�k<u$l��/�v������d���jwM��mwl�"kl):ò���{Kì���\;�zl�}1i笈t�nxT\�l5���X�s�W%���Єm �ۧ�Nݩ���HݛX]���A�n�p�����Ŝ>'����ѧ�pf:�d7mR���%�S[v��
���ͅ��K���!b1ԇ��ZukbwSNn�����e�^����#�3�m����\tl�\�ay����:ɺ�m�f�R��k�H�m&������Ͽb�:۹�r�^�u�h�9ّ�4�Os�-Tۥ��q�__&o-�`M��@D��xI1G�Z��Y�}]���)�vwG[�,jcǐ$\`��o-�`}b�l��	�Dƈӓ��M��Š}zR���ڰ�5�
[�[��9N�Kd8ٶ܀��f�����n�RB=���ƛ�.� 鎩�M7$�]zݻS��~,	�^0�T�����;.��8��ʙ��,�ͫ%�VG�D%bIj��G��r�[�7+9M���zX�ř<� �51�n= ��@��qh�e4]���vc������9(S�>�6�>,�ͫ �r� ��;22C��"xۘ���h�BP�7y� ��v��6�gUjUl���]�낵�z���k��"2�H�ř���brl����r�kcVIᮆ�l���*`}9nkX���"��4J�j�&�`���$�d�k�-���u�@�8��� AӦ���T�n=,��J!%��DBJlt���s�7��Ꚕ�9���m����x`��;j`}9n- ���
`�i��[4��hs����M��uĒyQ�k�+��������7)g��9}s����{���d�2Lx9�4���٠{�\4�Jh��h�Y1�j7�x��4۰?en��BI)�;_���>�w�L�ڶ��CdUR��U56g/�T�;�S��sX�iăG.G*i��a��D�n���ay��9\�PՇ�P� ��z]��.}c��51�	$�����r��{Ud��t�.#h����īq�ݍ18���6�iv�|�rdס���=�̖X��r9۫lH��'����`}ڨ�;%L��0,��8�U*�.z�����訪��`��4zˆ�w�c�Lm"c�!�vJ�{*`}*�0>�T`}��2y&0j`�rh�u��e4~��3ľ�@���F���yj�L�T`}ڨ�;%L��0g�f+@T�м
�c#̍'2#$�lf5ݩ�*��^5ΖK�T��rt���D��Mۍ9a��c9H.��!cv�K�!=�|���N�6B���ݻ6��`�=l;�D����8ӣ���6�:x�/����͌ Bv�5���=�M��|�1jy:�6wDqي�M�:��[.���C�m�gaJݸ��(������j�a�r������^�wq������#��s�^��w[:�c�d�t\<Ns8ۇ�E�ݚ��m�M��c���m�/��"��� �T�'eL�T`z��H����wY��Y�{�S@������뱩�ȣ�O)�-� ϳ]��u�g��S?v�,-�4��Q�<plRarI�{�Q�����T�'eL%z�/��`�V��o���U����/�,�L��hBˊ&Ǌ	5<X��xES�p����"�!������bM�{c�o�֚k�,5s���q$0�S ��0>�Q���M�x�&Bb"�	�&�w׻��B��^���ʼ����٠^�dǈ���d��@������e��NʘfNU�����D��Қ�[4��4��h�kRIm��8h�k�:!)�����Ł�q�`tBS����tힸ	��9��G*�v��yɩ�;k���g�i��[�^�g�+L�tOfݮ�_�=��쪌ب�;-L	خ����I�M�&��YM�Қ�j`���Wi��5j������|Xٺ���}�T��  ���(�$��0��_��$��Q0$Қ� �� N$�	�������4e	��SC	BA����<�d�����X�`�t�|=��,!���Ev���D
!1���*�����lt�ꈇ���'�E4�
�	}�����C3���N��,�U:,�C �0	�S��0;b���Y�!1Sԓ@;�f����ب�$�0?�߹�/��7�nf�7.��F��b�Y�G@l6]^��O\%�֐NFӒLx�&@JI=�~���ǥ�fn����s���:"��A��!����;j`v�K艓'��[ۗUH������y��������ŝ3�k��ջ���Jr�MQO�@������L�|X_����X~ �?��G���S�M��*N`���&(��M�e4	��� �T�;��{ܙ�#s���%�GV��'��Yv�2��.�.(��z���lӖ��ԷW.���!�r������3���	%LvT���Fl�\�Q��h��IIS ��0>�Q���M�x�&Bb&,j`������>�Q����ISȪY��.n���L�T`}b� ���$�4���2C�� cN��h��%�������ٸd̛�۹��|3�n�*��s,ڃmN8^�u%	�d^�V����۳m�\u[����Y�S�ܴ�۵���D���Y' t�%�Gk�Î�w9��ٛ��!^$���%�eC��6�����ث�M[o&�qٱWn����5�շ�t�ݠ��gtY8H/7h�ۍ6w.�^����W�72�K���٘x5���b�t]V�1�s,kDX������
�_��V����]�5d�Ƚp�h6�7��[ ���y��k��$� ć0�~��hu�@�������gu���I2c��&%���U�Q�vZ��T����1Dܒhu��=�)���;*`^��qi��b�Է|�>��� �0	�S��0z��A(�LnHh�l����>�)�{zS@�+�ؚj	��=�8�n�ۥ���<s'�����Wk�>k���ZX�4Y��Xiē ��0;j��Қ��h�;2A��&�?n�.���	*���ŀwv� ϳ^�{s��!�m<i�@����wf�:�P�ɹ���|X��m8hXa�ł���;j`^�Fץ4��c�H�ɐs�h}j`^�FlT`����S�ʰwf�/Zi1�����=��%�u�n��[����* U��=C�v%f��?��ب�;eLv���W��L�s��>z��T�'mL��h���A(�LnHh׽�*����Q��UUA�r�)�}zS@�wd�L	��&�LvT���0>�Q�vژD�`�d��@��4�l����>��E�p���y9�H4���rM�!����t;)�6�&�y��(�㋗&FHx�FLbp�=�)�[f�NʘUFٶ\���pXa�jKm��NʘUF�W��V�`�����`���[4�)�}z�h�٠w�*N`�D�Q�6㑁%T`v��vژf~���7gmL��R<y$������w��s@;mLv����0>��2T�i�D4�v^�;�5a��t�F�ژ�<��`�9-&��7 PJ1�f�^�h�eT`v����U��79�8�`���Q��+�e��{���$,N1'$�/YM�Қz٠��@>��̌�m���Q�Yj`���������1OoP�&ƄMK�X���u����>�zXBQp��$��[�����N�L;�ĕ�n�X2��h�Yl�Y����k��d�Sm�Ym&�l���ؖܖ�/F�շ���e켔�ݝq�]��,�x��gr��}�v�赧&�A�c�L���GY�b^K�����:�':j�m#�/I48�!��2�����V�0�f���B=�
���x� �E�CL;�k�Y�n���p�5f�˂kt
�{l	m@kW/9L�]O��{����=���>Tv�ZS]%�"^Fi�Z�����˹�N��'t�U���S;�>��W�m����`YU�S��f}�z�Ɂe^���䉸�m�&�z���Қz٠�Y�w�u)<��?�������S ��0,�� �^&��Q��ܐ��� �������4WqfObƦrM ��0,���T`Z��-��]��r��k���ķ�:6�8��t������x�'V�U/]NΤ�p���YUX��,�0	�S ��ʓ��*UI��L�?n=/T%
Q
!(B���I�A�7��߹�s�S �0,���l�LhD�i�2�77]�}�k��	DL������?���mC"�nH�;�Sʨ���Q���ﯼ�X~Na2F�q�6��@�e4�w��~ ��v�ٮ��+�	�#p�C��6��X�9��7��t�Ʌ�o�JѺÖV�dc�l*NQ4���;?�s��37]�}�Y�}l��[����1Ȑ�$�?��	/�{����F��fLq$D4�rM ��@��M>���|즀w[4z;8�h��-7W`v���j� ���;�f�}s�s2��O�4~��%��w��m����\���H���.��/&s�DJܗ:��>}s�Ɩ;-ͷ/6s�̏��c�d��Ɋ8hu�@;���j`}b�d��.�-ũ�I�Nʘm�����KV��t*p&H��c�5$�������;*`N�=H1g0A�\?��y��^��;*`~��_11@$!Q�$� MᶔBQ�{j�>�ڗM	�2葪���$�0?�l�_=�<`}b�����)A�Hش�GJ��]7^.9������R	ʹ��:F�yW02g4�쩁l�X��ϴ��������EI�$ܚ^���>�g��7���gٮ�>ŕ��M1J�[��X��%�0	�SY^0=�z��2Ba�d�4�Y��Y�u빠{zS@�m���d�8�&ɦ݀gٮ��
"7��/�}�����*�M��8��IY{h3���`�"a�,a�pt)0�H �K�)$!���:04&�A��`i_��)#5S1�t���o��x�%�82�C$��
ق`,cô�V��J�\t��Rj����,�,�*0��˚(=�&��� Ě��, q�e%�<]2ca.e��,0cAi���)$����6
A��Te�0X��᠛	�F��������FAPX��Lcea��folE��7�֦{(�I[�a�"04���Ve0�,�D i�l���z��"b4���F��b��j[�h��:`��F��.mv��H�h,َ���6/��^����`p͉������6#��F~M���y�E�K�'������?�_��]���	��Ž�( �f�z0���#��L10M�a-��y����`���k#F��[M5�����L���Y���'	"�B��-j1�L����8fY�G��#,a�<6�&�$aH����6E�f���� 0�[+Z�Y�f~>�~V� u�-�[V��+\WFn�d	ݼ�tj�h��IJ�A�&ȋ[- iР=<�������8��6.h��=� vq������^����K.�Yd��f# N��z;3-�X�x&���Ѻ�s�1�V=�ڐ��*���6ttrmR�Ѵ�ܛu�N�
�"ν��l�����"Y����Nԟ?o�' v��m6D�GSf���F5R�����M���<	-�K��u��B��#��@���Ё!4�sh86�9����z23H;U�_\"4s"�>ݖ�s��N݄.��T�b����5����Ƅ�ר����ip�oXœ����;�m]�-�kF��@�z�flT����WR�B���.#�yo<��
#�ظ;c���;eحWl��ۅ��n����d�k��\�x�c�\��8P���tx6���5��(rֳ�;��eg�JF%��P�U: ��0��T��V�8
�]�98��UX8�S +��raQ�Ց�q�7�E���5���ѷ�qc8Fv���n�2��7& v��\���y�13o� ͵�+R�Z-�٭۳S�4uI��r+n�t�[`ݸw �å�8����뀣�����|N�..x�q�%]��[�WMcX��+�/)g4�Jm�v:��vnH	q�T�'!9ƺݬ��Y�xr�K�,(u��n�ʛ��ҽ��h�6����Y1���$H�lO<yv��{Z՝���n��hO<6�un%���<����uF�	�x[�����7��OK'���S2�&�i0�Hm%�TT-�ݎ����I�eU�ܭ��=u�T/+RBm5�U	�eR�֞��*ٳ��h��9���lu0�5�q�g=\�g��q0gl�B��S��F!:RȐn�)3�Ȭ�qu�r�L�m&��V*�X�=Z�Bf)-�rp0���"��+�:�c>v4b�9�����'M�X#0�4�{6�1VE��J@tu?� 8> >�� <<�)���C�{֮n�07�������P%���X�H�n�$�pm(rj��6�` rc�x�\���/����=�K9�lq�tF �����ی�$��Ѻȃ��\�]�=�3�t���b{*��:��J����������:	2�@t�<���1t��O8HCj9��c1��7@U'���vlx8��N�oZ8�G����Ւ���5'q�.��]�>��ҥc���8����=����z�sd��ϝ+��"�uȹ#��ķ���%�$�x�튌YS ��0/e��� �.Z�π����(Q2���7;����j�7s\RG�i�29!�z� ﭚ~��]�zՁ��Z�?)�mS���S-R۰�;�����`}��Q;��@����c��lBN!)$�:۹�~P�3�������]�Fl�Z���ڮ`�a��1F��FԬ��x�p.z�.¥8�n8y!"&G�̆,Lɉ)3@��w47u��n�$���u��uM4��5l޷��^���8��:�+��D��f~�`~��V�nھP��˷�Ʀ$Iő8'$��ߦ����������8$Q�7iq&��`w��`ژ{�~�ٻ'�����MP9*��7v���j�:�4ﭚ[w4����lx�)y�^�R{N�ۀl1ese�Opsd�v���y�Q����xL�9��٠��vn�DG���V�sNmS����Շ9�&�mL	mx��ex�&��Q	L����IԺ���$�m��֬�͵f)IB��!"���`f��em4SHN��̶�:D�o~�}�&�mL.m�����o���o��c �q ?�L	mx���w4����bJ9䌞8�ț9ٰPoY���NpkD�nH�/hw����V��u���$�ݵ0%����� �٠}�B�d�'��#�ɠ[n��+�m��}-L	�G�F,�w�՟���|������0%�s@:�qH(���㙠m��7]���j�*IDD	X��͵`b���I��I���@����빠�4��17'!�,���3`ճ��=t�nI����n����z�˗#��5�`�rM�w4���[l�z٠\�\�̆,Lɉ&Ձ�fڿD$����`os�7wo4�uU9�91x&LRL�m���0-���W��V��ķx���I�}-Lmx��� �٠w�*N�(�$�M�w4����~����; ����_�A
#ݏ�pm�?-�n�,8�K�c<�헭[R�u�#q9[�j�˽Z� l[��Ǔ�c�ӣC�m��*�v����g�<q�h�'r�����7l<���r[@F0 :�����e<���\�5�<أ�t�r[��
ץ�à�^�F:x�Fܺz.3�^=�nz�ۛv[��,�h��<�
�R��g���D�ʈt�����>��|��lַo{�PQD���k������5f�sjv���8�9t�'	Em�uղ%�MU)�#M��W���<���}������� ��v�7_�%������V��S��:N�iStՀn��IL������V�fڿL�)�9�NfF��h��v�w;wv՝9�֬��M�J�<�G�X8��@������ ���>�v���Ë���n�,`w��`ʘݵ0-���o���c/�:�e:�\4C�:ȵq,[�=�n�7;��ΗI��Yn����;~��b�X�-�0�j`[+�{+��cS�6�H7$���k��T��w6Ձ���V���С)�3_L�
M�t���n��;��X}�j�-�4߭�}�RsxțO&�ݵ���V����ۮ���J{7�f�_߿8��#M��#���@�S�w?�voZ�>�6Ձ�N��Ҩ����N�Rs���n6�P�����y���Y�Uղa���q?��I��I��l�/ex��ex�/eL	bڳ���~����WL�^0;�^0%L�ژ�9�0s!�2bQ��>�)�s]����
!%vf��`}�֬�ᚩ�Sj`���Xr����`����͵a��IV��x�<��[�h��U19l�m�ٺ�IGv����|X�f��W���ґ&��	�"OTu�����rs�3��3&�4���r*��=@���$�q&��`vUF,���_���`vo\�4*T9��MT���o>/�DL�����`f�ڿ��
���N��:N��F���`�y�ٺ�脔)���Vo>,����NT���-SM�yyD(U[��;���9W�{�ܮ��(�&��VϹ���;�_�<�G�X�b�I�u�s@쪌[S �0?��~��n�乘z�����e��^�
���v:͔ñ��v�nS�@F���{��v~���7[�����~,7u�ٺ�%�7��X���s�b�L����u�o�������`}���IL����KS#u-�t�5M�os�3wmY�IyEV��� �{���ǳ4j]*i���L=�}�}�	|�0	mL����6�i��R扡��7v��ϋ�w�����`f�ڰ"%IB�\B��{���n������۪;n��n�;E����)�5碹�Ճ-���c�Yt�uS֨��.t 3�;-�׷M�uv��#�����"�/��TQƴ�]N:�	������G�̯#�s��p���9�U�i��2�'§i��Ŧ��7Da���8�[� �� SccZ�f�u�۷`�v�963��R�͗����݆�՟�w�����~�ն�;7@T�v�ĵ-����釲��[2�zHv��%�ہ�na��m�Lm8P�~�@>�f����ؾ���ĉ��`�q0�S[^0;*� �����m�2E1bq�9&�����٠u�@=��\�̆,LɉG1��U���j`Kk�sd���#��&&�m��[4��hu��?�癙q�	4Ӂ�2|�i-'^-��b\���m�]T�<�rT�J�o�50Y!$y$�nO@:��4��`vUF-��$Ww�9�h���$�q&��{��eT`ژe�@��TqQ�73�-��@��~4[S �0%�� ��.,_����sx�-��vZ����U4�}őŉ�����٠u�s@����u�h|ծ,����t�nn�x=v��eM[�v�¡]eݰ0Yꑼ�mI�$Q��C�I�u�s@�5�`�������[]Mᒷ�,�\X�쪌[S �0%�s@�u�����17 �l�/����?�C2K	D��J$ U�*э�`? �Hi?oH��E<GbI��`���LG'�)�Hb�XD�5D�0D��a�T�@���H�F*E��$�,�\<N�i�D��LU0�MSL e�K�`A$�T�k��q�C`:y*	��~ G�*~Qq=\"���� x���k����*���*�[v51!�8�Gܚ�[4��hu������I�y&(�̑-\I�,��Q�K*`���|T2x�$k$Ȗ%�����㝞��TXF:��u�����i���h[����w���|�^���j`K+�������	�� ��hu��,��Q��oaR���oXUM7`����͵g��Jg;����{_+2d�?b�q�4�w4ʨ�%�0����g%�`L�qa��,Lɉ)3@��M ���9u�@���R�w	�X�&&�JD�R�Z��p�|��mY������z+O��n�3�d��4޳@�ֽ޻���h۱)��L�<���&�˭��^0;j� �T��+��ģ�2Hۏ@����e4�f�˭zw]M�OQ�73�-��C�<W������l��mx�-����nji:�e�n�������Õ~�wەi N�D@�$�D������,�T�C�4�@���4��B�$!'�9Z�q.��jj���:5�?nK��ɖ6��k&�-i�ntrJv�D��s틝���,��d�I�Ƕ�<���^ۛ.�E7g&݊�3��W<i��y�*�����A�.�t�s�[mB�*h���ѓ�S��j�\-��+��XĂ^5����\��鹻J�����q���,����uӏDg=�ۂڎ�zcPÛ[<7k��{��=�6�uhӠ��ͯ�n�]=%V3��=����
��0���:�85Ë��Ll���^0;j� �����m�2D��`�z��h�)��4]���:�0S�,LɉG1�����Sl��mx��m�����Sp�m�.��۹�}l��o]�Li�y#�n&�o���U��	�&~�C�K���83�rH�����R���������\[�n�\6�|��<`v�Fm��6[����jiT̵ST�9����|[W��D/���v������7wmXfX�LA"i�24��4]��۹�{l���/��8�"bb�1��Lݒ�m�NA I"`}"�c�ҁ����۹�}l��[l�9u�@<���!��HU�\x(�ڸ:,R=�����&:�nEY-�7G�H�%<��̘��4���z��Z�z�hb��L�$��MLM�@-�0&�x������0/mkvcO�#�$rh�נ_��i��.� �W	�R�`Q���k߾��*�{߷ʽ��Ts�#�JdQ��~빠}l��_���b����o�M�OJ15�v�~;��'�y�g{���ݼ�:��&ǋ1O%2#$m���ݵ��=f����齻6��z��l���*f뎉L�74� ��vNnՁ��k�=����\W��#�Ħ,j`���9u�BS'wu�;����ۏi�N�YR�����V���ٳ�DL�������ڷ]53I:E	��MXtBJs�t�=�VNnՄ%�"�D~�S���>S�:�
`TԵ3OXm�`{��̼��>��ڨ�o��7�'lu�.o5Уۛ%���]vyqȻ����9��W��k�ﻻ�_Ir<^Y�"M��_ߞ���s@��M�mzwJ���9$i)q��w7��
�Q	U�������VNn��ď����ƒSS?�n�z���@�mz.��m��mq̘�a2jZn�͇�"S���`l�uX���9%	)�}�`b�ӛ�J�jUKET��l��	mx��	��03-���m���wl��ϦěM���A���4���Bܝ������W2=��f:7��t�s�6�[��j��"F����7;s�'.<��<�L�����S]9h��A��i�����{c��:6ܑq�aG ��7K�?=�y~�N��C��OQY��h�n�)�!.0J�I|���~�h�FS,�ԃ���NC��vϷ�]�nv���e�3?�������ѮXkKvYuvw�ٶ֮�]���6�Fu�x�c�L2��ވ�wwM4�e�!T�*�� ��֬��h�k�9u�@=쮹�y�`�j\�VۯK����UFO��:{ޫ36��LS�<�
r0*Jh�!������oJ��U��jcO�H��&����b����oZ�>�zXrJ~��w_Ki�)m�IH(��@�빠}l��궽�Z���o�^���"��c�1��l��f�5��Bֹ�b�Y�LNё��w�z��E@�)�S?�7(������U��]k���CszՀwwS���9r-7T���^�o�y�fx��+�;�ڷ�$v+O�8,JbƦ��U����u��=�ՠz�W�{_W2diA�I�Y�.0'ex�����l�`M��{�]s�"��1��>�ՠz�W�[f��u��9wn�d���((Ա�ŕu�����k��GWa6���=�#S$ x���Z��z��h�]��ڴ�]�cc�1�(�I���l���������=W��;�U&D�I&5HIɠw�w4�6ZJ��/𩈚��7;����s$��(���f�Z�~Z��z��%;�ߕ�gwS���9R�Kx��e����y|��UF��������͵gb��۔�������;әb�����̿��}����nsx�������`IUm��k�d	XL1'�}�s@��4�l�{+�cO1LɈ\X���0����'�������w+��<��I�@=�f�}m�*��{Õ����R]��EW�dDDY��~ݷMU��e9n�T݀}����DBK����wy��ۺ���]�`��dl�I���1,��<l��8�A�
�oap��Z�QV+��e�7RL	%x���0���vژ��-�iU)�?��կ�n����Jd>��`����ݵ}��gwS��XDF(�ӆ�_߿M ��4�ff%o�ۚ���@�_qdpX���0m94=	(���v�u�3^�P�L�wM�ί��,�sqɠw[��fk��>��`n�2!�	*D��D�L)�� � ��x>����9����<� ?)��ЇP��Tv"z�,��)(4 D�DC$0̤�$2IA0b�`!��� ����fl 0�4���`��xA�K2B��ZX�&�v$����,�2� �~,Y`
N!â1�Ć�nބĸH���(2L�#-�a2�xh3��N+�����hm[D�Ƶ0ՠ�� ��R���5�J�!�uk5l��Y%^U���{/etk=�.S��c=�����rb$9���S�;:�K�8�`�`X�V��κn��Ѱ�$�QJ���&c'f�[UOh�n�\�saIj��M@��JS�K�k�tăIϠ.� g��>�m�T�hun=���a����v�u[S^�����u8dslc�}�� ��#��B��R�������K��I�tr@8�w;�=��k/"i.؊k��\v��F:wO\7���ڢ�8eB{��=�،+0z�(
�2T�.5�:m����`W�z�F���ݶm�djX�vL�[&<N0,��yK�Ђl����M�y�R$9�v�lcr�����ܵ�J�uni&�J�uõi2g�{Y'T��-� �!�2'G���Y��� [%��kn�\哂��5�;lshEP-�Im�Q��/^�Sݪ�6��rE�f��v2�PmK�Yzݍ��h�`���3���꣝�q쫣�sÐ�u˵�M�\�V�m�pq����j(���<]�2%� �営d�]�p�ҧ9�p��`��1ͺ-Qr�LgC�6`v�M��ml��Rh�Ӆ١!�$�L�c�t Q��;{L��)�m�.0�8���p������
�L�s��6��1��|^n���]�6nv6��j��R�v�����V�㍗m�i�h�=99�I'8��ۭ1�q�� p[u�H�\m0sY�+�ݶËkql��R�
U��.�m�lt�1e�on�/�n�`�#t�S-+W&a8�kj���
�HS9�e[Wc8�T��`���Q�=U��2�-eQ�tB�UХWSǇhy�9-�=s� ��Sq:񴻭g�Y�v��w(�5.� �[3��Cq�4<t���mUW�&]�< )�m�*�sI�CP� �Iۖ�L���U��kZ�[�zބA:���
!*�z
��Aꟑ È	�UH�*��Y��k05��dF{m�A�]����յ8���rH����3�ʛA:�u7�61,�٢��|goeE�pqgL�9��ؖϱ��w7-ص�����5��k%'U���X{2����w!�ce�=!� 1����PZ7O\8 +!<��juu �jcv�ca�`����ʷ>@��b]��	q]dU<.�8�9�rd$�Lڤ6�'���ޖ�'������5�=:2��[v�aV�1�M �9v���`�-���{ݯ����{��u��\f�,��v��_�7{�X��H(�71'����j`^��%T~�������Z��79�C��JH��~�4���u��*�^��ҩ2'�I1' rh~��Ĕ��~V�>,�ݫQ����v��ALo#x�?�ջ��o���*�^�}m��w4{,F��5c���Z����h��/pX��t;w<�md��BIU;���S��D�UL�N�U�vژ��%T`w7��pF�h��UN���w�TB�	tR����Vw��gwj��������MJ)��t݁��j��ץ��g����3�~���k��S�bQ��;���v���ja�߷���6��$	j���&�`l��X�;����Ձ�e4�u%&<Y'�sRC'j8��v�u$h j�L�.I���t�eU�.\;I���q��٠^�s@��	/}A��z��~�ӚR�2f�M4��׌	9n�.�x�;mOۥ�Ŷ�j�GH����~���6sv�⁂;�Q8(��/{��~��h[^�0YQ� �8�?�y���{�`�y�����ݛ���D&&)�6����@�����z���Uֽߙk�	�S	�DE#Qz�p���m�����ݲ5!��gv��:�z���#K&,Ĝrh���;��@��k��;��ܧ��sIKTH�:���ݛ铧{��3�����j��&MJ��$H��8�����@>�f��ʫ���X��M���nZ�%R��i(���Y�[n��;V��<�?�������}��W�w}�n�h���8�@����v� �l��5�	B�N��T��R�6^���Ѹw<�4�U�Y���+�d���T�BALm
'�����~���h[f�}z�����׮dő%�4���~�P�K��7��`w{֬��V�ؾ�Ɏ	)��`�rh׬�$��=�g=�`��`}bڹ�\��3s�9�I&��`N��`���,�{�$b�5�s4�ڴ���;eL	-x��Oߥ��N}�9��8�u�Pf�uc���-�6���i���5�%�4�\bvm�O:Ad�ֺ���+���{Mv�L<��:ų�����`�'8�A�[��M�-��F�jx�Ȝ��M>}M;�%�pQWcd���@�g:	1ۀn �F,��F��w�r-��̞0ts�7�r,��c7n�u�}���u�[b*� MHj�
%#�Z�_�ӧNUUMKB��9�-��\%�7NT�rjmqkn7>��7c�{U��KM�m��h�s�gs��5���~�����@�o�cİ�/h��`nk�B��&�u�r���>��~S&����� �`n�Z�;�j���GZ�׬�;�"`��W��Շ�wt�{��ۚ�����k�2b�J1���}m�DD�o?�owZ�3�ݛ��kN�J��3$ƫ��C�u�MeY��;�qWbхx�:�r���7�x���`�rh׬�:�ڰ3�ݟ�P�Т�{�v{���5��i�&�u�o���@7��`n뾈����T�4�I���,`[�{X���j`Kk�)̝M�m��4�áDD��s�����:۹�w;V�m�����UT��� �w]���������6��h�\��?���%�,��H��\��qGQ��Lq�Gj�y�Nβ]�hn�Ď`� �������w;V�}m�СG�;����Ҧ���TMù�π�����S �0$���33���"Q���馥���Ӡnìo��a_�� B�Q�׾��U���f��?f�i�CSD�UM7a�B���&�����Xm����j�	s]*���M����I-��?�3�����@<�b�!�s$@�.ǎ�ܐCI��7%��5�%�]T��=t��Z�h�3�q��s�h�٠[g脿HowZ�5N��ln`����6����%	L�ws�7��X��7�(��J*��������ӘuR:��}�����'-�-��$Wx�\��h�`i��Q;�ߕ��]�`���DD~�qU���`n�J�jJt��5�swk���6�����3�������.��x�`�)�ĦLD��K�����J6�yq����Z��@���8ҳuĒ&7F�Z�٠[f�����B��Hn�t��7�8ja��Z*����u�����ݛ ��w��/BJ!U�s�Hn�ЦJi�:n��{֬�ݛ<�L����3����ql�N�Ht*���MXz!(����6�����vJB������;�ʚn`����6���I/$�"+}�?��{֬�ݛ��BI
!�ª����Cm��$.�v��.-�v�Ƒ��g�nJ�A1\��ܒf:Dv�J;8����h�S<X�uë�ݶmÇ�nč�	���W�]Rq����C�lp{A;�:�ȣ�8�d��,qc8WAn�c��3�V*����ô`��=�]����j�yc��:s��z�R\K"I8՛'��k�:�]�X��im&k?��{��{����S��b��eܜ���l�m�=i�����w`�	��� �����v.��#�n�7�����j�̭��Q�~�4l���<$sp)&��6��IL���6�����w舅'f�t����N�M\۵�����2�4�l�:���>��n`�H����X���j`K+�ٙ���ߖ�غ��y1y11LRM ��4�w4�j��f�|U�LM���9M�����ę$�O$�{Mm��H<ñ�e5��f)��L$j3Ȝrz���N[��*�>�'����p��%͝�5�5��[9W���u@�AY Q%�!%�����;w���fڿD%2l��*hM��B�Nl��v��?��J��s@�����l�cm�b���n�>��`gٶ���f�СG�V{�vx���i�i�Lt݁��j��Fk��ws��u��eR��]��kg��n�by��0½A���7l[b9i�!r�_�w�������댝s������ ��?��X���;mL	%x���
4�����@=��������/�����)I����ג�����)JR��s[�L54KUUM��!B>��p��'��v����2�$�#�:f���I�Fb�I`� z�t梖 ��T"P�B!%غ6�}]��w,�N�l�:#@D0,LL����ĄH�����H�x�P��
s{�&��$ښM������@�%��CA�v�#m6��^���4�.�<x�P�̪�� z0=)Nw[�qJR���ݏ%)O;���kz��ɩi�:n�Dy(��%)P���5D"S����R�����ǒ�������D ���n��̦T���j[j,�A	��s�R� ���������D#}�;�A�Fn�QdB�������uCu���L��%�#������v�ۭ�n�M����#��ZK��T{7����m����ǒ�������)C�{ݧ��JR���8�)C��}��f��l36e�k{JR����┥��v<��=�]�qJR����I��x]!��Թ��� �@�~��%)Os��\R�����ǒ��>��q"B��*i�*]S_��|��)_�0�k���qJR��}�ǒ�������	�HD&�jUy�s��ǒ�����浺޵e�Ӫ��� �@�7u��!B>��p����v<��=��)I�'{���������Ӯ+������b�Ж�Q��������9�_����_}�=��ֳ[����.�}��)JP���c�JS����R�>����R���w��N�jfj���۸�f�.B)����)J���JR�����B�BJ�B_�朹�t"���oc�JS���k�R�>����C������o�R�=��<��=���Ml��x�Z۬���)�2���JR��w��JR����JP2�^��q"(��n���D��Z��6��JR��{�)JQ���߾�c�)����)J{��y)J}�VA#�%%��OL��Q$��ܺ�M*��:5Ƿ6��a�7j^��zK�&��kV�<��������AQ#�n��*� Z}�.66���_9a67V�M ��$v�糌�6;,-cذbtm순�֤Ҫ]ú��Ά�c9z�9�	A�;��̒z9���O.����y�M�{;9GWd+l=5mՄٸ�YK� k=ك����Xќ땚���x��؎�K�W��K���-n32l7�6�ar̥*�篷�9{穬�n����m�v�������)�{��R�>����R"�A��k�M���U*i��o�%)N�_}�R�����ǒ�������)C�{ݏ$��0u)���꺦�Je�M9SNn!B�y����w����!��}��)��A����.�rQ-MT�j,����~���JR��}�ǒ����vn!B��E�"����)�-ff��Z����JR����JP����┥~��%)K�{��JSow�����S�ynk<��Y�� ��t���
\�Gc��u��(kY�-��j� �{1�k7��%)O}�{�R�����ǒ�������)C�{ݏ%)Os�s��F��s+[mky�)J{��y	�TC!E�+(!���K߾�|R����~��R���w��)�
7w[����.$��uM��!B>���(}�{���d�}��gA�F�sQdB��n�T���Ӗ��o5��JR����JR���{�R�����ǒ� $����|R��]�ä�Ԕ�M5��;j?"�}�qJR��B���%)K߻���)C�{ݏ%)Op�{U�Z��홺�;c���5.5=�.&��^4k;NM3$�q'/j���<�m#{ݷ��w�����<��/���┥��v���7���[��7�!,F�9p���jkY��y)J_��w�)J{��y)J{�]�qJR����I�*���[\�)�)�
j��n�D Q���rR��������P��c�JR�����)I���v�\�K�.jGN"Ȅ�BB����ԥ({�~��R��w��P��4����E�"�l�ۘ�
pU9┥���JR�����JR���ݯ%)Os�{�)JRzW�Nٛ������n��'%�u��i+Z�c&�RZ�g���<J�_����i���^��r�kc�){�~��)=�{��)�~�u�)J{��y)J{۽խѽ�{���0�k{┥'��v���$2S���k�R�=��<��/����B�(���A�xt���T����m�>JR�g���)J{��y!�*�){�~��);��my)Jy��\�&�*�U4�j�\B�
3wZ�")~���)=�{��.*� J�ā}?>��"~^��\B��3�����%���ڋ�?w��R�(,����)Jw=��qJR����JR�~���ݚ�T@ֲ��Ú��km�ƭ��}��]Z��F�9J�8�㛖[�{���ow����R��?w�┥��v��g�JS��s�R���������9�y��Y��%)Os�{�)JP���c�JS�}�8�)I�{ݯ$��1���4F�1�l��{��l�{�O����k�JS����R������j��Ӫ�T6�QdB����� �)=���R��?w��'��C߻�E�"��ER�M�e6�\�w�JO{�v���=���8�)C�}�ǒ�����qJR�n�Gޞ���{�5��u������nh�����S�-w-��(��2�^���)�ZF��
t��%�!ӷZ�u�2h�8�s��a;;�%x�p�8�α��e·��lH����n�y���c+�Uv��-�z�rr��5��C�Z�D��(���y�bs6\��a��;�Ըz�����jم�L��d�8��q��qD�l���uA�������דWI�7��i�ܴ'>y5&F��uL�u-����|�������o���R��l�5������k��8�)C�}�ǒ�����|R�����k�JS���t�*T�r:�sq"(��j,��/��w�)JO{��y)J{���B�S1!a��K�4�-MT�j,��/~���JR����^H�"$d�{���)JP����R���;���fp��f���R���'~��%)N�_}�R�����ǒ������D ���k\��T�9�8�!)O}�{�R�����ǒ�������)I�{ݯ%)H�];���������mrUa΋ps�sr��S	=���nMص��j勛�Tx6oe����������c�JR���|R�����ג����[�y��|[[�o26�G��%)K�����U�GN�)3��k�JS���s�R�>����R�i�ER�T�[e&黈A�n�k�JS���s�R�>����R�>��q"B߳e���#uT�������J�@�������R������c�JR���|R�����ג�������,��L�SNn!B��E�^��o{��D ����E�"�[�~�m�v�����HL�./BMӹX��k��rt����7i��]v0�g[%�+\^�u���5���<��/��w�)JO{��y)J{��┥��v<��?Oڵ�T�)Īj���q"B��q�������┥~��%)C��w�!/�Z�2�p��H��rR����┥��v<���)H��1�YS8�?�ƥ/7����)I������?g��5�5��Z�k[�)JP���c�JR��{�)JR{��k�JS���n)JS���ƛĜ��6H��4��<��|R����1����k�R�������*��E�"�NN� Rh)��U�Q�ۉļ��˼���1��=�:�^u���K�l)T�'-��li�n�D ����,�T��{��R��������R����n�D �ٽ-����-��5w��)O{�����~��%)K�����)I�{ݯ$�U�%;��k��D��U20u4ˈA�F�sQdB/������I߾�k�JS����)JR~���٬#e���5���<��/���┥'��v���?{���'D�a`dS�[����ǒ��'usaCR�J��j[w�!,��%)O��}��)C�{ݏ%)K����D Ifɺ䦩�M7!-�Ax����nL�B/;��m��0u;se��a�fn������%)O��}��)C�{ݏ%)K�����'~��%)Os�~5�5���f�qJR����JR��{��JR����^JR�en��.Jf!,;�����$�K�R=�{JR�����JR����^JR���{�R�����ǒ�����Z��)t��6�M�B�D!)!ow8�")�u���)J{��y)A�,��{�� �A�z[i�N���t�����?JR��_}�R�����ǒ�����|R�����ג�"���,���`1��O^[�+���9�\Y��C"Ai��?~ٵ	�@@�	2b"�]$�D�R�~PL�D0� �D�$f[ ЪyA$0��I,�Iѷ�%��ŉ�"�cJd�!�e ��6���~���� A?'���
�<1G�R�a�|_�/�7�%��0�)$ �1q�3-)� I4H�C�9�
���BL̝>�����iʹ�[G�m]EQ�9�Nv\�06ڸAu[U�]��Ŗ�� /*�U�>wm�v����ۊN�Y���i�F���]�v��	���{o@�`�bJ�͗����E�A
9n�	���u=�I�^έ���$N�� ��X�a �k���ZlqSv��2^�Ϡ�x��Z�K�[��M睓b ]:���2��Y�sn���{[�;F�����Yw��^{m`�fz�la��wh�-]v��:E[K�NM��T6�Z�r�=v��A�Q��;Dm�n�>��VC�8.���e4m��j�qvJ�U�iA��7fd0��N�|qO ;�e��X�25+q�#��k��g<�`�uuçg����B�;v�
o�.�n8'P�u�'����h��Z�lqط�r�m19�l��ˆ4�G��5�gZ�\l�F�m�^i�zU�e*��eW[cxe��g�	Ҹ�綐(�UҒ�zRnEcH���*���D� �J�jG�^��<&5�]u�.�	md-�C�]�2��pȚʶ�qnW[I��Аհ8�YL�.�]iqڭ�e��-���n���\�f����դ�H����]9gb ��;
ܢ:�����E(��겒i�G��o"��ʓ$���'�g,L%��=���`C������<�;,$<�^23�*���l�.L�R�x��E��ث @.ܨȉs�7m��1�ѦPg��ն�Ů��i��)��� �٭���+�FN�F����h�p�pV�����(��g#�����0�#q��ݬJ�q��d�eZ�k�lW[UP%$��z��c��Z�r�S�S�)���{T:մ1��r���T\�T�K�fs[������Қ�i�ջrg��I�2p���%�7"*�3��E��]G
�m>_	���`�vp�������@�P�,�Zɗ��zwh�V�޳-�5��~ ��?��(@P�X����|UU�OȂs����n�j�ofkF��M���aڶ�jx�+��vWZS�FҗX4;�ے�]�9�Y�f[G�n\JB����/K�5�� �� �=��{ <�3�!���:��)�x�e��څ�W�yq�.�JH<tC�������/��D��7[���S�8�ծ(dwn��ݩ�p����(n�lgs��Z}o�i��yH��뮧���w��}ޮ{�xv��炶��a�m:Iݛe�z��\	=�vi�vm������bΔ�u�k[��R�>{�v<��/���┥'��v��� 9�R������)J��ާD�M�P��M6�Ȅ���|R�����ǒ���u���(}�{�� $9)�=��{�[3n������)JRw���R����┥��v<��/���┥'��u�R9Nf[�SC��Ȅ��!
k��)JP����R��{��P�¤�!ow5D �Y:o*h���R���o8�)C�{ݏ%)K�����)I�{ݏ%)O��}��)C۾ڵ��I�+y�u��u;1q�Z���؍�����lv�b^���q��w{���-"��rjk��){߾��)=����R���w�� �@���j,�A�M�r�t�[ތ�������JR��{ݏ#��N����~!䧝��)JP�����R��{��|
�b��{߳{ټ��\�'Nfe�D �Y����}��ǒ�����|R�����c�J\�k�&
5���"4�y�����<��/���┥'���JP|��/���\R����������j�f���ǒ�����|R�����c�JS���n)JP��{��)�����鿿��*t3�觶��XgsvnKH2��:I}��!� eH?�{��������uÉSM9r��!B]��QdB��kۊR�?���y)J_��w�)JON��bȒ�F�Ng�y��g��[�R�?���y)J_��w�)JO}�v<��PXrS��ߍ�o7f���o8�)C��}��)~����h�v�A�8�rw}�ǒ��}[�q"(���t�jeM8�5#u��%)K�����)I�{ݏ%)O���)B ʀ�~�����R�]�޷-�Je�Ji�t黈A�n�c�JS���s�R�>����R�>��q"B߰�U&�MP9sN(�mmX����O<�qW�5�'����Y��r�{�������i�R7UIә%���6���)C�}�ǒ�����|R�����j,�A�wj�K�N�T�U9���>���y�!������JR��w�%)O��}���	��'�{���6[ժٚ�o{JR�����JR����H(�d���\R�������!B�?j֚��jB��N[w�JO{�v<��?{��┥���JPA�D?��<_;�߷�)��ݚ�*Y$�.��mE�"���┥���JR��{��JR!f�D �_f���ScuM:��}$���x�y%�=�����ۙ(�*v���-��AM5T7Q*�8��\B�
3sZ�")~����)=���R���wۊ�!���˗3S*iĹ���Y���{����'~��JR��_}�R�����c�>E!�N�}�7��Je�Jj��t�� �A{y��!���{�R����w�%)K����!B[�l�Ӗ�K��ېt�Y�O���)JP��{��)~�����$����Y�!owU�i�P���o-�Z�qJR���ݏ%(����}�)JRw����)��w��)JI�!B@��c��F`���wA�}6:x���[p�;��:�� #s�7��jn��j�����N�g&�:���۱śy�q��9�p�p�#kv��6�͒cvl:�c6�:�:�&U
�G�����v{b�sp\��/�D�Wݵ�x��r�u�sI���nC������G�o.�SNt�3��(�E[s��n��u.Ld66�n����7a�p������mR�Y��͈vê-�t���ys�M;`�yi�Y�\!q�f���R����o�R�����y)J~�]�qJR���ݏ%)O3�N��CRԅSN���!BY��E�"���)JP��{��)~����B�f�hԕ,�[�SD��Ȅ��{�R�����c�JR��{�)JD,�֢Ȅ�$�MU�J�N&�ͩJP��{��)~����)=���R����┥�}�o7f�,�:�D �Y9�W�!,��<��?w���)J{�v<��?�?���#����k��z�pϷIWe��:����m�T怣��r6�+��g��ַ�)JR{��c�JS�{��R����E�"Nn�� �A~͖�=��kZ7���ǒ��	BP�	BP�%	��s���(J��JqAD�>P����9�%	BP�$BP�%	Bf`�%	BP�7߶pJ��(O3�(J��J��(L���(J!(J��?k�}�<��(J!(J��30J��(H��(J���(J��;�~��(J��<���(J!(J��30J��(H��(J���ך���ݫ7�����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�%߻��	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'u߾מ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP���pJ��(O3�(J��J��(L���(J!(J��=��}y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�w�kz�v��kYl�k5����(J��(J��"��(J3�(J��J��(N�}�<��(J!(J��30J��(H��(J���(J��;��p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B{�����(J��"��(J3�(J��J��(L���(J��}��P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�^�}�f���-f�l���y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	߾���(J��0J��(H��(J���(J��"��(J߾�מ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP�~����(J��(J��"��(J3�(J��J��(N�}�<��(J!(J��30J��(H��(J���(J��;۹�7�h֮JV��Nn��z}�x.hR�%�z�q��<�Y{��gMQ�,7YY�������NJ��0J��(H��(J���(J��"��(J߷���P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�%߾�g�(J��0J��(H��(J���(J��"��(J���k��(J��J��(L���(J!(J��30J��(N���8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP���w�f�ozp֍����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�%߾�g�(J��0J��(H��(J���(J��"��(J���k��(J��J��(L���(J!(J��30J��(N���8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP�����<��(J!(J��30J��(H��(J���(J���oK�2�\P�7M�P�B�<���(J!(J��30J��(H��(J������(J��"��(J3�(J��J��(L���(J�}�	BP�%	�`�%	BP�	BRJ��'@�_�+���%	�0J��(J��(J����<�J��(J��(J3�(J��(J��30J��(K��o�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP����7�ٽ���f��޵�y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP����(J��<���(J��(J���(J��(J��(O~��g�	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	w���(J��0J��(J��(J3�(J��(J��3������%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP�{߳��oef�j������(J��0J��(J��(J3�(J��(J��=�}�x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�%߾�|��(J��(J��(J��(L���(J��(J�����P�%	BP�%	BP��%	BP�%	BP�%	��P�%	Bw���(J��0J��(J��(J3�(J��(@P�B+M��
i�H�sR�{f��-jT�'U�Un{��ڮx��۹n������֣{����ky�P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B]���(J��<���(J��(J���(J��(J��(L�~�~x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'~��pJ��(O3�(J��(J��30J��(J��(J߷���P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B{���ެݣ-�6f����%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	���o��(J��)�BD2{��lA�4>����"�(�>��؃��@H�(J��5�%	BP�%	BP�(,�q�SC���lm�ߔ P�B�(J��(J3�(J��(J��30J��(O�����(J��<���(J��(J���(J��(J��(O~��g�	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	w���(J��0J��(J��(J3�(J��(J��3������%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP�������{іo[֬���J��(O3�(J��(J��31��J��(J��(N�s��<�J��(J��(J3�(J��(J��30J��(K�����J��(O3�(J��(J��30J��(J��(J;߾ߞ	BP�%	BP�%	Bf`�%	BP�%	BP�Dd�W��(DBA٨Nf	BP�%$��Z��B�gI���M��\MS�R�����ǒ������)I�{ݏ%)O��{�R���L��k7��g�׋���w�ֵ�[OR�2n��e���v!g�^՗��}�l�;�[S]����J]��o�R������R���w��!��֢Ȅ4ݷ-�JfJd��k{���)JO{��y)J~��┥��v<��/}�w�>1JO��Km9qT����Y�!gWt�B(}�{��){�{�)JR{��cdB���Sm�.�������B�C�{ݏ%)K�{��JR����JP|������┥'�{���7h�j�jj��QdB�fn��A�n�ǒ�����)JP���c�JS���[a܈xOc���9�I�]���ud���<�=�c��\�:ͣ@A�cd�]�1�mˋtS��n0�ۮ�]��rX�X^Շ6c$v;]��˖��=�v[�2r]T�pTV���snKZr�2����@?�k������Q�+��V��M2�gv�1x�ph,�hȖ7<ډn{j�$tE�X��h�ce8�۲�*3�2����=1{��{���o�`��v���"Ӱ�b�9��a�r�L�l����y9�nӯ*:��v�)uf�߽�{ݷ��}�ǒ�����)JP���i�
'����JR�����JR����_��7��L�n�5D �_mn�� �@�7���R������)=�{��*>�9��i��je�M9��f���/}�w�)�@S�LR}���Ȅ}^��B�
>76\���9����mE�"���!BY��y)J~��┥��v<��=�n[N�ʚ�t2��w�!,�֣��ʈϿoﳊR�=��<�B37]� �AWӚ���2�n;;�6�S�jL�]��y�d�Kn �۫-�M�m9j�`�e�2ڋ"D/��f�)J{��y)J_��w�)JO{�j,�A�wjm��М��#��7�J{��y��| GJ���pS<Qآz���.���R���߶<��?{��8��$�bB�w���2H�KSU4ڋ��/{��┥'��v<��R2S��ﳊR�=��<��<��wc�hq5R�u-��A�J�����y)J{�}�qJR����JR��w]� �A�ֹ%˥S.��GME�R����qJR����JR��{��JR����JR���;������G�x`�+Lmv�tf0d�3���L]�w799�f�}����q��qu>�����픡��}��)~����)=�{��)����){���7�Z�nֳ{��[��R��{��R������R���wۊR�>����O��(��w[�ӤI5T�e7M�B����c�JS���n)Ob���0J�}�[7���%"���	viB��C[�`Q��Յ����7��zWZ֖p��q5�LS<��E��7���K��5� � Jbq�@�6"��� �U@�Q����p�]uA^�����
��6*��s����D#��w�!nf�m�ԔӚ�o�*�π��� �T�;-L?�ٙ��o��������"����ӆ�u�4��vn��ץ��D(P��V��.Q7�Гt�K��D�k�ėf�'��\u�T�9:��{J��Li��
U��o��;7vՁ�kӗ�B�K���;'�y���j���[vn��ץ�u�h�l�>\[ (����M��ץ�f�:"D)�7���֬�S�������\US,=	(S;���3{����j×脣S���X�OO)s%H�U-�t݀}����$�"{��|��� ��v�NN�")5����î���B�$aO��ˋ�b�6�:��ne�M)��Ȥ��BnF��?@��~��,��[S췌�u��Y�-���uv��ϋ�DD%!�����z[w4�ֶL�L�Y2"4�ژe�g��3v��x�������x�RH:�5SM�yBJ"'�{�����s@�e4��@�^,��Ojb�Ը��׌�{�����`]���& a#|������lz�<]m�t���p�<G0��Us���:$9�li䳩3�=Y�h5$�Z��)HZ��2�2[&��.�W�n��s��W�?'`�u;��J�n;qq�E�=W	�G��vL6\ZK&Z���ö�ڷ	�p�� ���Km؜�h�StfH�n7[1[��c,�t��v���Խ�����u�`�<�؆h��� ����u=��w��k���n�u�N�cWa��ݔ�Y�t����v:';��v �\�r"#G#����M �l�6wv��D(��!��j�;��&���TЧ��h[f�U��m��-v� ����$4H7D�M�k�:�ڳ�(�	L�Wt��s�1f=�ӥ2����ESua�;�ߕ��]�`�f�U���܉<C�MO�w=�����J!$��w?�t�uX����\� �&H)�Ĥ���f.�wDe��m��dc���k&M�JU�^��@��C ����m�[^0-���us��F0��NM�k�3��W�=Q�P5�[�����o�m���fO�x�S#�G�u�s@�ץ��d��vOwU��p��#):%Ӧ�*��脗�(�U�{�� �{�@�����h����!�1O����o��mT`��g/�H��fܼ�z���x�nΊ-���K�ɶ`�cm�^���q��{�q#ج��I%��{�`K+��S������.[?) �Hr6��r=�]���B�;��`�����ڿDDD�۽uM�Ғ�uSN��Wk���� ��v|��=��J���u�l���F�mŠz��k�:���-v���\b�SLM�&�U���d(�����]�`������S��Jt3����;������LOn]����7Nua��j��kW^n�(�,S��~�߻@�ڴ��@���W؈<��M�4U5`n��ߢL��s�:{����h����!�1Oqh[f�U��m��-v� ����5A4ӧNF�D%IUww��w���;��9]�h�H
k5��|���I�x�Y$RM �l�=�ՠm���h���H`�$m��I�z�t�.�gQg�����.�uU ;����#��$�9�����ɳ�����- ���$�0	mL	�u��u~Z�Y��Ŭ[S �T�%�0>��X.��#`�1���rhwY�����?���W�6�����wi�45M51��4��@��V�u�hwY�z��b��RB)�@��V��%������`���q	%���d��Q	(��O���{6�U0:��&՛l��p��/4�[+M�,P�<�B�k�A#I��fI�vyf�۶�!�wn?�ͻm�w��v�V�E�;G)���ͱQ�chN�[���m���Qn�v0��1�I`�Ӷ3M�<�l��݃z�m�� ܷ#�K��f]�"�<��3�[�A����(u%��R!Ԗ�M�;FL��ϭ��,hJn�3O-`g��G����֥�������i��.��E�<oi:�	�]��*K"�s������)�M9���; ��v���	/�uwM�|wT�UI4өl��IS�?f�_{Ɂ�s��-��2DY!0i��I�@:�4k�h[f�}�f�~�H'�s���95|o=�`ژd��Kj`^˻&E�D
4���� ��� �l�=�j�=�P]qD�0s"$n:�,�2��>��Q@F���1O�	�����L��!OLM�&�}�f�u�h�h[f��Y��0���"rh���}��g�߾ą9n��j`����v!�
H�cs4z�h[f�}�f�������$#�&9��h�į�ߦ�u�������v� ����i�B9��4��4��h�h[f�������\��Mv�T����O]��̼t���&�f]M.-���vj�zr��uq��S�����������{]�@:�.z������&�����zV��wM ���@�n��n�E�D
4�����U��|�䢔����A�,��|����\do�����rXfk�3wmX��f���L�w;��9�Ӓ�Jj��7vՁ�;��o���`����y�jĖ�b��J]:'g�q{44�����#�5�q���ᚍI#r!�9�1����Z,��vJ���w��K.g7Nq~���,��vJ�����@=-j�6��F�7$����%����u�K*`L��K7Q�sLKq&��`vr�`ʘ{�~����*�� ���߾�*���攘<C���rM=���h^�@;��^��>\u j,I�$i���2|�jE��8�.�I�ͳ��@P���	��D�(�$ ��N- ��hu�@�Қ�ڴ�uq�<I(�&&ԓ@$�0%���[�YS��d�7�d��hzS@��V�u�4�٠uvLph�Lm�C@���%�0	-L	b�l��Y��7<IŠz� �hzS�~���^
�W���"	I����DԒ�K�A2m,N�� �F �JR`���d� LhH�������&����zWa�D	M�B��!��0�J�DKJ~�������;���G�����c��B������5���&y5�S	�dv��WTg0O$�+B�O5�^�g8����+���@�J����A�r�`]�խ����ӱ;���������4�5�Ys]+=��2O+6S���v���QEKx,-��ޮ��T۰�nM���6�v��LH�۶E�L�q9:*��i�۴i��Y-\"D���/����^]&鲌��9Z�Jtt��U�v��y�Z�Un5�3R].Y[ew8����jj��e&ƶ�y0�J霌��m��đ.<�v�ɰ�09v�S�;h�{O�V���7�v�S7n��;�ﯠ��n��8�`�1�4���C�&��m�UI���[�gC.ӭ8�:�[vl�n;h�͎;f����u��mq�͝���-��ܮ'���Uv�T�y�#Lܧ[nV1�C9nț�A[[F3��ix�s�ʽ�H\���QV�*ӎ�K�e�s��P�$��z^&%XغS%z�����3J�nڧh8��Ma8*���.	y��^�U���]lcc��W��P�T�c8VM���إ�ɚ�=n���ˮ��b�!�v\D�ͺں���m�sRќ2cuMD�̭<i՝��|?|n��W^65�/B^W;I�ll�h�VA.�%��ţ��xqu��r�/�^JC�R4 v��6f�#F� �.IU���G,nۑp(.5}}����}����Ŵ \Ժ��V�Vx��Ms�f�n3X�]��z��D�S:��
�ch�+�B:�5����9���i�볻Eh�lHk��z�wd�Ggw^-��ю�t۷C���+� ����P;m�����V�wT��b,T ݝ�t�!�
�am�J��N����b�a::	S����6vش�a�n.��]���6�\�� +��&2�;�ޤ�[8*�U�l�nݵI�vy��NK=�Ѷ{
���m��/.���O�<�+�.4�9�<mr�a`⣁^,�hN.���m��,�%��*]����{�ɤ_DOA.(	��QS��Ҁ~UC��ߛ��v6M�'�3�v��1��k����rn&�n���	�]y����{)�g���~�ݶ�\a�M�=��s��x�����a[�^ˀ�ۛQ�X6#$��"@n�v�txi<�c],�"nX[s��뵮��������J���m<��5��k�\vyܾ�g�f�cd*Xi
���Nt��4��v`�v�gN�11��独}߭���+�a�1���j:�ɖ���cg��xJ��9K4��/Z��፲c"s�z���@�Қ�ڴ��h�вd��"�Y&D�`v�G���Oyx`{ɀIj~�ɓ�z�[E)�tS~�N���?�n�<�d��vuoM���7I�М�b��h}l��f���M��y��~�Ɓ�;�<�,I(�&&�@;�L��=_������'mL���-�z57,E&n+����p��F���L!����7B^Tuu�댼�Z����*0;j� ��0	-LM�,�ދv�kZ��ܫ�{��TO�IU��Q�(��<���;��`f�l�9�rds#Ʊ7<Q�@:���l�:�������kW1�O��^P�%U��;��Ł����3�נvwBɒbP���L�ɠ}zS@���'mLKS�.��Y����;;��4U��JlQ�&���;s�l����S�m���JjF���6��w>E�gۮ�37_���3��`n�M�l��Sb����w�� �h^��>�\4~}S��J3	���Я}�wʿw����z� 1�eEԦ
&0�9���\���|���ӊi��)i���:"(��,	�{٬v��$�0	'*A�b�mUQM��[�l�DD�w?���h^���Q]��X7���p�b��Ŵd:uv2N��ػN�un��ӭv�W���wp��rc�#�,nx��� �����f���M��Š���o'�I�S��3uߒQ2gk��ή�6�n���U&G�A�%�dNM�Қ�[�l�(P�M��`����ͺ��JiKNi��tݟ��N�����s��u�R�]r�Ȉ�u}Ł��7I��ɖ��u4��}���
��?�gl�hu����ƀ����#�8���1�vh���4�]zɻ��pA��:cv�a�E�Q��bn94�h^����Š��@�^,��<M�$RM�W�ʮv��;-O߿f�Yy�0d��Li���:�����٠u�@����*�Ɏd����n`�;-L��������n���U'�T��v�n��;���mw)���`BJ!~E%�b�k�[l>�ܢj�knh�)�ڤK�iֶ�=��>{|U�b�''iƎ�:�ƮUfQ�.��֩�̶�<�r$�n,Ղ�nI��9��D���1��XZm�6훩�"�9z^��v�ywlkcu��s���պQ�7p�M�'c+�N�q;ȦPյ��n@�A�a�����!�Ź�Mv�����Ӣꇶ��n*�w��덓_t��]�����v{X^q!8S�gU�lc�lz��Mv��]R�c�$����o��V�[�l3j`����԰Y��Y��W�y�����n���`�Ɂ�k����Sb�9�@;���l�>��hWn-��L�!$��bmF�3u������T��IL�w;��9��qT��)�`f�ڰ>�n- ��hu�@<ꎱcs�;��a��6�B�]'f��6����=���n5r�m8�`ɑ�"����}]��YS ����W�	�.^%�X�3I�q3MM�f滨��D fn�7ws@��qh���O��cƤ������Vr���ή�6���Yҩ2c�Q$Ȝ�^���ۉ�K*`Z���R�f�5f�-_�M��	�{٬�*`Z��Q�ݗ.�,M�E�4��
a0�0DBG�ȵ�C����&G[k�����e�˭�B�\�,���0	-L	ة�������-e��bIO�ڒhu�@��� �ʘm�X�q�9�j��݁��j��u�,�QITBP�FTd��{��|����|���;2dx)i��h[.�hu�@�빠v.�\��#f&狜X0���Ij`I+�mW�߿���3�@��e�'5��k0�v�C4�l�;�vV��v�un�;]�:��z��椘����\�T����S&<��0Y&4��:���>�\4�Y�������LO#sW��o>{��0	eLKSY^h�u��l�1�ҍ���w�� ��vۛj�$��ID(�v����ƁO	�����f�{�����X���%�\���iUT�5-6��M8�E;�n�"#���wNڌ7n-�z\`͗h31��C���QM��v�Z�>��S`���l���#L�)16����sX��%��l�e���!17���@-�4�٠[�s@��qh�WY&1��'1�ԓ ����W��[��-�0'tu��Fۉ"Liɠ[�s@��T��k���`|�����B�ؿս�|ʊ�;+��n��u�n���B\<hex�;�e�m�)�cgFm�p8r�3uڭۭ�b(��ۆ*R3ƭ��X 6�ZN�k���yX^;<�-l��0�=���2ᛞ5�ʚ�fV��g��z��cZ����m�P�D9���*nG��mt��w3��2�뛤Gl�m�Ūؔ�!��6-�76��4�z��tZU�%�8T��_����~���??��[c=t�����m�ؑ�we:���s[�zy�P�&��}"�59���iI廻�����Zl��Ij`[+����$.8�Q�1h�f�w[4z�hWn-��VA�h�RM �h����sX����l*����_��UE6�?�Q;�ߕ��]�lӻ�a�;���;6��PөD�2f�,`v����m� ����׌3߿��8��Y��\Q"f��>�]�aNz{���gf��u�ɱ:���kO8]_��,߀-�@쉁$X��rL�z���&D�87�w[5fy�|ff6t�s@��qh+k�;�:�ɏ#MƑ&4��;���>��Z����٠w֚��by�i�k������X�o��d�K��!�Di�Z��z�l�>��hWn-�T:��6`�E��l�p��P���㖳pPm�On$�=c"$틵;V� �4
xLRG�w[4��Z�ۋ@=�f��Y�Ǔ	�y1��4�K��[��>��%���7C���	u(m�$�Ձ�]�l��v~;��D��z��p0c �Y�q`1,pf#f
&�8?����5	,4pe��ͫ�� $fBR��B �� ��4���!�E �B��HH���`��� ��̤��DID1��:�b�	�0!߅����O6 耦ث�3�qt�A�0%�#Is�|w��s~�z��0#L5��^��e���?�)�e����JC�ߖ�2۳��"3�"�n���""� h�D@L�l?.�c�`1�tsA9+�M��EV C���0(/�GP? ��� �nƵ矷�=�w4]r�1���jxۘ�?ؗ���w��f�ID�>�6���6Rp暤꛰��`yFow����~Šu�@�]����di��+f�od8�#���˕��7)q��9;`�Ց�OȪƤ��#&4��>�w4���}��������l)�M0����|�=���j`Z������BUGwzn�c��JsR:�jl���0	-Lʨ��幬��^$LOL	��ɠ���ޙ�G���'����Pތ�}�����5��U&��m�n�,D(�}� n�; ��v���:jT�Rbn�ڸY7,��˲����\��a�n�͸M�hs�%�k6�])?���X��%���Ue���SN�U.*�����~�����`w���}]���Ud����)1�I�Ij`v�Fo-�`Z�tu��r&I�94����ۓ`��Ò����vgu̶�L'��&��'��f�	-LKS���*�%����a`������3z�[��Ek2ҝZ��Z�r���]�isu5�TQ�ظV���\�k1��n�N�n2��s�/W\�9x�v�ӵ�-u��ㇳ)c��F���8m��ˌ<&f9�:B�ѕ��'n�#-!��8����ݸ�t�N�6�N�.z{A�[0��lg#�ڍ�7��Σ�cj�IgQ!��v0e����ms��xx9�ػtjt����-����n�g��\�n�=v�Ы�m�a�}���Խ�j �Wc*�D����7�����Ij`v����sXw��lsRI-ES��3u��BS&wu�:���f�?N�8���5TRI��+�o-�g��t��L�y0�@D��A19��ۋ@;�� ��v��;�� �ҹ�M:T,mOs�w[4�٠}l���v��-�.�	���O�9�sɇ�ݭh��p�Ύ���GN^#�$��ܼ��ۆ�ȤǊ94�٠}l���v���f����C�8࢓"rhWns�P=4�&�P�]�^xg*�߾� ;����J@x<�����9��;���X��%����u�$���X�B!��s�w�� �hW�hWn-���
`�0&�&�ff���z�Wr� Ϸ]���~~0Б��"(C.�c����U���c���묢�a=cB^Tuu�ח�\���K��-�`��$��I*P ƞH(I��v��z٠����+6o��S!�i\Ӧ�*%UK��jl��v���������f���h���[ՒIRc�\I�I*`v�]`}ynk �Z��q�<��Y�@��U��$�	,��y g{��33]��;i�F���%[���5f�5p�N�g�9�K�^������v^�.�4���p����������j`J���XJ>g)��h����{�� ��4��Z�ˆ�y�̿��	)�0r94��������p`KS�'�&��ccrhs�k��{���M"!���)RL��v������i9&�����T��	yVw�� ��;�ٰ=+�I��n��e�Xb�x�c�Ӷ���2�7!�{OcF�ƙm�u��Q�5�t�R�������fk�>�͞��w>E�woP�&��BLy�@;���}V��v��zٿؑm��$�<qdRM�ޛ���=
!D���; ��v}�iH�M��d�^�����- ������=
!Nkޛwx�TԸm�\��j`J���XZ�ٞg��if&�֣I``؄�g<[b냒�8�s�ҽ�c��\�rMZ@�V.Ųn@`��u�����=�ln+����k�'�8'c����(�s�nG�(�s]�-�X�2k��kn:�ח���V��&����eP����E�"�5�u��\�l�r̻m��b��=jͻ,=gwe��ny	�t��K>;a��.RP�5�1Űc�73����{��y����]����vL]:Yy���ⶲ�T�&��&��<�os5��1q��q.�}o�����U��3���y0>�ӚqI����QT݁�c������[4����$��@d�ƞM��>�|� Ϸ]���2n�;�;�h��fG2<b���0����$�0;y.�>�\��H1(�!&<Qɠ�f��}V��v���٠r:�f&��܄q�k�i�܂�;�
c�O[=nm�Í���{r̵���(�)'�w�-�e�@;�g�(P�H����I��0~�ws�����Ie(R	(�$�T������4����׎b�86�ә��j`J��f켾�}�{5���V���<S�ɠ�f��t���v��z٠z�d���x�1��&d�^[��>��$��g��o��j���X冐��z]l�����к5����X�&�%)Jj�չ���8���幬�j`J���`����S��Š��@;��d�^[��-��A�-�!,�꛰��`}�����*Q�%���ش�_�@���r	�$i�E�I4����v�ڒK�,Z��y�cn��{�I[�jR��i������$�ߧ�ؽ�$�YbԒK���Ԓ:�ɩ$���;����c��	nr�l]��f�,�Wk�%v�`��.�WM�4dd��y���2�i�_|�J���ԒK���Ԓ:�ɩ$��n��_>����br9���fk���(IUT��i�����|�ߦfg6X�$���fOL'�Ɔ��Ԓ:�MI%�p����<���-I$������v����l��M�D�;��P�_ɼ���?~����󛙙����Lˈ��jD	B��J���w333��kN�uB�T��9�����,Z�Iwu���G;TԒ^�n/}I$��Cu��7#@�g'-���I;`(���M�rݶ�&[�z��rv�&uI#Fd�܋RI.��RH�)5L��ݽG�D$���f{��nff{���M��s#�,nI�$u�����K�߷���J���ԒK���Ԓ�R�#NL'�[�ORI}�����RIu�-I$���}I#��Ԓ]�U��1O	j6����f7o�$������GYI�!{n�=�$�]u�	D"3��p��Ivf��32��$�+{�陙��Ws33�<s����Q_�(����
"���
"��(���Т*+�"����B���� ��
"������Q_�Q_�EEo�QXQ�EE�Q��DTW�Q_�EE�Q�B����DTW���e5�����G3� �s2}p��  � @
           
     =*	H�(E*���P	(	U 
�RJ%(��A@  (�� P@*�J��$(����  h   
P� =>����A�2wa��@{�W'�W��n���ܾ��/)w} 4�ҬYJ͎ �^Cק'J� �)����wW�O�b�]�z�)f�_\�ڕf�{o��>��  �T   �R� 2 �)d�����*�l�bë� (�2j����ɧ[�]���+�s�b�x �ͩVl)� �=)�{2���/]�ݵ��u�� ���+w��z\Yɸ������  =�@   
(	P@ }ﭵw�ו�{Ƚ�nz���/p>�w�}���������Ϸ{����]�o �����ؾ�μ ��y:w���z� �1��]��Ү��/[��+}� s���w}�<��NO�kri�� }�    ���t{��m��[nMuN�={}}���U�뼥b�t��u�6W��  ֛  ��>��� P@�� @ @ v`
@ D��D �P    0
 �    �@� �n   " :E � � @1  � �  (� �m �   +�>�e��ru� U�)Y��[��Zrʾ��+� ��y���]�rx��nm+�-:o j��R�  *�)��*� "x�T���  "{J���R   ��#%)H  ��(a4<R�k�o�������O����s;���W��I��i^���PTTWAPT�`TTW�`TTW��QQX �����?��K�U��i� "E���j�%�Vrj�ĩTaH�aX�YIU�$�R�E�"�� �!CB��!	M�pIP0y��!+,�)�n$��R!��]��d�:K�@.��"0�R,Q���D#��8���q��e�$����+�@�i�^��*�@!3"ә�]4��a�熞\a���S�B8&Ń ��Ɛ�%�$)�HP����tq�d�p��� _���y(��?,	�OhHЅ�q�y>�L�!�B-O'��9���!g�!
B�!	)6C�)
�=��ŅF��x@�`�<9�F�ww8tQ�E��s�hb��(V�����W��B�|�6��L�fI.HR�
�C�B�]��w�9�80
)�
�Db���<`�70�BȐ�
Jfg�7��8���Ysh��9��Zf�ܐ�0�13w�	!V,'�5�nC<a�?>a,���R��(@"F��(��XN,)�����
���� T�$��l���ư�b���a ��܄ӗM�%"Q�#R#H�FH�k
���)����$V&�B�:��:�n�B]���� 0Z�����I!H�X�1ЉL�,"@�O4cB���x8 zpX0��
��wL�o�@�<2JD�q�MHW5��V*4q�B6H�����}B쨔�v%Wn�.��j!�V��D(�*ze4ۡ.P�L���7��d�0�7�OԐ#RbK�@����4���=�BS�X) RZK!���}�LW�Y/�l����F6���><�4�����ˁ��畖�3~g�t�\�.�/=�L>�����+�bK��.i�'�ĸhE��=�ː��V�R�^q1t.��z����K�3�	��u�Q��B T�`1R�x8J�1��_���I|�r��%!q!GіS!L#L4Þ7�����h�
���2�%Cp��b\�e�Є	Ya3�6[����-|��_$0���@��O�!V#F"P
�������С����$Z.�
x���N>���
���t�š����@(a�������<!$���䰷��a��,�_K�_7�.���GG��6�ˆq�\G���d癧���В
jr���x���7p=H��Э�9���$��c�V\2칒�W֜�^��i��`WN>B�3rBdaYw�y�Ƙ�.,	�XV��\6�B�&���7�.�0#��\V#�<�7�8c.9'��t�Zz{�S��p�xF�<@�\,�	LI�F,�x�5<����c�K�yS��dXLOD�`41��CE�t��!~�������/<e15㇇�1�st�x&X�!GW��+0 �`N#�`F!�9��l8f7a<��p9�
�O;�9����.'8��%߼a1J+��B������!\5!e&�.o��.^xK�yIi�hB��.�
$�ak���{r�٬,���t�M��v\1�!LT�$B��!\!5H��"�%��o�#�pxRS=!LP��3�<���=B5�w�82,Jf��\ E%�\�xx�a#����p�����d�S$�4�x��O&e��S4��S�ׁ�o
Y�2��w�l��B�ZF��s�f��>8�_�w�/���D���������}�9�ɤ�o��9���u���)�*JV3W��Lu#9}%/����]<|��书�p�!2!=q"@ 0"S)���`��
�K��.m�3����.s��B��3�=���{$���x���hi�<%0Ӟy��379�{3�3�ہ0��<��}���Lf�Hl�ϟ�>i,�s�xd��9�%9�<4�˓y�s�%�S�)c�B�p|ׇ����a����F��uF8�hj�)��8�(B��!re	�s�$��uB@�\0�
�fi�P�ԍ�5��	H�6�`p6�G70�!LԒT�w��Cw��
h�A�Q�`%\S�1�̛"R�Dэ$:�&���!P�"E �D���B)BH��S�a�L-��r��Y�z'F!\q5m!��nI
�o�G����	�ɑ��Ji��"�Hk�(p(UX��҅^ �F�u�����7,� �@)�t2R[�t7А"Bil"hJ����4&�B�8����$��0���d���e�J6�,�m7y��ӜVRF��
ēNhFD�sI%�I[d�f�e0,�7'%���
�6m�@�x����0)�K�7��� ����FBaU�(@��,J�HA�da�B���8� z� �|�$
���I"�Q�A@���� ��ԁca0Ra%���	#G  U�C@�p�q�)���X�-B0q׆�hb���S��HD���LP�U1��	%��$I"�lK�YaD)1�4�l�+���4�����9q���%��6>a�+��x�c
Ԙ��<��I(��������x{�$r��٣g<<}!XQ�q!B!�i���-!�t�2�+� 0b-`_0�B��IsSP��NB�DZa�8Cp�CS�#W�p�\�`H�#����ϟ�)29��)�]�y�{�H�z������:�q*�x�J�i�S���^xa�9*i�e�Fo���,��s����y�9�2���V4�Ӈ��z�Y�y����vs�`dB ����!�IoiH�$*F��)��L3<���X{2CIy4�a��{�1���F��l����8�Z�zt'�>�S)K��|z�ZƲ6�0z�BE�`@H�"D*qaC��K�X"� ��H3��I
��Y�(ˬ04�)$�(y����,�@$���|q���p��8p�x�w&q#��ɰÉ,�/��[��P�!V,ZӋ
@��D"$F����)��@� �Jfi�
�	��A� �t�<#H�C �s"HH���5$p�#6i,A���Md�4�	�e8L�'���b���"�����\��|Y �$$D�c�B�;[��Bc�`}��0eY	%C �,��G2\�B!�*B��I��,��>J�j@�JLC$fͰ�d�t�zu>�%
R< �x��(@�
f��p����Y)m�絀�{a���d���w���Z��M9V�@��p]P.8���t���Gee��4L9����
H�p�+پ{�LaR��W7�4�sُ���
k���͓��@��@��[)SS6AH]���顔���65_ �==�P�	%�No�e�7��Jf<9�#V��ye��Le��Я�$=J��X��ԈF��Rı�F�$���M�B@�$+	
A��V�$)���0i��J�'�$	�[0�I��Bd��иg����I�x���j��!D�O�8xA�����"��ȗ���,g<<#�Ŗx��D��	7��cr�i4�ټ!�>:��`M��� @�F
�HT���!��u�+HWP�"%\Q���
Ɩ�l�.V$
K�w�i���&
��+b��F�5���!U� �@��V�T�B�&��z�����������  u�H     �   h.�JYj�j��5�	 6%f�m�m&ֱΐh���m��\ m�ņ�c��o��:5� l�Um�T��  �f�:t�lܩ$�r��ll T�Vӣ]w����U�[<��f�Ә�9;b
���F�W+������X鐭�ت��UWvV=���u�g`��j���"�)r��ԇl�;6�v��^,�E���m�v�,��i�l��x6�m�l��[[z�к�  �K֑v�۶l�&� � 	:���� ��[R1�Z:R�e����.��V����v�����mլ�.	-���	 �K�M����EUs*R [UUUu@Q�*�R��L�z�6�;`MRIն�Knm�3���SԒ���m�N��t�I���r�{)����˻ iWMS׬�f� [BK%��!�UU�Yz��	�C����r��*��J���Ur�^��h
��*�d�] +倪��V�3`��]�7ee��<5	����E��lh -]vN��Hۉ`ݧ��y%Z;Nٴ���k|���e'��X*�8����n^U�J��m����$�{*�xRl\-��T[-P*6N��������V�� m�$�� e�dI&��K��   im�]�����q���@Ho7e[&˥��[[m ��8 m&�u���6ݎ�		 @Ү�I��d��m�B� e�h]�ܶ���%�;$ݞ�]�Y�Լ�A����k��v�VΌ�:@yڮtT�<p�.���u�+`�ֹ�v:�Ij�i�ħ<++��p�s[����]u�;�����P[]PW&�5���F��0Sui��&�R�	-쮸��J��lB1�x���Qض����8��J�ګ����6��j��)��r�]J���t�.�÷h�➗gf��]�:�R�#�Wf�z�\�-��U\����U�U���Z��5t�U��*��Ƥ��]�73� 6�y�+X�Q�L���U�c�v���`m��6�-�6��l�VQ;�O���;T���<Uu�e\;cY�5U=�UUYS[$J���U���v
�t�� ���N�+����`%�C�@H�hl$9�lH��`m�6�7  n�r�UN٩�cT�U�A�!+�T��kaA���  ;v��M�@�l8�z]��m�m�  v�3�GѢ� [R Ӯ�����I��-�������;�UU�`*�� m����Na���-���^`s���[l	�sV��� �ۖJ6׮lle�P$8۬Y���/]�6�HI�ċj@��벇�ݑ��>�`sE���	 �cm�Um
�!d���H].:D���m�j�`)]��+F�l��@��n�-�� 8�[۫�b�!U�qF�6.�0��M���d�ݴ��}�O�	+sPm��Ix [@ۖ�moP9��$�� m�d�  � ph-� �aƺm&��I�l$j�e�H�  
��VʵT��]U<��%�ynU�j��V]� �	@�-�o-��m�8 	%�p�i7$ �]� H ��H�� ]3l���V�H�t[���@UU2� �6T��� $m��JHv��ATp�Dv��SBú^����vݖͷ;k@[*�[mP%��+`A�kv���D�mv�耰�n۰h�l�۶�xp �fȑnv��oX*k]z�ސ		������O�7E�[@�[�ݶ�gӴ�u�Ͷźݝ �uv@��h���$�ؐ$��@�$I����ؐ� 6��mm�#��l-� p[@ ��mWE�1m$���ݶ m��T�<Ү���PN�� ]*F Ͷ�րm��kj�o�q$��vl8[]��쐶�sl����H���n@Y�J�����E��3E���Qc[�d�kX��M�`Uꪃ����� 浶�t�ES��5��M�јXbʔ�}����B�H᭕/Zʆq�����ܠ-�@[I
���5T�y�c;l�77',�'��XqmA���[ym$m�  nը շRUER�ɺm�i�B�����U7!!�)@� 6�	/i%-�[�mw]6�#Kje:e"�j�h<�X$[�\�Ā� Jă�+d6��'��j�ܶ�m;��ꪪ	s�]�;�R�]�b�mJ�M*�U*�m� 6�\��6�[��
���:j�	nK/i�8���؋���  8 t�[Vղ[h��R�U*�T�V��UA��U*�3%�L�F����*U!{f��Ve]K�]'Kl�	� 6�  ��κ�HrKl�E��[����p��5�\S�/Z�d�ڮ��U]�*��Ul��;�
���6���l�m�6��i $��	-�ϧ}~�o�m�  m��7U�Ӝ�����$8 �l ��:Qem[H m� m��� ��H$��2��[ aM����kW�l[Vз��� pm&� ۷a�@o0v��h$�6ۜ  �lKh�km���`[F�L6ͷ!l����*�u�SjU�� )@  i2=�T��
P ��*� $H㵺�d� ld 	  �h�ͷ` >�d��m��[R$�����6��Ͱ$    � m�U� pIj�ͷa�[v@[\
Sm,[�	 �㍷`  �`	 [@        �m�m�[@ �6�����0  D��rc0 ��I�t��  ,m�Ḱ �u ' �ͫpS!�\]%��M���,6[Dk��m�    �^h�1�T�ܶ�l   � H  �p ��E����H@���{ݶhz�Q�am�� �`�%� ����$� -�  ��F���l -6   {Mr�[�V��*ě�������` �v�� ���N�8ׄ�Wcv�c�۶j�T�l�	�z�6�W`:H�� �t�+�U���U� �]��9�[%[Mj*��n��߾<�.��Ҹn�[H [m�bڃc�@� �ٶ�����jP   ���K��	�:q�*������O�Y%u.A�D�Ӝ۰-��f� ��D78$&��L� ��}a���-��6��!��-��� 4^nʑ �ӎ�e�l�`� �� �`���6�z�k�M�v���&�j�N�S����l7m��� �m�`��,$H iÜ�:H,$��xI&�� "4Vؐm�nZ   6�@	 $�V�P l m m���hm�!�kn�M�Im-�2m�$ �    ���m� �^Z��'\�mUS�F�$ &�x�v�^�� �   �@$GP  � �d�e�@�����  � �� �"�6��M�l8@��8  	�l �X׫��� m���6�m�n�m��K.�� 	�j*PD"ɒU⌣!5mR�mXv�j[S҉:P6�$ 6�.�m�   �� j^�@r�3�m��4IM�8$6ۛl � m   @ �m����	�� � -�n8Ze��lq�Xf�k��ܵA^S����$Mk�����j �km�@s/K�!�d��a`Q�&;v��m     ���[@�d����;mS�	8d�  �� �$` �6�,4�4�b���ͻX��UO<�k�Nۊ��vxԮ�U��m�:� 6�||M�Ż;U������۶F)y^���Ӎ�� 5�knFFnl�\ �͝�sya��«��o�:��?�0 vv�I��e�	/��g;��'!d�&�f�ܝj�쒺ٺ\6�@�V��:� m�tY-������~���u.q��� y�E��m��gH m'l�Ɠljl��U9"����(�[���㡭�苷!5 I,���n�q�ꀋ n�ݶp��,Ҵ�Eaڠg�旈��T��E�/Z��(���$��m�Ѕ�H�o����V�d� 5���mm_kp8$��m]$�@-�^�����|�Dҭ���7/[v�崥� 8  ��f���,�v,]�]-�� -6 �V�e�ɔP��
��IE��+B�L�a�N�Jky���n�&� �;mo\H �m"ڪ�j�+cid9��X$n�t�m톋��k  -�  v�6��Z��f�ʧ.� ��� ����aۅ�-6��m�@���t��vbWA��U*	���t(���т����4�� �B�x���p5KvH
ӮyV�Ԝ�-�ԭ���n�m���6K�rg��PT��dP��$��+�|��S�U�`� �`����>�q?�s�h�&�
 j��04�HP袞�!TJ�&�uS�@� 8z�(� Z�|�zq| �C�*���Kފ@3�)��"�x��	"�"$`�D $���
�AP� R�	���>	G_��O |~AH#�Q�#�A�R���D�p�@ � ?qU�pU PD��A���(�	�:��� D���D�XD�d��b�����1�$���� �@�C�G�GA ���u��h
�C��� ?�z
�x�G�T9�b��*!�O�D蠇��"<R
�z����b�PA�z����j ���(�!��*�CT�UB&(��EP_G�u S���
�>��+��**+���"��T ��9�JR�U;�zɵ�J[��Ǝjά۳=�Ͷ�+�x	7�L��ۨW�-t�9��ݶ�z֎)�Y��YBIu���yŎ�8��lf��f�<�=��v�M��̩Wm��=P&ݪ6��/�m�ۥ:��8��˵�F�Q�����H7:��1ƕ�EP8���g��s��ol�nF�[s��mñ�� ��Ņ]�d������E����t1Z��Ck���;s�[r7n;>zC��{��9j��<�M��an&���65@K�]R^-�{<����(U]<����TQO9�Z��˺9nv�y��e�{p뀭5bؠny�`�j��.������9�4�d�&�N���O�.�W�E)����������z,�;&��b�;)۞$^{��zT��k�`�f��� �������1ͥ	��RM�fSs�R��i�^-�t�v8�]��N��Lһ����t�wC���p�仙-�-��Fk���i�8�m��&4�� (���76�î��"��0X�㙵���M+L�i�0y��ף���Hy������m�y�k�;��u���g\լ��
�Q��]���F7"����e˜%Ę/`��2�2ҝ7k�d sUUT�uq�*�G��[��ƲZ�i�rt<]Tˈ8&����]��%6��u���۞����,�o2v�fD�.|p�tN�E[5�i�gn�競�(�@��5�ι��HY�f�ceE�u��M<OAf�JD������P{%.E��B�;ta'@:�)[��Yą�[k�����crgi4�{N�����̻J�� ���8
������@�i���Z�%j��W�ڮ��sjL���	�ݶ]Xy�]>ɵ-���N �r�[\{�ڸ��.09�nZ�d9!#a�f��x�a�����<,qe��;v�%��gn:l<�ت�]�EY��M��+�n�A�N���� H��5�t᪔i�ٙ���������|��� E���!*D�� ����^| x!�O ����|�fY�ʌ��0�b�X^��5��(7:렀�^z�ҹ.��W�T���^�5'l.8ґUv��˽^����7֫��8Ν��7m��v�v��fly��`X�՜k�;j��z"Ŵ�7RD
�l�g��c��&��6n�l�&b�Y�n�\ؐ�gnA'6���=W�{*e�5IW[X�l(����J;�w���������AC�UL�p� �w<g���.wl�g�<��m7]$��nf� �c�_;�_�_UW���4���:��ƥ�%�z�"u��o}�y*@/3b@=W� n:[�����)�`ܖ;�u`��`�l�f�1v�=���ԔFs�X�6J��T�=-L&~�������fl �BQ��rX;�,������l�;�s����.��aMv�յ���t�z�˪�ӹ9�/fѕ����g%j�v��� ?�����$w&��I.�l�Iw6�i$��5�9#(��&���BK�6++꬟}T1�m(ZP �!���=���}�<����ἶ�|��9Ē�л����IҀ�r+I$����I#��R��mw}��$�͞��IwM�n�R�Bm9>$��I#��R�I.fl�Iw&��I.fl�Ii���Ө�8ԡ�$-$��f�q$��X���I.fl�Iw6�i$�jf�r
�BFIO��{r�N���=���#�WLg��\��{N�����*R`��Iɤ��K��9Ē]͸ZI%�ݜ�Ict��7Τ�JM�ZI%�͜�I.��-$��n�q$���\��ic36���$F҉��$��ۅ��\���)�}UR��$H�0"*T � �"Ec*R"V��͞���i$�36s�$v�=cR**O���ZI%�ݜ�Iɤ��K��9Ē]͸ZI,�M{NH�*8*I���H�M%��]���$��m��I.f��K�}��V���8�(�8�����V���qӗ^l.�v���:y�xջs��cN�3=��ٮ�<Xm8N��[�~��I.��-$��n�q$���ZI.�M�*S�&ӓ�I9Ē]͸ZI%�ݜ�Iɤ��K��9Ē[��6�F��6䅤�\���$�ܚKJ}�|�Y���$��ۅ��ܔ�Y�8T��I9Ē;�Ii$�w6y��~�6r��@�Ah��U�"�U���������0���8�u%
!�p��Igsg8�K��I$����I#�4��Ir�[�D$j:I��n�4rZ�7InXt�̃�V��'vēe�\"�UW։w�S�H����I%��I$����I#�4���6�[���$�����H��訃r�Issg8�Gri-$�����B�mՁ���i�EF�aΜ�L�j`eL�^0Y���`M����IҀ�rX:��,�T��W��T�=eL	Is�ǋBm9>$�����X��{Ӏ��X��Hi		��Vŝ�GzA����b�]nC f�f�r���^�AԈU�rM�W�)�Xt�עv���-8��T��V��N��x��;r�	��حcml�Yhڲt���żvz��7����+l糫��ۆ勥�dGI��0d���:6Lby���lp��9����@�۲�W9�2S����y�ӡ�ɜ�2K7kF�N�i���6;t�S-'&����s3e��W�F�It^�kt�-�Ξf��J�cB�mI*���3;/R� o�|����I*�����`n:[����*R`���͖��,�mՀs7e��t��7Τ��t8�`%L	��`���*`b;��S�H�������X;�,��,W�s���;Y�i�D�.`��0l��zʘ�T��,�_U{~���U*��I�4JE6v��,�u95��u��7%�F:�t�Iy�om]Y�i�G*LrN w��`�l�3�4�w6X�	��r�t@m�,���j��C�x�'��@$�;<X7=,��-��$sL�n��8�}�R�$�H��=���*`�e������F��� �se�{mL�*`n�F��[�t��ù�.��DH�2$M��y�@f\i`�l�5WM�9����>Rt�5�:�8.�u��x{Dz^;c�p�p�vθ��?wË�Au&�07b� �ژ;�,#��l�7)"6�NK���u5�^�HnlHU�H��qu�**O����s3e�sse��}U���M����c&$��$���.�Y�����s�I0m��zJ��R�9����`M�����m�`%L	�Q�zZ����3ټ�*R�4N��L(�\B�'=&#Q$Y%ԉեu�4����/V��{M6ߒ���*`���*`Iy���]:Q!�6�,��/�}U�RA�o��f論�ɥ���=����ϣC�J�p�R`��0��ب�=-L���~Ι�]�Kv̒��$���o��ā����z�"@ibM5lI$�Q�������I��}ݙ�a���s���R`n�F�*`�S ��3o��~��h��:+8��={U��,���ml���nؽ�B��0\U�Q�H`���0IS�q��rFT�1�,�͗꤃���sg� �f���6RnS�N���&�*`{b� ��0l���3F��8�m9>$���ri`�ږ��� �f���F��҉8���P�=��`�S �ʘب�*�"�b�w��=�3JS`��vA�ۣ�5�.Y����Vn�uh�n���x�M�LoW\��ݫ9w)ɭ�3��,zz�e1]��g&�f�Uey��q#J�܄���0Z�Al�nx�+` ���o�Gv=*��]��8"�X�SMÁ�F�ٰI�&2:PSc����]�lu��l��7�>�ҽ:Nu�='k�9��sO�i;�1\�$q*�� QTay��n칻�&ݺh�Fk<�Ag�M���S��PYխˑ�C��ո�dN�7!�t�8(�T��~�����ɥ�swT�;��=��)F8�	$�=%LlT`��0m���w6���Dm*��`w�4�nj�~�#��K �o��r�6�(�)P9�u!�z���=eL�T��,�={NIN�8�Rb�K ��������U��=e�`\�&���a]Y&�r`��5v�\\�ՙ�`C:�W��ri��M�5���D���m�������Q�z���=%LR��q���r|I%��ɥ��}�]RaٺK �we�s3e���WJ$H�*tۃ ��L�*`���*0,�f��>���#n�p���� �f��ɥ�s7I`w],{M����I�zJ�f~�_ǀ7��`�S�_Vx=b�r��F��&��:����h��w��������HN��Wk5e��.w��^e_l�`�S �vX+��l�EIJ��ru�RA����n{���sn��x����pT!��wvXwvY�r��c�!�~�)!(���x=	LH�HI#!����H��B4��$\� j0^վ"J�o�L�#1hJŹ0��.�ˁ
`@1i+��.(H1$d���H��Ɏ\)-�:�H�(E�JR�	IHJ��	a�`�#VB��,i(R���� :�QM��JJȑ�$�YIed4�V��"ET_@�b*���b����J � '��V	ED:
�('�<D ��D^�����W�O�
��6'ɵ������:jR�ےÕU�Y���37�^����<�,��|������7�up�rV�ə��y��[O�+��ؓ�'�y��3=����3)��(��R��Rct�P�a�����s�W/fp�u��9v��t�T����rU�H���K�_.��p3ޖ{�.���Ë�+}��:N�Q�M�`�����9��VV��}I�K�ɨ�J�r	��,'�&����T�=%L�%GzB���l��,fmՁ�ջ,����	ঁ�qTCn���|{�v6IJ$��r����`v�s]�s����rT9]���$㊤��r�.�p\�:��αmh䔬��K���eM<�g�:[���GBNK �we�s����f�X]Y���VT�I�N��i�# �ʘ��`o7���j`JKM��dCi��K��u`uuf� �n� �se���m��� R��6���o%L���=��Ȩ��ܛ��:n*�`���9���9��`]�a W+�� Zx�Bi�(3 �U5�;��=�]���rZ�۳xk]���<
d�� f�����X�c��ɷ]h�Z*�1��YWE����d��=0�.��s�E�T���Q�b���%;p��Uv���*��2`�Y<�s;K���u�3zٙ���Y�u�r�@�Kr+����&#�a�`8�!��9;q����<j���8�h=���X�2�o)Xðn�ws^ˣ�����_�;�mV=r���A�^�ʱ������r#���m��Gn��p�5%D9М����3&�Wsd�n��q�6B����(r&�Q���R`���T�7&=��B*%@Q9���X7vXs6X�4�7���9#(��C]I0[S �*`I͕&�eM����jF!�$��l�32i`uw6K �n�{O]j��)J2:���T:�R����%і�k\�qj^l\�ҷ.-�JGHLn�	�NO�rX�۫���X7v~�7},��m���h�P�؅ W*�"u��!4�k�Y����s6���:ݍH}6&�ȓ ��0��}��3?g9-��r^�X�K^�����q6��fl�$��y���=mLsgnw�3�p���é&��`o6v��j`��`���7S�"�q��6JI�V�{�^nܡ�8����%�R�:v�{�gm�F\�V07�;S ��0ISI�V��=�$e�$��,��,d���W��Q06d�Vs�Y���M�%�ff���K2��ꪪ#��@#$���$U �$�/�uAM��{�Xf�9�h�\M�'�4��Q�z�&�*`J�f����4tT�� ����}��U.��pw},fM,�<��
t���1�V;l��t<S(7'&�#���a�lyb�Wx�*꒷������???o�J���`���������q�H�xu$�$�0=%x�=e �f� ��l!NDTM9%��ͼ`���zJ���3eGz!�$a���c ��L�T�$�0u�|��Ձ���i�E(EI28F�*`J���`�x��3[����61��7�o���F�3ׁ��{cc��9b�4�t��ݜ=�\u�p�=�#rԼ-�0=%x�=��0ISԺ7W�&ӓ��36��9��,��,��,�jn�������헉�zZ�"�d�nƤ>���T܊X36X̚X�۫ �sT�;���ME���9ޤ��%x�=��0KS$�@`�P��[ۆ���Mɺ`���q��]<��qc�Cu�p�{nx�ٹ�wm�ծJ���[D����� 0�l:��N�v#@�3���틔
���>�m���p�`6�&N:�ջs\	L��)ѹʸ�?�}�ˍ*�4��iv��n��Lqݮ&Y��8��&�F�E���=���!Ƶ�8��/t4;U���5�M�x7����H�.4Ga���Y�������v�q11�K�́�[f�<�m0�`鎪�t�içv���u�ܺ�Ѻ�xIf�v��{aS ��0="��efl!��Dܫ �p�`���T`I+���-;ĺ�.g9ӝ`����J�{p�`w+*l��`5E6��3&���`�T�=mL��{�	ww��X�z���`�T�=mLfmՀp2�݅A�8�mG*����F����k)V7g���dlMlhūT�V��;�gz�0l�L������Vq��jC���
jE,���Ί��xtE����#�@�BASTUx��'s���{�u`�j�u�ש��DG��.�HwHw���4��
��$�vXk���B����,�۫ ��L����ٜ���2ߑވB�	qs�X�=% ��06J񁙛u`w>�.&�* 9SI"T�����e��[�������t���4Ma����c�r6Jv�.g9ӽB`���^06J�s3I`w+*l��`:R&��rW���o�������Zw�p�ЛNJ��Vs6��9���~���l�6X�۫{�������w�c ��L����+��^03n��>��(�*q�X3vX�^06J�zJ&�K�K;����n�Y�G]�+�+n{k����gd g���%&�j/���t�&�;��VrW��Q0KS ��۝��\1s�����W��Q0KSd��+3`�	DD�
&�X34��j`l��d�s����q#9Ν� ��06J�W�~��B D 6��� �����%������q��H�rX�۫d���`���7&w;z�;�&e�I�[3�ݜ�Ў�RC�J���ôB���n����87R:i�#�����zJ&�j���������BL�rU�s3I~�� ������]X�۫1��jC���$(�$י]�5$�|��l� ��"@�:Ktj/�������s6���J�zJ&�j`�;s��K�.w���06J�zJ&�j`l��I4��b�F%p � _Ie5!�D�q�Lv�bŋ��3qM���Xi�����w4�ٻ��v�HD�r\�i�L�`�^���03B	���H%"E=Q��d�4���J���i��B,� @��/J0aD���<M�4 p!�	���� K����i���
�D�H0�Ia����5T�q�*��!%��"��8���B�`c��1&cG�.Ha��R���"���VBZ�f1����ЗT4�jD+$h`B���1�	H*Ѝ0H�H1H�(��@�P
(Č�� �#�B����*9�a��M-���.,�Fmf�H$�! �i��@�0��V$)��E�D�Px*�~��$�����B D$N��T�HB�6� G���ԁ �B-`5�,��wp�������ޞ�׷3�6X
�i<ܷ��L���n���� ��q�,Hp^�\��7hqbn�:ax�9�Ch�u�/8�k.5�ۯg#cV�m��=)���U�vy7�VNwb�qf�Ӻ�����c���<�6x[�]�v��MsJa����iscs��2��F�f�v��c�m�y�M`��m�B2M&�ޔ֯dtt�=!��mn�;X�ݍ7<�`��'����9�u���GY�XѺ�ļ��-�giG�Dʋ���TM���dwn�U�f�9Iͮy��*��ʪ�g<�e8�Bn{M��
� ���I4.-���܇U��::�����I�btL"h'8���� ��"FxJn�U<������W\F��ZVn2��x��^Uj�(��.έ`	\rk�\�@�l��� �D���29�w`�'l��1�s.6�݋��v��rz�p*���8�;j"^X�m�1�Y,Ls��]q��t󦻰�;�vq��;�����
��m�Pm�����%��u��8+�Ҵ�V���c='
l���d)�Ss�,�N�:�=J�F�u<^v�Vۭ���n��Ū:z�&{a�W*�F/l�� ]D�]/eBKn�0 h��:��y-HH!�6�sk�i� �)�m�U�@ ��Sݛpm{��]h�M:ayE��#WR��.�g�5��N>��g�m��ad鳲�(����g�clvԃ�0��t��pT�2���Y�nHmr�; X�^�!�T�n����J�M�[9��6݊ݴ�êBYT֛�jv{5U;��ݾ3���i����՚%ڢh�6�"�s�kٍ�6r�pl�TK�ъ�k��̨�(#:h�B�t{*7��w�,q�w\e�j�[u����M綷BM�����,��S��rN��C��CD{pc��u�Ճ�iDp8�6����/nݲ��U�s�Il���]���\�R'������I
��m�����ρ� 8𮢃� �#��)���엖˚fn̳$��k'YR�Y��Wnj�mlm�8��`�Ohv�L��b9�q����O]Je���N�lpہ굧Ge5�	�����ZM��A�c�n�&��L�ݺC��8̝U�`����9��l�sr����:�Jｆ�*��L�m�����o�@���$j�����g���s�m�@W0�M���t�IQ�'���³����|	c��]6u�5�4��^��5r&����簗��t�WYw5eֻF��ެ�K�&�j`zEF�^07���Ԍ�*I�Ԗ�ݗ�����j�`[~x�=&T�ٓY��t���s�I0="�I^0I�0n��&HH�M�$�J�32�`�*`���T`z����s��ޥ��eL����fmՁ�]ݢ8�7 ���QF�q���חF��i�\�C��,��[��'2�������$�n�9��VfmՀs�l�;����� �t�$�<���樗H	�HH�� DUS|i������T�z�ȐfdN��v�_����&�I*���]X;
�����+��%Gz!`�,A���c �¦�j`zJ�ٙ��R��r�e??&�`D�LL��=mLI^0$�� �¦��#��m�ul��`��]�t�)��y1zzY֬)�v�VWEe\mG�e�س;����	��T�z����m{�V�Āg����	�䑸X��V�� �Ȑ=wN��K�+w{ީ�#��#�]�B�
�6$ٙZ��IyH�M,fmՁ��u�!Q��85B�"C[Ms��� Vdi ]�J���U�p뤷F��ȔN����:��n�x�=���zژ����.s���,�=r��Q�@,�6+I��ȍD�ד����8��9lp�33n��
�����������\�V0l*`���T`I6����׬��S�*I��,��,I^0$�� �¦̘����:�����$����I^0l*a? ����*�ݛ,��Rc�#�6��u,`I�0[S�W������ڹ��V�[�EP̶�W��%�T��jq��ջqӇ�-��^�N����P�=���zژ��`I+�c��ԇѶ�85B���ݗ着���������]X3+e��t�m5�D�ct����f�X��V���`��`���8�r"&���?�ww�@+1lH�2$5����) ���68�@�Dܫ �f���U�W������@f�Ҥ��R%(i5�t�� ��~n~�3H雙4�vf�fۼ��h4��-��l`��s����1�Ξy�]Ha�!9M�7 D�t�^%����<fcM@D �Sv�gF.t����|�l��6�������3�!��lzf�4�+]��m]������컮��!n��]�.1�v�
�@�u)�wOnw��']�zҡ=��QǑ��jC���K�-��ۻ��@wu�l��s1ڴf[���b���X�αh��nq7�
g&�f{o�ݮ��ᛝ�H�$�p� ������f�X��_������`f������J2�RK�W��ٜ�m�� �~ ��0[ʓ�	�H䒬�۫ �f��9����f�X���\$e ��C ��L����+��Q�'ku�!Q�%NQ%�swe��ͺ�33n���K���e7��9 n�c"�n2��6�;	i�-��m��������e%%%5�D�ct����f�X��V��%�swe�v��X���Tm�q%�	%x�����3��D�6ʘ�۫��_U$[��mB�	PMʰ��0[Sd�J�w;{��E(EBi2K �����u`]�J�֒Is�xlH�l#�P�ut�w�&��J�{aS ���m��߳��4�N�Ԝ]T:�YI�:x:� KLqR��\�ҳ�h��YH�Ongz�z�X��W��
�����u`sw[up��dTSrU�s�j`����ex���/{ԄtbL��$�nl�9��V}YI.��X;����,�h�9Q��'%��+���`�T���7�Lrk�:p���$�36��9�6X7vX�۫ �v�БP�Ѹڑ�)N��Q=�c/%�-��s��L�b]T6�)@�Dܫ �p�`��`s3n��۫{O^�e�J�i2&�j`zJ�$��06d����(�e6��36���ͺ�fV� ��� ��Ԙ�H�Lq�������) �ű �Ȑ���I�گ��-�p�;����H�2*)�1�zL��zژ�Q�$�~�������N��L�1�7��%���sl�!�x�����	D�9Mby��g8;�q/ o�|���`I�ʬ뤳i��$n�rX̚XJ�zL��zژ�goN���u����v	��	 ��ȓZI7���`wvx��f�� �8���zL��zژ�Q�$T`]���u8�)T�	��K �����u`fd��9�[,UU�_�}���Q��H��)3t��E�F�ЧK�V��Q't�Y��i��hM�5���Ʇ�;��T[Y��<X���#go��ѹ��n�Q�DoA��ח���t�˳\n�UЋ�m�m��ƶ��;tq���'b�3nX��i]���V͞���WU{g����j�6s�0e�m5J����1ҏ�.�T�N']��>�w|Cn��q�������S�&�&��,���&����ە���1Ϯøm�q[$�`�a���<�4�P8�e6���޺�32i`̭��ݖ�թ1ʑ���M�V�Q�zL��zژ��`z��t�H����m��9�[,��,fM,̚X��mHA�I�7D�� ��0="�H�����ٜ�۟+<�-�4T$��m�NK��K��	 ��ȐfdH�K���ӝ��Q�v��X���z�Y�@�ѣ����7;���e��q3��f�<�W6߿���`�*`���T`�Tw�1  ��R�ʙ�3N���M,̚X�z�8�(�R&�$�[S�*0$���
�2b�M8H��mI,fM,̚X;�� ��� ��Ԙ�H�Lq��EF�L�����~l~~�Y��u���0V4��W<�8��ݬ
�v����'%�T�]Q�l�����ʘ����+ϳ�j�`j��mI1��I@p��9�����I^0I�06�9j�zbA��{��v"@��J�.�%I�
�HL"� ��X�bD������F�Č!1P ̄T��`��x�A�_�]U���!&��0p"�a�!��`�
!�c,*Ha\�	!1"� !�adl*sIRHHC�Q������	HT�$!I��2b)'�Ej�ͤ!I D����:�+*�a	*��8*�؋�#W =@CEG�� A�U�Ϊ��
U�T��7&w������ �w���N�)%X��L�
�����+��%Gz#0X������L������36���}�Չĩ@rbjRJ��[�j�t�:�e�36��l�'����]45;��$a��`����J�s�l�;�Sd#�(��ڒX̯J�{aS ��0�����R0i�*��ͺ���{꯫��ޖw޺�7�����%@7J�K�*`�����3�d���1t�mI1��I@p��9������I^0�T��ҙs�t8��cU�0�d�i]q��МW��8�6�iҸ7&`:��2Rr&�T�m�I�`s7n�	%x�6L��zژ�goN�8	,�;�s9Ա�$�ɕ0[S�׌rJ���$`�;Ռv0[S�׌	%x��;{y���(U!BiS���UIw���;��Ձ��� ݅L�H]H0Bŝ;�$���`}m���	2�������pH�B$$F�F�  ��T���S��nf�ͣS`�����u�ԧN8";���Mt�ҁv{A�佳P���c�k�R1�����ӷnv�����v���Mf��nW-�M�nޖ��:V:�m�j�1q�N=��KV�9�^�֤���5HA�ݶT����2���2A�m�;V�U�-Ƹ�묭&�W+�Y��m֮�q�r��'V�v��{�w|?yi95�������;gꆋ%���ų5�,BhGM/27B��aVڋ����ߗ�� s*Fc�9%h�Oŀw��,��,wv������:� �*m��7rT�=mLm�EF��G$�17L$�n�9��VfM,��e��t�bl�IFۤ�LK^0$��v0[S �w��A$��'%X�4����ݖ3v�����-�*:�:K��a��e=�wn��z@��n:�F�ł��b��#�1	,A�Τ0�T�=mLf�Ձ��Kr��NH�T�$���$�������h@�L��������T`����b�\]H0BYӽ�I��k��Q�l�S ��0�&HH�n�i�*�k�=��P7k��;��j�n�g�����$%�w�R��eL������I4�:���#NTm9N1�N!@U��j{{9�y<���܍�1�ۓe�K�����-|�W;#����
�ؐ=y��
��5��������{�8|�n�rX��R]�UfD�z�"u��8�;�j�J���9*�����;�6Yu���`#V*DX�� @�/D_��~�n���;Y�Ϥ��"8��
�����k�f~���0=��蜑�B�
I��X3vXI�Y���/24�
�2$t�;�.�i+g]N0k��5�����9zzY�n�gh��iz�W!�9h�ݺ.��U�������
��$�̏�I�]��@3���d���Ɯ��̚_����7~ ߾�06Z�v�w��%�q,W{�$��$ٙki�r�vT���Ł����)�MD�	$���WԾm����}��J�.�%HbnP�B"�D��0P6}����w�/�ۙ��Fۤ��3v�����Un�\ ��K ���7l�?���j��y��ɯ%E�$<�Y�z+)�hFm �7���w����-]�c_GRRM�I�\w}u`��`��`s7n����l�HQ)���RWy�&�8�� Vnʐ*�%O�ꯩ#�Oމ�*�m9,��&��%x�7eL�j��F
9
N��!���*�|���RUy�m.r�v$4�9� ����w�IcI^0?��$�/ o�|��^0,�p+LOjSr��t�� �rt���3:v�s$�2t�욤�$�
�dq���tk�r{�
v��ڃmv�X���1Q�x��v[��p% �2:XƝsG�;F�X�P�Hڷ���/���s\1¢�Z ���1�k���m��m��n�<�.���݆ԏ8=�[N[���3�]w/*�j� ��I�K�V$�:��G3�]v�N{Aڅ�Tۼ{���3$㳳t��˝E�Hv�̎
ΐt�m����c������www}���p�$	{v�f�}���`���׌	%x���VȤ��l�(I`����謹W�4����H��� ���ԚIs��R��n?���m�NK��]X��V��� ��� �f=cUN	F�'!Hji$���� y� �Ȑ��Iw=�U�en��I
%1(7*�;���=mLm�J���\�>}��$"���Wn�*����eF�-��1C� E�;o����������
4P��� z�%HwjM{�]�ā����)��!�$�9�۫�����M6�$�^��� w� �ȝN���	�0�rJ�7vx��S ��0=��`m�{�Y��N�p��U%����{���n�Xz��ߋV^�I)�Mą�,�j`I���m_v�����\\X�Y%l�vB)q��n�1ٛn{p�)����wK㴻���}��'Z�i����bO�x��W�v��=mLrNގ?�8%T��`ff�_�H3=�`��,�v��;Y�Ϥ����`Y� �ȑ�I�$�iI&&��m���d���T�����DuU $ےXy.�},�z�����X~��K3ޖn�~�H@����Ӓ�ݵ�l��zʘ�Up���.��\k��:);����<�5��C����ny:��\�6Z���#W}��+��j`�����I) �8��`��~l3��Kw��;�u`b�dRJtS��@nF�07mx�ݕ� ݵ0/2Kq�$i8�t����3��X��{�{��4�B��}T:*T�k�&��;Y�X���P�J�������k�{��
�ؐ*�%H����kY/K!M%"��G�Q<���to"6�ι��)��ٹ��=sV]�i�[��nژ���ݵ���_�0>�߾I� �@J7$�wv_�H������Հw���}UT�����)������.�eHW���'�{� {���3D˄���I�*��}��3}� {� �Ȑ���w�� ���z�G�U���`��wvX�oI=�����騩�E$A�8t8�U:��. �G�D�`�`BH�`��$�b1"���
!�c1D� G 2�|X�3�v&"!�<
��DO��*EZzRY[h�L�FaVYB25�*��B!B�E�$��b1Hr2TBU� �	 �""$��$"� ��� ��KX��E�j,�`��W��� I8$�F$�`@��!	�� I�ʀ�I	$!$"�B�#F@��D	J7$$���"O8T�u�!	[`B��0#FҌ�$���� BIIHHq E���
�ww����/�촫�V<Z#v����J6i2$5�������r턼�Ӌ%\t�G��i������!�L��J��4`0������M����v�;�g���\�&ɋ ��,���:^�;I�,�yN�W R
Z����5� d�Z��7F]K-�u�ٸwG;j���Y���NK��^Cis�j$0��;��6{f��Z󝖳�%7<��jčDګg��޴O6­�Yۛ��1r��-��oɬ��9��
<h�vWMumn���� z�^ϝ���;*��+++U�����qgAqg�����	���gN���,��ݮvN:�[=�j'X9�'H�5pu!֦,�/�2]pH����Ԕ�WWH>HwPJss����ڙ�畷Qu^�q�	`�4����lm��ƻ 2�/,!:ַ(�v����1C�����uȺ.,�d78�s�e�f��7����;�dA=�ͤ,���/:�8�Om5O9N���ЪVm&�d�py7�k<�s��E�y���]�V�}�Ho ��l'g�s�H���wm$l��m��燶�N�6��ՃY-Ğ2�j��RD>(� [��)u�]��T*��۝v�8�Im J������`�������v`x�9x���pwW�/O.��uѤ�֊7d�q!́�T]Ca��caTܬ<rk�<*���ʷ<����n�r!>�B[�E��Nʙ*\�@��sS���qm�r������Ν+��>���@W�f�)u��T�=j,m:���k�Ô�U�HD�m�%���h���`�%-k7f�m�6�Hg�͋kq����)�-�li��Mڴ�����6-�&'�ɳc;q���vx���p<��p���9���5�]�V�e�v*/	rS
7kz����w=���WYGd2i��k����;!��ewm	��Y�d�L-� ��e�f�J��Z�2vi�T�Iu�����S.fۙ�&f�h��|RDD:�>�*?q@P���5�M���晔�gw7fVΥ���6W��on{`㈀�m��]�P�r��WXx-i�F��unu�\us���W&g��c���������Q��(.ݺ�;=e�۪Zx}Vjr��ޮ�ƶ^r��m�[��ju�9͂ڣ����M7X�K7��mP�I��o�Pl�ۏF-��	� �j��t�y��s�E۶����.hO�{��p��~��8"n���lu����gD����j���L����������|}E]�3�g1w�*�����`n����U}\@w=�`yV���H�m�QȐ*�%HW��ՙ�̉��o�2�_����P�J�������9ݩ�{eL�^0fʎ���0]3�Q�֒Ms�{� y� U^J������r�e??'t�(ܒ�=W� U^J�=W��ՙ�6����ׁ�G �]]�Iӷr��% ���z�d�2��f��a�_����G��(��YT�r`���Ձ���X;�,�͖i�&\$`7N:M�V;�uyMy&ڥi�M���y�U� ����J��@�8$� �we�seL�33������oh^��,��,p�R`�SvW�l�}��K��KUn�SeBE��ҎK�+�ٛ/�� l���=������Mfj�9ж�^�ڹ��z��t�<��{k�q�+]�W//�*F|ѱ!�]����/%H�2$�y�&߸y����M}$2��ܫ �we�s����sn�w6��RG����M
�D��
�ؐ*�%IƓ~���D�}i4�&�Zi��*@=y� VZ��9���Gy����6�O��oԤ��T�s���9��`f��e�J`�(�7&0=��`�S �ʘ��`	��~�j���\�v�4���σ��K�.c�
�unr�Ǜ�����,�N��=���07ey��/�}߃ͨ��dR��nK �se����X�mՀs���}�F��~�ʑS��t��v"@�͕ z�%I�����~� �ߥ�r�64��ȁF�)%X�mՀy���I'����j�x���<�^Հz��F��He5Q�V꼉 �^D�꼕 z�%H$�J���S��ɣU��M]��2��L�a5�ۍ��ڱ{%�PY银9�x-t���a����`�~Ll��^0l���b�o$qTr�6ܖ;�u~�����fo�]Xo�K �se��n��RJ@�(�IcvW�vT�=���׌�n�����*RP��`�l�wvX��Շ�fo�V��kͨ����I0m����vW�v]䓋E{��{p���!M7L˷r7zxY�Q�+k�d8�Ԏ��4��*v�7{Jw��wi�OsnR���ٶ�]6ôŉ/:�����aMs��1���;pW ��Mz9���A���g�6�e�u�2��V��/WH9�n�Z�4J�h�@7�孴u� ���5N��<.�ε�"��c��g@�P)�-g���k�;S�ط$�]����5�$;����\��v+i��D�YɊ����u�%�Z^cBd��'j;[n���u�������-��vW�vU�{�l���7-�4��8
4�9*��vi��������zX������ �f�4�BT�C�Ԇ%�0�S/���ʱ�V�,ƛh(L��U}Iw�������Q�nʘ�{x�W�g�W;�v"@�fJ�5���Ξ �͉ �we�Wk+C6BGRG#��!��,Bv#��2^q\)�W,E��y�z�p�q�-��܎�v"����@*�"@+/#�6��K���3~��~?~%GQ T�,��&�i�&���^D�Wy*@�����}�����jIN�p�GC�X{~Lm�j� ݕ0/3gnw�u&J�Jn��X{諭����V秋 �se�w���9Y�q��@���`Uda jm�˽����HY���������0ܡk
[.*�m�+N�n���yB�g��dvh�1�M$���f���F�r�U�U�Vd�i������`{i��6�P�A�,�ݗ�8]�ʐ.�4�
�ȝi��i>������⣌Lm�,�߮��f�"���W�x"�Ow��I'�w��'չ�eԒ�&(�9%X{꯾����`{� Y�!���^��:B���*N4�`��`~�����N����wf�Uwt*9$d�D��jsv8�7-��y�0�e�<'3�%��^Pպ;;Y��Q�3�g��I0�S�׌ک��������Kʳ}�q2T�St���2T��M�p���@/3b@*�����*��|w�����&�Iw%�7q�/���S ݕ0=-x�=�����F4��,=��UIf鹿fnā�̕!��k�$��iL^֒���&ڠ�*U��vX���������,�͖}��7�)#�	:a����cN��W�E�Օ��ƴEԖ��j�*m�#�*�11�$�9�۫�ل�UfF��^�{� b�ӽ%DB��w��RX�ݪ�v��7mL���?��Qs$��K�Mɶ˳4��C ���0�Sv׌ڨ����ܒ��I�,=��W�Ig����ݕ ]da!�m��]�ā�W�z<��7n������{��~�@{߽�@g3~�UfD��M'���&�Ϫ�t�/A�F8F�j�0���V��Ol���zx['8E:�3�ʘ����!�$x�f8ة=۰66p��S��]�"a1���;���]�vu�6��a9ݹ=�gSU#j�\+�g����qq�s	�֣�%79R�۳'b���3�;S��^vMfB��p��۴5mŷ-�vGi�n�8�{r�����ud]z�V�r��
R�[K�������{�o��/�_��n��f��Q��1�Z.��0���mL<d��J����2F
4�9+ ���`W*�Yy4�o�
��R��ӫ� �"9����}��}�A��K�vT�U����m���l�x��Ts�?.�u�I�Ɂ��v�0=͗�nToT�R�rK�ݺ�;݌$
�^vCSI.r�v$[�w���|��s��X�ݪ�se� ݵ0=��V{Ou(܌�䨝F!@�$䘊q�o5�I��4;{$WY�k��䆌���{�o�î�D�$8Vo��wse����~����O�o��rJtS���������QJ���!H!�K�.6����/6�H�H�^v�W�Wԑ��}ϜNB��$�s}u`w�4���R]Y�v��K �fli�S��*NJ�3�4�:�����4�$�o>���j���;���8GN��Cy������_�����j��~�w�k�G�nJD�V;4OU�X�.9�*�䝛�rV5[�{����{}�_YSn��/�q�=��;�u`w3n���w*7�)��4����wn��K�3w�Rs7���2$Y�w��'Ɏ��7%X�mՁ���f����PHA��D���ڇ1a�
$@��D�Y>B2�qqk���ȱ��1�!�P�">E8�M�0�W�.A�1~�"��0b�2�(Q��D��D"�B�@�4c��Cz���c����$'�=C������U=D �gj*� �%Ɠ~M6�1 VfJ�ax��aP���=UUU_����~v���`{ex�ݕ� �Z�������{�v#��̉�I�ҼߩP��������mG��H�	��D���)�a��*N�^Ш�Q6���|v��kt��:n��X�mՁ���X]�~�� ;�����MB��J6�I*�ݕ���z�=���W��߹��/|ƾ�QQ�(��`uf��;�,w6���sn��<�6� �A ��v�9W�^���T�[I�Sj�+� a�+���{��w�73�w6�7:�����&�׌�^07�/X��?}U�W�^�JC�9J1JQL3Z�m[<,�]���gT���+)Ƹƺ����e.��&:#���7}�����k�wvX��ՀsM�2TaL�RrU���z��p6}�`l���^0������A��v����ݺ�Ԗf���ś�`f:͂�R'T�RDH|�mr�w�@�͕ W*�s�{�`��F��9�mRrU����X�I�����{� z�%H�M$��~w���Q����IEwd�<�n{m(;=p:�ոܩ��p����V��a��s���(�Q�4�����]S�ё�f��˧a.����t�b��ݬC�n�v��n�2v�-���nK���kW[���mӳ�E��NC�rrr�,����K���u��2x4Y�.�����;�`�s���]�@7Lu�h���1�)��CK��{��H���e:�îe�D�zm���v2�u:�G!C \�*"��qu-��HcH����ߝ�s����wn�w6��ܧ�ڠ�$����0=��`n���z��?��7��7�H�(�JLm�,�߮�w6��Ԗ,�; �o����Z�t�)&�'$��K���X�|��͖;�u`�tL�D�:��`uw5��]����z���sn�o��D�B�̺v4[t\Td��.'r!�'�a%(/t.���U��ti���m�0&����y-�orr�Xn���ap����{�{Þ���i4&ۄ�oZH���*@+7b@=[��;]Ǭj��(�NJ�;�۫ �̉56�¯v$��RJ��ӼPuugN#�X�6Z��T��k����f��`{i��Tu�
I`�Ȑ>i���/w�*@*�"@���-HRR4 �]�n��mATRx띦�X��NX�l�&k��0�9yX�7n���{�vT�Uy*@*�#�߸^�;^�y:�n�H���U����X^dH�2$
��S���8��ΐ����]]��B��ؐVdIm$����o&�Ձ��u`3^���0n$��r;!�6�9W�����T�����,�zXj��J��*t�)$�6J�+��j`�S �����.�pk���\εrH&���N�q���q�ܵ۱L������k����nh����K���0m���� ��zƪH�N|�F�X;�/�U��$�ؐ*�eHW����k�6�s`�{�u��`�zX�m՟���ꤳ7�V��K���#�J��ܒ��^J�*�%H��$1�M��I��Έ'_}����I<=�~�nLٓ.w��B�*�%H&�|�͏ U�ā���XQ���i�!ʎTlIR�ɚq�-�;lmq�
�(�8�w+�.6^��uӵ����) �^D�z�"@�^J���K��u��ߥH�~�r"C��;ð� �ژ�^07ex�=��~��g�6��?��ڡRm�;����P�ܖ��e�r������q,`n��{eL�ja�~���~�0�~cU$b�>j�r��͖��ā꼕 U^J�!��k���w��;e^JB�F�6�\:k&���x�����M�L�9�.�D8w�r�6uoC�Kd�m/�Ѡ{Cg@.�{s".:�x-��U[����ay۶Ɲ�k�����s���"7`���њ8�AlgT�q9ۜ��ɺ.����h����v�Y�@ð�k&�x�l�;;�
(�]���
�py�^W�Olr/ ��/s	�ݓ�/��>f���g�hٙG��g`�n�`OC�%�r���$�l�^8������שׁ��$nN f����sn��6��9��`oi��#����J�ܒ����+��0m���������1�i6��rU�����w6Y���朗;���;�� 曢d��$�����)M��{y�D�^}�H��Rw6���׮)'�i�RhrK �wc�+���T��)�;WC�.���tLe�v*W�l�.��ݶ6D��B�݉:c���"U�V��BI:N��p���vW��*`�S �I�ӫ�ٻ��̦n��'����)@�}<�K �{���sn���zơRQN|�F�X;�,�ݖ~����3}u`��dmP7%������_�������^0l��w;�GeR��5$�9�۫�~��~�t7ߥ�s���+����kdQ�P����2.���.��m69��u�8��ڤ���k�����"u�4ۢ6ܕ�37�V��� �we����X4�%JuT�B�X�=�����ϾL��l�U�5��)�:R��$�w6X�og&� �����?*�����ܺ���K �4'�*�EN��$�lT`{ex�=���0d��8�r"�iS�;�u`~�w7Ӏ���9ܚX��M��r�JQ1�@:�V�$�@t��V��'�V�(�Z���*9�ơRQN|��`�l�w6X�M?qs}u`��8�aCu�� �Ȑ=WH��R꼉���8nS[��D��:rK��Ł���Y��;��`�����S�N�M�y��l��T�=���~�g�m�I �M'�ͺ$��9�.��9�#��X�=���0=�Q��ͺ�8��[�rINA"T�� �.��r��)Ä;,N�u/�7�	֎Ѻ)��
85C�X;�,w&�;�u������F�'Є�&�I,w%�^0l��{eO������S�ȅn�p�;�� �se�s����ri`���5
��q�����Ms�y� y� z�0��5ʼ�) ۭ�9>H ܖ����ͺ�=W���y���4�P�j-HRDH#Y$dX��: b��zy�4@8�1"�1$I"�I�!����)� F@� j����+Q2�
�.�!!��"�,�������0ˌ.k
`�B�K��a�����#0HSIpe!�LI(7eB	��j	��BAj��0ёWP���Ȑ�!�0$�@�`B,*�GE�a ��4`5V+�� ��E�,�A�8��C`@�A�@�$5E�R�y�ܒfn��ӷAS�2�x�Kf׮B�ʌ��=�=�bu�c<m��A����bHmۓqYh�u�b3�M�]�M�m�HH;6���t�ݹG�L;]�p=����"n֡���9f�E��0\��Wf�e�=m�Y�QW�ڨ�5��A����p���3�����-n�*��m��,xM�H�n�x�l�n�����s�^{k�2�oK�a�����=����n [���N�cVݜ��J���[��-v�lPV�S"�ձ�-q��C�jM�s���2�j�VU���5�Sn�ggY94�Vy��\�j��tU�uF�mp��+�Fj�3�L3�r<ו.��:�W��溴]P=����dmu�`�DsnY���%�����x@�7*�P���c��[���igf�z��r�㋥	�W6���L]�ܠHd�ցHq��G���)�c�5��;�8nwnB��1���2.-��5����:->:mͨ�L���rq,Zk�:�����p+�-�lЫ��!y� �=��EP��*��8U���+�G:����H�¸Yn���lL�z�@2�#$�CDAUUee.YV�!�n�Mn��սw��9�@Ms�ng�:�ex�;��j�X��6���K��Z�b8*��auYv�$��R�G��1>�5��y���]C����eo��vp�cCŎ[Ȳ@�n����λ:!��'vl�k��@@>Iz��� �����m�$l;����ZN�.����/<��*ҫ�.���l�b�b��sU-UV�	gftUW+�Sp�6-�f�d$�ޮ$��F��l��]��C��]bm,�g�N����&��u�l6ct2G����]�����)��\��L��]����!X���&�]h�ðb��9�s���+�� �3��]�i5��o��b�J^vl�]��ltJ���R���V��<$B�t��W�/��Q�C��T�8�S�A�`�|D�CQD��UW������2S��$Ol@]��5�ZXr��r���͍����5όJ�����ILv{Z��]�����n��6�=F��η��kX]�o�1�֎�.^;����M�9��n��=uv��H���l7,/l�m�]8���с��.L5q<1L����K��)d��=f�u�z���!��k��5���].a$��M�4�و h�i�2�9fȳ�������AC�^�)q���X-��Ӟ����#rVfwj�簵~��%H��R꼏�_&��^o� ^�~N:Q6�6ܕ`s��V��� �^D�꼕:�|�V��aB�s�9Υ�e�0l�����+�Uf=r7
cN���rK���W�w7b@�͕ z�%H|�K��͉ ���I.t;Ӊ$������ �se�s�����i�-�%JDA�Ru��F��*ǧA>v��Zs���i�ۓ�.�����u-�6B��Q��I+�w7�V��� �sg� �o��+5��T
r��9�R꼉Ʒ�6Ҧ�h��ډ7�u`s��W����H=��q6�I;Ԙ��`{ex����{eL�5�8�(����jI`s��V;�*@=W�!����*�b@1f����u�w����c�+��0l���ͺ�?W�UU]f��E*Sr�$t�F-�[-����˫R͓b.7���9�	g����w�V]�9R��i�] ���`�l�9�۫�ͺ�:�1둸1��&��I�{eLl��^0l���U_|�g��	P�8�`�)$�;���y*N$��6�14�Qnr$՛,����!NDF�t��`s��V꼉 �^D����I.�oԤo~c_G��('*�9��`�l�9�۫�ͺ�7��Mbc��RTmE��k�.j^��\\l�D^iS;95�tܓ$��{���gQ\aC�����,w6���sn��͖���q�IJS�6�`{ex�ݕ� �ʘ������׽^N?�b�rU�����w6$�$��
�ؐ*�eH����G$�X�=���07ex�s�`������'���wws62����&�07ex�ݕ� �ʞ������t�n��H[�Y8ˌ9�bNu��V'm�Y���/,������Q�]���1q��I���vW��j`�S �f=���ȅn����6����T�\�U�ĀU�āUy*u&�8�;�k��R��Q9V��K �we�K����37�V��[� �� �rXjM4�ʽؐ*�eHW��5&�\�f�X�k|8� p���$�9�۫S����^lH�2$.��i������w���7"b�3�K��t�����g��ډ`��+tnzA^�˵cmc�&�	�y�`�3��v���ܕ�v	����9%���`K:pnsu�k�v��p�b?Џ���kb:q\!�r�0��K���a��uN���q�`�Tmf�����[LC�=�5ڧU8�!������<�'&�Z�;�)Դ�[���s/nj{������Md�:�e&�d;mae���B�ɹ��$5ۓ��8B���F���3}t�=���0=��`���Ջ9�����K�T�=eLl���VV�H�A�4F�'$�nj`{ex��+��0	9�pX�3��s��u$����6W��*`��`�̓q|�Dm�J8X����6_��7��`{b� �2����F4�	�u�#�O8�2��Np��u͸^a�WK�p���g'��8�n�m�������T���F�^0�9Q�� �-�ff�$����抿��@��~^�W��*`]���uutŋ�s�]I�튌	��`�S ��� �ݭN?�b�n36��=���*`{b� �%��Y�$w�K�T�=%LlT`zM��;�4v�P#��RS���Ꮊ���=;��܋�K��a�a5�"�;�kC��m�y�9�I0IS���`�l�ůiJ�j��SN�$�9ܚ?��g8m�<`/ɀzJ��J��/��4�:Q���f�X;�,Uu�UW��b��>���K���I;��K ��=c_))
|��`�l�IS���`rr���z���z� ��0=�Q��+��X��AhR��*?[�����G�j�8�̗c��8mn.R� �7/b�a��E��s�]K�l���+��0IU�en֧�A��m���u{Is\ �f��xO�U|�sLԇ*R�pBGyԱ�l�&�*`{b�ٛu`wcm�0l"j�$��W��}�ߢ@����=w��2�L��m�������� � � � �{g��r��t��f��A�666>��~�|�������>A�����o �`�`�`�}�o �`�`�`�}�I�񛙓si�&���2aغ5Kj�)[ۧThƸn�^���8���q�{}�}������̗����A�A�A�A������ � � � �~�����lllo������lll}���8 �����K�L��]��pA�6667߻�x ��{�x �~�?N>A������� `�`�`�|v�ٙ��0�Jl�����lllo������lll}���8 �{��|��������>A�����~̻�$ۆ�3ww��A�A�A�A�������lll}�xpA�6667߻�x ������>A�������sf\6fL&��͜|�������>A�����o �`�`�`�}�o �`�`�`������� � � � �>����3rWI7vɳ[��nA�=n=uZ�,��e�3�����M�އYpB'�:�c�P�t	����tV�ht�D68�Q7��L��u%�q�ٺ,�tt)?��ۧ���h�vR���ѳ��62'�fR�u���[v�獜���n;p3[v��ٴ��$�N��J�]�U���;GcC�nGU�3Џ=�ӥ2I%2�B�m�-��5 �=�]���=1I��j냴ʫN,r��6���܄F�B K^�%�b{9ז�l˛���A�A�A�A�w���A�6667����A�666>��~�� � � � �������lll~����pْfI��3wx ��{�x �~�?N>A������� �`�`�`�}�����A�A�A�A�����L�m3&附�����lll}���8 �{��|��?��@29�o �`�`�`�~���x ����ٙ���v�]͜|�������>A�����o �`�`�`�}�o �`�`�`������� � � � ޟw?d�Y�d��ٙ� �`�`�`�}�����A�A�A�C�"��~���}���������� � � � �������lll~�����w--�t��ThٙG��g`m��'��*�O^QJ��	��^-��wffL�e)�3w��A�A�A�A������A�A�A�A�������lll}�xpA�6667߻�x ��w��3srI�M2L���>A���߻�ӂ�z�H�R� ��`AV�/�?x�A�67��)M'�4�8�� ��?&�\�m{���Ө6:#M�X��Հs��MM���
�ؐ*�4�axqv.(IBA�%X~��朗�鹿ww���d���f�XX,{u
m�1����=%LH����� ��0/4� �g9���Ѳ�v�Q����Ue��fl�of�e��=\qՈ���w{����!z�,�玤�ھ��`���*`�����r%��G��u`��`��`w2i~����H6�o��F�#���;�RY�뼉U���>%H�$�����P=�
��0CH:K��h�[��% ��)Y
9��(�`VV\�&ebRI�F!^LR�G䒌#)+*K�a� �%%ae)�SU�H�V�Q�D&S"sN���F b�RF�*��Ex��_EG@j �U�EW������uQK]KJ�M��.��$��R.OO�vfa$�6R�.���Kı/�}��yı,���ND�,KϾ�Ȗ%�� �3���jr%�bX����|�ܒm�r3sw��Kİ~�{59ı,O���O"X�%�}�wjr%�bX�����yı,O�TçK���˹�l7wl̙�3 �n�qsi7i��gP���o��?����~��	�\�٩�Kı?w���Ȗ%�b_{�ڜ�bX�%�wx� �&D�,�MND�,K��w��i�6�f�7N'�,Kľ�;�9ı,K�~��<�bX��of�"X�%���wÉ�Kı>����z��f�w��oq����߻�O"X�%����Ȗ?� !�2'~��'�,KĿ~��S�,K��>����36fL&n�Ȗ%��� ���59ı,N���O"X�%�}�wjr%�`~� =9������Kİl�������ܸ\.�bX�'���'�,K��TB9��۱<�bX�%��oȖ%�`��xjr%�bX�������J��&܌�P���0�
z��E�`��[�v킓���2�N�����7��,K�s�S�,Kľw��Ȗ%�`��xjr%�bX�{�|8�D�,K�O�vfa$�6R�.���Kı/��������(!]��,߷�jr%�bX����É�Kı/���ND�,K��^�74�n��!�����%�bX?}����bX�'���'�,�XdL�~����"X�%�}�����%�bX��陜�pٙ0���͚��bY��"{����yı,K����9ı,K��wx�D�,KﷳS�,Kľv}�ri�m3vۛ�Ȗ%�b_~��ND�,K�9�{�x�ı,K���Ȗ%�by����yı,Mr	 	"<�^���,�����il��34 �̼�&D}.8鋜�uغK���<G.v:��t���ٞ4d�;4l��q9�����o�:�^S@ug7.��':�/C���؎��>M.�e���*F�C������
b�J�5O8���b"�����멤65ܠ=�c�c��&r狖��7,�j[����pk<OBx�Knգ�[�J��Om�+�����?���������O\�k�:5s.�Vہ�vi��u9�:⫰��]����ݓX�G��rə��;ı,K����O"X�%���٩Ȗ%�by�������ؙı/����,K������]�r��2���'�,K������Kı<���q<�bX�%�����Kı/�}��yı,>��36��n�̲nl��Kı<���q<�bX�%�����K� �ș����'�,K����jr%�bX��߳�2�����˳3N'�,K?�FDϻ�v'"X�%�}�oȖ%�`���jr%�bX�}�|8�D�,K�O�vfa$��R�37br%�bX�Ͼ��<�bX������5<�bX�'���'�,Kľ�;�9Ƒ�#����^�N&��1��RB��Y�ڗB��K�\%�N.'0���7BSs�4�!�����%�bX?}����bX�'�}�'�,Kľ�;�9ı,K��wx�D�,Kӽ33�.l�s,�.fl��Kı<���q<���*��D�%�w�~ڜ�bX�%����'�,K������Kı/��v\�nI��۹�7N'�,Kľ�;�9ı,K��wx�D���D�=�����bX�'���'�,K���~?��is�];fh�}���Y�P�~���x�D�,K������bX�'�}�'�,Kľ�;�9ı,N���ܻ��s7.K����%�bX?}����bX�'�}�'�,Kľ�;�9ı,K��wx�D�,K��L���ٶ��m6�0���[6�яF!��6��yD�ԌKa��������wz�}��X�D���^����oq�{����yı,K�s�S�,Kľ}�w��=��,K����r%�bX�����2�ɶ�%�sN'�,Kľ�;�9����,K�{�x�D�,K����r%�bX�}�|8�D�Q��,K>;l��	���6]ݩȖ%�b_{����%�bX�}�wS�,}�:aȜ��|�É�Kı/���ND�,K�O�o��a6��)�����%�bX�}�wS�,K������%�bX���v�"X�%�|���Ȗ%�bzw�fr�͆d�n73wS�,K������%�bX~c�~��SȖ%�b_{����%�bX�}�wS�,K���߿����b�zuAER�t�og�"�xץZ�ϒ�ۄe�+Z��`�j���oq�ı/�����Kı/�}��yı,K>���Ȗ%�by����y�q���~~�~����e�>ﷸ�bX�Ͼ��<��șĳ�����bX�'���'�,Kľ�;�9ı,N���ܻ��s.̳-���yı,K>���Ȗ%�by����yı,K�s�S�,Kľ{�w����oq������X�A(�*��o%�ʈCb}���O"X�%�{���S�,Kľ{�w��K����(�{pѪ�9�����Kı/����˳&�n�.��8�D�,K�����Kı/����yı,K>�wS�,K��߻���%��{�����_�
lq]	3qX5ɮfY�"�m��x'^zѮݚ���.����fl)M�wjyı,K�߿oȖ%�bY�{���bX�'���'�,KĿw;�9ı,N�}{|��	��p�fn�Ȗ%�bY�{���bX�'���'�,KĿw��9ı,K���<�bX�'�zfg.]�%̳q�����bX�'���'�,KĿw��9�����ؗ��oȖ%�bY����r%�bX�vw����6ےfne�Ӊ�Kı/���ND�,K��{�O"X�%�g�wu9ı,O}��O"X�%��t�f��w���l��؜�bX�%���x�D�,K�9;�۩�Kı>���8�D�,K�����Kı5 ���I��� �c�N��=Z��Z�iw=h%{knx��m�秱�i9�����+7Zxz�e��7Z��gb�%P>�͇f��K
���c	�;!6��ӵcu�����nd��=t��8��]ήK,���V��\[�o5�,��� ��R�jq�cG��:���:_,��o2ggd�$Q�h��l�2�[mUڛm�&9���fz��:nWV6�����Kv���c�O�w{��������(�$�4�ܸ��9oGZC�,vQ���I�,�(>;K6'z��&B������{��,����r%�bX���|8�D�,K�����Kı/�����%�b�o����ǚ	E�U��{��7���wÉ�Kı/���ND�,K��{�O"X�%�g�wu9ı,K���ܙv��Jm�8�D�,K�����Kı/�����%�bX�}�wS�,K��߻���%�bX�z}{�3fl)M�7br%�bX��{��yı,K>���Ȗ%�b{����yı,K�{��,K������0�wf����yı,K>���Ȗ%�b{����yı,K�{��,Kľ{��Ȗ%�b~�w���h�uö�ZsS�us�X��;8�OMns�2��n��/K�z%y����r%�bX���|8�D�,K�����Kı/�����%�bX�}�wS�,Kľvw���M�.3l�Ӊ�Kı/���NB!�D+�2%��~�O"X�%�g{���Kı>���q<�bX�'�ӹ��q�.fne�77jr%�bX�w����%�bX�}�wS�,K��߻���%�bX���v'"X�%��}/�˹�3p�%��'�,Kĳﻺ��bX�'���'�,Kľ���9ı,O;�|�yı,=�:fmsv�n�̖��"X�%���wÉ�Kı/���ND�,K���8�D�,KﷳS�,K��DL����l���."+d�:�ꎫ��F�:3��S�krs���\Q�w\��6�Y�Cw���7���%�~��v'"X�%��~�O"X�%������lD�߻��$�I��ݙ��3aJl���I�{��"v%�`���jr%�bX�{�|8�D�,K�����Kı;�����0�t�!w3x�D�,KﷳS�,K��߻���%��/��:yȗ���ND�,K����'�,K����39r�.e���͚��bX�'���'�,Kľ�;�9ı,K�~��<�bX�&A�y�jr%�bX����n_7l�&f�]�8�D�,K�~��r%�bX�����yı,~��ND�,K�~�Ȗ%�b}�^�ݻ&�ےB ��B�Z���VE����X���Z��5��kn;�̙�2e��ND�,K�߻�O"X�%���٩Ȗ%�b}����yı,K��ݩȖ%�b}�K�r�Ge̦�e���O"X�%���٩Ȗ%�b}����yı,K��ݩȖ%�b_;�w��Kİl��陵�ۙ��2�͚��bX�'���'�,Kľ��ڜ�bX�%�wx�D�,K߷�S�,KĿ��ɗa�!�d��Ӊ�Kı/�gv�"X�%�|���'�,K������K����X�����݉�{���Kı,����3fl)M���9ı,K��wx�D�,K߷�S�,K������%�bX�߳�S�,K���ݞnd��fWT�5�[�X��Iēcv�=\l
Wv*v��y]��X9qt=U�h���U�������A�����Kı<���q<�bX�%�����Kı/�}��yı,O�;fg%��K�e�s3f�"X�%���wÉ�Kı/�gv�"X�%�|���'�,K������Kı<��l���&\ۗwN'�,Kľ߻���bX�%�wx�D�,K߷�S�,K��߻���%�bX���~�C��s9����{��7����~��<�bX��of�"X�%���wÉ�Kı/���'"X�%��}/�˹�3f	.��<�bX��of�"X�%���wÉ�Kı/���'"X�%�|���'�,KĨQ�U�\R@�E���� 0I���>@��H1�� 2J�ki$KBb�)�$LaO����E��`�a�K�St��
!�"D� �b��G	Hu�SȔ":!Ũ�0]�$ @ :sJD�R���`I@%}_W;�S�����n��!QIGe�=1��nz�\[�sl�	mλnz�Z�ud����m=�jӷ� $P��T����iK���m�6I8���N�niwMD�U6�'ci��g8sg��k�loG\�\FƖ��0�Þ�i]�7`ׯ���
��j����]���uGYT��ʷ���}���硂��v��d^[	��A��������i�����P=�e��s`��jM�n6�Զ��+��I9��;j�i��Ŭۑ2����a�0Z���Ɩ�q��V�C�v]�r��l�\q�ҋt�g��%R��`]�[�N���c�z��M��5l����8)[s�c+V�� /*�8��7/d�P����n L�6x��[nM��vۛ5mr�H��'=uB!��nMnQ%�e��ո+I���HV��ڕ�1���{p���Vϱ��7C�]�]&�;��S`����4�3
4���❞t���/�;u��*#�x���SΑ\�6�[\�ηY�۵%��WO`��
���5���ޒ�[m��U�g*q�B�U<gaUwn��z5���l�֌�R,�PJ��+4C���mKZƠ�󓠪,�نE�� ul X�i6�p�6�M��vv,��+%�����M],<͖��:�v��UU�m��m�������t%��T�B�;;=תU'j��ֺ-�76�]p8-n���-@G�^U8���=�����Z]Ol��R��=Ix�X��
�96vz+�kI�X�J`�ݖ���EJ鴉5u��bt�!�UPr��˵@U������;�Ηkv1h큠6��t��]��h^��ڮ�6�YhĆ����λv�n��b��4�l= v����V!�q{c�����m���cn��T��;+�nc�;�i��B��8$��2:��)�i
mʂ]���	f���&�}�~��q�b��?	��췶G��y��p�
�N��S�T}> �Ds�"'��uOD1@>UC��@<�}9>��f��le�&�g1�r���[���v�v{�NUմOEz�a5�
4q%P�ː� A�G�O�|sp���|2�����t �.�p
J;V9ֻn�Q1 n��J�c��n�91��-�mM��o,�ح�a�Xȩ�&�lt�jOG97�M�wmØ.�94��S�8cN���t5Wzc9D5<�r��* �Q?��T��;�}�9R�r��q�#tH��]kҺ8jX�0�On#��7\�7��t�`^K������ܱ���!�׻��bX�'�~���yı,K����Ȗ%�b_;�w��Kİ}�{59ı,K���ܙM�����O"X�%�}�wq9�H�L�b_{����%�bX?wMND�,KϾ�ȟ�C�q6%�gO��ffLͅ)�ww�,KĿ~���O"X�%���٩Ȗ?���;�xq<�bX�%����r%�bX����L��	�vaL���'�,K������Kı>���q<�bX�%�����K��E�3����O"X�%��������.e�n\٩Ȗ%�b}����yı,?�#�^��O"X�%�}�����%�bX>�����bX�%�������զuu�ؤUd,-�5ؘ燋nE��b�j�s	��:��]F�%i��%�bX�߻��,Kľw��Ȗ%�`���jr%�bX�}�|8�D�,K����ݸ��L����,Kľ}�w��? !� OȂ�)_"y����MND�,K��߼8�D�,K��wbr'�TȖ'����r;.f�.nn�<�bX����S�,K��߻���%�bX�߻��,Kľ{�w��Kİl��陵͛���-��59ĳ�� ���|q<�bX�%���؜�bX�%�߻�O"X�%���٩Ȗ%�b_O~���l͐��Sni��%�bX�߻��,Kľ{��Ȗ%�`���jr%�bX���|8�D��oq�ߟ���@.�\���#���jwV���j���%'���g�9�Ee{m���6fn��Kı/�����%�bX>�����bX�'����Y�L�bX���݉Ȗ%�b~������0�t�!�����%�bX>�����bX�'���'�,Kľ��؜�bX�%���x�D�,K��ۙ�ni�\�sswLND�,K�~�Ȗ%�b^��؜�c@>Z�C�1�2\�X �D�Q��
c� ��,K����<�bX�'���br%�b#�晴�ʐ��ۃRJ���ԏ��W�V�����۱9ı,K�����Kı;>�ND�,K�~�Ȗ%�b{����ۆ�&]ܒ����,Kľ{�w��Kİ�D?�xbyı,O���'�,KĽ���9ı,O�ӽ�wsv�.��p���<T��d �W�yhwR^�#T�.u�.ٿ��^K�e܎˘]�	77|ObX�%��w�ND�,K�~�Ȗ%�b^��؜�bX�%���x�oq����o����=]-B)\���bX�'���'���L�b_����,Kľ����<�bX�'~��S�,Kľ���ɔن��%6�O"X�%�{�wbr%�bX��{��y��B"~��§"X�%�������%�bX�t��ffHLͅ)�3v'"X�!"g�~��O"X�%����
��bX�'���'�,Kƪ�Q\ؙ�wv'"X�%���:f�&�7$����O"X�%�߯xT�Kİ�@B?}�ޜObX�%�w��ND�,K��{�O"X�{��;�w�ݗ��]q�� f����Zƌ���9��יc��8�P ��c%���ҧ"X�%��wÉ�Kı/~��ND�,K��{�O"X�%�߯xT�Kı<�����ͻ%33p˻�Ȗ%�b^��؜����,K�߿oȖ%�b~��§"X�%��wÉ�O�@ʙ���~��ێ�r��S3wbr%�bX�߿~�'�,K��׼*r%����>���8�D�,K���؜�bX�'���w.�v\���$���yı,N�{§"X�%��wÉ�Kı/~��ND�,K��{�O"X�%�g�gLͮ鹛�r��ҧ"X�%��wÉ�Kİ�#���v'�,Kľ����<�bX�'�����Kı7������������y�������<?vyy{f]k���n�v����1�";<4��:��(p��έ�#��z����C���u���We�0�.��gţ[UWGF�7
��;+4��8l%�\�GCaq{q��Z�۶5��1J���nrʲn�\�F���˫��v^eQm�3[Dn�CYSY0�E�oHA;8ѧ�Ã'-�帺a0I�.fe�w(f�0̈́�EG�$�5�F�7Hו�vj���̡Ѹ���ݬ��n�w;��39-�^�C���w�,KĽ��؜�bX�%���x�D�,K���br%�bX���|8�D�,K�O�ve�$�6R�37br%�bX��{��y��Dk�6%����'"X�%������yı,K��݉Ȗ%�bw�{�37L�r��&fn�Ȗ%�b{>��ND�,K�~�Ȗ%�b_~��ND�,K����'�,K�����0�4�.Kv�͚��bX�'���'�,Kľ��؜�bX�%�߻�O"X��� ��=�����Kı>�����͛�Jfn�swN'�,Kľ��؜�bX�%�߻�O"X�%���٩Ȗ%�by����yı,Op�N���yluըy����Ş�{�S���Sƹ�a�n�Oa�:Y��vfvV���{�Kľ{�w��Kİ}�{59ı,O=��O"X�%�}���9ı,N���ܻ��s7p�ww��Kİ}�{59
�/�A�D��E5Ȝ�bw���8�D�,K����ND�,K����'�,K��1�7����#������#�G���|8�D�,K��wbr%�bX��~��<�bX��of�"X�%�}=�:fCf�n˚q<�bY�`dL���br%�bX�����<�bX��of�"X�%���wÉ�Kı,���f\�Jn�Sff�ND�,K����'�,K����19ı,O>��O"X�%�{�wbr%�bY���������ja�����k:���^��nsp'�w5�&N�6�7+sW;Q�l�n�Ȗ%�bv}���bX�'���'�,KĽ���? �<��,K������%�bX���[����$�m���19ı,O=��O"X�%�{�wbr%�bX��~��<�bX�'g��Ȗ%�by��K�͛�Jfnᙻ�Ȗ%�b^��؜�bX�%���x�D���Q==��t@3�"yg��Ȗ%�b}�{���%�bX�ߩ����6i3sL33wbr%�g�T dL��߷��Kı?N��Ȗ%�b{����yı,K߻��,K���/�˹�3f	77x�D�,K�����Kı=���q<�bX�%��݉Ȗ%�b_;�w��Kı=��˙�͛�ܴ�z�M�l�`;]#��p�ͧ�Q/7TM.<u����w{����,s�$©\����bX�'~��'�,KĽ���9ı,K�~��<�bX�'g��Ȗ%�b_�~Ι�a��&��Ӊ�Kı/~��ND�,K�߻�O"X�%���xbr%�bX�{�|8�D�,KΟ^�˒��Jd�݉Ȗ%�b_;�w��Kı;>�ND���2&D������%�bX��n��Kı;�Ι��I�f�3ww��Kı;>�ND�,K�~�Ȗ%�b^��؜�bX'QZ*:!$M�~��<�bX�'��9���If]���59ı,O���O"X�%�}���9ı,K�~��<�bX��of�"X�%��>����9�s2�ԕU(7�M.���RG:vE�c���\�� ������r�֋c��37t�>�bX�%���؜�bX�%�wx�D�,K߷�S�,K��߻���%�bX��ӹ���l�f�ff���Kı/�����%�bX>�����bX�'���'�,Kľ��؜���TȖ'{��컑�p��ܓ7w��Kİ~�����bX�'���'�,�Q�Dȗ��݉Ȗ%�b_w��<�bX��}�36�v�͹��t��Kı>���q<�bX�%��݉Ȗ%�b_;�w��Kİ}�{59ı,K����2l0�dܴۚq<�bX�%�����Kı/�����%�bX>����bX�'���'�,KĨt�(���n��n�t璸x�e闭�u*�q�{f��T�r>�.3VE�HF�:p�o?�w�o�Cr:D��l5���m����j2f8լc��f��\w-k=���t>wJs�`��![`��v�t�'��6�G-Htsr���Ipࡸ�z��lp���ĺ94��cb�v3�I�rpZ��Mlp��x��hWs� 75��g1�����7!�����˲O<�Hu�f)\�\N�x�R��JS���c��+�\]ι+#�f�q�Z����,K�����<�bX��w���bX�'�}�'�,Kľ��؜�bX�'}7��7t�7lܒfnn�<�bX��w�����$r&D�;����yı,K�n��Kı/��w��O�W*dK���g0�4�,�72��r%�bX�w��8�D�,K��wbr%�bX�ϻ��yı,~�59ı,O{;�0�fݒ����n�Ȗ%��*�2&}�۱9ı,K��߷��Kİ}����K���$ș����<�bX�%��~����f�74�37v'"X�%�|�{�O"X�%������O"X�%�{���'�,Kľ��؜�bX�$C����iuS�7ny��n�w��%�!�y��3���u�s�Z�d��6xv�h@�^u�@�*��S@��_`�Nı,K�{��yı,_�ދ�IP���}����oq����}��qD�
�Ǒ9ļ���9ı,K�~��<�bX��w��"~*dK��s��M��\���O"X�%�~��؜�bX�%���<�bX��w��"X�%�~���Ȗ%�bY���̸Bf�Jl�݉Ȗ%�b_;��Ȗ%�`��xjr%�bX����<�bX�%�����Kı;�Ι��I�f�3sw��Kİ}��59ı,?!�{�x�ı,K��۱9ı,K�{��yı,N���S	��7&��5ݙ�ٸs�R]������y��7na"{vᣅ��`g���̳s.�Ȗ%�b_�����%�bX�߻��,Kľw��'�,K������Kı=��L�͛vK�7u���'�,Kľ��؜�bX�%���<�bX��w��"X�%�~���ȟ�*dK��?f�na�I��a����,Kľ���x�D�,K߻�S�,}�7�88��=�	$ �� ��D�B�|	露�Z$F��i�苄A"Ƹ)��(,B�F n�LP�G�b,@ ԉH2TzʱBK�b�H�`�b��M��K�*��y�Èqb�V��:�H�"�#B����!äc FHB���e��$�ЄHx��Z$�qI	jp�b���HHbE!	GLX�a��YR0�%�!��
$��ŀ���@ۂ�"��h>%DX ����� ���V��o���>�@OaȞD����Ȗ%�b_~��ND�,K﴿w.�v\3f$����%�g����xjr%�bX�����yı,K��݉Ȗ%�b_;��Ȗ%�`�����{PL)������oq�����<�bX��G>��؞D�,iR��W
���۫ ��n�#��\Fh�vu��z�C��h�r-�c=��؜D�/\��Jq�n/�J�n�#��9��`��`s��_�� 7w��=���i�C.a��R`���W�IS �˼��/�9���g�a6�$����	~�x�$�0l��zژӜ��NS4A�%X��V��� ����:�� �} ��?���U!(��1�9{��z{��\"���'$� �se����f�x
��R]���א��q�P�l%����搮�kV{a��"7;͢����b�:�r�/Z���+W�m����0=��`zJ�{eL;���]?A:�P�)%����_�;�� �o��s3e�r��qS�D)�$��W��*`���W�	�gnw�3�Շ8�#�c �ʘ���합�_5�����}�y��Pꃋ��z� ��0=��`zJ�{eLf
!�,A?}'���34��1s�C�̖�j���*s�ĳ�͌�\nm�8}��<6�G�,��������P� ��vm�z��]�vx�F0����u��ss�N˹��3ۤ���v9ķ5M�n��O�I<!f��`#��N����LM�!����\p�>��v:%���V�B�n�]W�s�6��Q�;
�]�.t��G�u��#o&Rzt�صЌ�>���}.;]l�q�����c4i�D$�;\�tK㬳Lz)j�1�M�]v.&�m�n�$������`�S ��03tKm�N2�n�6���uҒ��Xw},w6��更�\"���Xu%��*`����9������;���q��`ےX36X�mՁ�ͺ��Iw7����[�*�t���C�&�W�I^0l��zf� �v��n'�4�D�R�Z�6l#u�]Z�q��Ggm��d8g;n���<�;���0=%x�=���*`{e��1̓d)ӔFۂ���͗�4��x��m(I-IU�^��6T��ͺ��b�4��*U�fj`{ex���� �ʘs��:���t�9ޤ��+����T�9�����-�I8�)� ے�fm�Z�^lx�6$U� T���;CTڝ\�b�Q#YW]m��c�-�Q.6�j��[�b2��h��٫��ol��zJ��^0=%x�6s'j�n�(q�tےX36X�mՁ�ͺ�w6_�H��[�*�tF���,
��R뼉<�~LM$�&$�'�_U�v>�� ��� �bͦ��ԌR��0IS �ʘ�������6B�'ѱ8�������}��K��N����;����}�U���'W.�с6fQ붩5z�8u�<�'�q�5ӆ��e:�JQ�4��*U�f�=�Q�l�0l��7;{s�.���C��R`{b� �*`�S �n�7D��&�(C�ۅ�w3e�{eL�����F���q�qcr|9%�s���9����ri`��è5��s�o$��i�˝0٤��N�rK �n����}��@7��,�͖f�(��ԑ"'L���*^z���_<�F�GV�cn+l�ق�#�I����9ܚXs6X;�?}\@w}�`�[�j/�H� �#��w3S �ʘ�����G���_�ވ��I(���;��`����UU%����37����Ǭi�*crX�T���F�0�9͗���;��9#))�6ܖ;�K���N U�Āz�"@����i��!s��]�w֍��{�'�m��m�^q-�6�d�sǮ�t�pOk�)g�0	���m\�"�շ	jy��]�iQ��X�E[�I�h�us���_mD����ݴkb'�FP���hy�ۃV��R`�l��j�Eݘ�m����n8+OkpF�v��ֻy��Z^,A�v�g�u-��y{z�����^����]��s��.�g�����x�ϣi*耟��8sI��ۆٛ�L�L��Z�ݣ���C:K%������m`����g�I���@m8`�,�͖�͟ϫ�;���7��]H@M�'Ñ0l��zJ�ب�=%O�9��54�N�ĥ�%�ww���rig�6�8VfĀU�ā���Α�(�Qs��`{ex�=%L�*`�� �bͦ��ԌNRh��͖���N w}�`s��Vhd4n!|���zY�q��/]ѵ]��M�`4>h�	9ݸ�(����NP�b��`�l�fdH��_4�� �͉�]��N��e.L��I'�w��)�CҜS��� ��0l������ԗ@\�$�rX�M,��,����K ������۔����Ҁ�p��l�l��zZ�ب��K��<HAΝ�_��`�S ��0=�Q�l��m�;��v����N���8՘l�I�w"�˫��z3�uӬ=�5������[us���&�*`{b� ��0nl�7]-�FUD胤�I,w&��*`�S ��0'79�s�\��Iӝ��@=w� �Ȓ���i�jK�������i W
��� ]�	%�rX;�,��,w&���.��X�O_�Ӡ�*LnK �f��W��T�=���_�/0�SU���`�.Zά�y��^.�nR�'Y�p���iw6��~��:��A��M9' �o�0IS �ʘ�T���k9ެt$�@mIV�����UW�RA��K �o�����X�v���	���rF�0l��~�6_�0���!M��Pt8ԡ�$�����_��o=����ߥH��$%&��$�֤�j9y�,��22�6EN�$�9�۫ �f� �se�s3e�ո�kS�%���4R����q;��7W8U��uD���묉JJJJj/�IDbh�U�s3e�z�"@=w�����%]��T��3~���d��b��`�l��_RA��K����fl�7�����IPT��L������l�0l��7;^Ӓ2�8:I����Ի��U�f鹿s����]�zX��RnS�'J{ȅ w� N��}�͊ ������$��**+��**+��E��**+�آ���ʊ*+� ����AQQ_� Q��U# D� D�B $TB
�B
�B(	@"�(��**+��**+� ����**+TQQ_TW��QQ_�EE���TTW�AQQ_�QEE}QEE�1AY&SYu��,�ـhP��3'� an/� =                       � (	EA@T���@T�����ER(H�Q
� �"�) ���@�H
 U(H�U R�U        2  � %(� )A@ 4(f(�(�R��D�AD (�� PQ�  �b%ܟJ� �}��}9��s^{+�'J� ��+�w|��y���K���� �    
 2 �}7��㺥�3W[�w{i�� �r�e�']7�ί��g�� }>�>�9�7׽�� [�6]5ɝ���(t|�>���Ӿ;��\����X ӕrz�95֜���>�J� �    
S �W�nT�֜�{ۼ� �ʕ�z����NZ�bԫ� w��x����� ��oky��5+� �K���{�W����ꏾ� <L���ɯ&soM�{�W�<PP( (  "@hi�T�NvUw�畷���;�� ݥ��Ο}����m���r����ܯg7|: �P   D  {�� �٫�mr��rv���﻾��}��� {ҙ�﬷���ݼM=�3J����@   ����׹�nn�-\��=_[���� 3J�m��o{��4�����+�}�O��S�iw�� ��)J��>�H �JQ �@ "R��@ �PQ�JGf�;4���R�� i�
��J�Bz���*�i�o*�I � "x�T�~� d ��T�i%T�F�"����{ڕJT @D��JP��1M�	�]�?����E�����Z��;j�o��(�Q\O�����DO�AEE�EE��"#�H"**�W�?�`�[	g��Jr0�!HزH�FY[a
ڔ�L��	��� De2� R��F0���y7��LJ�R%��v8�D� 6L�H\�l���2��N;� �H�R��V%���1�ɉ����C>����4�<�9�ᴍH���!�Ms�'ٯ�W��B2���.�@)�� T�"D#H�!��}
\ւ$Xԍ l���@�����	t�!�Y�ޯ�3$�	�Ϸ�C�X�=�"�)"�d�
:`�602���.��In�S7�����a�s��횯l~o�u.kY�l����f�C�湼�	Y�[��C$�Bo��+~!��!X\�!Rܩ)�}�h�Ċq��GP�2�P���2li.��hbS$bQ�m�jMR�0�@���6�&�Ġ`h���L����RE��P�m�
2.D�<��A!fR�20�Lѳp(b�i�0�1,$)D�d�	$��%!&oz��.�ng&|��.v��s|�ړP�,IF�:� 5����3gye1	�a� C#�� `�!,P�c�j_���Ou.���kz��-h[�|D�¤�p�4}�!aq!�˭Ḓ�))���%ѩ�s[`R<0�1��6K&��e܆0u϶rL����?@�|S�1��e��m�$�e�h�Y���Ri�!�_}.�f���8,i���7��1�B D����Ұ��$��abG"�+
�K-e̺��<�H�	�K�S�g�7�r�>�'n�&d�r�7�$Jf�W���)��f�sZ�9�W��D�R1�!"�"��.h M/&��0K�B��@��$c0!�u�5��vw]�h�|�^l�ӟt���wl�
�w
p8K�kWE7&��	�35񼁳�.C�ى-u	�~��e��2�D@!�(��Sh`ei�.�"�t]K�#��7�㽐j`iٽ퓝��B�(D��I��J԰�L�T.���N/ɶ)����{3vs����ѶP��kK	@�c@�eR�h����4�
Y�&ef�;"B�S,Bn$�af�IF&k[,�)
J��*F�涱����`HY4�$�J��������h�#��[�Hz�0�HP!^0�i�Q�$!J��d�JE�)
I(S5�i�m�|#� ���`���Q�nf�),*%@�C����4��Q�[�"E���G��ށ�1cN#�� T @��"�GI�N:�)����{��
BiYX54�!z�].���R\���uo{�.��	^F��W#w��a�!����\�}�׉�P��`�
��)
4�T��*B����`5�
�];	�%Bo�Zhfk\	B61#BV$)��9��N�cC
�����7�ݔ��ϴ�asA.�|Fr��o����g�y�sLr�j�W)���3]0����ϴL��3뤚av�CG&�ۼ��8�i�r4��4��%ς\@��2I��3C��5�K6��+)�P�M���㤃!���04��i�A�#��)�a��f�M�h���L��g�a�H�0�V��I�kƘhވ�Ʉ�,ɬ`��ѣ|8�f�����%�S8�(d��w4�֍�XPqҐ�sa s���A�A���Q�k.�;�晌�t���;�}5�t�4!jF�\Y@�0�LВ0��K R�F"�X$�h���F �0��ar��]FL��_k�\�ϳ[	sCy����+��L1!p!LLX\��h�ٮM��4K�t\���ލ˚v�����ִ&�$����m���	��z�SwM��:+w��l8ic82��l�;��A���ݺ%1Ӵ�qѰ�.kG���@w��� q \6N<a\Jm.���y�}K�+L�8Hԗ8��X^as|��7���!�:X�@�o�SL���3{���p7�`:ٽ��h$75���o�D�B�h� q�����������;�>�N�����t������$S��
+� ���ΐ o��C�!t��e�4�0�φF�	��㌸hCg3_f��i�5�Jd�̝z¬Hc
�0J�6 $Q�Lk�!��ĸ�gA.�߉��?p9)+s�$�˜���%�
��MB�(K
`�+�jf�@+��Ѝu��+,((@�i)��Wa�p�#P�4�o��(d��B���34�]O��sDB��!!La\!	\!"�4X�40bP�T�\�,W4��I`\H1��4�#xB�)
��i��h�l`�)r���qLH\�l����a
��)�hF�$��k{��q0H�!HYr�pٚ#�Jm��r�j\���"\9��`��L��
�F�¸M�Ö},�3\�Y�L�K���9{m6����75���o�F���ȑ�����H��l�o��$>�`B������Jd0˚%���"F5������B�D�*JV�j@pѦ!R72�%!�RFG%��*
0��1ɮnI�tK��)�ƸF�$n�/>�>�E"Q�Hk��0X��F���"�Hh6mdH! B�j$ѵ �Z��,�2�M'С ����$��@)&��%7��@�"Q��@�� a C"H���CG�u�Jᡜ܉�K�u�����ٛ5B��RkI$�n1�p!��5�8�t�B0�B�����Ȓ��C�����]0��du��h��� 1a
0�
1��-LJ$D(�Ssw��u��
������1��
@:�,P�C ����"&B#4X`�
��`�F�!;R��H�%�@��h��#sF�8�F�H�E�-�p�@�ѱ�I"GD�dH�i�$�<��K�$bi��jb�H�T���E �;I��Ѹ�WB�.ǚ��\��5-�%�	.HV��i@��[�pồ}�x��Q��1��t@!��Ր�K�``��4�
H��7\]e�@(lL`�a�!@���IR0�0"F�h�� ��&��,�i"c6B���n)
a�u��BEh|�(0j�J��G+
�B�¬*J`@i��|��� �A��A���ֵ�`L�����n�Mf���I���2kSbB�.K�k焦���������j&�"nݺ6C[%���Е�Ih��
B[������f�Y��a
�RĐ�Ir�`Z,�SF�hkG�|�9��YJ`h�7�u�̎<5ee	njS!�Y�X�G~߽�F�.��9y߽��|�Y��j >X����i�R�4C|/O�HQ"�����!�5-��j3
cB&�i��Y5Ǭi��k���Ax@��RDc�f�e�H�FI���M��BkN�{��ȮűB'�X�	�`���@�y�#n�g$�FB\%�B^���P��[��#Y��aHf0&`^]l�N��q�8��8 �ͬ�5~��~ޤ
�JSGČ�(�kr%���WC�0�]�ݐ��6K��u��5���K)���8&�6L��5$	��1�ӵ�@�MXF;���$�դѠp�h8i�#\$F,X�v�K��g]�;��!L�BK�B@�,I&<)
e)0��Rh�6p��Z��@�;x�̓Nٓ)	\v��K�Ք�6p�p ���C��{��`�n�6��B"���',��%2%�l8���@1�0�	���(B�֛�cMB4�4A�@���qZ�4a�Zr�MB�"JR��B0�dh`ha�r!
b6t�b�0$7�&��w}��n���7~���~��  6�      �    m���  $     ݅H�i&��l-�"@�Ô٥*���NU�V�� �Mm���v�Y-I�q�ۧ(۫v�WX�4�@&��m�k�L���r����S���UeSq�źk��o�Y����I���}Ač�9�	 �m�6�&�� H �I-�Ԏ݀�l�ֹ��   �m�� �j� Zn�o8���[D�J sm���[V�H[@	��rI��6۶�[@�  �6�;Z���n��` l '[KK<�VU�⫗n��i6���Sd��F�`��4��vpH $ݶ,Ӵm�  	m�� H$d�   [@   5�  ?�>m�  � ā����Hj��T	31C����ݷJ����m�Z���F����5�[��'6�Xz�|�ۻ`�Y�U���)�ڪݸ#n���]��D�m9Jw��z$X{�|[v�`����BU�U�����V����n�o$��``�6��,�0|7�lajܥ:� ���i �I�il�� 9�림m���5t��d���#e�X�ݹV�:����棭�eZl�[C���l[�m���6��l�n��v�H�	$ ��bۉ��"ޥT�LIMd����7N��:9mڶhݧFضCe� m� y5IBE��� r�z��a����[r��9���j�C�pUUmP �U�.�*��뀥%�E�]طX���  �d���i�m� [zM�nU@m[QơwB��*�р-��	9� ��*�UmmR���
:͠�ہ����[*���I5�l޻�� �HE�ZN�8ְ6���h�7Eogen�hk�6X(mD˚�|�|8-�����@��y�č�� �m��ε�J���mHkR`�l�K�����Ҷm��!j�0�KU[A�.�m+R�5J�UP/l-��p��h6�T9jR�ت���9U��������$I��a�&� �� ��j������6�m�*m,�i/n����uە�iy�Q�u,p�����ݩڬ�@U�HI���m&��˵��rJ�Nؼ7�6�mr��6�-�����RJsj��;*�,�:`+���BQF�V�5v�Qej�;0ԯ U_�ϏZ�V��'m����N���j�하N�z��*]E��=z�d{5..���t�$u\��(�m7[%G��NN�L��,K�/&2�*֤�C;����( 6��S�u2Kz��tJpCV6�]��)(S+Q���l�$m��]X'&�J\]���n�p�U[@��2v�tna����El؟6ƦRP*��K�E.���5�`	8 6�m��h� �V��"]� ��ӌ:ޠǆ�j	m��� 8r�v��L  ඃm�   ���$�f�vݶ��p   �m�G��-��}�4��8  ��d��c$O��k�V $s��۫ku��Ā  �}zɶMs�C�mB�u�HM�@Am���V�A�	7&6�8pA��kh    i�s�5��U��   l�Y�z�� ��6���ol�*�+.�청t�U�Ԫj@IӡԒ� i��   �m�M��d�9#���p�j�@	�ݶݺ�We����u�_*tR�R��m�@�*��j���s!*��=+r� i0��`�z�m����u�Cm� p6�`��ZbCm�[k��m� m[�T:,�ݡ\�TRօ�m�Xe��e�oY�`�m��:N���.�K������YIT�yqS��@�
�uҬ���l���kd�8[\m�D�T	@�u�)� �B@�'dք^��� p�PRݕ�ZU����vZr�Z�g���v����qm�-�6��k���c�.�8 	�D��I%6� ��U�.��!]�V��������l� ��  ��  �� m �k�q7j۝�� �fۦ�ٿ���o��f�W4n��*U�VRZ��@k���ml��t�l��K*G�I�Yd�`� ��d���  
��码j��G���@�֥�ZBj�)��N�lm�t��e$t��J�R�J��-�u�4�)E ���ϟ -�����VV�WhZ�V�- �|[C��յ�؝������n���A�UU!Kұ�vڸ
U���F����UT;��:����S���m�B��iSi�@�Ivm�2�,0��[80K:����jV���d9��
R݆ܶ�F�M��v2���v��vS��azED������-�MF`ݍ��S�k���d�t�,��+��M 9m<.��(rtM��-�H/�  pqͷ`tm:Vu�������SU  �d���B�qoSm��8��>�߾���޷�n��/6��@I�I��[@   �� �k�>��PUJJ��e.��n�]	n8 $7Z�kV�m���7m��)m&�YKG ��z�oPVĜ��ݯV  �KZh�M���ݰLݭ̀A/Yl�Crޕ��� �g5��!�Nl�+��/(�&��
�ѵU[*��Ͷ�`�3M��m�ձ�FaĀ�k�U�w	�"k���ϖ$ j]nkM���$9���& 6ۤ��M&��@�k�6�6�hr�UWvZ�V����[V��m�f	���m� l �`i3m��� �vL�����_��]6�m�͎Kʫ+�WYc���������ڭ�L�Kkf�7RWm��+(�c^��d�sslm�e�gj���p��yc�)W��������7��@ -ɱ�l2;�v�l�`` �  �G.�å�w�`�d�VZ��l�Ӵ�lI"GXc�V��pI��p�lG9�$�d��H���KU��5H^�y��	ͫ���m�K.� �p[@�nH$�t��@0mR�N"�Y��۲�UPUW*�l�H.��9�A�@�I$�Vێ@��� �ZW:��e�q"i�+m&�������86�`��l����m��a۠�暪�V���R� $�ji{N�[wUU���\*�v�#�jm�؀ݶp$�T�v���U��� �UV���[���P �$�I�m��m[z��6݀	�-�-���;l 6ε���[u�F۳��>  Xp�O:z̫����*��`��Pk�m<AZ���zc�Wv�x(�6(8�jej�"��t�V��\��|�.�pԄ<�, 'cby��]�i��l26�ndS�#Kl�ݳ$�	 ŷm�l*m�gD�-���mZ�m �&�K�z�n6ݜ��7j�a�m�m]*�m�����UZ�r�T�e�[-�$����2����{vZ�j�^�[E�M��ҷ ��Ŵ �i.m�dI��&���WK��꫕�� *�[PP[4!r�٭�l�� $�@-�hp � �m� Kn�mE����Ŝ�`m�@  ��	��q��R�p��Zm�v�   8VVN
��$�V���`  �lA!"Y@ ,��jZ 8��!����ͨ  �ݹ�[���	 jm[i�B�m��Ѻ�Hl�[��������  ��p mU�(� H��W���֦��ۅ�'N�i�a��"�n�UU͕jU�i��la�8�6ش�so����Z�Y������n�%��� �H�m  �Cd�Zf�YYT
����g0 i�[l�.�U�A� G]�6� I�[~����6��"�k� 4ukRf�I3���D� ��[��R�Rҭ`��@����z�t[��Vv� ���� ��d -6�s��e�O�rϖ�-�ɇR��� ,�Q�/5U�.��m6a� �-�8sv�+`�olp�v�z�ZWg��Y6��ktIV�o��@J��++UUJ��Ү͖�km�
� [S�.U��	Tb�v *��` ��M��[���E��l  �pkR]6��on89���@m�� ���8���|9 $m���Q��7����k�[d-�p�i�H�e� p  -�m�z�YKr�i�` ݪ٣t̴��5�Hc j%gd.�    ���<qͶ [V�m��%�@U*��KU!5=j�ˮՍ�Xf� m�ut��`�]m���T�;5@C���d��N&U� n�L[vnD� H5�v�&i  r@HI  $nݱ�5e��H-֦G�v�݅�����R@ֱ%�V��kޖl5�J�f������e��I:�p[Ko��` ��Ԙ   �� H �٩u�5%���Me�5�dP4/�"/��
/�⢸����b'�*�UQ������&iA6�qD�l����(@�G�V*���P6��E (h�W���Q6�E|"�@�4v	M(�$PL@<T��8#Q:"� �P/O<t|��@:��(��B�¾A�TC�=A����uP:*qQ��z0Q�T �_�G��C`���/�S�)�|(��_�]���
D����,|"���a$DX�BYBE���HH�"B @�@�IŁ �f�^(�p>_"D@誘��)�`��~
���u��� g(Q4(�@�tP���A��GE�!�!$�v"�x���=AO"&�EҕT���8�S���� �A�/�W�S�OlبhC@��ES��v�!Dʠ�
 �� � �@O��h��� UC��P�EEx �
3��g���5�hm�i p �esb]-��.���qrK^�$l4�=]�1�Ε��!��6�;Wj]S�0
�����\��,���AWUU�,��`�����N;Y�.�^͜h%]��lJ��<�e�Ϙ�0b�v��;3�8�8�Mq�v���m��1�zԸ��O`�<��Z4p[J��GaS�B�n�z<8�Z<��]M�Ы�glLLm7U���ܷ*����zXD�Bzbٮ��;��x�l�R�'l�-�:�x���;l0p��j9ۗn�d�����jK��c1��𕋈�c���:�'n��!�#���g�R�� 
�v؃�U;9	�{���[Þ�&��ƥV�-jP�\��m�Z�ܘ��ٹ$��xѥ̵�t�&vAV`:�p+��wh���\N�����8P-:��m���Γ��^v7��u=d�3i����#�uFժt��晤��l�J� ���k�)��Ȇ9с�Y7aۙ�;.�<9Q�a0R����գn+S����Q�;D�+�<r<j�E�؄�^���4��$Ӣ� �䕪	V5�v�j:�Z�m�0�C�1΄�I��b��.�Y����ӷ���%��!�#J�5i��a���z���q�5��a�bev�E����@��ݺ�����d=�ܓ�c�h,��V,��:�+�m�[���bm����.��s)��]�r��y���m�kT����,� ���C�Z���zm<�N�������g�B����6�`�8��:4��\�nͭ=�`
���)���ٺ|��6 m���pl�k��"ۥ@��n@0��6PaAƭn��e��j΢8�3B��LV��㊺��"w���tnav8�����v�ځ$�\��t�p=����]��֨+dSS�a�e�T;-@Rqh�Ut	�:��!4�0�l��P.�ʠ+�`��*� ��N۩�'<�!��G`S!�Ф���U�>���{�{�{��;�ܒ+ �?�pQ���U?ؠ? �����@����ή{f��X^��4����Q�1�m�*ݺn^���rn�&��D=�u��l�ع��%��܎�n����4���WA�^V����@r���8�pg��y��ԻSg��κ�����z��T���Я.���Ѯ�|֒ޞh7Ju��XM���e.����;v�j��O:+v�w]�����v�������x�vD���ݗ�`����a��\<�v6P��r�2RfZYs:G5���>��h�H$��~�pI��n�����2%�b{��siȖ%�`���.nasZ�ˬ�&f���bX�'}�p�r�Z%r%�`�?~�Mı,K߽��ND�,K��l���%�b{��2�5�K�WF�nh�r%�bX?g�t��bX�'}�siȖ%�bw�͑7ı,N����Kı;'��&���4]f�Z�Mı,K�ﹴ�Kı;�fț�bX�'}�p�r%�`AX?g�t��bX�'>׽��h�ֵn��5.kiȖ%�bw�͑7ı,N����Kİ~�z�7ı,N���ӑ,K��x�h�Ս\�ʜ�bE�w���'.x�d�N�\q�5��:�M��Mr�x�����bX�'}�p�r%�bX?g�t��bX�'}�siȖ%�bw�͑7ı,Jw��s���S���]kFӑ,K��=��66+�*i�*��H�1@� �)�D�K�﹛ND�,K��l���%�bw���"X�%��^���f��h���.kWI��%�bw=�fӑ,K��}�"n%��"{��p�r%�bX=�߮�q,K��}�=��MMk35�s5�ND�,K��l���%�bw���"X�%�����q,K��{�ͧ"X�%���˛�\�Զ�4M\�q,K���ND�,K
�@����q,K��{�ͧ"X�%��{6D�Kı?�{�,�ݣ=�=���ɝ�I�=� 6� sjb�*ɇ���v��iU���y���%�`�?~�Mı,K���6��bX�'}��q,K���Noq��������F���&h��"X�%���}�ND�,K��l���%�bw���"X�%�����s�{�����{�����\�Vl3�9ı,N�ٲ&�X�%��w�6��c ]�
&�B,�`�=��Kı>ϻ��r%�bX���.{f�\2���h���%�bw���"X�%�ٞ���Kı;��iȖ%�bw�͑7ı,Jw������Y*�����oq�ߙ����Kı;��iȖ%�bw�͑7ı,N����Kı?
>�߿��~Y�.Xš����lvwi�/`�:3�c�l��ǃ���,����\��J�\ֵ.]k19ı,Og�~ͧ"X�%��{6D�Kı;���ӑ,K��_{17ı,N��3٫�5�V�k%��m9ı,N��ԉ��%�bw���"X�%�ܾ�bn%�bX��wٴ�Kİ}�ss���˭��H��bX�'}�p�r%�bX���f&�X�%���}�ND�,K���"n%�bX��}̹���p�ѫ�[�6��bX�'r�ى��%�bw=�fӑ,K�ｽH��bX��O�D�� �"�huD|�;���ND��7�����F���(�}�7�����{�ͧ"X�%��{z�7ı,N����Kı;���Mı�7���w�}��N��\E��$g�����kq����u�q�VW���k����֭˭LԹ��r%�bX����q,K���ND�,K�}������L�bX�����ND�,K���^���IQ��|��{��7���}�iȖ%�bw/����bX�'s��m9��TȞ׷��72�D̩�}�/��橆]]k3Y�i��2&eL��}�kI���2&eN���m>��D̩�=�oYjn&eL��S��6�}^w�Os��~r���Z�	U{�2�J,�;�wٴ��2�D���e����2&eN����}�L��S"f_{Z�n&eL��S���{5p���\��.�Y���2�D���e����2&e?(}�ߺm;ڙ2�D̿�kZM�̩�3*w^�i��2&eL�DX1(-�� �b�B(�P7�L�3V��mԸI�&�9��٩�ېؖ1Ί]�v�v�\�K5sӍ�?��o�ó�#vl��ձ��.�ݮ�]k	<����aJ�*V��h�v���֘��b�(s&��\s�vk�t�n�vx��qCɍmr:�Q�1�j�5�0���{j�i�&݃m���cph��u>U=H��-mh��s����M�$�۷�6�v�	��.����lAŮ4�f��jN:�jC�5�t�q��l=��gv[���,�b�N�̩�3*w�����2�D̾����Lʙ2�u��6�Z�2�D���e����2&eOw��.a�j\5tj�捧�Tș�2&e���&���Z����=����O���3*dO���e����2&eN����}�L��S#ߛ}� ��ӵ�U����{��r�u��6�}S"fTȞ׷��72�D̩�w�O���3*dL��kZM�S��r���������D��g�����3*dOk��Z���S"fT��Tș�2&e���&�fT�Be��{�ͧ�Tș�2%��˞�Y���f[��Sq3*dLʝ�}���2�D̾����Lʙ2�u��6�}S"fTȞ׷��72�D̩�MS�7�1���dY���_�@���6�t%�8��=��]�����y+��<�Kf�'{S"fTș���kI���2&eN���m>��D̩�=�oYjn&eL��S��6�}S"fTș��f{2��k��%U����{��S��}�������J�D�"�ڪ}�Tȟ���-M�̩�3*{�|m>��D̩�3/��i7�d��3*w_t�f�۪9Lݦ~{�����r��{��~H&�fTș�;���i��2&eL��}�kI���2&eN���m>��D̩���}�~X1\�!����{���֪{��t�}�L��S"f_ߵ�&�fTș�;�wٴ��2�D���e���S��r����Ͽ�/M�����=�}S"fTș��ִ���S"fS����~ͧ~��3*dO���e����2&eN����}�L��S"vkFd~��f��6�L#��6��;�-[����v,�X���ip�sm=;\QU�&�fTș�;�wٴ��2�D��=���Lʙ2�}�|m>��D̩�3/}�i72�D̩ϻ�e�h�ֵ�.��V�i��2&eL���{Y��~U�U52��{����dLʙ2�����Lʙ2�u��6�}S"fT��>�#��T�/���)�w�2�}�|m>��D̩�3/}�i72���Wb'�� q^��T޿}�m>��D̩�3����M�̩�3*=���'�ا�H���{�����r��&eﵭ&�fTș���6��bX�%�sک��%�bw���"X�!������J��%O����o's��m9ı,K��ک��%�bw���"X�%�{{�bn%�c��>��}"b���r�"�`x�p�;�׵���]\�\�v(�.�n��}�{�|���K�f����}ı,K��Sq,K���ND�,K�����Kı;��iȖ%�`ߺfg�%�]Kn�F�u�T�Kı;���Ӑ��$r&D�/�����Kı=���6��bX�%�sک�����,O���ezl6+ ������{��7��>��q,K��{�ͧ"X�%�}���n%�bX��}�iȖ%�bvN�yi��Xk$�u��kX��bY�^ ��Oo��fӑ,KĿ_~�&�X�%��w�6��bXP�1"��`���  �|(�M��z�w��7���{�>���p��R%$�ND�,K�����Kı;���ӑ,Kľ���7ı,N���r%�bX��-�ۄ�Y0ֳ35�&��v �s�x[Gd�4m��0A�q����mA�������֋�fk2]f����%�bw���"X�%�}{�bn%�bX��wٴ�Kı/�}�Mı,K�����.��2��Y��ND�,K�����?"	�B����'���fӑ,KĿ_~�&�X�%��w�6��b]�7��}��е�V���{��,N���r%�bX�׾�&�X�%��w�6��bX�%�﵉��%�bw>��\��ZӘf����r%�bX�׾�&�X�%��w�6��bX�%�﵉��%�����}�Noq����~}�~���Zf�w̖%�bw���"X�%�}{�bn%�bX��wٴ�Kı/�}�Mı,K@�!��{3%![������W��[��q�-	���қ�p��N�:x��z���×I�ك�k���ظ�\�� {�A��Sc�6�s��+h���m����j��/�gy;9vT��#��[�h6ǂTm����kk]!p�uur�ɛge/5�`�N ��ݶ:��nmŜ���91�N�8���觻k-�c����V焳�3�ωwACR���w����V�.�Y3k�j�/tS� �m����j�G�GN�m/OC��x���oq�������7ı,N���r%�bX�׾�&�X�%��w�6��bX�'d���m��k�*�w��7���{���m9ı,K��kq,K���ND�,K�����M��TȆ�?����kB�@��w�{��7�Ŀ^�X��bX�'}�p�r%��C"dK����7ı,Og�~ͧ"�oq��~�#��l<���}�7�ı,N����Kı/�}�Mı,K���6��bX�%�﵉��%�bS���e�a���f�Fӑ,Kľ���7ı,?"���{�m>�bX�%�}�X��bX�'}�p���oq���������j&(Vu�a��Q�bے�n#9��1�fn�ܮ�z�@��ww�hX\5a*}�7���{����6��bX�%�﵉��%�bw���"X�%�}{�bn%�bX�Ϻg�W&��i�f����r%�bX�׾�&��1@�E���R@�	�P��j%��{�ND�,K�����Kı;��iȖ%�n����~����O����oq��m9ı,K��kq,v�"dN���r%�bX���kq,K����&�a���j\-��iȖ%�b_^�X��bX�'s��m9ı,K��kq,K���ND��oq�ߛ~}��6�d�U>��d�,N���r%�bX~Q �~���ND�,K߽��ӑ,Kľ���7ı,O������h�fC5����\�q�L��,���qV���v/nn�A���B�@������{��7��}�X��bX�'}�p�r%�bX�׾��Bn&D�,N���r%�w������~�M���O����D�;���Ӑ�G"dK����Mı,K��߳iȖ%�b_^�X��bX�%;���nke�ֳ5�6��bX�%�﵉��%�bw=�fӑ,|���A��H� P���|�)
 Uڵ# ������kh��*D�4�� `HM!K*��cJkd+��F(�+��D������jŤ�	�`J`���)�hC�,'�.#�P�$+"�XU�~Q�B!$��7�RRB!��� �2, ��D"D�b8S"0"�R"0X�b`BI!$���,B0a%���R8�qH�SL*�#*ģ�D�#1���� I! �0w@`,dbA�R# ,X0�"A����Ib@$�d(����'�` ��k��mf �(��8��J <��ȧʊhV �H�ı//�k�r&D�,O���ND�Dʙ�?O�_�X\-T��oq���{��D��{�m9ı,K����?*���,K߽��ӑ,�@�D*�}uRB���kU�d�s5v��k������Kı/�����? ș���~��K�!�2%�}�X��bX�'���f����ĳ���w{������2E�'El봿��8�*��(��P,u7��"2�mf�<��u�[��5u��'��2&D�?����ӑ,K��������Kı=���6��g�H"_�ߵ���%��D��~�fa�5p��K��4m9ı,K����7��"d/���f�ʥ�����b�~�P��I]�ٕ2���ʒ仫���BS���`�J�>��>}���D������*�V��˛����I,����ϯ9(Q2>}� �(_߽�\�j~A�B�mQ_(��������l��x��E�jU*���n���$�>���
y�t%�B�_=�W ��f`�$��H�V���,mnZ�i�`wu��V�8�۵�u]tss�XcQH�s4׬�9^�@-�4�w4ۍ؛�1�MH���`M��l���W��y�ݎ�&���8��l�:��Ҥ.�4W��9}�ۯ�bB�9j�`K+�d���eL��`}z���'�8'�'3@/u�+ֻ���x�_>���K�*�s>��.����<�[a�\&�<�[nƦ����\kZ�	�qM��p�Yk����e(6�f��>���b&6�״;:Mѹ�T�k�mګu͎ܛ��,J�JKm�F:��G�>H���q^�s׵n��g�`w<\�=R7eC:vx�0h.zx�/�G]0jb��Ѥ3���C���|t�\�1�,Ҟ���S`�vy�y��SR�D*�Ț��Ly�ap��j�[˒e���]�۷S��i���>e���m�4jj���wq�?����lv�_(� ��,СL�}x�݊���������j�9DL�ou��b�
������!K�}X:�S]Jn��UUuD���(Q2>}� 9��I$�H9�Ձ�DDL��^ 'ܫ����R�nnꮭgB�����<����������7cȚqI4W����@��s@/u�[��'$ȁ�ŝ���K�K��\�*b<&n��.xu��ڂ4y���L#q�Hs�� ����׮�[����*���*�?�bEU��U��^,���B��I%vϯ@�^���[�o�;��F��ّ8*S3V����/]a�	)������4����1�(��M����y�,����Z�%���������@-�4�w4޳@�z���vY1(��d��$rd�o�6�\ѻ�5�M`�v�h�gkc��\h���17#=5��\������[/0&�S �Y���V3��Q'&h�f�6ʘ��Y^0n+�,\#s���f�������w��I%�	�O�j*�s�}�rI��nI��c�	�n<Iq��f�׮�[�h�W�r���G�ȱ&�rU]����9(��}�sϫ �x�����2c�<&x0�)�<��V
��n-ēRB��r�YN;k�Z��t1����-��l��[/0%����mc�D��Q�&���^�[�h^��oY�}ey29����.L�y��+�l����S�N̎LOq�G&��빠�g�� ��S
�� _6��щ�I���4޳@���@��z׮�g�}��6�r%1Ǒ8�I��,<�;)�c V�(M�6����⳧kAJ��Vx�X�6�J)&���^�U���]� ���9}�݉<#Q�Hs#�.�S�W��y�7֦�LZ��%#��Ǡ}z�h�f���^�U��z�ۏ�#q'�Nf�[/0&����eLY^0$����II�Erh���^�@���nI=��[�ph�E�e�m���.�l��1�\�m�V�z/u�.D�v��vފ�
b&2�_+���-�9��2;�/m,w;1���X=�� ����)u�Aɉ�p�;-�&�9�'z�����K�;ӭ����`�	�ӱ=��������U�[>�� ���s��*c���Omu��V��K|6λrI����Nh��@n�l�$Bhv��h��w~��{������ؖzu�=Z�#�m���c�ԓ�Λ�����[��].'�v�F����&�j&�+�z׮�7��
!~�s�Հs��j���UEMZ��\���`��	��0.�S ϭ�\f'16�NL�z��֦�*`z��[q^�b��K�o.L	��0&�S�W��ژ��nĞ��$H
G�r���>��`}�T���S{/-����ۼ鹤sYQ�v�e��N'N' PA�Qp�l��-[�[ncRc��x�N5�@����?��}j`M���,��Zr��ۨ���9}�f��N(y@�S �B)�
���g�߳=��&�*`z���kKqȒ�"�#��������ٟ�fb]�����y��;So&)$I��Uu�l�����X�z���.�����M��Lliƒ�=�]���*`M���BL�%���b�#Ѯ��)���'���zR�r��j�m=̫��f'16�NL�?����*`M���,���.[��6�j8�W��fg���u��/��4��s@��<nĞ��D��z=/0=exə����~��Z�0&����}q�7"Ć�94�]���x��eLz^`z��K�g%ڸ���]���l��OK�	ex�~~~_z�5WM��=�L#\�V$㭭[��$�q����W`�9���[ۚ�cm�0	�y�,�Y^0?�v��LRH�R5q�}�hex����6ʘ��J��	W-7�sY^0>��`M��$��3��dk��Q�&h������ܒw���& �U#��� ��T4�!/�%�vf, ��uZ�WR��UWo݌	�T��Yy�,������Ϲ�p����ll�ٶK����3��Ua��� �ɵ��-�I�����-����l�l����Ƭ`���&��:���${�ۚ^�zoY�^�q�0y���I9��w4W����ؽ}4�����mc�(�6Ei��9^�@-����l�y[�,����ս�{ur`[y�,�J�6�ٹ&��!��R]0�,+rf���XL�R$%�m����71��ֵ�Cr�~>�B$�F)#���AY���A�إH.�6ޑ"� ��4��؆4�0p�)3
�H$BBҮ%B1�L�&u1`1R	#����2�uh�=�F��"Fh
��:��v��0�icĄ!6Ŭ����H�i�ʡ `�`��?|�t?��0���`Så F��0�0@"L�P�B0dA�)B�#
�"VԔ�����T��
. CKi-
EO�M@��33i?�f�@ �m^�6��t#;3u���#<���y%�	o�ϛ|��>-S�M�vL���H�UUK�Wjێ��]�x,&`�d�X�p�����d�(���cyH|^x��u��8=e{VS�Em��z�`N,\��ųҁ�v-�xH������d�)%��;%�8�f�\ԍ,rpA���ŉi�|8�����P�Ү��'��̕�*e8����,,mYl��Jf�sݎ)� YwktS���h�4�jݼ�Mah{u��N��fn,R;;O.�Sq�m95I��l�8�Ҡ1sn؋����1��9-O�M�X��;h��ju)�զ��T��<�H�M-�p��%M)=uE+�]����9�f����C���`z�J9�ڜ�745v�IAk���nx�t{Gk˳�kW�ʎݍ�mJz�lV� AYb;C�&+j���|����̳,�jx��Tv�M�1!Å�լK�2�~Y���C��mn��{gd.L�!���Xj��jE�#�9�^;DN�]o!�ˠ<H�����	G� h6*��@�jj��k�(j���\7n�`[�t؃9�˷iM�Nv6Q�״j�lE�V�� {!�"͌�e�j��l��cB1ѱQ��z�4]����F9�	�u���.L�Bv�CX$6N5�S4m�Ni3XL��v�%���4U���4�`�vrm�.:L�\����7.�N�c9j���KtRpg�xC�.	4� ��M���/Z�$n���;�2��-��>̌��rU�t�9%k����Rؕ�U�2�W��ŕ:�kI�'T�7F�	�:����E��������E[�q���n,��[�j
Nx�����J)G���0�g'!�4�b�T�
[)�`�h�RB��vL����k��J2�2�S�n����U�nM�:�W �M��.��825V�R�9���n�Pt��'�Sˍ���<��`!��n,�Z�F�R���MR��<!�����S@��^�P6�����C�������;�����^`9��apQjݷ-J&������;�K�6���{�]�(�9Ee��E{q��$��n��{bi���ۖ�KK:��Q8�yJNXx^	Zu�����I��%�\@�m��v(�8�.ѣJ=	gmp�����kx���)�q��c����v����Z�;v�b��b�ñ��l�!MiO\;��vJ���{�O{��ݤ�7H�uoR`'���0��p�Ѵv��]�q���c�1b�+���\��~m���~sI^0&���>�� �[�^K5q�j[�Wv0$��y��M���[��w4��Vc���ℓ4����n����ذ�b�>��UN�q&�B�8����^����s@�z��ݍX�N7����%��~�%x��eL�o0>�:���q3D���;�`�&㑋��c�.3�mWh��ͪ���5�ݞ�7 ���W�	�T�>��Y^0=mi9�+�D��m�}������}��7B5D(��&3�������w���>��&�LRH�R5q������+�O��7vJ�6ʘ*��;�		.H7����$�l����ff%�����?F��ڍ9���W�	�T�>��Y^0>�/ϻM�j3VVc<��k�wħ<�9�M��L���uk5�Nŝ<����l�u��w�k׋�(�j#�	�ۚW^'�Ӊ5"HǠ���5�ŀn�ŀl�u�	%
ds�T�0nE�E��/��4\��BP�"!(T9�u��w�=�uUh�wVU�jfj�%
%�ߖ �V ~v��z�@>�u��D���I�3@�����7퓘��$��u2b��f'�&1c��+,ɳ駎�V��e�w<k����f�@���ɀ}m���`I+��*`X�T\��-\�7����$��W��٠[���qa��4���$�l��?~�������W���V0�6�P�f���z��x�x�BI(��(P����^u�v4�MH�)H���4��`I+��*`}�w�[��vh��5��r�oE�t�p�r����ێ8M[e�A���)#Ƈ"�r}}��I+��*��?}�y[�'\Iv.�ʲ�L�Z�7u��%
"dsϫ >��4�w4�]ic�D��I�3@�eL�o0%��I^0>�Sd��F�"R= ����]�����U���W�m�87���)&�׋ �P�I%��/��~�`��krM��H ����R��E����n��*a�a��j��l�e�]�nQ���l��]WAÔ������u�{+��:U0nM�݃[U&s�ܼ�[�l����Y㰫��P�x�('�,�]�s�GH��3�v��Ɯ��%����ʭ�/��:��<�^��m)%³�ۯ����>|@�mc!epJ�z����i��k�ۡ�ݎ��;i[l�ǥ�[�չ�S�~P4��*��3D�Mk5&h�!E��.�gG��n����em��u�%Ӯ���x�8��ڍ92�������9}k�ͻ�J?Ho>ŀ���Wjj��˻X���tDL���x��X���|�7Yԉb��@?��@���&~�����^0&�����ob�����x������I^0&���?��@���n`�G�$�h�^0&���>���W�I��^øz�v�)�<�O82�q/7�n���f�ݣ<û��M)ͣW&�����������`z��~��hl���)wR��!!�D�z�m��?~����s@z�,e��
!L�먪�*�ʥIrA�������I^0&�S ���[�*�f��1$r�݌	%x��z� ?6��$�_>���U=t]3��qBI�+���ٟ������ۚw]���*���dc�ȤS�p�K���}��2D����UhuݻnK$��g��`�7"d�(�#���{�@��s@�빠r�^���ƬǊH��r&'���W�	%x��eL�o0,�q�1<�Lq��Nf���s@�z�5(���q	$��7����`6�UY&4Ei��9^�@?��@��sC����V�f��Y�L�$$q����}m���`I+��*`}L�\��[3\�/����uF�
7KJ�;����v�8��qef�dö�i(���`I+��*`[y�Kq+�.��đ�Wv0$��m�0��@��s@;�5c#f916ℓ4	�T�>��Y^0$��AE�:�#IEz��������}}���}�r|��G�NNw�s��'o�ƬǊH��r&'&�׮���s@�z� ?6� 䣶ɓ�*՗E���v��ؤ�W-����X�Y�p� �ӹΌ���ԂxろLs?���s@�z� ����]��n���"Lh�$�v0&�S ���	ex��W��}Rc��R8�JG��٠u빧��~J����_=�m��1�mrA����W�	%x��eL�o0	n$���\bđ�Wv0$��K�X��x�x�	J�M���O��ܑ̫ӬqP�䮼�1OZUa�v���7mpɣ�u�����;�l:[l/���������W�ܞ�G=j޺qr˖��؅@��1�:�1�	˱��r�V�`˺�٬l�#��<��d刻Z�wFN�b�:m�w`8�m�u�gj�&�m�٬�U�ⱺ�y��u��ZFv�� �A���tm���m]��%�o���S��Ngڙ3Yu��2�j��+*D�粫��Ҏ6D�vz�㫎1�j�ֲ��y)����qBI�����٠u��$�
,Ԫn.Kx\��L�o0%��I^0&�So�-�)#ǉȘ��^��w]������4�.5 �8�S��w^,e� �ۼB�/�~X����r$�ƈ�M9�+����h���7u��9B������sVR�F���5��ݲ���
=Y�9f���s�un�uVNc�B�9�!��`���������	ex��W�	�T��T$���ū���sY^>���d��)^0>W���l��u��diɌ	%x��eL�o0%�� ��2Fc�n(I3@�z� ���Y^0$��AE��B���nj�;�0����W�	%x��eL�_���vzv��=r*lk�X���#Tʁj�;^�\��#����\���-.�z�`��`/]t$�����x��Ɯ�����4�h�w4VT�>��Y^0=min.;N�Zt��MZ�6^��ͻ�T�H���#<
�@X�`F�֐	�C�4~RZ�:�hb���mN!j� v	� m��4�CLk)
	۠��B	�H�"$���*
�!�cH���P+$�����HBH=F5R1�p��R����10`FE#"���^"�O�����^/�j�N ����B(�'��|;]��]�|`�������-�IB���ŀ=׋ ��k��V�nWb��v�r`[y�,�J���α�F�Ʊ�$�:��`I+��*`[y�BL5^5n.���V�k�m	�^m��u�w+Ҏ.{r����m=�M��Ǎ����6�ӓ4�*`[y�,��\��b��Iv�����eL�o0%��N��p��n�Ŏ6�Sq���`�ŇDD$�[}� ��Հl����x��7#i94z�h��h^�B�~�߱���@��sƤIE1n����`]��}o0-�����L�#�
6�I�RF8F�Ne���k>��dx�x�\킔����i�����@/��޻�����9�D�8�q)�_���^0,���0>��\.��B������`Y+��*`�� ��S�*˱R��ʫ���
y���/_= �[4z�h*�:�$�916�rL�*�^�_���w4��f�!'V%j���/��'�Lu%�D�A��3��a���D�q�$�l�#�9��j;��ɛ͐�nOlQ]c��bGu�g8��;�n�\���ѻ9���hv��m\i�uQ�1�FiS��h�x�4��u���ή�ؗ�<��:N�:�ͶY���c�������d���ˊ+��Z��l�����*#�t��p��/;Y��^;Jd3lp��MP��e�,���µSf�L��E��v�m-�HI�$�Lm�;�&g�n�` L�F�3��c�A.&v�����0-���^0.�So�-��5w,�\��s�^0-���0z��K�����ҊcI��-���eL�y�l�Z��\�cPQ�������f�o]�������>��&��j'1��H��w�r�}�~��,��Xɹ%�	6z�c)u���s�p��nF��I��i�U�ݍ�۶��P���l�u�l��%��`[+��*`��[���]��M+*�� ޼YK�$�B$%Z1U~i<#�}��u��nI?���[�s@�U�\d��&$�rL��u��9L�>ŀw>ŀ=+^&�X�bq
8�>�7�y�=�����@������צ<N(,jF$����,�l��[/0>��}'8���J��s	ɰ`�孰�u�3���ڮ���,��������+v{T�]S5k�ϱ`^����(�!��o���s&I�AF�s4
�W���x���΅
d�k�j�Z���UWu73WX�����¡BV�#�US�@�#��{��|ٹ'����@��+prLLmǄ�h���׋ r��%
g����UG\ݫ�R*��Wk o^,������޾��w4ϟ\�IHAIܖGS��-�\�p]���:1�	�=���Ѷ�]Y���1ɉ�"�f�U��޳@o^/G�%P{��X���5^��U]Q4Z��� o]�$�L�ϱ`ϱ`^�@��cVc��b��4z1`�Ň%
&zy�`s���UV�E��Mͪ��D(��}�`<�7$��}����b1�A\_!�-��3@���8����h=u�t(P������ o^, ַ���	����a��������ڇ�wL]����ux9�u�᥺��w��>7�y�6nY�8��=��[ҙ�[�s@��z��Xۃr`Ɯx)&�oJf��D$�No�`<�����BQ2�=�!�y�3@����*�^�_���)�ʫ�X��LMI�X
"��}X��x{lX�3���}���\M��"�1�
8����]�8_��� ���J=�~�o��w�f��`�z8�[�E����t:Z� ]��q�h�r=x�.ÖW6����[kj�F�t���l�
�J� �\�c���n��Ɲm��6ڎ�h%�DAǜdh0u�6�;i�;�쳰փ��s-ln��ɧui�1Ѹ/��Ga���ʜ\��׷ �1���lr���s�@�=���Q���p�y���v��o�|��n�K�s�����2j�JB�#��r��6�|��6�]d�Z��Z�q�	[<1��tB����NZ�5sd�7vT�����%x��eL��`zι�v�U3v,�Y�	(Q�I(UG����?z��س�(��5�eT���v�����h^�z~�h��h��h�;Sx�c�7��{�g��=ϯ �w��׋�Q�ϫ ���pnLӏ��-뿴z�h^�����I-��+�mWu5fz ��5�p�:tu���c�ܙ���[`8�\v�亭��"3/Q�7j�T�iYUw�w�`^����DB_�;�d`zyT��%�f�.�Z���z����«�zA��f^ �yz�gD)��Z*�'"�1�
8�޾��w��o]������j�x� ���nM~��}�0�ذ/]`t�s��7��m���H�$�ӟ�z�h^�@-�4z���A�,�bp� F����F!��غ�sxXݺ[�����0��[�?��|����1�(�Ng�^�zoY�[�h���?�v���$q��� �y�L�ϲ0�ذ/]g)��_kMɍɃq�$��}��z�nq@ڄU � $�߮oy�!~�4���T���	��C��{Ͽ,��V 7��=
��ߣ s�ɯF$�"�G!$4
�W��/z��_o�ޔ�-��Q8�����6����i�`þ>�(V:�J����7n:�)����z"�18� ���M޻�@��4
�W�r���1�p�b�Uw�7�#?�L����:y�`z� �۪70xID��s��oJh=u��N�׀w>��7u�L��Z�W6M�Tݘ�ϫ ;�^ ޼�! ��HJ	��O��>����@��M�#�)n%#�z�Т!/{����{�� ��������S�%����qJ����N�%���ݸ<q��.er��k��4�7@�H�� ��0/]t~�;�^ >�T?)1�	ŉ�f�oJo�?$yz��s���b�Q#��U=tMUҹI7$4/_= �������g��=�<h}�7AAc��z�����׀w;�`��D�s���Mzc�&A1Iܚ�)��)�9z� �x�I%Q�BH�!#	A HH1"�!R��$D�H� J��H�`Ad#"A�H��$S��E��,�1R�V	) �	"�EJ1�B���b�r
m�p>W�R��FKjVQ��J��*
G��b$�4�
��>X� `B+!$H���G4��JV��(y���$,B	 f�	j��h��dHCL�v@��I���$# 	�b�.U�;Wxy!�5�]�,FA @!)5U�d��,)	
0�2�jo>����fۛl mKvإwL	ͷ�d��k����]K�S�R�ev@�N4��a�.:砦|��82<5qeMtШ��UMZY��l -�m���u���7��F\+Ƌ=]כ�7i�]NLn=d� 1�U[�ga����#K��{��7��gq���;�ᮣ�q�b5�q�7e�����=����u�.}���n-������t��(]]ԹM�]�:�'�g[��B��d��n�VFӳ�5�y��+��T�� �s�RY���v��'�.�lR�޶.w����F��5�g0@�7'c��;�����Ô�a7�azvB��!Tk�n)�΢w.���-ps�:�i,��
ӯJ�u�Ӕ�!V�q��[�!;n��2=�J�t�g4`�)@p�Omv�Ź:�ڍۙ�;`��m��*��6�.�v���F�ɞ	��Z��V�H4�vI۪�I�ˍ;i�//Q�a}0F�g�J��"Uli�·�S��V{�:�7Ca��䎞��m�m��#�r���\�@Ks�)=��3��S�7�/O���x�g�\J�ݞ�����)&3r#�!��WQ��c���oz1<K�R�(�6��ս�J��S͗��U1�3�43�s��y�'`���s�f��ݭP�:��k'1�/nHv�ec�t8����؄���C)2<`��`����s��&#�TdqT��]䜬���Z�����ZR�E�r瓷FRT�{@nw@��`Wgf���Mme��kϘŵFj��A��l�ؕcPv���j��wM��EݘK@�tmab�8�+ŭ��鮣Z�m���֎�C�l7Lv���I��wTp�ӻ+m8�����w�V�X�DG�[Sr���;c���M���N7(�9^Y���Mm�r!��\�	Ӥ��Ft��y�l8���vy��歓Xؠ�8Wi&Θu�U�;kt�ٝ��r��L���
H���IZ�kZֵ�YsYD6�QE ��P6�U�;US<��<�v�CJ*�jd��Y,�5�����7l6���ym��m8�	�q����0$�a�s�Z��Ϯ3�q��b�֫��<m���gn��́%��j�H6�G2�X�6��-����/n�Jf�#U�zu�Z5Wb�8�A:b{�¯���]�(�ڇvu��Ve;�%5�Ѭ��cz����keҗ\�1�.��ώY�/���'.�th��wz� _;c�uι�K�x=��5qGYYgkѺ���ڛ�ȼdzw9�+���|�����R���n������X ޻�I/��x���ic�L�"���!�Uz� o]��`�:!B����Nd�(�q���@=��[ҙ�[ҚW��?�]i������MJD�<�`����u�ВIL����_{������3@��l��[/0-�L`����M*3�H����ʝ�:ӛ��¤��w:��v[��9������|b��r$�p,��/_= ���-�L�-�M���
W*��*�uu��Ԕz��P�$�bJ=�>�ۗ�{�� ��z/��9?D����4zS4�هDD)��}X��xͼ���/#H�R��^�|h^�z~�h��b��������̈�"���,��u�t(S����}��=�f��~����Euv��]rܙr\er�qF�(Z�:�x�=m�ƺ3R1ۥh�n�"�nf���������"%��O�Հo��SUVUU�Ut�����F ��0�n��w��dr�:)2C	�'�޳Ɓ˭z/߳���p���O���w��=����U\j�i��,I��!�����z���^�o# om���i�aP���7�[�h[w��oJh�נ_�������N`�]�h�ʹ6.�lzz:�K1i�E�}��[h�ljLx���mɠ}m���)�r�_���������D�'���R`�\`vٜ�G/������y�K?$u�֓&LrdLQ��4
����l�>����Jh�ڣ�2GS�%۽ɀ_[�[_��������~��X�l��{��rO������4�ۏ	$�>���ޔ�9u����)hl&���SJ��ʸd�g�=܋�T�l\���\v����{��۱<��L�ǉ8�����g��Z�޳@�ۿ�U\j�'#��7$0�n��!%2ϯ �����f��4��7&	��޳@��3O�^��4/_=�ݍY��~���4zS4zS@��zĽ��w�<�s���)15!��)�9z� �x{lXDlG�D&��y��c��^�6�+۬�j��Ϲ����s�y����e�F��u�^{Dh�e�=���t8�b5�ۃYP����������&Z��-�鴪F��p��/(����ڹ	4��%:s����-�˚mr5�0V�]lt�$�ѻ�g��������W�vNCT��3�0k��z��gM<��uS��-�NwVS��*2*jK����C¬���jkD�\ֳ�`cWF�S��n��Dv�F�k>���q=�:t� �r$ɓ�m���y�����b����sw]7J�]�������� ?���D(�;��n�h^���1#�g�ۃ�	���r� �w����&\�6 �n���lcx�	�I�ٙ�^�U�z~�h��h*�5c�L�&0/]`�����s� ��4�u"�cq�rMLn
8f�Vg&r^���Z9�N��<��{L/��{q[��MU� ?����,��<��B�_Pz}ެ������VU�weM]��g�E���{���n��w�	D)�{���M"�nQv���Xs��vʘ��������,�
�W4M�Tݘ�D)��Հϯ w�3@��4���Ԅ�6�RV ?���Q�����9z� �-B��,cSڟ�#�in˝��lk�!���6�j��`�q���%����k-]"�� om� {����\�D/��ޚ}�l�Rd�<Iǉ�f�{��铧�V v�^ ��r�QJ"P���^��U�Ҥ]U�wf��z��{���
�TC4 �k�ס�'��M��u5nLq�{�g���s��;��{l��S�ϫ s�R���j�F�q���h�ٟ�/������@�z����Q�Q�"I�ì�`�c�e��
��3`\{U�88NV�M�R(���qE��ڐ��Jh���6^�興_�;�`ϲ�Z��Ș�mHh�W��߳?$U��_[�`�ٜ��%Gw]zn�Z.캴ۉH�/���@�ҙ�u�M���ﬨm�䘡�
G�����{�xX�|`^����D+J!/(�*P�dBKw�X ����ݫ�R���5V,^�0$�W>��9�Հ7���m���߻,�:������*[:u�v.s��x��v_.K� �Y����Ts��]v`^��6^��ב�BQ�B���\m�5nO�qh���7u�`�ـ~t��D(�UW���cn5�$IG��{����)�Wj�9^�@�ʣs������(P�K�`uwN����3��m����}�7��"iF���?:np��/%
u��_����5��nI�
�H"}쟮L���.�.�˜[��4sۂ�6�Ξ��v-�wC��'1��i՗�]��^-L���Wm�.�xrO�۷&�R[u��k]t5�..��tRn:�hi��I� �mQɛ�dN�m���.�됙�3TnՀ� �k�zmѺ�gi^[�8��̖�b�q���t9Ÿ����W��G]�1�r��E �<�������{M��z������{��v��9��.�����pr��&�94�v	٫��餻K9�Y�l���FMUU�\�{]`��0{l�D(��C�?yhw��ۍ�0�7$�@�瑞�P�d|����6^��B�J%_c~P�$1�N<M�4�<h�ڴW��;�S4
����$x���0>��`M�����?�?~����ˮ6����I'�Z+*`I+���uUn�'�o^[�C�`��m����>|�q��#�m[t�\6��W��<�vh�{��~|�>\��}�g�w{# ׶�����<����W4L&j�Z.\ӹ'}�zo�Gb �Tڋ��r{�o�'o�߳rN�^Fz""ɼ�.j��SV\����ݘ�]Ӏl�u��!L��# |���U9�H㉶�qh�W�wu����`yB�^J+}����~�j�j��ՕWvM�`��0BI��?�Wt����-ˑ�S�F�E��[Fs�{N:כ��i��o7�V�:��bn+o�������f��'''��=�x�?��h���;����Uq��H�����v��Q���Ͻxw{# m� s���tXp������v��y�$��&fq�O�]+�F@v1@�bcID�Ԅ4�[V��+V1D��`AJ�dF,`��~���< �A͡��6$H�!
#X1!�0RS|]@J&����"�V
DSL*f���B9H�b���!1- ���"<xQt/��"$P�D�`�,����T�Sh8��U>_�O����J";��W���J�_�����w=�7Z�Mڪ��)Y7vT��(�	z!%]�� ���~t���]��ssV�E\ܫ�EM\`�`IDz"7��O�}��7u�`��R'h�5b��ҒFʄI<��˸o+�Ku9�#����_iD䉼����J4Ԇ��]�@/�o �בВ�����9�뛕V�n��jIr]��^`I+����F�Z����f$}�<��NI��m@nM���0/�Q��V� ����ĕX�ՊT�]*�����ל`uwN=�}����U �X
"p"& AI���䞿����B�Z�Xr\��Un��y�$���m�B��]�s����EZ.�sw"���-s���}>�Ђ=��m��v�g���#TF�ww�}�6�5�Li���{��&�o]��_�S@��z��4�����Ի�ב�
d�w��ϫ �� ��TN`�qE�Ls��~�M�ΰ�IL��� �}��~�yST�K��U��MMف���S�ϫ ;_^ ����3����E9�H㉷���]���w>���w� ������~��W����;]p��n��6�d��/��shDb���l��T���#p��v��݄�B�`6_'l��=�m�!�87	�fv�x�Q�29j�Q��Cg���u��� ��uptR熊�չ�du�J�ժ�:�#�Y� y��N��2�{v��5���:���3�9]nr�x�۬���ʼ����ڹA�3l�[[�2��{�<���S�%���)X �����RtV�7�[��F�F�u��y>_,Uut����m��~����`]��}/0	n$��9C$���3@�t��U����h�س�Ъ��O�O��7wJ��U�wf���`�]��/�d`���6~�m�<��I&4�z�K�}4����_�S@�z���px��9Swxz�0����t������o����lsn���f����72�k&��V<�ͭs9����gH+��n�f��������`]��}/0%��`}:�M�C�1��i�����?g�g�IR��Q�Xu�����������s	"�&�JG�r�^��^F�"e�0<���m�5W3wk�$��w�0%��`K:�	�T���~�ʿ_= ��6ׇ��&�c����m��C�}_�sϫ ׯ# �����&3�I����;.�G˫��vT�\N��Wc��O1GWhG���O=Z��6^��6^��5��򈈏���U�~��x�2I1���9^�@�# ׶�e��IB����*���WvJ�n�f�� |�# ׶�$�\~��3�uz+k�>�U�<�d�U3W�%	K�`y�`/]`y%/�~�y�\�+V��������0	�T��eL	e�Σޝ��b+��m:��$g+�������"��;Ş��0�V\H�{��{����]�eMƤ�U��u뿴�)�r�^��z�I�)&7���z^��}��~P�����}X��Y�
!L��T���8bĜhr~�/��r�^����DL��Հw>���j���n�+����l��6ʘ��0���~���
���)�z��A/�k����w��P��"n=���%��}�? �����?l�*���7l�\t3�]ש/:QַA2�;]ӥ�%�rsq<rAc��z�w���m����%Т#��w� �z�19����G0i��^��*�נt�u�=�bϢ:�Ts�&UQ4MT̉<�yw���r�w�v��>�4�,�c�Iq6�=����)�^����ߗ�{�@����n(�pm������u1�,�0.����eL� �w�2x�Lf�Ɇ�MI�e���y�N�j�v7NW�ϫ*�q���m=����&�sj�r��ݍr�N���Ӷ��P����]nvlk�=�J湴�X|KmA����n,��V&���\�s��MV����h]��ۅ��sd2��1˒������ܧ���Pu�F��f�6Nݰ]8�����C�؀����z�f	�d�r6���{B��۵��a;<سy�ѝ��ns�{Ms�́��Ӹn;r����n��n�=���z6֏#�,Iǉ�g��<h}k�9^�@�ҙ�UUƝ1�Ǒ7!$4
����W�^뿴�)����]q��%5G���9�Հ=ב��!D%2��N�V �kUUuE]��E]��U�B��%
��� �u����`/]`�*r�x9�9�@�Қ_Z�W��>�w���덛0j90���JD�\`�Y��:
N��kv�t����y����߾�x~Z�y1�Ɣi��*�y��W�}zS4�)�}�4ɊI�8�qʺ�6^�ƪD$|�D.P��gd`�x�9}k�?�]i7rH���)Ɂ�+���u}j`M���UUK*ʱR���*�X�Q�Q
�������r�^���L��u�NJR�n�l�� ����<�B�%��������hzS@���*i�5d�Bܶ��=�]1�r��C��3�u`�|���\�ӌQ�n�'���z׮��:�����^�k델��ȱ�H��� ���΅	B�;� sϫ �}^���kf4F��ē���)����qU?�S0�t�����D>W��
�s���3rO��߷�@��Zo#�pq�jCC���_=�_=�]��u�M�LRLWE�M�������DD/BJ!w��G�w��`/]`�X�M)���n��#r��G���`����֬n���ㄜ��iպWM��&6ԉH��)�^��6^�䒈_����ܪ�x�*�Xj��.1�,�0&�Sm�0%�Ş���>�S]R���
���˻0<������J)���X�|`��i�j'��L���W��:��7$ﻯM���eA '�C?���z�����1��zY������eL	�T��d뼇�Y�MV^��j8z�.�l:�>�M��nܝ�'V�=E��\�4����0k�f������BI(� �� �_lM�q4�MHh�W�r�� ׶ŀk�fr�P�M�V����i�ԏ@���@�ҙ�u�M�����ZM�$�"&�JG������8X�|`^���DD)uϫ {kÃ�<�p��Jh^�@�z� om� �ք��
R&0$�	:����(�!�DW�H�� �dH�@	A"� ������XT��.)(����1A�<�(b���|��������4.(J%0�K�	q*V��#1��p.J"5#X%+F�f @^l��ā�Z�@�&ACA���FI!(TL�`0RBa��'�˻�'���~6��@�m�� :Ćؓm�l�WI��b��CkLi�
�ٹ:�Q��pu�Uz�P��n�\�=�j�ᫎԭ�B*ٺ]�v5�k4� $Pۂ;]-�'[k���l�m�@unW��r�1��x�W���˻B���q�KS�#=B�W�N��W'��q��4q��y�jcjb[Adi���'�h�b��`6e�BG ��v_&�0)�b�l!usf�E�ꧺ�T�lt:U����5];�cX�Mu=���Y�d-,\M�:1��Gv�l��<����͏f6Xl����t�vOXx���/5ޅ8��]���^4 �6W8�!�	@�ڮUڪC��]������d��-�W���nALrs��y��$�Z(��f;4`� �<�Y�s/(i&Ng\tJpH�� 2�{sZ�:D��jd��s�L�S���1v��]�V��D�:�ӫis"�"@dZڎv'r[R=X�lH�����]5Xύ���C�k���t�Q�Xf�"L�OLu�͸�֚;9^9���cq�tv���$�4��LS��t�HJ���J�}(Q��Y�ɭ�9U�WQ���x�Z�x�	�D\��N;qd����kmR�J�b;��R�Ԗ�0�����v%�W�d,[��r]�.̜+;mֹ^3��mH�0D9኶��2���΀#�"`Q��X5��h(����N�`�e�nyy�m�Umь�!I�5�N�9�\q
:��y�y�����mӲI�'6�n�ɸwQ6�6�\�Q7�����V����D���G�C�܎�&n{N�H���VIն��^��v0t���7E�.�XmL7�}t�˪Xgf��e,�E��hӲl�I����wj�v9���դ�*��"�+��.Mv�v��'KX�Kۥ�k��i����Nڔsʭ�;��4��TL�i�*�tON^���;7N�a0/�v��q����UUK�������>;ܯ��QqQ����@-ڞ~04@� g��h�����sպ�.�^mSm1g�N(�ú�^� �'Ov\q4�m�1�k�X����W���<�!�rݷv�ڃa��7e��d�s^����'�����픦�Y�A���8-�k��G�<�Dsݴ÷I'&�8L��Ω�G��㱡u�\��e^-v��E	E�5�Y��
4��=obF�X���'�Iħ;vm��k��5�%�V�]���`���34e�Z�+�u� �ע8��v.s��츦��g.K�m�lrcR3q�I$��W�^���� ����"}A���z_*O�����"���W��-�L�5� r��tBI)���*��
�W*�Cq����@�Қ+���W�}z�[1��J'1$����W�|hy�`/]`yB��|��`ϲ�G��J4Ԇ���z+��z���]��[��LO�D�i�˵��;��kZ�NŮ;��U�s�<n�3Zz��{���͍�I26�nG�^�z^��@��s���3�^�z޾֓qI$��5��Z��;��n���`�E�A ~�! �����Gv_>ŀ}=ΰ����
!)��}ʪ�ッ�8����__nh�W�r�^�׮��������H��e�e�^�X	%
_>����o�pX�!$ȓ�@�z��Ҙ�x�����D$������fJ�����y��p�i蛍`�i�1vm1^�l\ru$��;��w\�������lFo�C�������W�	��0&�SYq5���5����:���9^�@�z��Jo�?~����}�7��88ҍTլ�>�e�5(U �(A
/��(JQ	%
��[0z�`}Z�9��#j!��z+��zS@���IzJ+��Հo��S5W7wwrr\��Ɂ�:�	ex���SU*�:���)�s"r%r�<	���ظ�y�;my����Fǎ5�z�%��{�����+<ٳ�8�7�/��4
���_U�^�M �q����Ȥ�C@��^���Z��:����~ď.�oȐJ��.�\�]`���vه���e��4.���k�H�ɑc�Iq`vـk׋ s�u��%	B_(QP��_ߧ |�VU�T���nj�3v0%�F�Z��u�d�0-�#s�k���Ɣ �#��|�����:۴�W-�˜]<�҃H�7�	�͊���_U�^�Of ��Ɓ���T��wj�䫫��]k��DDB�9��@��ƁWֽ����>������DN8��@��Ɓץ4�fg�ؗ�{�@�w�@�_[���Ƣx''&hrR��N�V���(Q<�~X}�kј���H�$4
����O�����X��`
!("
o���]��
ܨ����.4�l���V�����9Ϝ;�R��m��OfN\=p���%m�$ͻ[s۷���:|�k>^���k˻*�۰�]0.T��n\��h���]ك�=�Ӡ'�qw)X�=�s͝�Ж:�K��㋪���8h�W��
G#��;n�9uq� � �&����;��G�����МWg���`ݿ���ݾl�0��]{��n��SN�'����Ӯ��O|ur�s��5r���c{N���'$�q��q��Z�^,^�?�H9���;��T��\�wrI.���Σo�L	T��u�d<�F�sNf�ץ4�Z��u��+����,�٫�廽�w	��0%R��W�	gS@���7�dRd�D8�@����$�-�ߗ�;� ����?m-N�I�g�VN����9�@�n��[K��3�/s=vN��mU���P+T���(��������u}j`J����q.�j�0�5l��ܓ��7Q_�A��(Y��߫ }Z� ��ŀکv�NG�"�(G�ֽ���]��Jh��m�8&I�7JG�J����Σo�LT����ɑc$����>�w4�)�r�נu}V�W�\�"p2~O�I�k,�Y{9���E�9�^I�@�r<�m�Q�V�x�Ei�II�^��9}k�:��@����>�v&�9��F��4_Z�ؑ|޾��:�������9�I�5�=���]�5
&JL%�(���|`_u`�WRm�#M8�R-��s@�Қ/�zW�h��q�9#M��`K+��Z��u��+��{o���gIXT���*n]]���L��\N��6<Tr�=�q��p��Dū��7֦�]`z��,�}1�P��&F�Q)���[ؑ�̀k׋ �wf�!$���kU7j�]Z��]�%����<`K+��Z��V�׮6�5"��R	)~�د����={��nI�g}w"�T��5P���~y�^�}z�M�s��(�Nf�7֦�]`zΣY^0=�ر�v"��F�.�8�8\8���U�lO6��,������G�ϖ�r�j�3�|�W�X����W�	��0/���nIhi��h^��^��/�zW�o�1#���7#�$i�njv0/��x���SU.�=ex�:�iֱ9,�8�$��ֽ��8�^,�Q/�~X�j��J�h��Iv��r`J������7�^����ϳ�m�X���H�@�9�a�7:�������Ûn&�)��n�Kt5D���˽�[�yv.��)�9���M�����x�٭';K۷���k�����[��/[4V��;��y�8J�x;��ǲ�_�9ә�:�pr`;s��Wl�ʔq���kU)��[�1ɨ.����v1ƖR��Ӟ� ��5:�8)"��.�#�w������|��#V���t2�񋱝/JNɼ�n/b����n�+�:�#'a�<��:iV��>ŀk׋ ����%��}8��4�x�Y�JL�:���9}k�:��@����>�v&�H'�Uk ����5ֹ��BJ<���~�b�=���s@��,KȤ��q���K�Y^0%��o�L�tI]��ԕ5us7s�|���<�/(�����|K�� �Z� >F��b*��Wr#y#������]/��k�����n{qk��������x�,\�jė$.�`K+��Z���@�����tbr<YqBHnI����D4�F*�"A�:~T?
������| �A�A�A��~��A�A�A�A��~��� �r6{�������ut,�O��w�����w��A�A�����b �`�`�`������A��@bA ������<��������lA�lll~׿sS�h�j浬��؃� � ؊�=����y~��yg~͈<�����k߮�A���߽���\.�Mf�kS-�M�<�����{��<�������f�A���ߵ��b �`�`�`������A�A�A�A������!Wk7fR.0Q�p3%ܓ:駹|�:��h��:չ��w�{���|��ؒF�<�������ٱ�A�A�A�A��{�؃� � � � ����lA�lll}�߸lA�lll{����Lѫ��]Y��ֳb �`�`�`������A�A�A�A��~��A�A�A�A��~��A�A�A�A�~��؃Ȉ7w��n�w���������
�"df
�y~��y~��yvy�0�b��0ʝ��0h l`�Hݸ��h��pX�����"��gG��� �E�tF隴�D̢aL��],3 q"���:2�!XX0F�K��Y��B�
a�l�@�X���ք�A���Y���4R%IF4���>��@8�/�	YFT!R�X!HV��E�).2.+0a��2*$��{�8��)KQ���<# �
��"A�
��AشE>|��C����N���<:N�? ���A����؃� � � � �����A�lll~�~�ff��f�a�5�3Z6 �666>���6 �666>����y~׿]�<���#`�����b �`�`�`�}��?L�3XCWY���h؃� � � � �?{�lA�lll}�^�v �666>���6 �666>���6 �666?��?�p��MkWY��Z�*�6��2P鍉ˋćNs����h�/m�k�f�X͇WCL��;�����w��������~��y���y~�� ?����������lA�lll����˚�f�E2k5���]�<����{��<�����{��<�������f�A���ߵ��b �`�`�`����fg.Z��S5���F�A���߽��b �`�`�`����ٱ�A�Ull}�^�v �666=���6 �666=�����5�W5.e�˗Z�y��&A�����y����v �666=���6 �66
O���>��~�y���5)�&��Y�Vf�Z�lA�ll@���~���Q�?w�_���l��`�X�p�r�P���'=��-�d�����gv��p�W�[M�Śr�H����=ex��ul��*�Xl�Iǎ87������Jo�g���z����hz�h[�:19,�H��� �z� �Z�$�L�}� |�Ɓ����C�d���7z����b���@����:�����z��4���1c#����:���?ٗ�|W�~��;���h�H���I#��E*?���#���cR����s��):���ɝј�uw�[��l\(��L�� �8��{
u�����>�C-k\1��<��eD�I;κ�.��Q��l�;�L�ȳR�)vԄ;K��)ӗ�L��N�+��7`��ZS�H6�R�e�#���ی�lF�GD�p�4��F��k�4lv6�S�p��)��A������͔#o���>q|#8��ڻED=��z %ԥ�m���3c��nq��j�囒yn'�E�II��?Ɓ��z:�?�!G�ϱ`�eMR��j�n��Ļ��*`J����`K:���`�̊L�Ɠ������:���߿fbW�x�*���/ܥCn7H�������%��� |�e�����F�xԉ�mƇ&hz3 ���~�>�^�X��j���jV�u����vVv����m�����.)�;ˑ�^����M.7^�4�/]`�\����� ���j��͇WB���~}>���s�;�(�%�>�ŀ>w���� �kU5�H,dr6�Z^���n����3?%W������@����'�d��HT�����T���`>�V��s�m빠^�X�G18(�73@�z���X���k��n
�٫5�P�8�0�N��k4݋b��L�M.�<��V(����/�9�*��������t����>��y%�A�>���q��CN8��@��s}��f$u��4
�|��ڷ��+|6���ܩ*�`��`/]a
"�	$B^�	D���vN ��, ��M:�5wY��wq�݌	�T��V�Y^0=��h��nĜ$�����>�n�%���׌	�T����L�Qe���<ĉ�n��O��z}63f��V��44�!;N�Jrz�N*�l�7�X�����x����m�0=����}�$�c��iI��n���z��Z^��ץ�y��Q�1�3@���X���k��־7���&jK�����	D���>ń�w�ٹ6�=�(��@w��{z���m��i8�R-�]��׌	�T��V��.r��صvv�d��މ;Mv�g$<�I�rV����݃��n�ڱ�iǊ87������s@�eLEn�%�� ���LZ�,�w!ov0&�S�[�	ex�������d�d��Gz��Z�x��L��ŀ9�Հn�j���W�ۋ���%���W�	ex��eL���>���O�ゐiI�^��IC�}_�}O� ׯ�%�C�`X�B�oN\�?[r]e�g���\���F�<ݳ��,��n�����m�Zc]�܍����e���`�F�v)�sq�;���F��H\�te�h�IãOo�|bI�b��5)`i��s��щx�9���`��l�Ց�;�[��l73v���f6�k�X�OWg`0�X�nͷ�t�<���;�v�t��� �p�xU���m�̓�3�n���]��u�u�b���g��\��I��m��v�n\����\-e�lN$������`J����`K+����&�drA&���_U�u��,�l��}7��.K���]�ݬ	ex��W�	�T��K���F�x��xۍL�:���9^��*�X��Kqj�-\�n�ڎ]�	�T��K�	ex��W������b�r�-���rx�F˂�^�+T�vx`��F��nѺ�;rm�9.�_�����`K+��*`Z��N$�x�$i���w6��?(�
����,�s�]k���U�<rG�% ��4�w4_Z��]`z���(���v�5#y%���7֦�]`z��,��^���#�	4H�@�����s@�����ДB��k�䛪�V����InܾN��N��K�q�[;��\��p�+����6�6�q���q)��ۚ^��+�� ���.�4����h]������z&�]`K+�-��H�,��9�+��_U�6����H#�A6(�������`K+��LW�up�ݚ���]�`�\����5�ŁСB��|�y�cN$�x�cqhz�0%��o�L	T����bڎ��u�뮛�>k�3�:kj۫n�[��ZI^96�ź�U�Xx�����������|o�L	T�������	gvv�5#y%���7֦�]`z��/]����d��M9#�:��@���Y^0&������$�.KtZ�n�k�W�	ex���S���B
�E�A׿s�.䜽�q��n493@��s@���@�K�Y^0I�W�,5gn��ɒ臡�<"c�i�F�RbҜq͎1�GK�t��N4���x��j9�/�zW�h^��^��/��'jL�8��U.�=ex��W�	��0&��ӣ���)$MŠ}z�hz�h���_U�u덽O��An����`M���*�X��`^�X�I�8&�i��9}k�:�� ��ŀk׋ Ց
.���@� �H�� DI" D"��d� ��B,BBʙ"� D��ZU�ƒ����$ ȡp��T�B!e ��P�j� @%%t�S�]� �H�*�,	,bA`� �>2��H3ĩ
�h@�l��"�H���|�$p�ĸ�5A�A��ڲԶP�6l0&��`��&
0�0�J�	��U�Ԃ@�0	 F	# �I�T��9�kZֵ&��֍��  �z�Ζb�.�BD6[,[t��}2��<u�B�w���%&Y�[����3Mv�nl�u��Z6��f��@ג��Tl=a���!8m����ګ��K�)B���c�q����rq^y��y�m�"�6ۥ�݉�@��ż��\�]ٞΟa�ݙ�1��[tj�c��I��D��$�k����޶G����F�[��̑��d�)t]cRu�z�!o`ڇ^�<��W\le�g;�vZ�U��˞�nD/&KVt	���̝��Zx\c2鼔bU7] 1@^��1�s����'�[�Ǥ���Av_
�N�st��,�lU:]֪���8�v�&K��[Ge���uX�s*���UR�f�;%�Τ��v�����
z�Xy���6���xxd�B�ne",̹�;hĜcw:x�[b�5a�ŰDP.�&X���T��h��[��B�v�� T�gst��̚8�ցր9sl����Ɇ��9ݫQ[Ѽ[��S�ڵ��܍����vT5�ƃ׮g@f�'c!��vS��zZ�y���9}o��Nutm��nf^֍[���]�l�j�ˍsvڧuJ;�2����c��,ݷ���d:'8�-�a�ѓz�H�l�YzMϊ�牮�>q�.�� ͍ok	F���nr�l$<��)X�;�~m{���9=]��Z�i�v�pt	IV�z�4�-&_��>t�<��������p�9�.׎8<ٴ� ��:��ɚ��/�5�q�8����c��z���8�<��ڵ���,����[���f�k��,��\.�1n�J.M�͔1��Ѹ��c�P`�T�W9��8,�98N�z�ۧ����@�ye1[qY{g��p�}����;*`��3[F[�Q��4kk��u�c#��m�[j�:f�&�WQ���Rl*+�[o�i�:8jU�q0/�����@�2���`���tʪ�g�@�]�M�@�UU*R~{����iF(#��#�|��]
��� �G����	�AO�E��b*�Av�!��{2Rک�{7;m�l�9��=m��n���˪��#���͢+uH��]N���i�t8z�� ��7��l�`N3�ţq��U��gt�'��/wll�<�ȥ��vu�0��͔ⵏߟ)�@n.�M�]s�3�Tq"'M�z���t��1�;m�V�ܩ��s���/H�/Q��r��{g�5��Oc�v��N�C��nġĻ���{�����s���j����xÑ�@#����@���whǱ��h6�m�2drA&������}z�hz�h�����n7�i�q)' ��ş�#�ذ;�X��9�(�f6r��8�G�NL�=���s@����Ц_S��7�b�mT�]]N,[ܹo.��Z��u��+����}}��V�zQ7&	�r=�k��(�}�~��X��� �U��mZ�PKs�eݎx�\Y�/��:���+��:��Kͽq�Ѯ1Y=6��Me��z��,�}j`J����U�Jn�ʲnʙ�X�x�WB�V��J�B�^IG�9�Հw��8�^,�����"pM��ә�r�נu}V��빠u빠}�YbL�n4�D���н	$������ذz�`?Z��Gq��i4�8��@����%��o�L	T��=���L��I�ռ\�ѹ�</WnA��k���Ů�pf�����曃N<Q��mƇ&hz�h?7X��<����Cy�, }ʦ�N8�<jG�f���^���Z׮�׮�˸j�j&��8�nG�;���{�ٹ��v*�n�d C@����H"!�l������9w:<R(<qG ��/%	DS�{�w�ذ���e�z^����H��$���u빠y(P���W����>z�`�dڔ*�Ů&d�����.�����{>9����]��~��{��|�q˹t]�]�����Xl���+���`{=e�2A��#�E�r�^��?~�H�}��__nh��Z���Ӎ�4�wE�����ŀk׋D(����t�z����F�x��xۍL��g�����|�p���)(���B������>:�=��f�ߺe�C5�d1U���]Z�?m78�D'\����,�]���;�"�c�&&�(H>�ME�0N�qAds�PF�ݭ��\m����V�ra$p�E�r�^���w4�w4@��4��H��E�8��׋=2>}� �k�p���ДL�ϓoS�"�"�Bs4������@�z����>�,�0�#pONc��Sm�0=�^0%��g�X�&F�@h�����z��w{���ϱ`O��jPB����~����]n4�]��+lV���r۱���'o<�{s���\^I��Y��VQ};u������]���v�T��EݺN��㴃�P湳P;uV�k��/�ԧ;ue�ѧ)��Yƌ֭ݐ�N.1;mu�E�C�a���;��[\��6�X4�mEq�:F�8�y�X�j\@Ν<c�=���bC�.�M�L�;)�������W]����>v��8�n]Օ3{&�$�&2d�q�b7F��qV���:SA+v8R���0i�����빠u빠r�נr�^����4����hrf��^,��29������>z�`��:c�35��3@���@�z� ���^��.�����G*����^�XДDN��=�F���H��)q��[4	ex������eL�������ڻCD=�=mt 	@\�p�����u7��)&��d��xӃ�"��H8��^���֦�*`�����xK;���Ը[sF�_����C�)�������o��׮��V�&F�@Y���Ɂ6ʘ�o0%����V�~�(ӎF6�"R= ��f��W�o�L	�T��}n-\�yp�$��sY^0=��0&�S ���o��~��[�ѩ[��[Ods��u�1������)�8�-�&خ��ۚ��$N7$����@�z�ﬧ�������*������17����W�{ר��W�o�L	�	+�7���E�]T����ـk׋�$��p����w�}��䝾��rN��ƞ��	!!��}}��.�����zץ4�K�H'�H'�%����Sm�0=gQ�,�m������)&���xns����=�M����TH���&��������|� ����H�����@����׮���^�~�(ӎF6�"R=�Қ^��	��0&�S����r���X���u빠r�ק����@�Y�@;�Ӧ9&1�9�4_Z������0JD�$  �@F@�� �h�����'/{1XDܘ��M��W��>�)�k׋ ����<�'ܲ���I��U/)"H�7O��{���5�gO&F�躳�wĺvβM)ea⧞s0��v�߷�|�~Y^0&����eL	eũ�7�xXwq۽�Y^0&����eLY���Gz�A����	�I��*�y��W��K�g���s@����d��H7�{�0&�S�u��7ֽ��Q��m�D�zץ4z�`?7X��XZ���(Q�b��ŷ&nB�!������Kڧ0�n�}`%7V݆�Cm<�u<F�w���a�Z;Q�=hh�#��tc�!�!���/`�9�G��<3Z��X�ۭ�l-#�c��χ̮+O[���p�ۋ����b���6�9�Nl�1j;a�6�A����@�Nuc��ǁ`;'<����h�sl�D�׷�m\���ɧ�%�X#*�n�ߞ�ww�w{��{����;춻\�%`��N���8:ݫ��Լ��[�{d���q�TAE�3r3��X�rB\@/��}j`M������4�I�x�NG$��ֽ�S#�}X�0z�g���XT�nLM�&�z^�zץ4�w4_Z�]�n��H���6���g脧y��ذ���J"�\����i��8���Nf�׮������U��}z�h-���.��ض��ƒ|�B�S�;9��5�e�0�r�m<ue��^�Ua���m����������==0=�uZ�r՝���ܘl�����~���	ey�r�׾H�X��q����dJG�O���Y^0&����eL�����.ū��,�}j`M���Қ�F���ǎ4�rL�6~n�Q	�>��o;� ׯ��/�)�-��0s�����c��?-��./N]L�l��ǃ��t�8�56J�!k��-/�����u��7֦�Lm��I<c�&�zץ4�w4_Z�W�����ċ��i��8��K*f��>ŀl��`$�D$РH���>�|����Ra��"�U�х -�6�p5 E���O�<RNq��J��!��
G3&5-h�ґ�P�c�Z&ÀF7��"Db�&J$
�*Jh����P��غ!aIb��H
D�A!�����Օ�0̂B����B"�VZ�B1����C4����m���;��c	�F��T|�qO?0$��A"@8OT�(��"�C���HB�k0�QP��
(. �������S �U�AC��D Q(��n~��� m�XݷER�"y$�x�s4?���_{�@���@����:���>����27��"�=e��B��}�~��Y�HRB����q,K��tt��e�f��e�p�'�����p�=Hu�r�8��kgv〭���;dV��3��������ow�߮ț�bX�'}�p�r%�bX���f��L�bX�����ND�,K=ߏ�ے��e�e�v�|��{��2w���"X�%�ܾ�bn%�bX��wٴ�Kı;�fț��QO������[�oq��������y����r%�bX���f&�X�%���}�ND�,K��l���%�bw�������oq�ߏ��B�t-f&�X�%���}�ND�,K��l���%�bw���"X��!����P#E#`�T�����L���bn%�b������<T��j������ou��{6D�Kİ�TV>���O�X�%�쿿f&�X�%���}�NG��7���������[\a뮛�Gg�$3pm���n���n��C/8�q���@��#l.j�Y�f��4D�Kı=�߸m9ı,N���q,K��{�ͧ"X�%��{z�7ı,Ow��Jf�5tkZ�̖�Ѵ�Kı;���M��EX�L�b{?{�m9ı,O~��H��bX�'}�p�r%�bX�m������g�*_w��7���{�3��m9ı,N��ԉ��%�bw���"X�%�ܾ�bn%�bX���~�ꦂ�S�����{��7���ޤMı,K��m9ı,N���q,K��Ȟ��~ͧ"X���~?nJ{M���-����ŉbw���"X�%�ܾ�bn%�bX��wٴ�Kı;�oR&�X�%��Ȭ�k��ɑ��.f�qs��d�R�[��7v�;!u�m��OM��K�]����c�����>q�;�=V}n6\D���܂.X�h��f&2g�l-�1��قM�r��y�ݦKz�/%I�2H�겶=;q�R��m�Z�P��^�c�/	����=��C� ;Z���s'Tv���5��/��<�d�-v�d�E�O/�3ʞs��&g52a.Ve֦MSR<�xD�״�맰��b���q�*8:9��%y�d0�ff�u�ND�,K�_�f&�X�%���}�ND�,K���"n%�bX��}�iȖ%�bw;�/�&]\�h�����bn%�bX��wٴ�?�PH�L�b{���D�Kı=�߸m9ı,N���q,K��}�/��ֵ�3Z���fӑ,K�ｽH��bX�'}�p�r%�bX���f&�X�%���}�ND�,K��70��af����jD�Kı;���ӑ,K��_{17ı,N���r%�`~ �߿sR&�X�%������kV��kR�m�ND�,K�}���Kı;��iȖ%�bw�ޤMı,K��m9Ļ�ow�~\���j��\�/Mr��aOt�X/7l�Cю;v"瞃ip�:4��M�MkY���%�bw=�fӑ,K��}�H��bX�'}�p�r%�bX�e��q,K�����.MkZ�j�fk&��fӑ,K��}�H��@�� ≉�@J�&D�=��m9ı,N���17ı,N�����oq�����>ܔ��/"J����%�bw���"X�%��_{17ı,N���r%�bX�﷩��7���{��??>�~�7<��Q��Kı>��f&�X�%���}�ND�,K���"n%�bX��}����oq������m��k�mf&�X�%���}�ND�,K{�5"r%�bX����6��bX�'�}���Kı9��]]f�����n}1v�s�:���7���S�r��L�݊7�y�WnJzh��+?=���7���{��oR&�X�%��w�6��bX�'�}���Kı;��iȖ%�`��2��5u,ֳV˭H��bX�'}�p�r%�bX�e��q,K��{�ͧ"X�%���z�7�eL�b~���%3ZԺ5u�p�捧"X�%�ܿ�f&�X�%���}�ND���`������7���H��bX�'߽��ӑ,K��ײܚ��jɣY��k17ı,N���r%�bX�﷩q,K���ND�,K��bn%�bX��^�˓U2΁������oq�ߟ�~[{�d�,K���W����Nı,K���q,K��{�ͧ"X�%���8���O�(�5o3�8��9{-���6�ݭX�:�kv:���諒��e�MffjD�Kı;���ӑ,K��/����bX�'s��m9ı,N��ԉ��%�b^��.z��S�fkWZѴ�Kı>��f&�X�%���}�ND�,K���"n%�bX��}�iȟ���,N�e��2��kE����ֳq,K��~���r%�bX�﷩q,K���ND�,K��bn%�bX�Ϻe���kZ1�ֲ�f�iȖ%�bw�ޤMı,K��m9ı,O��ى��%��
�Q ���߽��iȖ%�`��sye�k5�ղ�R&�X�%��w�6��bX�ʠ��}�����D�,K�~�ͧ"X�%���z�7ı,Nt�t\�Z�of�S8+�\s�nl��%6خ�ώk�1�2W��N9�E���=���7��,O��ى��%�bw=�fӑ,K��}�H��bX�'}�p�r%�c��~m����ON�T���oq�X��wٴ�Kı;�oR&�X�%��w�6��bX�'�}���O��}������Tt�!4�3�����%�b{߷�q,K���ND��!�2'r�����bX�'���f��oq����~}y�e�x�m�n%�bX��}�iȖ%�b}���Mı,K���6��bX� &HM��XB����-���Wt\�Su��]kFӑ,K��/����bX�^I(D;�Ր�!I
HRB}�aSı;���ӑ,KĢ��/s(q�K�q[dsѝ�L)q����U�Qf��E����N�J<{�]�d�uroBa�vdq	���v7&2/��.]��v�t/�n�vm�i�����8����4���.�Ct"X�\t+U�Q�İuF��`]�2��x1������}:��%xnv��mZ��u�1��[��{8ݣ�/�lVm�7��FWUFNy�+]mFe{��Ͻ���ϟ����0�qD>�u�6�'f5��k��3v��y��7#��g=+\-�i}ߛ�oq���~Ͽ{6��bX�'}��D�Kı;�����A�DȖ%�쿿f&�Y�7�����O��<�Y���oq�ı;�oR&�X�%��w�6��bX�'r�ى��%�bw=�fӑ?Ǔ��q�߿y�/���|��ı=�߸m9ı,N���q,�"{?{�m9ı,O~��H��bX�'��s-3ZԺ5tj�捧"X�%�ܾ�bn%�bX��wٴ�Kı;�oR&�X�%��w�6���7���{��}����ӵ�/�q,K��{�ͧ"X�%��{�5"r%�bX����6��bX�'�}���Kı/�N�,���d�ɚ�q��&J��l�g��8��a�ظ�%�Y*�L��@��w�{��7����Ͽ)q,K���ND�,K��` ��2%�b{?{�m9ı,�^W��l��-�����oq���m9*lH)�ȀH$v
�P��ı=�^�Mı,K��{6��bX�'}��D�Kı/z{&z�MSu���֍�"X�%�ܾ�bn%�bX��wٴ�K�"{߷�q,K���~᷿��oq���S��k��-*n%�bX��wٴ�Kı;�oR&�X�%��w�6��bX�'�}��w��7���{���'��<�,�ND�,K���"n%�bX��}�iȖ%�b}���Mı,K���7��oq���������3���F��{@���8�K�Lt�\����cc��v��9��|����5wJK��&�!~!I
HRB|���Kı>��f&�X�%���}�ND�,K���"n%�bX��w�Ջ����=���7���{����bn%�bX��wٴ�Kı;�oR&�X�%��w�6��bX�'d���ʹ��qEK������ow����m9ı,N��ԉ��0���?�T���"}��{�iȖ%�b~���17ı,N}�{2��f�V�f��V�iȖ%�bw�ޤMı,K��m9ı,O��ى��%���$Ȟ��~ͧ"X�%�}����k5.L�]ffjD�Kı;���ӑ,K��/����bX�'s��m9ı,N��ԉ��%�bxϼx��M���mҖ������0 �ݜ�Wc���׵��)�5�Ƌۭl�w����,K��bn%�bX��wٴ�Kı;�oR&�X�%��w�6��oq���S��J�t-/���bX�'s��m9���,O{��"n%�bX����6��bX�'�}�}�7���{������dډ�eu�ND�,K���"n%�bX��}�iȖ?�U�Dȝ���bn%�bX�����ND�,K��70��ae��v��$)9%�J�]������"X�'��f&�X�%���}�ND�,
���������q,K���~�Zf��tj���-�ND�,K��bn%�bX��}ͧ"X�%���z�7ı,N����K7�����Ͼݮt�(�c�"�p;>5�˻]�H�u,�� �����Ej�ti�d�.�u�f&�X�%��w��r%�bX�﷩q,K���� %�MD�,Oe���Mı,K����#��V��=���7���{�?>���*ș���~��Kı;�����Kı;���ND�,K����x��"i���{��7���Ͻ��"X�%��_{17ı,N���ӑ,K��}�H��bX�%;��#�tQ��U�=���7�����wu~�Mı,K߽��ND�,K���"n%�`3"{��|m9ı,�~'�_�^��д���oq��N���ӑ,K���߹��I߽�I�$�r��BH$�� ����������(���QQZ"���Ȋ*+�(����(�������A@(�PA��"� D�,B�TB�UX 
/�QQ_����������EEh�*+��tTW�PQQ_�AEE���TW�DQQ_�QQ_��PVI��O�	7:�` �����\#�   �           �        >��E PUP(T�B��  E% QR��R*R�HHR(�R�
��H
$UJ��E)U0   �  (  $  ������t�]{���s���}�� �ʌ_}�;�s�p��ӊ�>�z<i�w�I�N  /W���   �PD@�@  " (�
}� � � �J�l   @� � T ��@%�� �   ��h� $i�(� �����  &�@��@ H�o�{>���מRݞ��c�Yq����rWq� w�b�f���#�ݷۼot�� �  >��  � ��|�{}�&�ӗ�^�#���������w�s�Z�Z�g.��(���M�vU�k�8�r�Εp ��G������q�;۽����x� >>������ݼ��ۄ��:W| <�      1 
{��k��oM�ִ�[u��U� w�q�����\c]n��w _{�kq�v��g< �{k�$      ���,f�g׷�� �=�X��ݝz�y�]��MG�  < �    
 @���u��o��w/m���rt�� �/=^�]�����s�7���>�� 
{�|�;t�|  �'���X}��{��맾}�y��O{y�8�0 ҙ��{O�3^{}�'�ˑ> =AS{IT��  ?�iU*���Ǫ�RoH��  D�*������F#CO�2Fԥ* �"$�JRHL�hx��	�����O����mH9�ڊvݻ��D%	^����PTWAT��(*+�UTW��AQX (���t��X ��$XP��Y���(o��-�л���iYp!#dad�y)�11d�u�</��%���JI7�L�d�X?�)���R>؅�a"�4=���6< \$Ӓ6Zf��rB51�BW8m���$d$$H4�)��������@��B������)Sԍ�呎��a� �1�fH`1�Ս�T�#D"@�rd��HB���\FP�\e�qy
sp���c�r�	+
�ˌ(A�+.o'�� TĈWP�Л��LQ�I��\cXR��sS��i�6�>	����%��͐�y�(t ��|<�K����+�0ٚHƜ3?#EԆS�I'	0��X�	s�$.o(�(Sy3��	,.���]6.����l�60�`��cM��!L|<�^�_4"e�/�B��[�˚��#!�	��I�(Gs	s��5�&���1�1���IYVP�ژJd.;�$cLӕ��a	�l�)-��+4e����VV����%���f���<X ��H���U�noᒰӌ������#L&i˦�����sx��Rn@�١���%�P#��L���g',,#�/8z��9�I�����&i.l����&o)|y����e�no��6��'�Y}��N�C���0�]Zv�j:D���\9Ä�{Xw��o}�WJy��y=_χ'�d3NB������
�-0����*�*V(��
1XDӛ��D�ՃMx�B�D� �Q)���J��H��p#R�B1bD�#�
L59ā@�F\�)$��s�������ً��0 1�����&7ye
��Ӈ�Ж$�&o#8T��5�71!s�]i�aw����!� pӁ
��=X���@��|��S	���|�{�ln�!�2!��j]v��Ò�lI���hH�q�d��nMͰ�G�!H]9c�+�
Aj�X�������tX`B�q��zO����Bc�r8{�Ӂ�+���s���i<1�G9�ayp���w��������<�<%3N_F\�xo�s�K���hK�at�B�x�椦jK�����y���<��3�r�c
l� Is�0��p%�1�8$,����&d<��IL0�!���-q�.e�7O!s��j䌠Ss�no �R4���wJfː�����S���,��h�HJb`@��ar���T��# `P RC�4%S�y�	@�]���h�y3�~?1Rs��.h�L)�(d)�(J )��52GN�<%�A�ᇇ!\5gb��8�
��ZJ��xs�=�~�wK����9�<�a�g�~��q?)��D���8l�I��8y̴?g����5%1���+R+y�$�[�����1���k4p5�Jsǁ.2�.a�
q&��1�B�I�rp�g0%`L.�)��y7ɛ��)
iYnJ0���+V0 I�?Y?%�k���?Z��% ���4� Wxp�|���
��ĲSLÚ0��s��(`��n����3x�np乼�LS#q���8�0��x!L��F,R4jB��хL4�lX4�l-pu�sm�9bXB�x��:P��	��7zn~,��ɗd�g�!�����M�H2�9[ ���Ă�>���q��B)Xw�&O�/���*�aP!J᰸m	J.����BR��#�B�o-�y&��I9L9"���j@�l
0��
k�Qn���Ӂ[�xk
���$��Z���<�asÇdJƒ(`f�9q�BIapxO3xK�g����7���ԅpLJ�D�D�����$��#b��C@�L�̈A�#�$
���@�Ɛ�D�e0b��s��jqa�P	VP�������C8�=����#p��sF._<���%�{��Ҙ��1��1e�!w��F4uy�
n0�p�o�����q�p�fz�BVxˁ��0*)3Nh~�t��L�'�.BJJK�+`¦#
���p省 B\7��������~`�<?$
�Ʀ)
I��+�3����8�:D��+��|?��o����P�)�DI�A�A!MS���R�A�N2���b�`x�M����~�<$�]HшL9�
;�f��i�<?@��)��d.hB�fp�n�zSɞ�ZaHq��L�~fi's��g/<<��o���W�y�\%�)&���p���q���4�<�*D���`x�	sN_�0y���D��i�xR�N>o�����~�L!r�'�H��?'<H\e�R���IsN/��2�'0�.�����?kvp�L�&��c�6\/%2����6HS�$�n������3|e��sF%$ėg<8o�s�ۧ9s�~����G��������`�^(D�:��%�=�"re���V-2#3>��k����L 7-9��l���1y���} ��P��HE�HH�p<�=���&P���x�9�$J%}��|��/�_�J
EQ���R���E#��*�k�a)�������EZ�q= �1!s4�!�22���M`ɛ�!�8��0��4�B�Ɔ,
�h�t�����0��tx{���IL B �ɓxK�d#e��a.M�䗉.$���_%1 VHXW!L�5�0��)�\��u%�YM��&��[����9ᦰ*BˌnJa
�F��K���Owx��{�!�X�<`Szg��n�:2O2$
��R6$5"��H�)��K�����|��SR$�U���G`�HFR19�B�i��p=b��F�>
�"D�*H&(�D��
��`�xh+���B��+���,hfJ��<B4�^&�#� �:���q4��
�2�L�!���A$(��"��Z���)����!����8�@�@��,R74�N0!���H��J01�S�h�(���������a�i �E)��.�䜱4�
0��)��ĭH�#!��X~a�4y��,�X��Á�,[�0�=��N䟥���|�HPp�8xk��u��H������]��OߓĞUM���*�@�C�.3Ie�C#^[	y�&����a���|<�iōmM���P�X�$�
S�2��o%���㧜8�xx�x�~d�j@���B������
��MH�L?Ùm��0�q��0�0���&C$��LS�8�H�BPӏ�y��l%"��*�
J����&���Nfd&[��g��� �"|w�`�=�	�<�+��=W�X�H��c�d��?�b������!-�����$w��5�$5ńR\�|��g��1�����r�s<��M��
HB�	dt$�l��׉��x�Č�i�<$Z8�3�ф*葹6>�T�����M�����-�����h�'�
D!B��#MF�%3YÒ.�dn!��f��ͬ����#H�@��cL�ɶ��S4!S �"���
��@�aJ�	#*�f��ZD����M�S	d1b4 �H�����Ii��8�HB���R�q�\5�V`���21�@����0!L��� H�"�!B,��J�w�ݔ��$�G�K$�Za)��̅M�C�H���2>�#☤i)9i��#�qd}��ɕD�x���fuM ��!�+3\}�B{B�I�!��$I�$�b�O�Ēp��`�����Y1]IV-�B��s�1��0�Hd�Ր$0q�&d ��s��Јd$<,��?����A"�7HxR�)[y�(\H��s5�`�-7ÀE�
D�`hi�:$H.�D�B���_bW	FQ��.��d����ZL��2���绻��M�-�����n��ۖ�W�}��ur�����j50�YTȵmpm�   m���JI� -��� �]i� H��[@mm�n�- m�( $����p  t�L�����l�ЭJ���b�$��^F!�K����j�ey!īJ�tVfH�+��k�����U�jWy���ʛ[[��  ����X6�v��{����>��lB�9:m��۷h@-6��&�v7Uc����`�[M�UT�s�d�<��7Xam�  �m"YE�M�bۑmn�׾>[@�&�n��d� �ڶgK��n�` �`-��.��o�e���t���t��k�l�!z�!��a��a���^v���m�l 		 ��I8H�`����Uy^Z��#���-�l�:@�Nr��G	sNڶ�hmfvl� �M�Ԁ6�;�$>�[]�J�Zăd3��6:�^[�Z����0U -�#�f�iG �ח�U�kd>��3�]We�% 	-�p��ʭ�mS��zU���m��m�I� ��.��١��d-�-��Z���Ӷ�ۀ6�@  �S[v�_$���%���t�d-��� ���B�m6탂�$�mQD��%cz��� m��m6�@qκt�l�{j�8 @� ��h�! ��M�� �~��m��  ml4/k�-�f� �`��֛[�pm�    	���`dgN��An��� ��\�ڑ��ΐ�[)q�hz\�ҫJ�j�6��[v*�8P��Tc6�ԫ������#!f�N:&פ�֜m�!��I�iW �[M��1ۯ�荱�`jy�j���n8j��v�(���-�Wy��U\�jGl� e�]��c��	qU^�mm m�I2ICI�GR����-)J����l�۠ �B�&ݮdúE�0`�����������T.   8 ��8ٖI��Ժ)v�q���m��媫᪌m���2������v$�%�N����UvٓpU��4�sC�\J�Lepz%�-��A�� �N�9ݧ,�R�:UZ��H-�L�m�]5���[I��m�`ַ'@$ !$f� {D�d�&�n��[Y�m�:C���[�m���8v
b5�A��mn�*�����b���*1O/F�N�����m�L�`[mif�8����/!�UAA�҃M�� .IR3�� 8 �:^�m�8�e��y�W�m��/(rN�mm���f� [@Hp�hH8ԻV�$�R�bB�s��kkl -��e�Ih4�@-�H � �BO7m��5��n۰� ��� ���� ��� m��mt����I%��8�� l .���ۚv�V�%.sm��Z:8����l �[Al�m����J�m�� ���:;:`$� ��$H�$m� [�h�m� $6�M� l�,�� ���¶�m�%4Pm��0m'`���bU�P:�g���\�' xy��m ��wXl5V�U96�At���I��Ԋ��6]�v�m� M��-C4�Y8� ����Ս��A:�ʵuu����Z)m�D�im�H���k|��O�^����*x].��hN)j�e��6�C�0�(���&��[xkX�n�� p����l:����WK(��  �JIoJg]�J�knւBk٩��I��  m$�[E�\C&�H�Y;I$��6i&��vl�� �-�n��e5���u�ݭ�"��YV��g6�@���h!̶��$�v�g��l�P  ��4Psh�Bh�I�~+�̬k8� ��� -��m�e[h�b���h
tuU�p[UU)*��T���@���m[�8 �v���hࠥUT*��2�\j4s�'�z��G$�խ���M��t��m�!��U啩nVut�E�W6]jy�/5[�򰶭�z�m&`gI���P��i�P�UT��^���]$��eʵԫ<�+ �t�n��[���8�^���?�|��U������g����7�jR����6BTU�َ)j����]F�ݔݒ���X�Tki� �]�s�@�k���n��dҪl m����N��VF�7vͶ90��WR� �2��q'm��Դm�d�,�E6����ݻ��$i�m������.Q9K�*	��+UUJ�qj<�UVq �S��^T�����Ғ�	�K���m�  ��;k& %�ZM��l�6�2�QÙ�+��^j�z&����W�O��PY*���U/C�^k�Ի=UB@ ��h�m �U@U*�[*�UA�t��/[���m�z�� y9`t�J�۹�E��ՠۀ�}��H4Idm[�� [Nm�m��b��ڶ����d[Y H�^'�ۖ��`�F��kuI���]h m��g�L�^�u�9������Y�iWj��+���m8p �����r�����m -�� p�����%�I6��m�����,ݱ[l���9+�-��[*����Mڀ���h�2��h�����Ŵ  m�Z��G;v[V�	  մ   IK if�6�q?7�S�,�j��^T��e9VY�WUE 58l�I�m������֚L  ���  9!��Zn[r/Que,��m��7lA&��A���P'U��,���`�$^�8��� �p �$m�6Ĕ�|��~R����Տb��V��*�@p*��^&rp/�]Ul<&b��N��tÀE��쾓3�$2��#��n1VҭE���Y9�U8 �VV�F*��� �u�,� ��r��m ڶ ���F�#vI'H��֜[�ڹ�&u����H��iY��J�++UmJ�U&.�0T�C�v7A�1��ưP&M
����[���V����V��`W&�ں���y}U��K�:*�[�6�-� � �^�nʫ�O�@~J�*��V�T�ҜH9��@�nj���ڞ\ભ��m�ۀ$m�$�(/V���m�$��#aV��j� (@x$A��Y��z��� m����HF���-I�A#�� b�m� %Hpm�ui6�m�� �,��v۰ISH�F@ �l�l@@ГeYˉ ����n�H��nͻl�m��p8��X֮�N��@	gm����ZO$�q��V8�0H�u���u;��6�HH�u�-����m��Am8��P  ӂI�[�C���t`$mu��F�۴�.(����%��e�j��4]@�Wm�J��}�F�����&�k�[l�8DB�s���Y6  .��Hm�o�iА��m����kh   
]\ҭ��{�KU*���m�  m��޹[uk�6�e�M���m[5�.���:Hqm�ٓ:�v�Y��6Z/Zm�    9��hN��Qmr�˲�- @��� �v-�AL�H9�UU�Ji�%�	V���Z��屶� ݶ]6�>  �K�� v���� �J��� �6�%��Y˶Ȑ  k&�L`-�Y�EPN�kwf��q� �� �D� ��L�� �g�Z��U]uα�mv�p �lm��ve�͵M�$  ��N�afI���zVUU���Wl�ݩ��B��U�	T���ǭ���KL6�ٶ	K�  h�ڶ��fضMl���WV:�*+�ee]�Ӓ
��5,i�Pz��m&J�Ӣ����[�`�V�@5���m��i.5�0 ���6�����}��`[@6�Y�v�l���U��Z��q��VZ3���l0;�n��������v�Y�lE���ٶ��n���m�UHL���*躠%Q�VTv��3���&m[-�b� e�� ]��@�k��p���ō��[D�pn��CIi�@�UFRwj�<݈C͌T�q3�:N`+�V�� �[r�[&�m�v�2�@ -�&�-Z�R["D�JA��^lm�6�8`�ZV�6݀�� 5����w+l %�D��[wIz�-Lh��ݶ  
��i|�Q�j��Ea���i6��v�b� �`9$�� �R��^� =Bi�s���;��ʄN�  k�FM�mmt܌8H�C�kN6��[�mj-Șn-H��m�H �ׯ0��  H$ ������;�QT�v�**]U]O ����xj�I ��T�R��g� ��Q�!��鵻gAu\I��c��)H]&�H�&�  8�$��c�6ݭ����V� N�� �`*�i.y%�Hݦ�9�ۀ��  $��]UC���ʻ�R�t$Cm���  -��^��� �]�d�m���ws�UD(�@~W �`?�A5A�����Q�P�
���'���@�@� O@< ����?�� 'PSAC��x~US�<
�OAG���q���#�tT|D���<L_U= ���'P"��� *��\N�ު��(b#�P8����}P��W�'��T��'�A�)���'��&�	�� @�*"Q�x��#�`��*�>����@N�(&���DW�T�$�dI,X)�D� �����F�	a!0�H@@� D�$�dHD$!#$		��/5E*����=D(�]�? �@�P��
�D|�8���T࠸�(�?�@�z*�����<�0G���4��C�>x��!�< ����@��} ��cPR#ꇩ�? �D���@W@y�U �&���T��~}]ODP���=U}8��EC��.,�~��⨟�?�
�����O�~���\��9rKM�iq��n'@pH�,�⤹�-v$�\fE��řM�n�6���݉:M�j���ܜu&ۗ"���nz��Ë���'m;r�jn7`��x9��)�@����D��xQ\�ٹ�-sNl�dϢ���@v) x^�҇
ͺ���{i�[��"	��UUm�M�r�6y��v�.��w8�Scc��B�K����;`!���N�Ҝ8Ĝ�NⰑ�62�rFy�^w$��Uѩ��%s��%�q����,����:wku�_in��6x�6�G��<�T��nN���݆Ѱ��-Z�m;��4��j̦n�c=e u5Ok�N�kuj!X�;�\c���;�X���	���7lvx|��/j���x��av8���VYkQ*�Ib"^Rj��ю^lٯ��6nݭ��m�9���y���p����KN��m�Sn�:��ȠZ�<<����ź]�x���qQe�[�$+;)��\�:��[�[���v.��l�J���u9L�iœ�2Tƙ;,^�b�]�';9!l��%/67
�3q�8�ɳ`*|����tq�▌T]3Ǳ���6E ��e�j�L��=��@����0v.�m���ct���r[���x�ǭ���]r��PU�B�����Vi����=���nd�)=�88US���yv��4Z�|�%��cmvq���05۔v���7l�Vݝ+��D��Um�"� 7W�`���6�={r�/�K����[���R��-�n�g+�Eʙ#��j�9W4��Wv.L�[ď���ch�z	l�v��88S��#��G*�OkBY�G�ҦΥ\nxŵK�Z��9�(�"mu.A��W
�&��A�0)�RC�`�I��s^[%�RH�M�	u�m�%�cRFMr��wO)��vj�.v$0�<`��<���i͜���lN �Uk�ڮ`x�۞���سv�w2ۙ�ݰO��:��E",�@ � >T�P`#_UO� �gS�"����A^����<�n�7sm���r�Q��۪Yi�����/N��s�7,Fc�v�;�¹����3w7[RHe�݋Ѽ�u����`����ΨW]�{/s��;�^������C;r�/��M˛�s�.I�f�u�r�����n��n
[Vy���Km��
�����/v�u���e��
jL�ٞ�a�a�������s���u�����x�㭌���r�� <�9�PvL����0.���j�R(�*E�Wv���f�Ȱ�������+���?�%��N����躩�� �ۼ�I(_(�To]�9�o�,{�SP6�m�N�m���@�:hz���^�%���ĕ6��0�p�6�"�I>����̓��Ӥӻui���@���v��X�I4	����7|�h��=;��]��iy7�d�o	Iǵ��p��	p݀`�*���E�v��X�I4�nh�;LM�i�I6��p˪��*�(�F�PH�Q� `�P�>���J��ـ9m����`��t���ݪ���w�� �� ��E�vk� W6��SV�6�M�f�������4z�h�%��:im��i�������p�;��m�E�{�����!&&�!Z�<ƻ5ۊW���G:�Mɝ\<��,p���f-c�&�C���Mp�~0�8`}�`�Ȱ�[����i%M64����dX�#�;5�]��8��:V��t�N�f��, ��Nh�@�# �5�Q�A,�b�AO^�����0	��ove[v�M��B�+M`m�@�����@���.Z��cmݤ:i$��;5� ��o�� ~m��B�_7���̅������������F/g���u��P���pJ6�N���k���'N�,MݤZL�G� �� 9$xf�`vT��պm�IҤ��^�4�נz�MH�{h�)�t��CJ�X�#�;5�L�)#���4	�|��x4��a7w�|�ـn� ������\�D~B*E��)�pN����<��oʹ�ĕ6��0�p�6�"�Iٮ��T��M�	RTX�ɯN�q!���K��KX:�c��ۛF�ey��w��>@73���ߛo����ͻ�>{l脣�n����[�cM�4+b�� rH��p�7u� �� ؤi�cmݤ:i$��=c��$t�"�����܈�:v�bn�"�f��wr�Ȱ�G�vk� WeK�M[�ݤ��� ����:!%?wu�y���2I� 3���A�R�a�Oߗ�,U�Fvy����vݡ5��v�=�.�V�X*6�s[����@��m�ϴ�5;�ä8c,����m�{;a������Mg��Wl�\�D�ݝ�ˇ1&�/�x8ř`��^�pҼ�3�p�;ghw`�c[]W�y�n���r�+$�U��s�+T�#��+���&��n�p�����W\����T�{C;<���+���#��ŷ9�=���V�p�3r�d�k�h��K]��z��;�ǳ�E��㙢��յlm��i� w���;5� �:{�A���>yA�x�hM��:hGM/[��k�&��M�i�$�6�ـn����v��X�vQ֒��O�cbi�ـm�E��<�\0^��0�pi��M�m
ح5��<�\0�p�6�"�?W�����i%la���um����V�r��۫�z9�{-�V�f[U�瑟ͷ����`�p�6�"�;}�`-���;l���f��Y�}�gE�K�) $"z�'�ʇ�}����$�����f�b��+��ܦ�$��R��T�4�נz�MH�zp�C�uv�44�5����y���`��m�E�oM����bv[o �� �P�-$����9|� ?6�~�����Cj��fU��q�=��-�Nu���Y9n$�'W	{,G�sM�i��^i��@�:hz���^��4lwv�+t�:m'i� ��=�UU}v����~0�p�;p��M�]��U
����n���0�_DBP��$�B�Y�g��`_:�5Ӧ�Lm���ĭ6��p���9˴�K�jI%�k�RJ���'��\1����bԒRM�z�S%�5$�����������>���S���c�q[y5����f�/�����Y����#�.��`xy�Y�nx~~ ~��~;� ~}���� ��E�$��N�$���i�1幹9m����|��T32��o���o{�x�.��l�g���WsI�/���&���RJ~��Z�JI��RJd����]���$���ƛ17����bԗ��s�qam��I+���$�m��IO$�!`�ւPE	��E�$�a���|y��<6w�%2]�RI.�_z�^��$�d�w�%3��X*�c��fL\��lއ�<�x��)Y'g�̙)�ٻm�h�h�T+�X�ԒK�Wޤ��:-I%�6��IL���� ����H��.nQ������/=U����d����S،�����|�IZ����k�6$���Z�K�m;Ԓ�.�$�d��I/\tZ�Isו+Ǎ7��`f3�I)���IvJ�Ԓ��E�#��;&ӽI"p�C�|I�ck%�I$�%}�Iz�Ԓ]�!�]��و˻�*������_�m����c;-4��闛���ݡ�����-�Ź����D*O.�	�����;�C�J��'/V���ut��U�Z��i����N���>;u�7<�d�9��r۲�0-��؍�q�M���A���7�`�Y�s�gZ�	�u��sӖ��m\�]3���ڷ\=����wBs�lI4`�KY�uG �v�yy����v��I�?�S��sU�y���7$ݙ2�W/�������,�����l8��Zz(�wC�M���Ŭ�m��DٌU������> �iޤ��wI$�%}����4ى���&��KD�$�w�%��ԒK��ޤ��u-\��I.�mi&�c6�nf���m����m������P3'��%�$����RI+VQ���m���1c�jI%�k�RKպ���$�oP�V�F]ٱErݱ������;+\��y��}� ?6� 5뒉�6�r���Z9l���{fC��2�'�����w���m���$������$����4�נv�@9����ܷt�.l��}�~�Wy�9�a�|��-Z��@99�X]�bn�Wi� rH�E%�U��hK��'���x4�ЛznZ�	#��$�� ����i�[i%V�w�n�ꯪI�W ;�y��K�=�}�/
��n�ӻ�m���k�j�Ӥ���{\덥'FdvHb�@\��%��ݧBt�t�g �{+ 9$xnZ��}�hGM ��F�|lm�����X�#�]���� �?�̬b��)�7v�ؕ��Ȥ�	��g$C:�BF@�����$$���t��΄�0�2�3�b�J>#��>)
'���%0	a��D�!�%%����"@����U%��G<X%cN��#0��B���0��c.J�!�c��R�8�c��EX��)�P��(ꑄHBI���KE*T�I"�c�H��U����I躐"$��(@*�$��$B~#D�m�	"&���0���Eu�V%%�F�M@�?���P=H(��� 5@OJ	芇�+��(�� >�� � T��u ���}���<�N��o<D�zy��[�ۺwv��w�Ϫ��I�0�b��@����R�����po.��5m�j�t�BO$�V{����S?uwN ۾:�%	-~�]�R�:�^�狞v�W9�i'�9��A<�+�5q�5����ۯf���A����������?/�������G��L�w�`~IO3�߭M��.n���n� ���s�L�I	���q<�bX�{�ND�,K�ۼ\G�/%�WP��$.�'�W7aw�3��wn'"X�~`dO������%�bX~{����,KĿ����yϐ dL��Ͼ���bX�'�����n�3M��v�s��O�Kİ{߸jr(G"dK��﷉�Kĳ�@�o�\O"X�B���TDT1Uy����y�EOs�������ٺ�V�k��{��%����}��?D�,K
�}�}S�I��w��H$������O?����r���uX� �r��;��獮�`r�nG��ίS��\�f�M��3wx��bX�'����Kı=��vq<�bX������bX�%���<�bX��ӹ�M��LͲ�s6�r%�bX���;8�D�,K�{�ND�,K���x�D�,K����r%�bX��Ӳ��svn\�0�6q<�bX������bX�%���<�bX�'����Kı=��vq<��TȖ%!�a~�72�.e����bX��3��}�O�,K��g�\ND��T�Dȝ�y��yı,��i�"dK�ﳧ�nL�7&�͙�]��yĳ����߾�ND�,K��>�O"X�%���"X�%�|�{�O"X�%��=��l�u��:C�;�t��!��銵E?������td�)iL���#Ճ\M�������q����u$�lг�+jl����gx��I�Z5�G.ݞE���ff��]�ީ��G�؛����v��p[^����][c�cY��['N����m�0�狭�]�< iڛnvL\eMʷm�v77��j�Yn�v�k�*1ڽ�������|�|۪������v'�d:a���Kj�ܶ`^����TC�,Ua�b+�QK��7���{��������yı,}�ND�,K���x�D�,K�^�19ı,O߽;�l�vL�w4ݻ��8�D�,K�{�S�,Kľw��'�,K�����ND�,K�}�gȖ%�b^�&vm˦��ݷ2�sMND�,K���x�D�,K�^�19ı,O}���O"X�%���Ȗ%�b{��\��M���{�7���{������,K���y���%�bX>����bX�%���<�bX��ӹ�M��L�-��nbr%�bX���;8�D�,K�{�S�,Kľw��'�,K�����ND�,K����3�WjV�X������B�H�{vZmKt���s��c�^ӹti灷�w��X�%���Ȗ%�b_;��Ȗ%�b~���'"X�%����Kı)���d�˲乖暜�bX�%���<����� )�R 1�EC[�,Or��br%�bX���;8�D�,K�{�S�>Tʙ�ﳧ>ܗL�m�ٛe��'�,K��/�f'"X�%����K� ��p��Kı/��~{�7���{����1�����54�r%�bX���;8�D�,K�{�S�,Kľw��'�,K�����ND�,K��N�-ݓ4��7n�n�'�,K������Kı/��w��Kı?e�s�,K���y���%�bX�����~33v۶L����=�4��8�wX���I�h����x���/.��f�ݛ���S.i��Kı/��x�D�,K����Ȗ%�b{���yı,��59ı,O{���i�]I����{��7���}����Kı=��vq<�bX�{���bX�%���<�bX��ӹ�M��L�-ۙ����bX�'����'�,K��{�S�,h��� �,�=�Q"f������%��}�'�,Kĳ��u9ı,J~��zm��7.f�[�8�D�,K��ND�,K���x�D�,K����Ȗ%�b{���yı,JC���d�˳0��暜�bX�%���<�bX� �Ͼ�5<�bX�'{�}8�D�,K��ND�.����~��7�QWS���v�kha{CՍ�l��囓5��\܀��ƹd.K���6˻�O"X�%�{��"X�%����Kİ{����Kı/��w��Kı=���n�ٛ�nasffnjr%�bX���;8�D�,K��ND�,K���x�D�,K���ND�,K��N�-�L�w4ݻ��8�D�,K��ND�,K���x�D�,K���ND�,K�}�gȖ%�b_���6�ɻ����a�4��Kı/��w��Kİo{���Kı=��vq<�bX�����ND�,K���Y�6n�˙7r̹��O"X�%�{��"X�%����Kİ{����Kı/��w��Kı/��۶�n�SQ7jݤ�秱zy$�P�l%8|�nضm��y��JˮZݖ����|��{�����y���%�bX=�xjr%�bX������%�bX�w��ND�,K��v^�nn�˙���'�,K��{�S�,Kľw��'�,Kĳ���r%�bX���;8�D�,K��l;�n��r\�sMND�,K���x�D�,K����Ȗ%�b{���yı,��59ı,OONe�e�n���.��<�bX�%��wS�,K���y���%�bX=�xjr%�`|�"g��x�D�,C{�����L�b���{��7����y���%�bX=�xjr%�bX������%�bX�w��ND�,K� �D
#��9&4�n��&l���n��\���|�����+v�N����AWh;�jҎܽ�]v��{GYf8ů:����h�/]D��=��|nЩ��ra&�g�/>�:\:�������E�9�"V���hֲIq����^��M�u�o�RO��Kg��7�b�uE�m���ƞ�v�[r<����p'A�j�	�j%�3L����nI��&e���z� +�~��\r��;q	X�/��馠�*�C���΋��:n�N�nؖ�g�nn���Kİ~��59ı,K�{��yı,K;���șı;�����%�bX�߲}��t����w0˚jr%�bX������%�bX�w��ND�,K�}�gȖ%�`���Ȗ%�b{��Y�6n�˙7r̹��O"X�%�g{���Kı=��vq<�bX�{���bX�%���<�bX����ɦn�&f�����ND�,�D�{�Ӊ�Kİ~����bX�%���x�D�,	,K;��"X�%�Oޝ��ۛ�r�i�����Kİ{����Kı/w���%�bX�w��ND�,K����'�,K���w3nK�fJ�n�n����^�m�.��-X.���&g�%9��u�nyMյ%�
׻���ou�{���'�,Kĳ���r%�bX���vq<�bX�{���bX�'���&vM2�wL�n��<�bX�%��wS���$�'*& ��X�^�#�"��&ı3�����%�bX?����bX�%���x�D�jX�'��^�6����s�.��r%�bX���vq<�bX�{���c��C"dK��}�O"X�%�g�}���bX�'��;�l�vL�w4ݻ��8�D�,K��ND�,K��{�O"X�%�g{���K��	�>�|�q<�bX������1uSX����|��{��Ľ���Ȗ%�a��}��yı,O��}8�D�,K��ND�.��~����t���m]����î�%Y�ogk�V�Ѱ��l\�^������I��i�Y�+W��{��7���}����2X�%��}�gȖ%�`���Ȗ%�b^��w��Kİ}���7wi36˹�����bX�'}���O!�(G"dK��Ȗ%�b_����yı,K;��"X�%�Oޝ��,�ٹs4�����%�bX=�xjr%�bX�����y���POF��Ȗwy���bX�'����'�,KĤ;�웹vf2��S�,K(D����Ȗ%�bY��u9ı,N��;8�D�,K��ND�,K��ӓ�e�n���yı,K;��"X�%��}�gȖ%�`���Ȗ%�b^��w��Kı=&^��6n��6�]:�D�Y�W�vv��6Κ��q$	Z�b�/1v�Mwf�l��e�wu9ı,N��;8�D�,K��ND�,K��{�O"X�%�g{���Kı<������7M��v��ݜO"X�%�����!Dc"X�%���x�D�,K����Ȗ%�bw�y���%�bX��r}�1Z��NF���{��7���������%�bX�w��ND�,K����'�,K��{�S�,K�������ZUi2�|�~oq����o�{���bX�'}���O"X�%�����"X�ɫ��@rUP>:���?D�>���%�bX=�{36���&f�s37wS�,K����Kİ{����Kı/w���%�bX�w��ND�,K��{�m7t�#��JI�J�뎷Nݜ@�'���1q�g��7[�9@���V�E��m�����K��{�S�,KĽ���Ȗ%�bY��u9ı,N��;8�D�,K��l;�n�٘\�sMND�,K��{�O!�G"dKϾ�u9ı,O��}8�D�,K��ND�,K���ɇM3rm��6ۻ�O"X�%�g{���Kı;���xB�9%Y
���\,!I
HRB�?z�������ow�~���e�<�*��,K> dO��>�O"X�%���p��Kı/w���%�`�]�����u9ı,O���6ۻ6黺n�ٛ���Kİ{����Kİ�#�{����ı,K>����Kı;���yı,H�����"��|�`|Jc+��4�LH�1X�)~ёH`@��Y�� ċ�!�Z�%.��S�,�UZځXl���e�Sx��W
��\���kE��@�F	�-�� ��sm+KH���P�(@X�8�$�S}T�����	�+�-+4�IFT�R+FS�) ���~�L �F�i�C ?a
<p�ID��$$B��HT0�D�BCA�FP`�l�P�0^�Q�	"�bD���s5!"ũ�G�E�A�4���*(��.$�(B�0�
`J�
���@��ˉ1��D�$�p%�f1��Q�T_s]
cG�0"�$BRD0�����ff�f�wr���5��m �m���9�����0���ԁ5�mQ�����n��`��/��h;<q���m��n���f�#�^n�V)�HJ���ϕUm��x�!E�E�ӝmm��D���,�S������/�~f^�m�^�F��#�s!sQؑkg^خ��#�;�UW(�\��:��Ʊqol�����\1����9.��+�Xsv83�]>z�����/d0�D��:Ŷ5�����uu��ݶȹ�ss��u��q���������b�p�F�q�n��=��i���ơ��i�ڥ���n����]����]@�6��������f1mg�6�r����g��vV��Lef���] =���;mvssϯ�{����i�#B�O,�&��;[X���n�פ륵�r�99ܰDv66�+)��ԧZ� ��d�L��XK����z ��,��c�99׋�ov��qt�lpX{p��U8���E�;	ŵ�3��wV�r�>�5�Olݰ`�+���c���w[��+��m�zZi8��}����jv6�<��P��n6��H���j�t%��u�'��;k��'@��L�m�PPt�ͺ���=ö��ںH)�l������x�� g]���c��mԩ��:�vg;���ش���+�ܕ�خ�1��T�أuM,���3n�mZa��`'�8�|PUc�m�j�wY��x�3�xn��On2ԌU:G�[l�K8�J���.p�����AZ5��k�۷X�6� o(�ݳ��N�<�W\�)^���$�G u��|��5�-n�m��;8<�����m�ӳ�ґEq؀}/v�]�SUt�.���I����okeT���WK�3p��vz0fB�'��}�v�^��7%����b�,����ۍ�W#�Kd�s�����E�i���Q��֎6;jN�ݣAeCȷ9D�ڦ�W�v�ڍ]��/;1���L�䤚�|����UO�?��&���@(���!�����sdݹ��͚l�.���d��&�L:7z2O�rr���y-'=i�ms9���/O9{6�:��\J��h�/�'!�;�͝���nӌ�=s�	ٌT�'l�>n(����mh��X�v��gny$��W�'��]7p�k���/:�L�t�x(p�d�Չ��1l�6x0g��a�%d��v�1��_>|1���çg\vk���v�pg8���zo�?'�b�M�&��a����Gu��\�x�ie��N�mF}ޗ�����Z����X�%�}���x�D�,K����Ȗ%�bw�y�����dK���^��oq���}���_�ҫI���yı,K;��!�?�WblK���8�D�,K�����"X�%�{���'�>*dK�i�fٛ��fM.ff��r%�bX�w��q<�bX�{���c�C"dK��}�O"X�%�g�}���bX�%?zv^�.��˙���'�,K>`d���S�,KĿ{����%�bX�w��ND�,�dO��>�O"X�%�H}���2�w6f��"X�%�{���'�,K��O��u<�bX�'��>�O"X�%�����"X�%���z��xv�Dr�0���=�2��l�l��b�l^�����pm�?5�s��n�
��Kı,��S�,K����Kİ{����Kı/w�ǿ7���{������k3eyLUx�Kı;���y&���Q@P?�ȞD����jr%�bX������Kı,�{����#�2%�����n�ۦ�黙�7gȖ%�`���59ı,K����<�bX�%��wS�,K����K=����]��-�Չy�w��"Y�"g����<�bX�%�}��r%�bX���vq<�bXȈ]���������$.�����ɫ�����*�wx�D�,K����Ȗ%�bw�y���%�bX=�xjr%�bX�����yı,K��l�w2�ə�3���Zl���\B�hm�j�W�ݷ�l�v��=,f�e�
�^��oq���}���gȖ%�`���Ȗ%�b^��w��
3�L�bX�}�۩Ȗ%�bSޟK����̹�anl�yı,��59ı,K����<�bX�%��wS�,K����O�D2�D�)���f]3n��ݷ4��Kı/����<�bX�%��wS�,j*)�U0ț����'�,K���Ȗ%�b{��
t�<3wsd�7w��KϑX'�}���bX�'��>�O"X�%�����"X�BX����r!"����ssvf���ɒ]��$D���u9�O}�MNı,K���8�D�,K����Ȗ%�bw;;��mۻvfm�-����ڻt��>M�+vM	��$;����F�n�uP�n����͙�8�D�,K��ND�,K���8�D�,K����Ȗ%�bw�y���%�bX��rwv[wf�����-�59ı,O;����%�bX�w��ND�,K�}�gȖ%�`���Ȗ%�b{��ݻ.n�ww2K��O"X�%�g{���Kı=��vq<�bX�{���bX�'��|�yı,{���f��I�4�����Ȗ%�b{���yı,��59ı,O;����%�`x�� �Ȝ��7S�,Kħ��e����̹�anl�yı,��59ı,K�{��yı,K;��"X�%����K�q�߿~�kȁmBK��s��ڰ)P8:k����S&�R8t&�vx	�v�7VK��ٛ�暜�bX�%���<�bX�%��wS�,K���y���%�bX=�xjr%�bX���0����6K��O"X�%�g{���>P9"X����q<�bX��}�S�,Kľw��'�,K����{�f�ۓs2d�wu9ı,O}���O"X�%�����"X�%�|��'�,Kĳ���r%�bX��;�6ۻ6黺n�m����%�bX=�xjr%�bX�����yı,K;��"X�%���y���%�bX��rwv[wf���˚jr%�bX������%�bX|��]���۩�%�bX�}�?�Ȗ%�`���Ȗ%�bzǅU� �wܷ�ܗsn�n��=�0�v��Ss�r��B,���S�Q6�t�xֹ��ڮ�C�Y]z㗩�)�HQ/f��ٗ�]V-\'�u�Cv;\`�ָǣ�.��M��p-lnl��l�4�Km�:u������9�f�ݫ��}y��㮸x��u�l���g�˭��+�mv�)�Xw�8��[��p��v^�,��ݞt ����p�9�r�iۏ<V������
�N[���xZi�����ܱ�n7h�s�ܽ�\ 9y���q��d_g��{��{��Թ�=����oq���?��u9ı,O����'�,K��{�C�P�o�ı/�}��O"X�{����o�.���u­W����o'����'��#�2%���p��Kı/����<�bX�%��wS�?�ʙħݟK��m�s7$�6q<�bX��}�S�,Kľw��Ȗ?��,��S�,K���Ӊ�Kı)�æ�tٙ�7m�59ĳ�?}߷��Kı,��S�,K���y���%�bX=�xjr%�bX���:a����l�7x�D�,K����Ȗ%�by���yı,N����,Kľ{�w��Kı;ٳ;a����陥�؃�=�g��=�vZg�Ű�f7JY�8��W7�vm͹�d�wu9ı,O=���O"X�%����"r%�bX����x�D�,K����Ȗ%�bw�����+����w�=�{��Y�����"r���v&ı/����yı,K;��"X�%��}�gȟ�._s������V���Dkow��"X�%��x�D�,K����Ȗ%�by�y���%�bX��y�'"]�7���o�}��J�&U�����,K����Ȗ%�by�y���%�bX��y�'"X��L������w���oq�����e�
����bX�'o��O"X�%�£��͑<�bX�%����O"X�%�g{���Kı<��<ن���7m�6�O`�vsB�B�n������l=�f�a�t���ͬ]b�E�=ߛ�oq��N����,Kľ�����%�bX�w��ND�,K�ｼO"X�%�Hw��4��˛7IsdND�,K����Ȗ%�bY��u9ı,O;���<�bX�'{�l�Ȗ%�bw���xf��ɲ���yı,K;��"X�%��w��'�,pA�E
lM���6D�Kı/����<�bX�'����i���m̳$���Ȗ%�by�����Kı;��dND�,K����Ȗ%��$ș>����Kı>���6ۻ6黺n�M����%�bX��y�'"X�%�}��w��Kı,�{���bX�'��{x�D�,K��q�����.�%��]�.1ӊ��ƛ�����bCڴtd�]�pݸ2<�Z�j�Ҡ����oq��������yı,K;��"X�%��w��'�,K��{͑9ı,N�{���-*��V�{�7���{��7߽�ND�,K�ｼO"X�%����"r%�bX����x�D�ʙ���.���u­W����oq����߯Ȗ%�bw��Ȝ�bX�%����'�,Kĳ���r%�bX���izl��s.f�3oȖ%�@ȟ}��"r%�bX�����yı,K;��"X�U���E�/�;��>�O"X�%�H}��M2�3f�.l�Ȗ%�b_{��yı,K;��"X�%��w��'�,K�M����)!I
H]���D�ՒM��Y�G�k�[���[xn�kz�0j�ɇ����7s�uU����w�����d���ND�,K�ｼO"X�%����"r%�bX����x�D�,K�z^�4��nl̳$���Ȗ%�bw�����%�bX��y�'"X�%�{���Ȗ%�bY��u9�ʙ7���������e��*>{�7���%���sdND�,K����'�,~HdL�g�}���bX�'��~�O'���{��?Ϯ�X
��H����"X�%�{���'�,Kĳ���r%�bX��}��yı,N�����oq���~����kLJ4�Z�{��bX�%��wS�,K���oȖ%�bw��Ȝ�bX�%���x�D�,K�M	�÷����d�G]��/^jm2�E�����e^:�6�{@Q��WFu7�`0�{pQ�0��b<��b��j�ke���+z�{����ܑ.�t]�p�����B�jÈ����;�Ѻ6���yZ8x�{l��q�{sӂ�.���j�4�IJ:�g9��;^u�0�7V��G	��u��'1ѱ]Kk	<
�Ʀ9������l�����޷� |�~�<?nYd�a���a�4���{�������;�nƵf���֜�q�6�)�wrLɥ����O�X�%�������Kı;��dND�,K��{�O"X�%�g{���Kı)･���̹��\ͼO"X�%����"r%�bX�����yı,K;��"X�%��w��'�,KĤ;��e�ff��.l�Ȗ%�b^��w��Kı,�{���bX�'}�{x�D�,K��6D�Kı==�I:a��wwd�n��<�bX�%��wS�,K����Kı;��dND�,�?}����%�bX�'K�3Lݛsfe�%��ND�,K�}�gȖ%�bw��Ȝ�bX�%���<�bX�%��wS�,K��PC������B�/8ϫ'nc7Lym����/)SD:{9�uE��{]�Ӡ�;6\ݞ'�%�b}����,Kľw��'�,Kĳ���r%�bX���3���Y�Y�Y�_b#e�M��nЬ���,Kľw��'���blK����Ȗ%�b~�y���%�bX��y�'"X�%��w�{v��۹�ws&\��'�,Kĳ���r%�bX���;8�D�,K��6D�Kı/��w��Kİ}����7wrLͲ�fn�"X�%����Kı;��dND�,K���x�D�,K����Ȗ%�bS�����ܙ33vKsgȖ%�bw��Ȝ�bX�%���<�bX�%��wS�,K���y���%�bX7�N��ɘ���97G5�x�쵌�Ͳ�tE5�-:>�]d�b�\𛮹.�ٶow���oq��﷉�Kı,�{���bX�'����� ��2%�b}����)
HRBi�UD�WWvwy�
D�,K;��"X�%����Kı;��dND�,K���x�D�,K�z^�4�ٷ6fY�]���Kı=��vq<�bX�'{�l�Ȗ<(D�x�vH0�!8�z.W��MXT��x�a�+�x! U�.�S����	<&�И��$!4Q4 �@���A*������T�Q��! � r z�X�`�G�@`�Q�� 5��=�@�LQC�=(��:���� ��N ��0N���@8":(.�DqUJ���UQ5ES��ӱ?D�����%�bX�{�wS�,K��Ӽ��wI��晻�svq<�bX�'{�l�Ȗ%�b_;��Ȗ%�bY��u9ı,O}���O"X�%�w7��T���f��|��{��7�����Ȗ%�bY��u9ı,O}���O"X�%����"r%�bX��S�:A�a'�#�]^^�x��3�jCd�ِ�A��v���8�)i�Z�&n�Ȗ%�bY��u9ı,O}���O"X�%����"r%�bX������%�bX>�{�.���&d��fn�"X�%����Kı;��dND�,K���x�D�,K����Ȗ%�bS�����nK33vKsgȖ%�bw��Ȝ�bX�%���<�c� �"dK>����KĒo8�_�R)�JnDժ�VUYV���^�v��	#��9ϗ9�s�RM��9��j�><m����^�$t�$���k�'=��l�MZ�v�vؓ���^n.�Κ���t	Qq��8����:��9rmf��������'�I4�נ����֒l1�7�o��H��� ��u� 9���m��i��X�0�G���H�I4	r⩦<m$�i
�o�_U�}�<H�`���<��I�m�Hui$��$����@;mz�k�9�ӟs�,�
E��D��{4��ɻ�]��Q�ی��6	��gI�[p$�[��Z�ꊤF�F�sR���>��g����nֈ�	�
��uN���]��#�s^���= �:�(�t<�k����5�����loGg���K�2��<	���7e�aۦ8����^�6�?�|��Y񇶈�}�	���Pv�!�K�.wchUR���k�/l;��,hͮ���Ϝ�s���޽����OUػLz�i��.�7�gghp�nY-&v�^L�]f;s���ʜ^�C)6i�}�� rH��G�n� T�,�N��bLL-3 9$x�k�$����@���5x�O�6��m�m�@�:hGM ��]ڹ��N��%bm���I4�נ����֒l�ٍ�6�H��� ��GnE:M��M$���Ӱ^��m�;��R��z���$��%���J��� 9$x�#�7u� ��b��cM�I��!6��G�~O�?EOU*��?�O��� Oߟ� ����m���$:��m�u� ��=v{}�����e�Ϛm]�&��3j�\� 9��z��C *W�ez�	�-10�f�_Z��נY4	#��9����&m�+���_$��6{VB+�����5����[���^�����>u�Wh�@7��� ���{�X�y��U���;n��m�u� �� ���$�=��g}^~wvح�7M�\�ـ6� 7xL(��	J�� D@�]TM�! H��"#��-�����7��`�c�&���&�J��� 'dx�#�&������ �^�lm����I+m�����G7�~�|`�����3�1l�S�4���ˇ�d�Rmpq�l �:����v�u���N�!n�v]p���&���;#�}_r���'���6�I6i��g�ꪹ�������l��r&�jɫ*�j� 7x��xt(����������|i�>1&އ�����EV�޼��� ��f�!ZQBD`N"���9��y��x{�{��N��%bm�u� ���}$� ��� 9$x�H�S�m�V����4iD��n�a��cL�z2!tfA6���ɉ�m���_U,�x��[����v�8���	� rH�	���F�I�j���IWf ?���(����n��7vٞ�B��Qޯ�����U�RV������M�w\0vG�sc�i:m�	�$�x�ﾪ���� m� �n�9(��3�w^ &�T����ZM��f�����π��o$�����JEϕO{�)����e��8r�kPSu�����Ӯ����9U6xͷDm�j)SqXṒ�\�^���+�G	��)c���\�:��醻O-�:F\�=���9�<��A�A�lN�������`؃��g<���d���ݒ��^�8�)svHܕ9CX�ø��V��J������ƨ�����Cgi�,��0�N-��cu�X���w���iܨj�qѵ���4�/S��^v#���Ӳ��	���g�>����㎲��t'L����<������G�Y4	#��9��j��>1&� ?6�?��zD%T{��`�~0vG�����앲�؝$��+[o ����;#�I�Q�wm���鶝��W�_U�3� {}��ͻ��%<�q�|��j��f�4�f N���G�M�wm��B��_R��T�vU���4���l�7+��[��Ѱ���yJ�Y#)���w��W�ڦ۴���Z��@7��� ���{�����xg���t�hMUU��vٍG�	B�	�a//�v< �窪�*O]_���V]��Zf$~0vG��<n�`JnDբ�Y5eXMY��
g�����xղ�=UrL�J�N��5v��c�]���G�~�s��$�� N��m�����9[�M�����=�g���(�i��uNZ��������|��>7��V �� �S׀n� N���G�v��M��x�x�mhGM ���$� ��^z����ZM�J�]����ـwu�����_�Q	���!DC��w|`�l�5�T�i$�*V&����x���7u��}�U�}�<���i:m�	�$�x�`���< �������|��e��zYS;�6��ez��4�SVm��&9�ָ�붹�.�2`f����@;mz�k�$��R���:�Zbai��#�~H7����~0ݶ`�عM]�ڹ�&ހv��	#��$t��^��ݫq:M�Ӵ�Am�n�`��g$�����D�T ��S�;�}ψ���%�u��i<m���ـn� �DBJ{{����xݶ|�}�?I��r+A'�xr�L7����YmřѮ�l���]{<�4��D���4�4�נ����I4�+�퉶�&��j�x�#�}_B^�=�~0� �n�СD����n�m+���Zm����7u��]��y�}�< ��ur��M�v�i�P�[y� v�^ ~m��'��0�^���t'L����0vG�m� �m���0�T@�B�F�		$��d�=�Ձ��0"��D��Q�� G�F0�`FI�+`�	�H@�a,�)D�ai�Q�)4=���� �
b��0"!�[T'�	RST�@�(��(�F���t�cGP��!�x�*$�ӂ(� q	IRZƕ+�� �p�FX�l*PaW�O^,"���gB,��+��`��<@�,pBH�'j�D;��*�C$�BE�E��% �1#$I��$`I$�1P�QbPphFH0#���H:�� �0!��b$a!$"��A�#(@($�ь�#  ԕ�� H a!0v��wm�e���*�,�c[T�qtl�1��`A1,hI��@6��y:;v^�Tv����u:�p�c�9�]�6��ж�"b�D����l;�8S�H Ц�eݱ��)T�gr�*�F}N�pɶ�Up��ry�UbY�e�"�n��m�W �rv*j�%9n�V���1iZ�s���^���[lV���vˎ��u�t�v̺��$=bx{Q͗�􁝻�W��M,tpd��p��Gd��vG��v�usN��i���le�eܾ�(.��0(��d��v�V��3T7dm#���*�pW=n3�j�Y����I��nYum�h�.i1�w9�ּ����9z��[�bP����7\�`:m�{��u�lg��tl�s��l�tM pu멥�ܝ*iձ�喷�m��S��v�7�L���-��[�هF�mq�=��*�<,��<��x�[�:�¼n3����vN�t����=�.�kg��1\b
퍲G<��kak�k�v�ʘ�z�6�t��exg�Ӹ}��I×;Le2��8m�J��������\.���s����I�]���v4����򽫥yZ�f��`��#���^m�{X�8�*�J�' I�f^����Γ�N%�wn�����%U���;�Z8t>Z	(w<�jv�-Y�W%�k�Cۣ���1���Mr��j�B�5�����%.�[puv!��ź��L�@S�s�\�Q��ꜰ�2��u�O���\]v(�*�
��@��p�5Y�g;l�qہ�f��;T�J`(B
Ƶ���]=���a���vd6ے���k%[ 4v�#�F�n��]6l��I�ɻt92\9�H�ӷV+zw��a��ܰNv�%ڳ��)�K��-Ʒ<�G�ͣ��#�^�[��kvU��X]�)��u�l��1�V7^5�4��	�rT�1��Mg�\��܅���l�9{��4�Mx�FY�jC\�K��hݗ�b���e囈ba;u��&ӭS\<p{��������P:3�����^�����"p8�>{�����s��p��<2jI�kql+�v��뇭�x�Jp�\5)�\ݯN2=���Llk�'(�v^�u���d�[���t�ͧ�;v�-�=f��J�q�˞���)�c��I��v���VS�2� !]��fq���<��h���,��W�e,���(Yۊ��nNܗF���w.�kX��ڋp=g<��[g���K�ɸҞ�������6נ(�.��9��dz���u�>�-�p��	�ф��|��\�6��X��$�����,���p�U}\�=���%l�~N�`�IX�6�#��$t��^�v���>�w[?��O���hqrb}$���~��ֽ ��GM��X�6�ˢ����IB���� >���7vف�(P���`�uqsE]�MU�R�����^�dt�$��}k������ɍ��MF�6��g���H�� �؉�G�]��^�ꃞ�������~|D��+���Zm�H�`���< ��$���x�m�,f�$vr�C��� ��q�}�o�?o$�~��M� �ʗd�Cc-�L-3 �� ~m��)�n��w��6����ؘ��e�o��]����=#�n�꯮����%l�~N�`�IX��x�p�=��<p��< ��ݶ�Glv�m�m&�6P�H���o-��4�Ӝ����l��Y�����.�&�7i�� �� ���$���W�����?���~�v&��hm5n�f ?������n��7vٞS#�^^wh�ڴ��I+m�}�<n�a��DR!���>s;���y���n�m+���Zm�tB�Jy�� m� �n��n��e�)�i�;m���w\0�~�y����7\0	}�M�4�����s�%���-c9���1jdm�4tk�~m|>�����Z�v:t62ۤ��8��� rJ�#��$t�'�ǜW�4c1��$���^�dt�$��}k����U]��U�'I�i��Am��?��0��Ty�׀�z��;w37M��ۦ4�l��rL��y�$��H���P"�x#�y=��0	�&S�4��Ci�v�0vG�r� ���`���"�M���3 C�']!=N���ڀ�.�m�ټ�����M̚�qR,/*U���{� ���`� ���t�i]��BM�n�g�ﾪ��H�`��x.H��e�)�m���Zf�$t��^��m�����vJt62�L�	� rH�	����� �Jj���ؘݺe�7�����I4�נo�~{������ܺ�b��[/c��Ҙ.��t	�.�%�ɟ, =e�Ьl�[�cl��˞#�OY�˦;F휛\綫�'r=t��p]����Q�[�9mpZ]��=�c��6�vs:��(�t\q[n�+�l[/[�8yY4q���n)
we��Y�cNv��H��7=�ɶo�қ�MӨHz�S��j�#-�6���Iw7f�23M�_���t��g�ݧh��c7;U�03�N��sVG4���;��S�7L+-�g��`���?}�߽�w�~wv�'V�tƙm��g着���������=
&O��䫫����ջm����˒,'�]�07u� ۣv��һ�wWbI������� ����;#�9#%���V��	6�	�e����I�8���˒, �ԡhJ��i�B�[n�W&�J�Q�%��^�5�^��l	J��q�B��`�w�n� N��\�~���(Q���Ӏ	�zd�U�&�U��4�ץ����s�,<���vd�@�og>Ug}�7�K��&�-��I?_��M[/ �� ���ݫq:�˶�Vӡ&�=_W�}~�z�	#��<�$X%GݺIն�;�ӫ�wm�DB�S����{���������O�\2P���u�<�:r�������Ͷ�*�o4�DYВH�]Hr�ʭM[�ـ�<�$Xղ���_Wܰ�?����[mZM%Jն��۬�k�wm� �n��!B^��RF���֛M%i;�k ���ׁ=�����D�"qDx+���n��c�;}�X[�����v�`��p=��-�� ;{� ?6��OG=x����S�v�6���<�(IO�����wm���ӻ��렇<�������Y
n
��e��&[m^ۂ���K�p��p؋���6���u`�l�7v��P�H�׀=j�G�����I�n�g�����#� >���?Kn��!z"UF����f�N���ݶ�� ����#�9rE�n�̈́�v&ݴ��jݶ�%	D���x��Հ}�l����(�!��� >����矾��}��ڮ���I�T���˒,��W�}�節I� �����Ҳؐ�+�sQ�-,�^��RiɅ�i����[���#M[���i+Iؕ��7\0�p��w�!$�Hwu���\�f���˴�0�p�	� rH�	�l�B��y$�P'���®.j��Zf ~��<�$X�p�7u� ޚ��Z��5w4Z�f��9B�J~��y���0=/{� z��Q�왻����U]`=�`����$����> ��^�[u�}�

�(���a��k��.��s�òhw�Ds����g�&�H��s�6a.Jd��lh�=i��WON\*S�����nq������(9�ͭ��gK���K�e�m9�*c>�ڬ�,q�¯G��`v�.���\k�l�'n���h�nă�nܕ��Y�Z�r�s��n˩r��ֈK�8옴��x�O���Tq{�v�杰n&�e�d�+��9<�rM���r��x2t�m�V��1vyئ���ә�/K�ǳ��n��$��n�Ӷ��_� ����ۯ%	%�A�|`>;�Uv]Z������0�n��!%2}=�Xn��7vٞ��P�Gԧ��UM]UU]U*�6�������`$� 䌖�M%i;���;��n� ~���BJg�� ����mU��M��L�7u� 9�< ���p�&�X�B-R��mN���t�;N�e��<b�]8vm)sf�M5����FӖ�&?��4���y�$� ��꯫�XI��J�ߩ�V��:ai�y��y���"TF�D?�x?���>�0��y�P�F�7Tr�]����$��?�a�ꪫ���x�{� �v�7wn�e��1�m���0��x��x�Jz%O��� �~?e;v����l�엀zO����w�����'��P⚳c�a��@t\�n����n9+;�8��J�	=���Z;����|x��¨Oa[o����vk��������Zlm4���J�o ���_}��_�QTwu��~�������SW3ht;M��L�7u� 7�<;U_?�_���8C�D��ȡ"D�:k�DR�c�@�}���*�bE E�D�0A��G�c�F3�<`H�bB`�H�d�(��ł��8�|��	a�1�� 
�?b���\���#'|E��P�Ą�x�'��� �P�D����L��P�PuDU�:��og���䓺� �i̍XU��Z�	�09DBQ䒪��^ o���>{l�7vـ?�R\�wrU���d�]����IG�D'����;��`�����S5qE6�f�ٞ����a�Վ{7m�s`zwV�u��ɰ�uՂ�&��m�}���n� 7��!/�OwV�.��3tӻi�m���w\0{#�9rE�vk�z�������e�;M��C�ـ}�r� ��w\0	\����[TZ���꯯����7��ӒO}�{9&�@�ׂ)�#��uT|�����'{��7f�nf\͵t�k ��w\0{#�9rE�o��������ߒi2�At<\��vL��^�Nc�6�ͳ��6�]2]��٦�f�0�P9y̧�t�[��ڴ��=�?� odx.H��p�
�w)���I�Ai��7yСL�OwV��wm��� �6�Lm��i��$Xf�a��#�}�n�۴Jl�m%m:*��=
!N��0���w��������ת�Ӥ��t���f����/{��OwV��f�D-�w{�߿_��gt��nx�����"<d�6�S��7n٣)���gh�A�P���A��3vzI��Tٶ���!��`�^!��[�mu�W%�t��D�Мn9As���fԎ�
GY����MWv�<Y�kǜ��]����e,[�H۷Fy����N�f݋b2X�m�o\��mm��e8�#ԧ���9�(�;m:������繏��5�T���6:�Fx<W[���m͙�[ՓgEױ���=��-�jfmO�I??_���U�4H�I4s����b�v�M��$Xw\0�p�l�?U~�#}���m�i��'j�&�=��n�)���x��Հ}-Ԧ�m���:v�&`~��&x��y��"�;���R�S��鰴� ���UWW���6G� ��E��v��'���]s�kl$�k�<f�n('x�͒�EхY�7Rf�]l5�m�m��:hGM ��r&�[�m���wK���'�}��x
0���(�!(K�]
>�~�0�}x�n�����'��cM���@�:h�n��
&~��[�0�ǖLҶ��M4�m� 9�<�$Xw\09DDKo8�;�Otܢjɪ���IWw�~��`Jky��w� ~��o����&8.t��Rt�6y�딎L����Jڻ=��jQz��m�&�˕�t�k ����͑��꯫��{� ���z��C��c�i3 �� ����[u�}�lΈ��d�鞦+O�i��i���<�$XUW���}�|/H�vGM��@�K8�c����UU}}^���?�`~�����y�T�~vӻ��Vӡ&�H�I4�נu[s@�&��`�%��μ����T�݈�|�6�(��v���9|����{�>s���[4�9��$~0�#�9rE�wu� ��c.�4�v�m�f sdyﾯ������w�����#�S�7)ڷV�MQbm��{� ��?W�U�ܑ����x�5-�m�i	;WI7���@�:hm�C�|��9�߹�΂�¨uQM� ~Uy�w��E��S-�Э:v$��n��
!O����{��ݶ`~l�\ѝ�.�������u���H�������&�WF���B��m�ߛm�X�m�����BJ?��%�w_������;n�0��˒,w\0ݶ`����CeO5352	U�l	#�w�F���^�ͨԲӡ�v�&Ӵـn� rGx�m�B����`>;,�WU3r�7�M�@;mzU�4	#��$��I4� !=7�ޛ�]�se�G^F�`���z�	D���ή^�*D��Ϋ��Ӆ��9L������+GY/^HtZKx��ċ45��:;n����s�nqQz9+����&�N7=��'��F�;sx��c��,u�.[��mu�-�f�������[K�.��^��m��ҺW!�k���d��jp51ۂ����04����7)ͫn6v6͉�W�ez ���Yz�v��u�C�vn��ٶ0����%W�n�cC����G�/�t%�e�,M����n����#�7��m�m;HIںI��n����#�9rE��ꫳ|�h�2�*j��UV`�� ?6�DB������,H�`vT���m���0��P�/D(��{׀l�ެwm���4	�q�lYƛO�7�u[s@��w\0�G�muEBT��;�n�������Ơ�ۣ	찅Zy�rи�&^��G_���|#�Lb�"��������	#��v���nh��*q�4��ۛ��O}�{9�P:���n�_�������6v�'V�o�f�v���nhGMHـk�-�ʹ��5%]"J��(�(�����{��w\0�G�ocDm�]\�W5*��ݶ`Q�!ww� �߿<�$X��Dm�t&�M�i�]eX�.��g7s�&�Z����n{`�J��ӰV��I3 �� ��V��$���
���617̰�� ?6�9(������w���zo�NSe�m1�M��"�=�������UMO�
@`��ET�*Evz�tO�Z����~��n�۸�e�v�ۡ&�?}{&x�$�� sdx.H�mF���6�Ӥ�l�7u� ��}�BJ�����{Հ}�l�6X�[�(e��:�nָ^��nxv:�9�GIubpzv��g:H�T�[wge1����~�� �-��>ݶrP�~�m�u+��S�n�X����9rE�wu� �� �����}�}vM�G�v�v�Zi]$��6G� ��?U}�U���<��y`�Z%;����ڴ��n�f ~�� �-��؅	,"�	yB��	}�K�
!}��� '�L�]vX���c4�נu[s@����m�߿k˓]�����K�p�Yn��F�.�7òػf�3!���u��Xz�:ai������`���������<H[^N�N�[�BM`ݶ`�l������Y��L�5�^�RliZt�CM����l� �����	��HN�i�j��f�%3������>ݶ`z(�rg��U�K�;�ZiU�6�\�h��@�:he�@\߹�}s���X�d
A������!�!  B@��,HB	S(�X<5�3E�#X�5�V�i@���J�H� �0#�iG� _:�� $o����0 &�,h@���K�#q�c
��2���
a.K�LMF\� �H	��@�A�E�!Rb�,X���B, @��"��p�,XD#����M��I���n�0�9Y�[��0q[K��B�4jLr�T56ήv,Kl�Ugu2�ÒPgU��z�.=���&iz�Tb�C�%�c���vG�I3	�d�%�W��6N�,K�<�a�^1̻�;u��!��#�K��t��nM�:�-�R%��}��Z {um�V��ä���6ۡ�a�q�8�.��Ц�NI#]s�T������C-�2�ZӞJ��{XɎW�)`zZ��l܉V�Gu�`�B�;6烀�n�cB��e4 �ۮ��lٳ�k�%\v��L�]m��P� ����N1���pm���T�J�scun�j�m�OQ�/6Y�*�U��Q���Y��k6�2Z��vo;n��iv��kD4�8���=mk[F��7v�ƪ�f�5"����v�[V룒n���cr�aqrjn8�n�]u⢤t�n!c�۬fS5���(e2-�^�n��Yc�'m���7WiL�#��9ݹ�ݲ1)��3n)HO-�l�
��Tm�]NN�9���hɸ��<7:��{g�����t�K���wn�2<��ڹ�<��^��$�z��\IvW��"�m���b������p\��94�!S���;���z�v��c�y���va]� ۂ�=���m���牞[�$�m��ʩ��sX��z	�p�y��ؐ2�2=*K7�s#&�kc5�ѻE7��h�:�i�v)�
U'�cn��gu��Q�	㞇�c����W��g"(����T�O��������l;�µC��it��lLAk@<�U�Z1;���\`;���Ō�����)����m�`�dZ��מEF��l.SXv�ػ(]e8!71#�<�E��۶�t<p&�8�E:
8�1X�78鷍Q�e�����M�V�sn�X�b�t�:{8��)�T��wN��[��vݳ`y�4�x���[$�p�Uv�n�e�������s�^��;s�-iK����9@���U=D檜��}@(q�:hpF��C� q^���AO9���M�d���92���E�\�\t��`�f8�K��õĽ*v�ckkm���=S�L���k<�B�A�A�^�٨�<f3��*��r)b������b@�Mj^_<d�ŗ-�F�;m��΁{]XMZ{1Ɠe�<hd�y��f��ɷ>xc&���m���!��x��u�]n1�:�uY"x��$��F��#��h6�92�n�
��]���&ٖ�7��f��[��e��
�;`Ѥ����n�q�e`J]3nիM+��]��w\0��%�I%Pl�ެ��4yY7w3S5t�ZL�7u� 9�<�$Xw\3�BQ!Þ��tM�dՕa5f |���:���zGMH�_��xؕ6�酦�?}�}��{�X��`�ف�J���^ �&닺�&�f���I����`6G�r� �>�g�TZ˥kc�����7�E�@���NL�ő���zlOo���������7R.�hi��I� ���\�~���#�vx�2�!:N�M��l�l��ь�F H�I#  �X$�B F ��P����Հw�l�7vٞP�!U��*��V�+v�.�o ���Xdt�$���k�'�¶�6�,XҺI��wu� �� �ʏ�_}_U_W��o���vۻwm�ē0ݶ`�Ӽ��� �vـz�\���s����t�'`痴���6^���ح��Վ�]!��i.��
͜����wfK�&������\�`�����a$~0	����6$6�:aj��9rE�n� ��f ~m;�B��#l��vӲۻM[��X���7u����D�@������I���s�9�v�����I��6`��m;�?Kn�<��$�*���0��.�$�ݶ��v�0�Tx.H��p�7u� �بv���V$�+s�[t\,���ŵ��Yݏ]yyb�(uͳ�w�w{��b��cC�v�H�N���{� ��w\?r��^x�4y6&���4��m`��n� rJ� ������������*)[|�}��� ?6����S?OwV ۾0�2�S�"�V�� �˒,	��g$�C�=UP�E39����^���6�:aj��9rE�I4	#��v�W�ZeTY���&��jI�ݙ��������;�D��фg�WlܯgM�&��P2]�~m�o��ݶ`�Ӿ���C����>k��j�N�V�m;M��g��ﾻ���}=�X��3�B�D*�{ǲɚUV���m\�ـ�/^�[u����e�~0	#�lU)V4:�m4������ ��f���P�G����������lM;IZi]$��7u� �o8��r��?Kn�
�����"$��=ٻ���˶�2ܷ�����)v{s��a��9^˓��WJ����Τ��٫8G-�Ԡ����˨-���']�c���nk�l�E�v�m�^c��ۭ�t5[�؞�uėIs\�0����ú�v6]���a4������&���:��c����c9�P����娯Y���n�o�7+�R\���nv<=���sm�]/F�����1�Kxn0k'�n�	���s#��H����tv�GF�:�l��8��d�v�8�!�D���+o�o�߷�`�Ӽ�����A�|`zg���m�vZf rJ� ������@�'ˎ�g�>0Y��\�`�ᇪ��� wޯ<wKj�c�ӻM[��X�`�������}^���^~v������N���7vـ"IO�˯�OwV����m���'�}@�IctdN�Q��b�OO75�IK�.���]���K�����ӷN�f rJ� �����儑��'�yR�[�n��m!Zt�˝�r���8 �TMQ�L�w��'���0�Tx�4Dؚv��ҺI��n���~�;�W������-�ۤ�lV$��n� rJ� �����w)�6!6��i��y^��m�H�I4	ro��׭H����u�V���klgMvշ7M��8���9�Vs㛫.�.�.��ۚ��@�:hm�z�MR��i&��i�w\3�]�G� ;�W�˒,�Q�i	�j�6�w���O}�{9$�w�w�����|*��W�Tsm{� ݏ�̈́�]���m<k8�l�����nhGMH�lU)VН'i4�N��9rE�I4	#��v�W�Nb��xcc-�.����G!�9����vz6��(���ؓjY�C0��r��m�~��w�7u� 9���9rE�v)hR�ڷN�Z���n�v�û)09rE�s�G��꯾�m˹M&�����i��y��V��=#��$t�/��NSbCI�[��=��_U�{�X����{���=��h�� $+����UWّ�q��-�Fݴ�V�X�@���@;/+�:���}�?Iw�$2�P;�=��V��,�Vͳ�\ܤ��J:M7��{n��>v���;�g �?��˒/ܰ�G� ���eګN��M*v�0{*<�$Xf�`�៮�yW�y�Н'i4�I�xo���;5� �� �ʏ �ƈ�N�V�WI6��p�7u� 7����}��{�X��B�[�n��t�ZL�7u� 7���9rE�z�Ms��8�*O��X��������vc6�����/a�s����p�9�i�cb�"6m��s�s�fv�9�=Xb�٪3��q�2ͮyv#kN�K\bp�'��8vӗmہ��v�4E���Ǟ����v�Ps��۩�\��Pyt�l٭fѰ�|�~|�qm� �����9�8��,�Ȼ=q����׸��'��=J�9��e���w�mV�}�N����r�/l"L�f�we�s��n#�۾u���}R�iȅ�L�d�jπ9�z��۬���P�H6��O����!�݌�T�˒,�:hGM ���@��x����M]U�j� �� ��fԒQ�Tz~�� �����9*LbC��v���M���@'�+�:���z�M��v�ӡ��J��� �ʏ ����脣o��|�_�wm��ڧ7USVg
�:.�7g\D=6յ���a.��v�J��dM̚�Չ��,������>Ȱlp�7u� ���X�4Dط6�˛�l���'��{9�B��M��(�W �T�D�C��Q���0;ܫ Ss�Q��ꖅ��:wm�դ��?ou�ÔDDL��t�>�0M�2���4���e�`~���Rz��^����M�t߮��ćiۦ�'K ��V��]4#���%�h��+*��،�;�8km6�9���ūT�zn݆�p�Ń�����|�<|���"E�|���7\0�쥀N�/ ���$:M�i�i4ـM����`�np��СL�w�LҚ�]���+��0��V ���[��	x�P���M	B��;�F
Ĉ@!
��	��I����(B�a@� �"q3x��C�+*����))
"�*h�v��¦�D�F�<"d\fE)�M��a�,Bp�)� ᤢ@����9
����HSX�e��8D� 
c
-)&a�̠ɊB�'�XIHIQ�T0���VYp�X̗)Z��P��P������Y��W��Q�	�qP�Q�T���>&(#�P=@G�����P=9�<�:芟�P�c{�w\0H�*l���NҶRI��'T��oc�7\0=U_^�OR�&��ɱ4�Z�ڻw�oc� �m��������I%�K��S\e�6�I�ʱ(��PŰۃ���<vU����&,��b�
ȋoͷ�w���X���D$��ϯ� N��M�jݖ���Q��K�=c��dt�;y8��6f6���� ��� {��:�S<���^x�lj�0��iX�w�������7|`��x�_�DrJ;��������]P2�o����7{����N>A���芆}���x ������w���A�666>��}8 ����}3m�ܻ���2��3���ez7/87I�.�h']1�CM�ŵ�f]7v[��&��ۦ�ݜ|�����o �`�`�`����ׂ�A�A�A�A������ � � � ������ � � � ���a�733L�r칚n�A�666?{�}x ���&A �`����8 �������lllo}��x ����7&nm˗7rܻ��� � � � ������ � � � ������ ؃� D�A�w���>A����;���|�������Y�6�n��33g �`�`(�?w��pA�6667�~>�>A�����ﳂ�A�A�A�A���ӂ�A�A�A�A�{>��.n�wr�6pA�6667�~>�>A���������?��`�`�`������|������>�|�����A�"�����?�L�4�L��8���^��ruh�p�x'X.�G]�#\�ɺ�9�x�8��s۝�,�8fvV8+S��띛���\7W���!�"�Nv݌�]�KyP�۱jI+Eѧ+N��m�/K��3`��v5�?6�����í<i�e\=X��Z ʐ�kkyݍ�6�4x�p�du<;(��R����]� �]��ՂD.�o������|����4���B���ȥqUvd��2f
����8�Js���n�f��ݳe�n�A�lll���?���A�A�A�A���ӂ�A�A�A�A�����|�����ߏ���A�A�A�Aｳ�g�&nM��n�]����lll~�y����lll~���pA�6667�~>�>A�����ﳂ�A�A�A�A���>ۙ4��nm���ݜ|������>�|�����ߏ���A�A�߾�>A������N>A�����O��n4������ݜ|����� ����?���A�A�A�A���g �`�`�`��{ϧ �`�`�`��{ϧ �`�`�`���p�ٹ��f�˳34����lll~�~�8 �@���ӂ�A�A�A�A���ӂ�A�A�A�A�{���A�6667�{��6̳����qR���;/^�.�-[�P�Z*�q��o�!����3��F�F~w�����666?w��pA�666?{�}8 ���o �`�`�`��{߳��A�A�A�A��~�3��7-ݙffl���lll~���pA�#���
� y �`�s�� �`�`�`��;߳��A�A�A�����4�ߙN�V[jݖ���Q�~�Xz!D)��|`���ը-��i]]�Y3j��(�B��[�� ~��M� �ʏ ��U&�iX�V��;5� ����/�,6߻���۪-eК����	�vm�a�\t\7Bp:�BA#���X��=����t���5���&�M��?��/�/��,7���;��]���v�v��l��N�(S'N�V����3�B���yו6;I:nҶ$�7�z��Xf�`bQH�����0�x��S��ӵj�j�[k�׾�� �� oeG�K� �>�t��b�i3 {����{˯�;�X�m����������6p穘�л�痴�������f�7��G^.�&�mn����g &���	}ذ�p�'u� ���Se�m��T�/�~��&M�|`�����x�l�Rj�4;J�Ҵ�ٮ�`�Tx��X�U��lM�����L��_TB^��߼`?/^ ��u�0Bq1�$U�
�pS� S=��0vv�'V�i�M�� �ʏ �݋ ��w\0���Zeg�UV���c�6�m=�	Y������;7dA����.��hV���W��������p�'u� 7���;��DКv�Zm]�m`��N� oeG�K�ŀwU�b�]�j�:V�&`�ـ�N��%=:���|`�̦;M����f oeG�K�ŀvGM�:h��x؟m��7�9�]`�-�~���4� Q� ?Q"�"����*٣/6�r��n��Y�v�r���a��Ђ%J�E:,�N��;�t�+�s���h�N��ɳn��fƁ�t�y���<��<��;M��lF���&�tq!v�psc�\_���|�½�g�����m����X����	��j�ڭcs;lT:�)�r���I)Ts�s{8V=`�q���:7jαVnbێ��ll�feٖL�㊦�������d���B.t�3��&�ۛK��ݧv��G<^�.�s@jLv!�n^�����m����4��ו�z\�'�����bv�3 �� �ʏ �݋ ���v�ӡ��J�M���/�ٮ�`��T�;tյlI:o �݋ ��w\0{*<���M	�jզ�ڶ��4��ו�z\�=-�3�&�9�ɠ/k%��ݫtv��/�q�rV	�]��7��
ȋo���@;/+�*���zGM �JS���mL�l���}�RD�.h��@�����^6<m�hY��
�.h��@����y^��u0t�S���m5�wu� �� �ʏ �݋ ��n&�Nŏ�h��@;/+�*���zG��_Uwf*G���i�Յ����ѯK�7I,ɗ�����@���u����]����f�=i��i�M�� vz��	}ذ�mr�lt��TU:I�Wn�X�7����4	�������r%v�;V�V���;��ou���� DX"p�z6w�9��O��w �W��]�+V�0�`5�x��P�%:�q���<�e���mL�l���c�;��ou� �i>T�wmSj�'M��Nu�cG��bi�Vz-)���7eG%���']Zt�|q� ����@�:he�z�G5><���1�6�H�I4�� ��׉�x��v$ձ�f��͕ rH�H�vR��,|km1�٠�;�ͻ�>ݶ`rIbI@�(DD" D*t� m�|�rI�����>ccĚbX�ށW���:hGL �ʏ 7uEWM+E�ڻ�I�'[f�M�G8�U�9��+�]q�Ӷ,�k��vjL�"ӧj�j�[k ��7\0�*<_dXb��S�t�I:IZL�,���y^�W���:h$*R�ۤ��M�Zf seG�K� ��M��^NA�^6<m�hY��
�nhGM��������5>5�i��bM�$t�,�� �i� ��� ��,ID!@�
��� ���^��O�F�(;� �f(R�B,��$��+���0Ȳ!%cP�����t|XpI���	HDe�,� A�����T�il2���"@��)*CR#� �\C��Y
BB�l8q�2,$H�$	��80���
�:,��B�J0� @�
�H�ёe%�	�� �b��R#!���C ���P�DǊ��`�LiLĄ���!.&� �ڐ0�2aB
j�~`Ԃ�U<0Mq� ��B�*��$"�`@,���A `<Ԙ�7�B�GT%�Jw���^���3.ir��i���lXy+v8:(�KHT�R�-��\�zթ��r��i��:v%�wTm��zX熍@�^}�P8�q[s�J�fӷ����E���[|�d�ɀh]��n�eAθ�q��8.zu�M�C�Cs���vp���H�T�h6�W6�Ll��E�����K�6Hu΃�ݶ�S;��	է2:�c� ]+�c��;8��0�6�V=�@�Ҝs͗D�79Y�OIu���[\�W�u�y�GFv2����B]gB�m )u#�;a�Q�<�8���͵�EG;�iM�geڜu�(�%�UH^G��%�4��Ўj�mnI��Il��:�(;'\I�=I�
mL���'Wvi㦙��!�N��� p��+�H'���� u��]d���^�r[�\�]�����8|ړRm�G�^��5�g�1s>�h5�;oe�a2��(��۷�b4��g�n�:g�ۉ-�c��֋v(^�����j��By��ܱut���I�$�M���;�����p�vf�ӳ���5AGu�n�ʛ"i�����Y�9ez����nv��N.�ܖ8�3�:�ixв�fqJ�h�8�FӁ�mv�5�@�nxy:퍥n0عL��7G�����v���k��s�K��r��������l$�ڇ���z�ÃvN�C��Hrpi�.���[WfM�<ga�f7hT�{S��H�gS�ۦ����B�����.֚���:9�T�W	��xe�J�͕@�1ֺ�Z���p@��c[�d-�D�Z���dy]����V�\; +0z�q�;�0�2d������\�#�i-0[O,��ͷD��چ��ʂ�i�z�Ġ����ɺ�jۯ*���-zC��ӷ4q�n����;~9�6�ݢ��mԯ��<Ļ�l�ptM1�Kv�w�J����t���9�	���ɖ[Wm�Q�!���\�25���E�������8�:8�:V\����w��ww��
� x���Dj"��_PS�p�>D�� �}SDW��˹�e�.��d�RZ�l�N���㲳��������ݻfҝv�!�����t'.��<km�ָ�.1�@8�Ev3!�p��*T�b�ga���7+����m��5YC�[����>?7�x#u�	��\5�����\�]��OA�O]��zbn�c)�����v�.��C�Vݸ�p�a��9E�ҧ[[�7\�S�K�k,�B�l�C��{���������ujRѢ��7�=���sƍ:V�/U����u�up��7/��uLֆ�KI�@�u��	�Q��"�&��	��UiӴ�v�m� 'eG����d����9�� {���%�UF��z�`�65m[N��?\��`u��}W~���o�� ج�JE�Nզ�ڶ�7\0	������_U�o�������4�t��f7\0�W�_����={<�	��m썧t��-:�n1u��u�]�n�5wi�tR9ɛ���>�Ηx�\��\�3.Fߛm�����@���dt�/���99�xشٻ�6ۆ�$����s�
>h�(\�$��"|We��>}~0�Ӽ�'ʚ��4��4�o@�:h�� 'eG����n&��BM]��Y�興KТ!*���0��׀�7\0HLeڤ�4�n��l�����W�Y4��L����R���.;;7��[h��s��B������7�4��յ�i�������� m��%
?H�����z�����եm�n�`�����	ݏ ��%��li*�UEUY�?�ـ���I�IA�фE?��j �Ab�Í�����
�%ܧm	�I4�`r�$�%U����>��vـ?��@���\�lO�m��q� �����K��?�� 4� �}N�¼�،��3�h��p����tZ�-�O`:�{������ǾC�W.��|�?�`��wc�7��bv��ui5mݦ`�៫꯮�����l��&��	��T���m�M��*< ����_W�Uw$~0l~0lu6�ݻe�uw��Q3�����?�فq����O�D���>�I;�Y�g�K��$4�+m���~����l� �^x;��6V��i��S�R�t,�7��]�ED�8��^9Y�M�251���t��f;��*< ����`wj]�vН4�@Zf ~z�璙�׀=w� ��fy%6mJ���6[�6��M�}<��a��l~0���w��bt�S��1�6�	��OGM 휯@;dx쫘ݶ$�ZM[e�`�p�<�D��u� ��^�m� ��I(�.�����߶��:ɍ`.5tj��R��dѠp]��=Hp\��F��qY�%9�ݵػ#WF۹vz;��sA�i�7 �6#a��Ƕݕ�,in���.�/.�'';ۆ�{�K�ʤ=��3ϓI�mmv0&�ts8�[�+�۪ݤ�qsl%g�3�p�@��m�e��t�#�k;��g�x�it�\��s,R�*)��$�D��sݤ��D!1�����������6�Yvy�2�\/i�;s���9�h]1�CѮ�j�r	n�X#S��O�����^�=4	��w����ci4ı� ����>H��Ɓe~0�j<�Y��M��Е��=4	�����l�@�"�)�;�j�$ZL�7���Q���?�
^�
��� ���|�n��i&��� �ڏ 96<{��\0\���J�0e�v�W�x���W��,�WH�1u2[`��T3�v̑������κ�st�Z���O<{��\0�r��'�9���M�cBm��Ӕ�`(� ��A���o��9 w����M� ��s�ē�I��c4	�����l�@���d&2�Sn�M��m6`z���+� ;��N���������e��[-'M�&ǀ~����&�� 'v��'d�P�i]�M�I������A��G˅��x����ӇM��C+s��!�+M�w\0�`&�xɱ��Ȕ�4�ݫt�i3 �� _NW����:h=yR�i�캪�j� ��;��]�P�C��.'!�#�@���{��$�{��rI��Ч)��1�I��o��}<�	��4	������G.h�|i��hM�z:h��@;ez�+ݶ��O�uE���֖���7f۪��Н���V0�y�-��*��+r�ff3@����+��^�=4�:�Y��x�c��6hl�@;ez�t�'����WˌhM�7��ހv��	��OGM ���Ȕ�4�i�Zm�~��l��|`��*�D"�P��Q(�{����y}���6]�v��0���w�� 96<�������w��w�8s���Xwg����qi9��O-l^����q�c�&���Ќ�@Zg ;��v�"�7��w�� �mhS��j�ۦ���� ����]4�nh�.]|O�>4ۤڴ�ٮ{0�Wr��X��� �*�6۲��i��`�p�"������:h�u�����ƭ�ـm�E�v�"�;5� �{���xj�����!	�h*|o��ͮ���9ٓ�eoVW����\�2�����e�a��\������;N�����u&�S7FK�s��[8����p�����"v�7m�j�v�O8;�t\h���Z�Y0�[u$ȧ^��];{qIn�{k�����0��>7U��̈ↅ���)��5fv F �X�u���`�' �Ӽ��LT�ݚud�Ϊ1�n�.i�M>��|�9a�-Y�xy����h�):��3�7���C�Ê�&뛳�1z\s"�%5�f�'��?����\0�p�6�"�6+"R��e�6&�k ���\0�Ȱ�ȳ�vK�"^�v�˵I�0�~0�nhz��=c��r�T�O��UWA3V`(�R�{� s�Հ|�فВ���y���
�]�J˫*��5�m�E�~���}�o�,wߺ����l�f6��\��ԯO={G[N�9�x�v]����^�5����tU��,y�%���8hR&�d�l.ci2��i��`�p���U*�A��s�� �?7X�m��d�Y~wv��m6�ն�0	{�,��ٮ{0�̦��i�6�N��Xo�,�\0�8`}�`�Ȕ�4�i�m���p�=����%Ｐ�dX7ee��J�ӻu����Mv�[�w��7	[/�p٭����r%cI��4��V��f��o�,��ٮRT���tؒmXZf�������4z�o��P)��-Sbn�5�mＰ�píN"�x�c(����!Y#=Hq�Y!)$IV,�	F$�	 ��Xb���_f�Ȁ�$��H��
�8�
J�����:�0�B#0uMZAH��Dԉ,��"Ā��R4&��HQ�eVD�Rx�Bb����hH1�S�1	H!
�� Z��0F���UԍY5�&C�,���Df�^f`%�0��4b�!Fb�]z�0��
?�����%H0[�@�-�BBJ�x��UQQʉ�*0b*?�P�P�F ��#�:� S��=�g$�^������S[���I�i��U��x�7|�`}�`�Ȱ�\��am��4��0�8`���}��6��Xf�|�~��I�}^��ض.K�NN�@�Ϸ�7-��K]��c���nz��p�5���CV�l�6�"�;}�`������~0	��M1��bmX�ݦ��c�>{l�7�`?7Y�BIy(UC�//��&�-!�I&�?y�0�`}�`&ǀH�ȓ��i!:ZL�'����� ��YϹ�����2���P��`�**�><���'$��Ƕ�l��nfn�	�0����	D�ϯ����7���������tv%��r�d��:�GOZ�W�t��S�v��K��nn�=f��-5��y���ou� �� �t��hvۤ��ٮ������^�� 96<v1��[b�M64�w\0��x�#�9�� ��c.���cV�`��8��x�v�%
�(����� ��즘��m�&�N��G�s]� ��f�ֹ�.Dz���w{���������4�\���mB87�z�}	�+��/筰�R���"w$�H�vȒ9z�q,d��	�IQ���'i4�uΩ3�}�^�K�� �ۺ4�9{x�Ӭ܉����;/V���c�����I�m��;0�T9ݹ�݂�ר*ڝ��PYN������/`݉�ծx6$�������p�������Q�kJ,[&v2�J]ru �P��3�)��L�ëv9��n-p��=hlrؕ�s`���G�3C�]4<��uҭ_�o�k�`��wV��I���'B�ա�Ui3 ���}_}��vlS׀���lp�
�\�&�i&�Wi�ul� ��������?kkB���TƘ�v��6G�sc����BS��N�r�x-]�i��hM���h��@��V�vH�v���6��Lv;cI]�Q����z�ڷ:[���r\Z�K��/i�|��a���blI�w\0��x͑���sa1�iЛlj��0��y*�O@��?�9'~����~ߦ��{�)��ݦ�m!6�w�����h��@��V�nrek)&Ҵ�M$�x68`�p�;�e�6G�n�dIЩ4!�Ui3 �vـt(�]���>��?k�`��ᗍ�Q�X�:�&��{n:v3�5�N"N�]y3p��K|�v��&�0<<��55�,g@�/�����h��@�
r�'m1��;�l� ����f�ֹ�D$��9�l�Ut\�ګ�n� ���}�l��i��*�_��	1Q*!���;���c�;�.bi���j�li��t�=2U�����h��ı�wnf�ܻwvrI�����O�O���������7u� ;��D����y�e�Pӫ���Z(�v����)t���ّ����p�en��)3�Ͷ�����c�\0�p�6�"�6*��I��!�I&�ٮ�`}�`$w��!D��NN��R�����5V`���"������:h=yR�c��v�]�`}�`$� �����OQ<�Po3�g$��Ol7���6�l��ss�I�{���O�D�������l��`��z��I*�n��g�7gdڴI<uh���`�銺]֌ka���m�gE\�*��~�}���7u� ���}����'��6�ݤ��ƙ�n��� rH��p����}Uvvx�2�:m5i�hv�0;�X��xy%�w��6�{�)&�;M��J�v��Iٶ�wm��D%.���ԝu�*�i$�M$�xf�`�������K�y`$� ���߫�QK�N��i��0��i���s��E×n��b⬦�^`|����هf�Ʊ��X�\v�*C�wWVLt�5���r�y���#��y�\�����0n�|�.��cr��\�֧v�1��̨��	�s�m�6C��3���8�.ٸ���[j�k�]o]:���ta�nM��Wy::+�9�]��6o$$����ق2����|dZg�F3���ww��;��??�v��R����%�n���EB"�Nr���+Ỷ���1˴ɥ�6�C`��f��o�, ��+���a��� V��w�e��V�]�`z���^��4	#�����ĉ(�S�6*N�j�V����xf�a����#�K�y`ݱ�����hM��:hGM/[��k�7an7m�۴�6��0�p�?}UU�[�. w���;5� ۄPT�Nm0l��v�u���:ϟ=��6���Mŉb�4��A-�3\�e�'�����ͻ�>{l�DD~�m��ت��nf��ܹve��I'��w����F�eV�0�P8y?w����`}�`\�]$�V�餓��>{l�7vه�"!L�������	�t6ĬlZL�7u� �� 9$xf�`vT��ě�ٜK�E�s@;mz�t�$����>����u�$sv���b�,�WYwb�ug%\�<�ƈ�@�<��wx;|7_:�I�M��&���~xf�`��m�E�ov�(�C��'e���p�$��^�4�נID�i��ĕ6��0�p�6�"�}�}[TU���dIHbT	���	���"��rB�I(�U��}��{���Ym��t�wi��v�0�Ȱ�G�vk�諭��g�l�RM�i�i�bv�5��<�\0�p�6�"ͷ���蝾v}r��9�"��){F+]���c��r)NN�:U�Jc���w�3�]�ei�I6��?�`}�`$� �m�'ClBn��ZL�7u�=
"��u`��x�m� �i��j�cV��Wi��dX�#��}_W�{��`G� �ѶS�ة;i�n���:!Dz"*���x�_�wm��(J!I|�B�+����epZ����1�6�X�I4�nh$� 4��j���I�;M�;��nH�0�P5Uj���YCG�^ɺ)��V��*m��`��m�E��?UW���P?u��7�_�fj�]\ͩ����0����(�����|`�l���ɳ�I7i�ݤЭ��X�{� ��w\0��`�;LM�i�I6�?U}��L�I�nlX�������t��W7d�w34���wm���7�����?�PTW��TW���?�QEqD��PTW�AQ_��AQ_�A ?��� D� @ ��@�$TB B�B
�"  �� ���ࠨ������ ��QE|AQ_�E��pPTW�AQ_�E��

���b��L�����A� � ���fO� ��~             (   �   ;�  <���� 
T����A(
@�ID�*  �U���E 
J	@
 �I
��(+    `4 (  
( 0�
{��ry�{<�^��ޗۼ{�� t�����5�����Ϸ}��=����O@�0  � 4��=��g�UL�����s��>YJ�Խ��O��Nv��]���q�����J�� �    ( 1 j������l�ݵN\�n}��Y�@���<���˻S]��m���j���4w��{�:K6� �&��|�  A���  �   �@  =` `   ��� �  7P� ��F j�� D :1  �( ��y` 1( M� f�@� (��m� � Z�  =���� >����|ޥ�R�[��Z�` =ܫs����o}��[��m�y:�� �B�@  @(� 4���n����W�W^�}o�/�Ǟ��x }>z��w��O'^�<������M��ܯm˾7�^�=| ��j���կ� zO[�x    "  ����}�G����iɮ�ɥ����x   P  ((P�=�ڗ>����|wv���ӯO��_M���4}�۾�OO->���<����}��O'ݞ�Mx O^��]��>@��ک��Z�������-�U��/g�)^m��y5��ɫ��=ԫ�OPT�Ҕ��!����T��e3T�R ` O��j� hتT�(�  E?Б���   ��&Ҕ� �➂t�'��g�������rv��������*������U�T?�U���*+�
���EAAS��G�`���g����_��z���1��@��0*Ʃ8�
�B��jbHBR�r�1H��"��0 ��Q#L3d5$)&)�`2B��Mw��4$t�xld�&� H7a�v��B��0��s�Ǵ%��/	,����q�a	�<�zA�1���K�#�]�BF�~������x+�H��I?,&�@��?��o4r5"X��x*��*��nn[B��,?SxhfyX��P��R��hM�0�L @�䓁rBٓ�Ʌ4�Ri3=0��k��&�ۤ'	Hc�c K&�:y��}�G9�C�iH�B�XhW�f��K	5�_7N_�g�!.H�Hl�Cp�\�L2�(�0l+����i�x&#
c2"BJ�[Ysz��q��A�@b/�!		��V5 �(E{�c���<fs6BN&�Yǰ�c�4�peq��7���wz<����h��ъ��C�BI\H6	E�M���0!L`B4фY)J��<�a»�*J�5�4Ɯ�2;���a�#'��#�+<+�%8��(K����2�%IJ�<�%�E]��p�4�CL]k
F���t� B_5��a�CO%�cF6aH˹�$+�Mb�HP����p#
��@�	��Zc,%��HI��y�.J�����J2�
��Rh@��!Y�3 m�(`A�XP�P� �D�hE(B�e��v���H�<aq�p��@���6�.;�%sNX[��6���4���tC�\�p�
7��@�)��-|�Jc�%%�1�	 a�cYXJ!-����s�����k&�B�8i�P� �1j�$X��F i�B�F+�+�)
�9�7�sɆ\�a@�e�J��*�硆�H�X�Q5H��P" T1%ɻ�����O<����T���$8\Hf���2$d���l\��SSR����T%Q��4�bjo'����r�)���.i��e����m�5��BP�2�+�A��67	@�N�k�� �I8�Hi�渑$��!�W$)y�D�	9 �"D��k)^�o!�e�79�
@��p%�NL��p6�-Ƙa8l0�d!.$(@�#�t��S2�u�)�#$�{s������p�s�������D!�W�{�B�	��@�����	u �(hx�J�I�!x�������SBF#"Ѝp<B%xr_R\5`�������_Y���́1ʙ0�.$����#cd���xB������bK(���$�)�T�M��aq�\0Ú��D�p���ń�nf��k
��L����*�cL1�T9f����	��g��VŌXB$X�"D�R��%�X��!�j"��4��	W9B0��\�@��eͬ�B6��6�)$���J�х(J�6�,�HZSH�)B4(`B�I���l� ƲcX����+F����ch��8��{ ��k㬔��w�3�%�h�QL*E�t�3K$+S�X@��-7��ܦK���F�XV���K��� ()Z~X S @�C57�8B2�"Z�d��.i��IJ��B�+B�����p�5"W7r�2�35����<�<�oV<"�Y�x6G�k�D��4��F�cB%Z��z0�+��Q�1�����Z�-P��{�^�h��0�6}w�K��H\�<!t�K�#ʘ\ILI�d9�(�k����b~�/��<�ć1��u��D�<�~,.g$��\e<�<汧���{�A(��"��F���0���q=
�B�	w����g��3�K�%e2��%XRQ����	�g�$�S���M璙<䒜Ca�nl��R�����+B+��i;���X������/�K�Ќ�$*Ff��.q��S�q����!�)�U
t^��^u`�>i�`�Þك.��������ĉ�o�\4����\�>&\֘p�����TÝ	���x~1#ほ�$\Is�`�K�HaRZ:��	�[̹�\��=������K�]e�qq������?n!
�!���F2,.K��E�[m�O3�Mp��?�<�eR���/�~P�<Ѕ�99'? xy��y���F�w�(��g��!]��`f˜B77��b�x��ƌhs�������
qS^,�i�G���|᛾G�� ��tOG��1��A����~d�/�#��J�+���%CHÇ�=���_ c��<��=�ˁ)��n�܉���$�@<"@�$��$��Ė_IwsA�V_I��s�߿~a�`A"ԉHD"-`A���1�:A�:i��J��
ĉ7ԛ��!p�-�B]�?RZ�@���q|e�.F䆛��)�.l�B�wI�j04"�#Lb�LH�\a	�SS<���2-�8�\v�r6��Ӟa��r!4�d��xV!IrS�1С��<%�
�
d��He�8Jy..	*B˄�x~��'��5�M7<�)�%���y�<�=��.�t=������W��������'m�Q*���2��8�	��U������B<�p�@�c\�����ip���㿳Bx:D=L��������Z����H��Z��$#��h�(bk�j�H,Z���n���H�k��|��C!L ��r!MaL�u#L%0ы04X5�40cr\�?3p�)�Ii)���H���8��g�t�H=9��sȓсc?h��H_9��F0h~'��I���͘~p�hƦ&�F�*Huq`&�B����qŔ��SdHB���w<������L���`�,���!\gP��#�C����a줅��6�<���xL�"AMH�G�@�������F��̉.@S� A �0�� �`S �$�#	*V8B��/"�4��r]��hJc����Z��B�HR� ��f���C����O%\W�!L7
1`p��13
�9��L�	|p�0�p�cZ�d�Jf���Z1�.�k�	�-y�p�n��5�%1�2FFK��@���0�))�ƥ�!`W0։�1�`Ywr3-�5ԍLr�rK�$J\6�L_�*f��>(��U�:-����k^]l�>��Hɼ�U�w%��'�.���NTu-}E�����P�\Z���eC�p��WV�Q�V�u(����U�����r�*볙Q��\˕���K��u^(�B7M�t���Jח�D��� B��.�NN+������v*�r����Q�k�rr��*?<�:�����:H��@�r��E()+)r�hf�?HR=8x�i�l��b��C��j��0����	P�6C�ᧄd)�����4�C�����������q��)��L]4y��6��7���E�$��&:s�˗yM<��9��2\+濲���,q���"A��)p=x��D�S�XRLOFB4p�##�t)%p��.Jl�����8B�J�D?'���iL7���'&�9�=��}�,�2$1FE��L5ps]HTq��#	%p�!B4���SA�P���`��0]4�@���ĀP"��BBL��.��zν���_�t��~@           m� �8 �`  $ m �����"m�H���Z����#R��'a��mI�܀    6i���m	4Ѥ���UPFRBb��A-�^>e^VU��� j�g��M�m�  �kd��:�   -�����KHu��e���l����I�^bu��ۣ���θmz����<�ô�����-��#Wqc�����]p�\r��2���[H<��^!d�D����3��@��l����`97\�V�]U\�U-�0�am$Q�ѷ���Z�aŴ,�e�`H��Z���-rݗct�{!ĭ͚N]�fҒ�g�{m�[U/<P��S��`	�U;\���4��k��fz�.�  ��5���C/C��M�ޒ�6ۀ	j�.y�U�CH�Uu�Fy[a۲�;�UUUƥb�Ymv۰��-�j�`��  ���ic��tI@m��D��z�K(� H   $8	r]�qa���m�m�r�հ 8	 [����mԻksv �[�#�rڶ���2��)@mZ۰   [Vݶ �  �e ��h  ������uԒ In��I��f�  � p 6�ÎpR�  >��]uC�y� ۶5v��_�}�ݾ�6� ����pjI8��tRv:�Tr�z�P� ����*ʵU]*Ԥ��엛�;9|��B@��Z������[E�͘٥ �S�iP��Ts%���P���֝Si�;%���+f��-Xѣ{J�N�]-M�C�B;0�-���m�yvWvn����`
�d�[@��u���n�Kz������m  � 9����+�I�p�`$�,2e�[M�`� 8Z���l/Z��m�  ��v����mZ-� [d$�p    6�ߏ������1 ݷc�m�i)@���L��c�U��Y:�4$�7�Ӻv��rܫ[V��Q�d�}�_R�(K�N���Ue�ڗ�5�m��98�[�[P`�`�i�+�8ȓR*�V�ҭ�/.�Q��Z��HD��]��8�`$#E�6�p�K�VV�T謣U���_V�i �� H��  ���M�m�NZH���UK��mxl���8�aǛ�)V �L���YmکMR*�.���-��IQ�kUK�{ym��t'7T�4 {jV�^vٕ 1��Ur�R��ͺl�6�f\�Ii& /]1�I�Ή $�/M��_&����n��a�\��4+���c]kd��m�A�X� /ZжȒ�^�!��6��k�c�&�	���Z%��6ٵӵV m���!%(-� 7m��iz�Lj�m� ��1��M�\�eZog��mF��zݶ ,�E   �[d׮�`x��t�    %�vZ�_/]��T�q*�*�@m�`6��� ֋iWn\ͭ��h�n ��l��n��ۛVͶ �zCm�x��ڷ��6���,�����wV��(R�ɩ^���ꮍm�R��/)��eV�e�lm:+n��}��Jܬp�z��tmFxQ��-P�%UUT�gg�%���-�.�	�k��l�m�t��@	  ���i���phH4�7  H -�Ŵ�ki�\�&  �v�t�v����+hN1 �*�]V������l�����p8qčN��`�v[C��a#m�P�Z��!��,�uAm�l�Z�ړb#m��q N���u��� �IfIv�	�,k�ʫeZuGd���veWf8�h�n�\ۭ���IY�`�ɑ���-�n�l�`6���=j��eg��4�B@�_6Bn��Z�
)Yٻl�ˎt�v� 	 ��km�l�[Wnn`ڳ���btUULkp m����d���`:�%�Bںl�)�l�Hٲ�����4�mU.�X�]���Яmm�ܵ@@*��TP�-ܫ���bE��]�ĵ�T�ұ��i����齙 ���D�ml@APR�U++�Gf�d���Y[��Ӻ�VX
�����aݮض҄�� [Rn�f) �ꪀ�U�޳�Fq�Ԁ ��j��"Ω@7nێ:Z�ݳm�� o���M�� m8����M�,5�  n� I����N�2ɮ��`  t�V�-6 ��|i�Àp�m^�΍�H'A�����I��(�n���n�[�m�o\�-���z�	�� -9%���S; me[m��n� զ�]�Ն ��3�hmZt�[mrM#m����'V���ͫlB��l�I%kB@ 8m����U�]�bQa,�[\�8K*XV���m�C��P�m=6� �-�9���Y�l&\�m�j��e��ܛh'ma�� pmm�λ e ���vkk��e�fڂmUOZm��4Ͳu�HH� V�t 
�H)p�T��  $M�l� �brÖΕ��Jԍ���	-����f�%�I~���ڧWe�퇝��k��v���jv� )Q�q�,�bq�S��T$7K��R�-�U���Lq�������l�*$�p6�P ���t -�Nݞ��֫d:��Gcn�඀ �����Z�� �j�"յ�xs6U����j�媪�
۪� ��)�;s��0N�m�c�}s���WM���+nP[e��j��{O����y�PsH֕q���.�-k4�7 m:-�E�`0-�R̍4��5��:J�k�4�F�Ř�j�&vvj�R�%�j���
yT��y[��˵��@e�7�؍��������y�e�3rm�:\Z��L��$�($	-�nH�`�l�G����� �J�m�қm����2n��p��<\|%�h���L��]���`p�e�#�ݤ��6b� �` s���Zk�HEH-��d�e� 'n��  ^ث�V��Y[A��0l�  []�l$p���2P6�-[t[Z-��v�CӠp&� $o$5(	 �	$��� 8�m�-��a�W���	VP㗲�Tq\m�bm[$�8 �]٨�m�$  	 ��ݶ�˰ �` D��m�7k���	/C�U�{U��Hn�6I#�@�[@6���í��h     88t��۴� $����[CEm��d��mh2p6Y*B�	ڶ �C��pm��m�Z�U� x#`� �J�6�m9��RKM.�%� [@�*�ZR'vB�����Z��X�R��y���wd���Uu���������َ��Xڶ��U���&�[ U*�,�@U�������5��jUڕ{k�!PV�,�����.�sI�� �  m�   6٢�� ++U����ҭ++*�U   � �� I��l  -��� h  m]6&�8�� @���,�` �j�  '   �� -����m  m s��  ��� �    8�뱀�n�6ZmS`  [[�|����O�VU�cb��8�ѵO<��IUk`"��Ҥ�UU:ݍ��pu��OHT+�v]X�g@x��� �  �o 6��l#�]i��[wZ�3 �6�l [V��Zl6���� �h ��unm��H�� �`   rڥH! �a$�ZW2.�;dbc�49f��8� $ ��W�� ��n� [
��ͪ�I0�[B� 6�lm[m�8mmb�`l5Z_������$�k�ɷ ic� $  �   Z�	eٶ�m���`�Uj��(
�UU*�m��	mͲ� $��h��7VҭU+���nհ[ն� ��Ͷc�-� Znz���ೄ%:YV�-�V���Bafv^��܀�ش�23m�@sm� m��`Kd���ݫ`�ɱ;�
��y�1Ȫ���U�j��*U�Z��^m����n�*g�`�Z����UW�� Iŷ Hh��U�W�����t��
� n4����rXls�Zl�fH8�.�]Y��npM�mUW*��UN3�]��6��{4Ҳ�N�qW$@Kä7�YW�jԺ�]��pX�
�U��Ò�+:id�  �
��l�j�r�{:E�UDJշK奍���l.�q�km�l�%�q  R޴mU�� 	=*^Z��Ζ�&�pl mƶ������v�tW]V�,�4�rYN�mfE�ɵ�׶�H� �ҭ�I��v��[ �m�6�K{ m����\��g-�:CH H �	�����%����V��@����[BD�6�Z�7�{��w{��U:��"�p�b��� V�G�X���x �D㯈+���τ"�!��A�O�`��qZ+���<A^� �G4`���A"�C��A+�}Q��4�����0OT����}��B�q@��T=���JO� z���"t�ʇ�(!�EA�0E��0�U@�=�B�Q�'G��<N�w�D�U榢CC��0����A^*TT:(� 1 � � T ��z��!�P"D ����Q�T����q1$@`�X2B!�0��!"HD�  @H��@�$��$H�� `* �� ��= 1 ?t�U4k�(>?�8�
#�@z���A|@� 8� ��3��OEQ� ����T�� CD���= Oދ⧪+�~�W� 芺+�A�T|=Mc����Q��@ �.#�T<�����R���)�G8 �@Q�������E�₫T=��:���!�D����E8��E�*A_�!�����p�C�*�~?���UUZ�h	[���n8]�T��u����Q}�ºR�=��n.�D�2��m.�q��X;h:��f�uk�⍗����Cb�L
�Ԧ�g�^��nKLq�5Р=v�\� �I��[9T���fRY�j��� ����/*�Qܭf^�lv�ڱ���&��r�R3��������p��lsuvv�qm��6yv�Uڪ��;�a�\]�8!é(AV��e^6,\<�x�+ؕ��J\˻=���{&KB�W��l&�j�9�V���aR��M،��)][pa��l�'��;;/F�s�Ft=�u��&t�K�8�խ�l�ӌ4��7`9-ԓ�[|��ܫua�nw�2��u�v-�b5���:�`���j�r�[[Vla: P^��e���$t�� {l�gY�u�@�#q��@,rc�h�����z��+8��eq�8�Kv�k��2�;&�tgc*6mi\\i����>�\hA�fx���y8ڕy�n�M���������ָ�
��u��s8Q�F�:��V�!�+����f���.�I��]�:�]Dm�\�`���.���V��N�({�U��|i��T�h�]�s�ig<�;��\�.�@��	d0�-�jg��I�Ͱi�p��5�U��J�K�L�	�`#M�\:24��M;&&�.#������}����hp��v��3uټD��7L�[^��f�h�u�$ӱ�o^U.��m��J��c�y���'b{�Z;&gĵ:*Ц�]$In����kKd��Uכ[�dS��]@妪��5�PΫ��ܫH\$��4t�v�l���
�nh6O(�ll����(k�(�{'e"�eLL��6�v(ymɷg���c�^h��ՔiݛW  %C��sۉzG���ݮ2v�v�c��+�h�ŏrm=H\�j�hΊ�M=I�^�l�KK睻j�j��<'[.u�]%Ӗ�6��M+�;n������H�R$�c��0�@q�=�
x'U<0O¸��h�@'?yo-̚Mɷ6]&�d�Qa�X8���"�৑8tTr��ծkڈ�7=<�CE�g��l)���@cu�\���:!nر �{\nv�9:��i�p0��7�^�zÌ�^��5��1��+�
�;��<@��a�L��a����:\[�tn�n.-��v��dj:�g���Vճ�7]�[vm��ܭњ763�Cuu���T�u!�ٷ�d̒�L�8=��dOg��L�;��9|��N�G��Y�zu�X�m����_����@�}x��Τt8�e6�ܧ`s�4�}_UUW~���sO� 7_^�^�X����X28!�p�1w5�{�,-ͧ`s�4���I5IIM@�R; ���ұ��=U���:c���Er���Ӱ9ݚX����͖s֠G(��TR�:�9�`�my�8�k�e�;lh̛�\Y3ђ��U�:�)ܒ���������`��8�6�����V�
�rH�6��I=���s���T��P0hb�*�`AP�AG ��_�(�����~�g[U�{�ـ]�zH�R:M�28��ݖ�Ӱ;ݚX�����Zi��8�8�6��#3�Ł�7��;��`s�=5Ԏ�������f�>�k5�{�,-ͧ`z���^i�$N֦j�k�Fku;;mn��l��VР�%�N�ڧ<����ͷ���}�vD��Ε�ؠ�&�y2��%%5(�)�w������vfmՁ����F��hJ(ې�6������I=�������",��,$  �AE(>*^�I%iB�_�l�:��� �\�ԑH���vfmՁ����9������v�b�v�
�rF�j9Vϵ� ~m��^�X�X(�߿���g��r\n-%v���<���Ӯ���:ْ+o]�\��𹻳�ͨ�S��X�g�7�L\�X����׽1�s�E(�6J�(�8�6���Hm�/��Aξ� �w^ ~�%�˺EZ��r))���V.�"G7vX[�N��GFlc�N7mI*���u��w�~��V��(H�\�"�#P������OP�U_<�r��<���MSP!��zH��ұ��{�ę�o��劉������2X�v�����x-AGS��a�=7Ont�8�v��2�0zy��v�g���	%�@��p�E�:�)�9N��vi`b�k��vX[�N�#v�V�R�I�$��x���쉁�+�B�2���(�t�5v����si���,]�v�Fk�(�6H8�����v����_��7���~�w�OD}� ��)�O���ߝ�ӌf��0��Vūv��c��v4`�I��	{�������H���Y�|@X;�+�V�c��n�9�z����7=n�1ln��	�I��l9��Q1Ky�65[	��D��vK��nMq�!G/gc�9�˲���B�c\�9sU���kk�NÅ"qi�I9�M+[���n%�J���	�χ�v���ib�8B	�S��ruq�������qޠ��r�-�N"ipQu�wƮ:zԓd�*p]�)lZ���\v����GC������x�g�s]�s������v::7c:qȘ�Q�X����$���:���`w�4���J��R��E��;݉��+�A�׽1���ɒ���nB8�rX[�N��vi`b�k��vX�j-��jFG$NS�;�A�{dLvD��ޕ��~��¾�^x�cS>���
3��-\U�N�`�w/�k���K��^eIz�mH�?I��ɀnȘ{ұ��V�dVi���m��I'������� ��<AOȾ�|DCl����;�O��� �5Ҏ�pl�q�I���+�A�{dLvD�;��i#��"n��9N��T�wܫ �{��9�����m;����8��UUwk ?y��9D$�}����}N��ͺ�5n�D�DG�F�4�s�.�����ӧ�g�ם�����Vx�����RiG)�I`��`uw6����u`b�k�7�{B�F܃q��?K֫9(��w��ξ� ������j��Td�IN��vi`n��s�����T�\�o$�_��{�*�j�9#R8X�5X{�,[�N��vi`]�{Ju#�驂ŌvD���+�A�/zc�_��?*'wb���J�ڜ�a�n��qs���[/��Қ��.����F���l��,K�K�+�A�/zc ݑ0�`�����'"r������_%	L�:��w��>֫9(���R5��N�r(6�n�o��w������v{�K ޘ���4������Q	(�����*�=�l����?!*�K!��DC�u����`gX�{Dl�9�i�`K�+�A�&t��"`l�S�&��ɛ���/:Xl���[�����P^:m�lk�nV\�#�
v�ؠ��:[ ݑ0%Ε��]k�RRF��N��W���a��L����7u��^�N�Z�WH�Sy���I\�X�݊	3���3](�G�)���ͧ`w�4�7^j�iw���7��(It܍�v{�K�{�|���KV�U�����H����ꮨ*Հ]d�&˺�.�N�Am�Z;�vQr� s�����I">cF�v��O+�=o�+�]l�8��y#�f�kt'%��t�S��ia-#�UzSP����Kq��,��%��|3F�!Xz��ok�qU�In9J"������nLl��7`֎4����U�;]�)��R�����RMv��	:}��Y٠�{<h���7�r�����a��l̶nm��3*m:�v�,'C�E��c���������{]:-��q�N�r(6�n��X{�,[�N��vi`���j��r��D�+`�&�ұ����L�o*��4����F��q��5n�;3,>��"eξ� �w^�j�8�J�Z��+�X����׽1�zH�[�N��i���@TI$i�'q$�f�;I$����$�[�RZI.�oNq$����o��\C�ȷUv��j���X�ƴ��lML5�+S�ӛ���s��yQ�v�Iw���I$�6���]�ޝ�ZKTۧi$�kQ��GJH��(㓜��{�L�j�� ���9o7���ʒ׻l��K�ݜ�E��(J��NF�Ii$�ݽ9Ē;�Ii$�{�9ĒK��%���IF=iө�ڍÜI#�4��Iw���I$��RZI.�oNq$��Ѫ��$�!$%��]���K��U7�꓉$�=~9Ē՛t� ~��ߟ���߽(	��e��W4��Z��9�zIކs�m�ٲmF��/:����݁�nAH�rw�$������v��KVm�[i%���q$�����S�Q�Srʎ�Iw�zs�%�6��I%���q$��ڎ�If��_�R�H��N�Iv���m����|�������	@��H��bB#�a'�0d�֐$���a$dc�,�ea���"����dd � �c ����_F�uL��"A�8��$!�H�L/��"��2ڐ�J�YH��@�ݠc&2�0J�F��`@e�A%Uh��Z�@bB�B����*²�(>��<��bo&a�b @b�0�b7B4�\%1_�{�?(A x=I�ќ��h�!��(��H0@� �LZ# A#R:h 4@<pP�"���@G� �?�� ��@��T )� �����4O�C���;�s���o���O<�	��|w�9����MJ�BZK�UM��zs�$��?}\m%����.��ʪ����)�I%��o�(�I8��\�ޤ���Tw��O�3��ޤ�����I%���q$�}_}�o��V��\n��^^x�挼�S�!u����xģ�����N�����X���f�����u$����s�%�6��I%������̉$�{�Ii$�IG��8BJ�mF��$�ܚKI$����/6���Ii$�=~9��_g�W�_���pj���9*B8KIq�����K�����I,�_�qz�~[�e���a��	:�r
OTR\�z�B�����Y�~9Ē�ޛ�3�S�ſUUWǢ�"&�������<� �����})Ԩ�)�"r���\����x�RK>�?]/WB]�zs�.�4�S�$��^�L1�Ls:.�n�^��X:&by�G�0a�ɴ�����t���j���������[-$�>}�zw�%���KI%����ImfӸ�S����2�7����`N��'GL��I�k*�YYj�%�06�0'tt�U]ȣ��ݖ.�E����H�qI%����N���nH��e&^V!	R/31%L	::`dL�"��X�I�	BMђ]UY5wU5��e�aՌa5��"g0n:�C��e��f�WP�n`y�w��{jy���p�{F�����~��GE����8έ�\�[��C�dK�0��l$�8��jڹX�ѓ�$��i]�vӈ�ꦔ��۰G�WM����unu�Y��Ύ����X��<mv8ogHKY�F�lU��N݃=.c]�k� 働��P�ru��uJ�l�Aj� ��s�M�m�t�ܒ�a7N�0J�j��Y�U*76.e�w����5�e��@�R��RW@=���:�vKs6�q���ߋ ����&�7 �cwyТds��x7عB� ���B������+ν��R��SqE$����o�`]��(_�����
�[�w�{ƪ�(T��%#Qʿ}_}I�<`ou�Q�������o���}N�N�t�JTN�ݖ.��`nf�XܚX5o���
NR*O�A���[m�"{^�x�׭V!\#��5�9|�����*�����Kwd�73n��M?�@{=�`{���#���$ڊM�I;��ʀR	�B*$�s�X���ۻ΅	L�ґ��4��*�&������ ?7xt%��{ޒ��ﮬ��jpj���$��T�&ȘrD��:`I�� �i�`�PnAH��:�vKs,�x����:"�}�l.�T�pk�59Ru���s\[]u�H��#3⋛��F��DuG��Ý��~$�����w�׋ �� o]��9]���I)$�G+�{�� ��� �͖�mՁ�Y��*���M4�#�`���w��y<QM��DDU�DD_�����0�l�ҙE]ҫ��X� ���:`I�� �"`ut�$tI*H�q'%���u`z�����g�,��,�kZ�M��k5#d�v��u=��؛ktl��ƻ`u�rZEd%Ɲ8BJ�m�%XܚX� ��0'tt�킩x���,W�%�`dLoD�����6��:j�&�7 �crXnl`N��ӣ�6D�ەp��e*IR��Ę�:`t��M�0�~������{,i��ڔ*I�"Qʰ:tt�&ȘN��;����u�ʅ�q���]c���7m֭[p6i������/<��V'����h�K"JM�l��t��:`t��{�Y&U�	,��V�ĘN��;��L۫ �����iH�T�P�F::`dL�D���F�iӑT��rJ�3sn�{�,76X{��{wܫq�/'� �q��%Ll��t��:`t�����	EN�n7�;&�4�l�r��	��d�˧n��7ϯ�w۞'�89�;����Y�{Iӓ�r�'mc�6�c�wY��H�3v�ڍm�q�ph��b�;6�.�N-�c�C��k��iް[mpa�����GDn�<tv�୬v㷗\Z9��\�#�uōsF��mk����+[�$!���9�R��Ё��-�y9^q���Iր�8��[q�;��ߟ�R�����c�s�]@���ԧ% D.l��=�]�F��䳩�pS��ⶔ�K֋�u�Wd��Uw���x�x�z�B_}��zX�KǾ��2J��4�'tt���� ��0���V�J	��"Qʰ3sn���,76X��V�fӸ�S���Q����w^ >}x�X�x��l��J�#��(��3se��ͺ�3sn���,n-�M���7#Q��=]c���z	�U�e݋��[�$�n�Z��YB���%hX�����0N�`����GF=iӑT��rJ�N���砐Q�P�=��`�@��0�Q�Z Q[C@D �G�|�7��y$���w�gsn���kq&#��9*�?=w����J��ذ��X��V�I��R6����,�mՁ��,��g���N�gE�WEڹ-,�I����������|�t��w����I��
Dr:d�16��5���+�uize�2r���x�[q�i1ٵ��79�U������}�K �ݖfmՁ�Y��*��4�tԕ`��~��!����b�=����L����JewJ���]]����7u��T$��"�}Icݺ�n�8��#�:��V��0;�:`oH�zH��Ύ�zӧ"�*$�qʰ;��V�}�N f����ͺ����5*(���뎲�Np��Q#��F�<Qڸ�"�]���BXn�$��}�������"`wtt�ޑ� �e��+��f$Z�X� ޑ0;�:`oH�zI/R:����)�d�$i�`ff�X��a���x������3V��]��Z��"u�~X�� ��x �PyD
("�������>~�X��~�qT�MA����� ��0>���|���L�0=:e��^�<��P��#u%����^��qN��Б)u��}����sW-��~ ��x�X��_/�z�߾��_�~#��D�J�)���ͺ���W��U�ŀ��^ n�y�&OiHu�.���D�N9V{޺�n���~���{ߥ��{�Ձ��-n$�P�j4�ݬI)�wu�wu���`r�=��U�{P�/TI��Q(���`tD&�~_���ŀ�w�J�	D}
��	!R��x�$a ���| 0Z�1c$��)	!(硬.#.06V��� BJ��ᡢe".K��\T��	P��pM$�5V%�\�Y�)�!W�p�E @��cf���oD�f�
���v���f����;���fa
a
c.hC@ hl�@ F$���!#0��a.n�dd"�	�9�jB������.K�.����� L�XD$�B%eRT�X%��8��bH5
�2�£*K�5F4��	"Ơr����$d�!+�
��ⲑ��X`rX�$d�P!T�!*��ܒ��O�~F��P��#`A��
d�[��c
��-R`1LO�@��P��1n�CBV\�J�C�"1H���aF%aD�IXT�����a��b$H$) �������ff�U*�B����#�m���[���T�f⋚��=���Q����p���=g�,�tkdG�n�[Z��E΋a�ⱞۮ�Fyٜ�9f6���L�v�1��w,��z`�L�s����Q�������eBs�6cS=�HMU*� m�x����h�uS]���ݗHMýi���39,JMR�od:	y۩�3�9��Krn:�]ͣ�Hny`�
��13UT�h�Wcm�Hn:�l�\�pWWەm�Dz.z���d���tt,h���ۨN���˵���Y]<�	mg6FN�\l�M�؞��H⫀�%����X����T��a�� UWA��m�����p�i
W���n���ƇK����t�#=����ۭ����;<�Q�T@t��_o�xG�7�r��V�kb�u q�Y�u��&��S=�'�����)ڻ�m�i�"P�a W]֩ٝ�+�J�QS��xl�k(�Il���9��74��TbB�5vɐ���ZR�n�=�z�,�Y�ƍ�۠��1�4�m�m�[�q��Xr�ڍ��^�tf�W�����;13iڱɵ���FMbP��=*3��qù[�[��4�lvt�!UOaD��q�vv�NH5��u@�lV�!M�d9� �67
6�f\�h�N}q�4���g.�-�z���۶�� �l��h7L�ڭ�]B�[�`ݸ�iy�}�j��M�.�nM��P�Q@�IUWkI�@(�v�ã�gi�V탋R�S�,��=k�����-�0ۮ�i�ڸ�5�O��d���$v�X���$yB����Z�Nb[��g��(h���4�j�c�j�:�z���ؐ����j�w:�W��Rkm���:͝�m�����J,�/��۩4#<�6�'ʪ�ݹ7l�/�kv��P�9I6� T(����n�bG��kX��ȰDc���(�nW���g�լ����p:x'� Ed��,ѩ��wGg��w��1�l�c�պ�7bح[6�[M���:(����:�y���D� 8Q�p�� �!�ײ�ۛ�r]�u��n�)v9�ɞ{7I��nv#���9�@��m��AI���k_�����n�����s��¶��&�X�.Ǯ��o'�k\��ˋ���/=s�c<#.˖�q֊��d����[$8�K#��k�Ë�=�����B�m��l�����AkV�0��д�.��r��<�����"�n3�k�u^�{7E��I�n�N�{��]���];<�M)!Ζ� �I��:�Ҵ�AI���>�{��>�;���n������X��|�G��u�NGah�MZ�Uw3uk ��,����B��߾������7u�΄�H��|;��:j5Qʰ�ޖ��â!)��b�wb�Ѳ7JT���Ujn���:D����}� ��,}_%�{��ņ����Q8J��I%���С�w����x���i��CV���Y�$-��vT�m&x�t==����z�;gj���ܻ����F�Eb�>��L�D�:H�����L	��y��aB���RJ�n첾��d���O��(���O�g� ��ŀ6�,�BIL�蓪�L�(7 �Q�`��,�۫;T��۫ ��0	]	�VR��,1b��0;�b�o ~m�D(IL�w^ ��z�
�r��"Qʰ7wn���,wvX��V�n���%":�i�-9��-�y��Xrsf��jT�h�Y%��=1ȪS���Q�� ��� �ݖ�\������ŀ�'u)R���1U�X� �D����$����~�����Xo��*����I,�b�oZ���脢�5���n�9��͍ӑH��i�*��U�˻���wu����׊��w#��6)�)%X3��.��`w��Vn�Ձ�2iMT`��1W�u]�:��[������l��Q����e�dȍ�I:�r
%���,�۫������J���YJ�T�ŉf$�����GLl��t�0&���RNT�Qʰ3wn�{�,���$f͖�mՁ���qT�MA��suk �� ���u��iRIDZ��:�ջڰ�#u�ӧ$��)#��:H��:`t�� �"`z�%��H��t��yy㳖�p.��F��+�h�����sl��il�ܩ��;��N�����������t,��9��&�r��۫��_}Iou��׀=׋ �;��\�P"�f,���0	�&Ӣ`N��Ӷ���b5����6�(�rXnl�'tt���� �"`���VR��]uwWw�=׋ �/$�}�}����^ k�x����U	D#_������<֒�J%/&��5�"�)�L�#5���	c���eJ�Jra�P���nb�v��K����0�.�c"���b�D�d�\�`���J�Iv�sw#�����3�צ��H-�v䝰AW1��͜[=�;Ta]�<�E�/7V��G!s76O�mt즻8�wi��ۧN�C�v��r]2��&�ܴ��q�AWE���sp�=1�
h��n�^��X-�^.r������ܘ.'2�_����v��\p74w�����X ����w�	,�z���`���NکN��MDI*�7���}��$�^��,^�Y�)��j{��T���թ����ϯ {��С*��� �{����GQ@�J�#P�K�o�,��X ����w�~�HY��r)M8�X��V�{=����X��V�3t��29T&�B�Ա!��l���r��\jAQ�\��N���9���[q&�$��~�ߥ�f�� �^/Т�v�`h��534���Ss7Wx�]�$�Ī��x���`�w��B�O�V�]ں�n�RL����GL�D�:tL�h���I9JT�Qʰ3sn���,[w��BP��ߖ��f��Z�SeIWS7V��n��IF���u���7v��9Z�岜��S�'"661v㵮+v$�8%�W:�Ez#;6���	���9%')G���,�۫6GL�D��Ӡ���IRT�-	%�n�ŝ2>�ŀ���m����Z��"��ӎU���u`��e��������wn��o��M�P�TRRp����,7vX��V���}ʰ=�G��$�A�)D�`dL	U�0'tt�&Ș�v��q���PNH�M�
1ѹ��딜b�1�UgR[t:ӷ�7�kI^$����wGLl��M�07��7�J�r��"Qʰ73n�{������ŝ
"d�}3YR�R��,ł�T�>�Ll��;���V��[��9%')I���K��o$�w�p䓾������z %uNq0%��YJ�$�*W���`N� {� ?7x ����vS�4+.�� �%�k��-=��Dd瞻�]P�z�x�R�b�-t�3w�m��:`dLl��;��tVD��Ib��%Ll��M��]X�۫�}I�#���N�۔�����׀=׋Q	L��ŀ�׀���I	RYkbI�;���x�����w�?�ԩ��6�+���z:`dLoD����$Q4"���ޖ�)�ve���v�2�T l�DƴE�s�m���rTpe�n�uu�������ٔ8llgg�g�-jݬX5������Si�6��"G]�]D�<�常�����x���OX�ka�x��s�%���._��9��m��<�X���k�7�Մ]Fh�ѤV4��[q��E���mX���kb�sg�g�g�ދr�����$�v�뤷d��w��'���g���UK��uk<v	y�nu1�f�5[���\һ��^�0�l6�s̝s�d��n`�`z&z:`���Pt��)9JH��l����u���۾���ޖ,7bu	%8D�$����7���"`z&n��Jr(J�M��X�۫ ��� ~�x����`z��EP*��-�T�6H�މ��#�ތ����߲��u�ӆ�n\�fl)`��O�:�YZKW#��"@�DNm����KΠ۔�Q�������ݺ�7��V�ݖ��7�N�I*6���,�ۧ�^+0����"`z&V�Y?Jt���9RU��ͺ����l�37n��6��R�8��D�X� ���:`v�t�6��KFVV$��+V�&��0;�t�����;����q��i�S�8�q����u�w�)C�R�������l��k�5�{yR�,@��B���`wH���� ٻ?UW��X�J��䎥A��J��0�&��0;�:U��z#�J
q��U�w���nn�!P 0 �dR#��a1H)O1��"A!��X��`1!0�$a�#�$�#��`)�A=`3ҁpOA�x�� E(�$�����c))V��j.�@5Y�H����@�
�ဆ� �R����yO<���u���C�z"N�^�,�O �p��P�P8���� ��*<LT�u]U?'@�} 3��E�.��*'��?
/��}���Ձ��Kq����A7)D���ztL���=$L�����)RIx��&wGL�P`��g�;���;����n�t�A'%^.3w3���N�1�&�V�y�mی�U�˟Jt���9�U��ɥ�owe�sse���u`f����M2) �"`�wGL�P`�����ԒS�Q�`��`ff�Y�P�^�� =�ׇ�HRBڑ��.�.�͛r��ݩȖ%�b{���yı,N�w��"X�%�|�{�O"X����[�7��6�"X�%��{8K�t͛�M�s3sN'�,K��{*r%�bX������%�bX���v�"X�%���É�Kı/{7r�۠�6٢ȗt�iw&�����r�J��:]�g\��Nd�\.���ZmS�,Kľw��'�,KĽ�;�9ı,O}��O"X�%��n�T�Kı?d��gl..f�w&f�Ȗ%�b^��ڜ�bX�'}��O"X�%��n�T�Kı/w���%�bX����d�M��nn��ڜ�bX�'}��O"X�%��n�T�Kı/w���%�bX���v�"X�%���Ng]0�4�f�q<�bY���o>�9ı,K��}�O"X�%�{�wjr%�bX����q<�bX�'{نs)��e��6�ʜ�bX�%���x�D�,K�����Kı;���yı,N�w��"X�%���ĄJ6��	d"�!E��J��"�w��I3'	�f��|K�,�("�\s�:m��5��=�����r�+�ciݴPѧ���g����,�WOF�=�n�0:�ݤ��,�!)8طr*�g�ڥ���jv��Y� #,��e���L���u��;[;��z{q��6Chi8��X��X�3`h�8[�ҷ���y����ܻ(���E�#a2ż��8��������}��}�ͮ��y�x(�c�q1Ib�-�#qP����牪�6�����\��pvr��n�?D�,K��>ڜ�bX�'}��O"X�%��n�T�KıR���/�)!I
H[R7uEՅݪ��.��ڜ�bX�'}��O"X�%��n�T�Kı/w���%�bX���v�"X�%������3fm�f���Ӊ�Kı;��ʜ�bX�%���x�D�,K�����Kı;���yı,O}�,��.d�ni73w6T�Kı/{��yı,K�s�S�,K���{���%�bX���eND�,K�N��t���m��fn�<�bX�%�ݩȖ%�bw�{���%�bX���eND�,K��{�O"X�%��0���w4�.���ć:hh�1��I�Y�Л����I�z٨�'�K��]��kIQ��{��7����É�Kı;��ʜ�bX�%���x�D�,K�����Kı:~���3I�n۹�Ȗ%�bw۽�9
QO�S B�|�n*�*��r'�%�����yı,K��mND�,K���'�,K��{0�8f�f�ۛS�,KĽ���Ȗ%�b^��ڜ�c���>�~��yı,O�~�ND�,K�z^�����4ۻ����%�d��ߢlA>�~��$D���&�$�����'�,K��Y��dp��&�#�}V}H���#�����yı,N�{ʜ�bX�%���<�bX�%�ݩȖ%�b�O�������Fj���qq�C���O<�y�u����c��;V��vm�c๳Z��?'�,K����r�"X�%�|�{�O"X�%�{�wh|��&D�,N��xq<�bX�'{�,��.d�ni73wv�"X�%�|�{�O"X�%�{�wjr%�bX���|8�D�,K���"|)�2%��O�ٟX\6\ͳv���'�,KĿw>ڜ�bX�'���'�,x���B�W��I�-P0V��
��=,ND߮�J��bX�%�����yı,OsӸi��M�ٙ����ND�,K�}�Ȗ%�bw۽�9ı,K����<�bX"g�϶�"X�%����3�d��i4��w4�yı,N�w��"X�%��s�~�x��X�%�~�}�9ı,N��|8�D�,K�����m��ekM�f굉�G%�M��=�N�D�X#Y�z�L�2u�'gE��"X�%�{���'�,KĽ�;�9ı,N��|8 �L�bX�v�ҧ"X�%�/�]�a��f�ws7x�D�,K�����>P#�2%��{��Ȗ%�b}ۿJ��bX�%���x�D�,Kܳ��ɹ�L�4��f��ND�,K���'�,K��{*r%��,2&D�{����%�bX����S�,K���g	{n��6�ne�Ӊ�K���������*r%�bX�������%�bX���v�"X���X�T�@���Dz	�����zq<�bX�'{�+��̷�c����oq�����x�D�,K	�"W>�}�<�bX�'���O"X�%��n�T�K�q������� ULV���暇��tݲuЍ���������j�߾�����~1p�s6��37|O�,KĿw>ڜ�bX�'}��O"X�%��n�P�I�L�bX��~�x�D�,K���7d�i��33v�ݩȖ%�bw�{���ʡ��,O�w�S�,KĿ{����%�bX���v�"|��TȖ'ǿϝ0˻.��n�O"X�%��n�*r%�bX������%�bX���v�"X�%���É�Kı;;;i�˲a��3M��S�,K>D��}��<�bX�%�����Kı=���q<�bX(�2'ݼ�T�Kı/���7wL�n���'�,KĽ�;�9ı,?�=�~�q?D�,K���T�Kı/��w��Kı5a�!�ܛ�?���+sf����O2�A��1"���\:]+�)\��!��˰�u�S��6�ή�E���l�%�+O=�ꋵ%��vԋ�=��7�\/Bj���5�C."CkQnP�64���W:ܼ��=��׬].ᑶ��u�c��h�X�V���Gl%�rª�I\�L�X �(a�'d�[[l'\���f�٬B�*u����~�s��텼��.ۤ���{9tgs�}s��݇�Ju�.��)i�/�{������Ft��]�1}ߴ�X�%��~���yı,N�w��"X�%�|�{�O"X�%�{�wjr%�bX���p���3n�&�]�8�D�,K�����(!]��,K�����<�bX�%��?����&D�,N��xq<��"TȖ'����L���%��͕9ı,K���'�,KĽ�;�9ı,O}��O"X�%��n�T�Kı?d��gl..fٻr��Ȗ%� ���w>ڜ�bX�'{߼8�D�,K�n�T�K���?}����%�bX�gO��I����37m�ڜ�bX�'���'�,K��۽�9ı,K�{��yı,K�ݩȖ%�b'��[�36�f�)s-�f�6�ݞ����i�\�뮰pkys��ؙ���������2�MͷsO��Kı;�w�T�Kı/��w��Kı/��v�³șı;�����%�bX�O�̻֙&K�7f�ʜ�bX�%���<����;ı.{�ڜ�bX�'���Ȗ%�b~��ʜ��2%�/��a��f�v�n�<�bX�%�s�Ȗ%�b{���y���DȞ�w�S�,KĿ����yı,K	�̗\�K�vnn��K����ߎ'�,K���J��bX�%���<�bX2&w����Kı;���.��6�ne�Ӊ�Kı?v�eND�,K����x��X�%�{��jr%�bX���|8�D�,K��'��7&\h�t'J�4��ޗH��g�.5$�GY�����&/3��|�N͝n/��=�%�b_����yı,K�ݩȖ%�bw�{���%�bX��w��"X�%��'gs;ap�s6��37x�D�,K��wjrr&D�>�~��yı,O~���Ȗ%�b^��w��O�*dK���i0�svff�S�,K����É�Kı?v�eND��+�@�b�R!Uh؛��}�O"X�%�{��jr%�bX�?t�u�ܛt��w4�yĳ���=���S�,KĿ{����%�bX��s�S�,K�&D������%�bX�O���ͦ�L�fn�ݕ9ı,K�{��yı,?��{�mO"X�%����'�,K��۽�9ı,K�o[�3m��nlf�lek k\]�
�p�ŃZ�4�8^���i8/�����}=U��_��X�%�{��jr%�bX���|8�D�,K�n�T�Kı/��w��Kı,'��2\%�n�2��ݩȖ%�b{���y���bX����*r%�bX������yı,K�����Kı=�{�^˦��l��w4�yı,O���Ȗ%�b_;��Ȗ?C"dK�s�Ȗ%�bu�������$/it:��WWa5{���"X�%�|�{�O"X�%�{�ڜ�bX�'���'�,K���w�D�'��QB��_bwo<�9ı,O2{;���˙�n̹���%�bX���ݩȖ%�a�*{����~�bX�'����Ȗ%�b_;��Ȗ%�`�w��6�2˷��W-����ܽkS��'e���K�\��:�W79�s��b\_w��g�ı=���q<�bX�'�n�T�Kı/��w��?DȖ%�}�}�9ı,N��ɟ:i��n��n�O"X�%��۽�9�P�DȖ%���oȖ%�b_{�mND�,K�}�ȟ�S"X��I�3�M0�.�ݛ�*r%�bX���}�O"X�%�{�ڜ�bX�'���'�,K����ʜ�bX�%����ۆ7I�]���O"X�|"g�϶�"X�%����'�,K��۽�9İ>E���y�
HRB����EPM��%˻sv�"X�%���É�Kı?{w��"X�%�|�{�O"X�%�{�ڜ�bX�%�4`� ��Ј���"H�"F��K�&�"D�d���$�2�HH	$`��ES�Q���p��1��:@���E$"l�*D�$@��
���F*xH +h,�: �h:�$ �$���!
��(H$)�+(!XE E�BV5�\H��iD����z��T�+����!i)!F�����W�W�Հ1B	 	�E�;@y���x���F*DE�����yĈ{��I	�Æ"�"�2B��� �P�)FH�1�	���Ӥ��;m� i��c�I:8켭�MR�69�I*6���Xc����ٓ�(ض���+\޹M����s���՞�z�vn.t�+�uƷc�3�B&囔�Bd��g�KQ�wg��:���UF5U��g�m��*�0��]J���0q��U/8��g�X�]�j8+�ů�NQI����W��[���ˢ�ʺ��O,����-�ؗL��k�%.���]�I�,��$m*l's��іx������W��[���C�8M�֔��.���P	A��ƴ灌:��%�{\s�-���ΗqK�ƑM�l"�T��;MU�z�����,YiM��M<��)�<��km��Z��3�
�6`<d=�<5��Q�p"ʫ.��;�\�Iz�L9�N՛S
�`�YH��������)�|Y�bm���^�H�O*��*��6�'�Mr�D��3,��S�kfݞ�	l�lnC��m��n�+�'a%�s]jx�*���)���}�X債�p���<��3d��۲���@��\-� �mma޷<'�Rv�ل)8�;;���emWk��S5u]�Xx�r=;9���l��U{n���N��������N����3Fҝ�q%�yɕzZ{�
g�k4��d�[���s�Km*F�'J�ȕԴ�mt�.H\4�j;n7$�g�ͮ9���qs@Vʻ[z�*�9�ꪻmڍ��.�	��Hm4:vY/&ׂ�2zH�i&5SDqn�+i�廍�u��rh᭖r��D�=�m��+ʍ!U�ҧ4�`��4�F�7A��lHG]����x:"�66◳�Zr9x��8յ�k؛��� *,���Q:%�T�ԫT#c��p$�y��\j��5�=r��%lfմ� oXR��n�����kvc��Z7<�ӫ!��«ϓF�S�\��
����,�z�:W=,9�)j��D��zqƺԶZ3�g�7�2t��l+UU�uWl�����kR`9ras7r�s&nS32�(�?�h���@G���������8�"�z/�]x ��⯃��ٿ��enZd,�5�r���չ�v���.l�s�cF�����[��[$�g�W���!�,dפ�oU���:��g��Tqs�n���=��\ڶ��8�a��H鶖:��5�v�cl�Q�xrOoo*�9���:٤W$�E��j˱ѥp!�1�Ik:�6��u.�}�&؞�Va�+*��k
��@�!.զB������{��}��F]��UG�.�e7Q��v�q7h��WP��j��W6x�}�t��v>��MZ�Rn��[ŉbX��w�S�,Kľw��'�,KĿ�����V���,K����yı,N�7'�l����2����S�,Kľw��'�,KĿ���ND�,K�}�Ȗ%�b~��eND�Q2�D�=>�s>��l��v�˛�O"X�%�}�}�9ı,O}��O"X�%��۽�9ı,K�{��yı,K������\�ݹ��9ĳ���;����yı,O{w�S�,Kľw��'�,K�T�=�}�9ı,N��s>t�7&�ٛ�sN'�,K����ʜ�bX�%���<�bX�%��wjr%�bX���|8�D�,K�s�7�e��N+�8��x�9���[#p�Z�GuÛ�^w'h���}����w��[G?G\�qgvn��%�bX������yı,K�����Kı=���q<�bX�'�n�T�Kı/�����0��M2����yı,K�ݩ����	���Np�T|Dؖ'߼���yı,O�w�T�Kı/��w��O쩑,K	���3$�]�\�77jr%�bX��~��yı,Oݻ�S�,�a�2'���gȖ%�b^�>ڜ�bX�'����͒�M�8�D�,� dO~��T�Kı>�~�8�D�,K��wjr%�`

!s}吿��$)!oGU��*�ݙr��l�Ȗ%�bw?w���%�bX|�s��Kı>�~��yı,Oݻ�S�,K��~��|۷�e�� �Y��v�\Mr��B0!��$.���EŷAW9��=ab.�?{���D�,K�ݩȖ%�bw�{���%�bX��w�����M�bX������yı,O����6C77ffnۛ�9ı,N��|8�C�9"X��w�S�,K��=���yı,K�ݩȟ�S"X��s>t�7&�76��8�D�,K߮�*r%�bX����q<�c C}W��\G�����ȗ}��ND�,K���O"X�%���;L��L&K�7f�ʜ�bY�
��{����%�bX��϶�"X�%��}�Ȗ%�b~��ʜ�bX�%����ۆ7I�]���'�,Kľ��ڜ�bX��~�~�q?D�,K߮�*r%�bX�����yı,��m�˗2���^��8ٶY��R������l��k'5�{yR�R�ظ��Zh�}���X�'}��O"X�%���{*r%�bX�����yı,K�ݩȖ%�bw��	{.�nn��.��Ӊ�Kı?v�eND�,K��{�O"X�%�}�;�9ı,N��|8�D�^�{��7���ӿ[iۙ��Kc��Kı/����<�bX�%�����K��lM�����O"X�%���ҧ"X�%����2u�6��ܻ%��'�,Kľ��ڜ�bX�'}��O"X�%���{*r%�`q5EY�*
�(p ������'�,KĿ��͐�M�ٙ�����9ı,N��|8�D�,K�n�T�Kı/w���%�bX��s�S�,K�� _���Lϳ37l̒�nn�sG ��7Fjʙ�-���f��l��s���Ϲ��8�nM�nm��~ObX�%���ҧ"X�%�{���'�,Kľ��ڜ�bX�'}��O"X�%���;L��L&K�wn�ʜ�bX�%���x�C�U�L�b^�>ڜ�c�C"dO�߼8�D�,K߮�*r%�c�2&~:_��p���4˻����%�bX��϶�"X�%��}�Ȗ%�b~��ʜ�bX�%���x�D�,K�{�s&a.��%˳sv�"X�%��}�Ȗ%�b~��ʜ�bX�%���x�D�,K��wjr%�#�Gս��Z�G$ �d�����!,K�n�T�Kı/w���%�bX��s�S�,K���É�Kı ��ȓ��n\��3d�&-՟r���@���UMwn�g����۶�'��_y�ݰ]�^28u��Y��ۏ.��:��x�X/#���-�n]��J�s��6ô�z��Ӻ�x���l��<� �67g��ntkv�iW^J��$���ҷ]�ܑкi8J�	��)�+d�tv�{v�*�z֢�doa=�#�d�l��ۍOqX�k���D\���M�{������r�>�4μsی���#g��'��\�!J�r���lJ�Nsd��Nۛ�.]�͕?D�,K���8�D�,K��wjr%�bX����p>���ؖ%���ҧ"X�%���s'�m���t����%�bX��s�S��DH�L�b}�����%�bX��w�S�,K�����'�?�*dK�w�6C77r�n�f���Kı>�~��yı,Oݻ�S�,h�lN��u9�	�ݪH$������r幚��I�>��ןJ��bX�'����O"X�%�}�;�9ı,N��|8�D�,K��v�ͦ�L�f��ݕ9ı,N��|�yı,>�w����%�bX�w�xq<�bX�'���Ȗ%�by�{3ɤ��l6��QY�L3�\�nD�XP���D��kQVƲL�����}��oq����{�wjr%�bX����q<�bX�'�������7�M�bX������K����n߿����r�	i����,K���'�� `�Ȗ%���{*r%�bX������%�bX���ݩȟ TȖ'ޝ��d��n�i��ɻ�Ȗ%�b{ۿJ��bX�%���x�D�,K��;�9ı,N��|8�D�,K��rw6M���-˻���"X�|��2&}��oȖ%�b_{�mND�,K���'�,K����ʜ�bX�'㳼���s7r�7x�D�,K��;�9ı,>U?w�~8��X�%��n�*r%�bX�����yı,N�������72t���1��L�f6Z�L 
td��M3x[��'n&aswjr%�bX����q<�bX�'�n�T�Kı/w��� I�&D�,K�s�Ȗ%�b|{����ܛt��w4�yı,O����G"dK���oȖ%�b_{�mND�,K���'�>�A]�ؖ��S��M0�36nl��S�,KĿ����'�,KĿ���ND�� N*�TLP!�,N���8�D�,K�n�T�Kı/����.]�.�ws7x�D�,�`dL�����Kı>�~��yı,O���Ȗ%��"g����<�bX�%��o�s	�3t�.��ڜ�bX�'}��O"X�%�����}*yı,K��}�O"X�%�{�ڜ�bX�%����(%<sm��F��krÏ(wQ>��O\=[��:��ͥu���4����<�bX�'�n�T�Kı/w���%�bX���ݡ�O"dK�s}�d/�)!I
HZˣ���]]��f�fʜ�bX�%���x�C�c�2%�}�}�9ı,K�{��<�bX�'�n�T�O���ؖ'O��̷����n��.n�<�bX�%����9ı,K�}��<�bX�'�n�T�Kı/w���%�bX��N�!�i��s7%�ڜ�bY�*@ș�{��<�bX�'����Ȗ%�b^��w��K��C�T������<�3�S�,K���κa�M��72f��<�bX�'�n�T�Kİ��������Kı/~��Ȗ%�b^��w��Kı;��y�Dr=��XIn+X�l</,e��GpRl������4�&��s��i�R�"X�%�{���'�,Kľ��ڜ�bX�%��x$�"X�'�]�T�Kı/��~ϲ����w3w��Kı/��v�"X�%�{��'�,K��۽�9ı,K����<���>�"'59İ�r�e�&���ܻ77jr%�bX��￷��Kı?v�eND�,K��{�O"X�%�}�;�9ı,O�{��.I���re��'�,K> H߯>�9ı,K��}�O"X�%�}�;�9İ?�Y�3����yǍ�7���ӿ[iۙ��ǻ��2X�%���x�D�,K�G�Tk�}��S�Kı/��oȖ%�b~��ʜ�bX�'C�cR�w�%?x�(8����\˗���c7ZݙM�c����l�r���Ѫ���W(�m��%�a�'b�(��mh�ʷ�<�]���cm1����#��)+�l����x�Hu]X��{�ڸ�����Si0�gOMrJDg���sk^�%��V�X�7��-�jh7�چ2���,Y�]�uV�`{cg������nѻbvn�%˯�Bs���3.�ɰ����4n�ƌ�5咃=�I�v.9Y�mF��{ܥ�<fB尴��_߻���{��7���}�9ı,K�}��<�bX�'������șı/����<�bX�'���3I0�3ss.�sv�"X�%�{��'��H�L�b{�ߥND�,K���oȖ%�b_}��ND�TL��,O���|�]6鹷&n�Ȗ%�b{�ߥND�,K��{�O"X�%�}�;�9ı,K�}��<�bX��{N�i�&f�͛�*r%�bX�����yı,K�ݩȖ%�b^��w��K��@&D��ϥND�,K����.]�.�ws7x�D�,K��wjr%�bX�����yı,Oݻ�S�,KĽ���Ȗ%�`�w��wv�ܗM�Mʹ�s�˵�8Ӌ�b{�^���p�gS����������1�<�Ct%��w�{��"X�����yı,Oݻ�S�,KĽ����P'�ı/{�mND�,K���}�%�3w7!nL����%�bX��w��! $ ,@*�"�ʦ9bX����x�D�,K�����Kı/���x�D�L��,O~����7$3sw%����S�,KĿ����yı,K�ݩȖ?Ȑș��~�'�,K���J��bX�'�Og|�w&l��ܻ%��'�,Kľ��ڜ�bX�%����Ȗ%�b~��ʜ�bX�]�����x�D�,K�>?��$�4��̻m�ڜ�bX�%����Ȗ%�a�~��T�%�bX���}�O"X�%�}�;�9ı,O����?���a�[�usf�bN���o%-�Нts�9�N��46'��wg����ٺcsnf����%�bX����*r%�bX�����<�bX�%�����Kı/���x�D�,K��w�M0�f鹳weND�,K����'����M�b_���Ȗ%�b^����yı,Oݻ�S�,KĿ�e�;�.�L����O"X�%�}�;�9ı,K����'�~������~*��b��@���EKJ0b�b� ��p��H��B�0@���$5M��)�O3(�)�� L�� �C�,�*����T��X���a�~Ŋȇ�4`,�$A�b�Y�7$����6[�x��Ob�	������*�
~_1G����1�� 
q��*�G�N�b"p���O�<���S�,Kľ�����%�bX��or����n]���9ĳ�U?�hlM�~��'�,K�����S�,Kľ~�w��Kı/��v�"X�4���ك؅�#T�俫�ԏ�	b{�s�ND�,K� ?�k����x�ı,K��?��"X�%�~����%�bX��훓.����ݷ[���ԇ"CM��ދ����g�.�������cN��rBf��n��iȖ%�b_����<�bX�%�����Kı/���x�3�L�bX����'"X�%���~|~�Nl�%�������oq����v�"X�%�~����%�bX�����,Kľ~�w��O�2�D7����׫l�s2�ﷸ��{�K��x�D�,K�{�"r%�bX�����<�bX�%�����Kı;��g\0���������'�,K>��;߳�'"X�%�{����%�bX��s�S�,KEE��6�� ? 	��A� �"_w��yı,_���6�a���rm�"r%�bX�����<�bX�%��������$)���~��y� ������?nkVw62�9Z�v�\V8-qgNp]\T�8^k�_k@��{�~��<��b����	���`��GL�$�Q�ZӧNF�F�#��;��~��;�,��K ����׃؅�"T��9�4�wvY�������9��\$BR4�a��������0	���7z&�(07��i��ۑ�	�`��`{꯾Y�����������D"��(�ܯ� �Ûĳ
a�m��'��Ոg�D2֣��{�&�GNR���N����m`�췶�{�6Уn�[�;Y�i��oS�M�.y��ݷ3�������[�]r7@���໣�i�y���tF�v�]��0�{F�e2]�5��g��0nG���C��ʹ����]E��Fv�S�k�!��+��vs;sg���Ϟ���uNS����r
��v���֦κ��F���Z�N �.Z\h��BU.�@��v眧mD�����`sri`���W��`{ձ��N�*9rI`svـ����]�����EP�.���R�5NJ�B�3~��͖~I,������Q�bt�9)�jF�a�Uw:|�t�0=9A�{dL�f-iӧ#R�j�`�l�?W߾������K ���4�1��q��7
(���u�������J�l��)lP��ů�?���
rD�&�`sri`� ���D��3��bĲK�nl�y���z"�@?H��e�$f�����sd�;��I>��o sri`w�D֛Q�������x�k�9%>�|`���>N��S�)�Q$��6XܚX:��r����� �N뢕"캻*��� ��ـ}
'����� ��� ok(���n���9*���@�N�V�[a���a.)yܜ���#{�u[�y:���C �ȘoD�7z/�����7�<X�_�t�9)�jF��l�{]���0������j�iӧ#R�j�`��`srifU}J������]���GvaUws*f����J!O���� �n��_}�%���|=<�Fԑr��=�&��0މ�����?�W��~���0�$�:�h�nu�Ѧ�r˞u�Hڞ���K��ww��k�RW˥x��}>�Lw�`zr� ��,]�u��t�9#n$��{�K��D$�Os�0��x��y�
"�ܝ�|��!�F㐰;�,�ݖ~����G�� �w��[*݊�*�wj�f���n�}��{m�#""#� N���x����ql��:Z�'N�����nK ����$�n����|`�7x���O�NDᕘ��/)ʹ͌�Ү�����뜧S��պ�*]���-�Ж��m�[l�?=�`�7B�	|�D%��}vV����*I�n7&���� o���m�GB�
��,�U!I6bd �{��9�ps��ɥ���ZmD�m�����͘�����fB�
g��xN���E7)�q$�;ܚXܚX;�x��x�Q	ZIW���D�U�M�P4�q[��4;Z)E1�4���F��[�y��q�]�/j�m��®v�=���u��7�B�&M�\�ٳ�e��Y��T�ȃuj;dr\A҆!n�b�g�6�NN��[�{'F���c��w+a��F9�V�/nF��8뒓���z��٦�n��ms����#���\��\�֔��\�.y��>���?J5ʙ�㊞ ��vn
Ѧ����l�3��(�rr��{������V,�Y�8	�_�"`�w��r�T�T�MT��q) �we�o���m� ��ٝ	)����iR��Sj��� ����fB����g� �{��;F`�t��NTMB;�J��QM��~����n�{�,W]c؄Ɯ�*I�n7&��"`�w��UY��Cq�3�k����Ҝ�7�P&w������.�)4I���쑤�E���?2O���;z&�(0=9A����^e�3r�n�6��$����yA��(�7]�{������Jt��Ub�If`,I���NP`� ���kp�~��#���p��UK�G��7��0މ�_v(07���B�J�]ڹ���0���������_����XܚX�h�&�¢#M�F��˺�r���I
*�<:��5d�M��kj��܉ӥ$�)���3����ri`sri`��ј-*nS�PX�w������/���ɀv�LW]c؄Ɯ�*I�n7&�����x
��	���G�<�P|�����|������=��߷�O}�~,h�5�l)�"pn�.��&:|�������r�y������*䚻����9DGТ��?z~,�ݖ�<�J:�1��)��L��� �:� 6�r�5�;M���l�kJ��J)Ӕ���#���ri`sri`���B� =}x.e�E�E���*�ZCӔ�D�;z&�(?��UT��Z�z)�U$��JB�;�������;���=����J�w4��%V��� ������� B+EW _�����o$��wE�t7)ʉ�G%���������9��`��`w�F�n6����K��L8��7P[�q�S�\�{Z�ON13�:!uc���	�9T���,��Հs���;���U��<X��|�'E5$CX��0?�{'O�w���������QDԃ�NK ��Kw����=�&�]L����Uyw5H����(S���� ����Ks},}����D�DM8X܌��n�}��{m�(K�!
J����B��B��dN!��"H�Rb�#�xpA�B4 @eH0�e ĖP�ijD)+� RC�y@�!�.��N��XF$*Ec@�F�<XP? ���q�#�I�J���R(�	�D���F+  3KRfk0�).$)
E�����q͔�MX*��!��2�Y� �X��p ԚF� M=#Ǹ������� �Dt"��s����wwwwwwmؖ��X�yM�ث�fZ�bvN�UK�I<�LV�K�������ٙ�W+��5�g��ns���];����蜭Cc��Қ;k�Tap�^Miz;3����7:I�)��P�zk#H�����h������Z����Q�uJ�(j�@vˌVûs���d�7:��ə˝�OL�^iq����K(6�¼m��7��f�+�+1.`�j��᭡.:�����s�����ѹ�)8�IN��\���f;Iڹ�wl�۫iyӸٛ�vA��lH��lXk�hqΪ�u2˭��h���K�l��Pbm{pu��)Ke�gph$'vݕ����A�vz�.ֈ�Fa��� 7L��h
8(�;g�Z�pV�Ц��\t�m��0��۵mv���t�W���au+�����Ju�RI�X�Z
 j�����:�/c��ˡF�CY��n�.��eK�z-ƚ9C���pa�s�r��L�sn)5s;�"�T���Q᝞n9�Cs���0=mN�tpǳٮ$	:%��g��k%��y�xΑ�Uյ vs]��{[�6�;�-u\��!m�l�W&-nD-��5*dܱdc�*�����kr=���vs��ƔA��h5����b��V�����wM��K*��V�+\n���=�ڴ��NQ�;d��V:�fyq���v�������K;��E�vS�W+��nK^�ت���N��3�-���\\���pclaVӵ��wN�nw �IlӅ;q�0 ����W8l�l�8u@T8�u`�z8��P�Ӷ�j8��ڕ�4���@7ZI�ƹ��+j���%�"9�	2-�V�Z��,��lTm���*��xHij]�<�I@��m=\���IF���PسVv�-`ݱ� �-�زT.ۭ��8�Wp6�8����ʍ�Q4�"�!��3�Kt[��q�3�6��u�Fx�6@)zY��[Uc�:U�=��uu�ڠpN�S�r�z #�]�TX�x��8!��P"�AZ���
����fgi3r�&Nv��E��K�nI�2]�rc��W85�o\�(M���P��\<��v89��-u�	��ڸ�9ܙ{N����׭dnm�, VI�iQ�����}����czN�trc���)z�֬�ظ�EYƐ�x��� :�����*:�F�ƤӘ��k7�M�9i^�M�¼Ż-m�GWc^���ې�����rA�;C�&�n߽۽�{������������2�wJ������ka��E��wgf��f䆴�+	cU��MT��q) �{e�gse�����В�(�Po���+��T���j��$�;z&�(0=9A�{dO��U�A�n�4��r�j�`fl�`sri`���l�9]u�br5*f��Y��DB�s�0��x��x����Y�~,�u�p���!���=�&��07yA����L��R�v���q�S�`;i(\�hD���#v��{��s~����Z����*�Ixt�07yA��������+�j���NRr&�K�ɥ�U~�H!$#F���� �5�H�����/�� ?}���]�(P�L���E*�T�"&�,�g� �we�s3e������1T�T�MT��q) �u� ~�w�{�l��	D��� �a5��:t��Jr)%�s3e������� ?y��>J!(�9�E��t)���kv;s���˻\\[{�]n��a�ں�Z�*���8����NTMH��w��`~ݶ`�7%
?Ho� ��N��4�iRN�p�9�4�wvX36`��3�
d�)>�	�"��K��3g$���}��O=����
ԩb(�%	t�n;� ׷��m�������Ҳ�L��07yA����B�(JV���~�_R���V���]�L�P`{�A�{dL��06w�6Xȗ��ө��n��j�n�D�mu$����us�z�)����v����=��2X�#�l��{dL��07yA�ݬU6)�U$�q' �we�7]���0۶��	(S'K	N�擥�"�Xw},�&�~������<Xsޖ�3��7)ʉ�����ـ~ݶ`�7x�IZ���@��C37�o$��{�۲]�sw.��)f!����0މ����}������4��MqT��G[%�D���x��j�F�.ۏ����c\Ͱ�I�q7 w=�`��`w�4��}U�ݞ,͞I�>L�)q
I`�w��(�&�0s�0����}�6g���NRr&�Kw��`~{l��2{{� <�^ �[t�"�G�B�˻���;���fl��	/�T�~��˥_�+T�U��5s8��0?�^����|0=ܠ�H���4�R!,������3��bڵɒ��X���Q��W1v^��z쩏VN�(��B�;tA�O�8�x:\f�.ݠ
r�]XsJb�ج�!<W�[�9���ݵ��ũԽ����n\5L����sx�F���%�\�����ś����Hܱ٧���h�{Liz� �d4���(�RS`KAR�4UЩ�O�v�]�[rmۮ�G-����O��ǩ�5�i����7#X1ָ�v3v�c#��4�8^���D�M���N�(�)JE$��~�{�K��O�q����e�y4�r��J�&�(0=ܠ�=�&���䭐r4�'Q�X̚X6D�=�w��+� �
ň�fbĩ�{dLwD�����,�扵)E���$�fl�?�Q�8���0����l˺��N'���������rn^״f�t�=�\�Ѣ�q���FeN�����z�m�_����D�=�T�Y+(ʻ�sl�ͻ��O=�{9���(h
�D(T�}A�� ;~��{m���SaR�5RH'p�wvX36X�M,fM,X
��N�(�9I�{�&�(0=ܠ�=�&�f%��n2A�"rX�M,fM,�ݖ�͖sT�M:j�r�E\]Vֹ�t%����]T���嘽��(�&��m�tN���ӑ�I:����d��9��`��`w�4�9���0�.�� ���>���{�^���yVz�Dڔ��	q
I`���~���rp�F��!������ �論��k����$M�NF�(0$��{dLN��*p��'*8�R�mՀs���7se�����3��P���(#Q�۶$o(�6�3�Ф+��j�';����\n��:��N��$j9V��� �͖{�Kw6��4�U�bt�(&����y�2{i�z�`�m_BJ&C�f���n2A�"rX͞,�۫ �we�n���ܕ��Q��)WUfB����Ｐ_�^ 7��"<�S��1Z�!�swo���n�	�8���RJ�wv0	:&�(0$���&<J�`.�����������t��Y���^u�͇CvW�ŵB7?%��)��''@?~��{�l�׋�����J�]b)b�I^e+Ę�������0���H�{H�R�Iʎ"I���oΘ��`tL�P`l��Q��P�
5�����7se������T���*�<h*��:��lq���w�{�l�7�l�?O�� Q.��w��2m��T?2�+�ݎ%��Vs���h�3�ͻh61Q�;1X��sy�l���&m�����'�!��UE ��W���8ЧV���{M���P3���F��:�t9�Om�7ZXy�IM��۩���!��6�k�|ػY�M����ƘH�3l�T�d�V�;��Mt���m9y%�����i��>��1�o���n_�m5���P[6�0���{ߟ[��Q,>qs.�J�)��\Pù�J��m�&t��x����չ�ݨ!6YՕ���{|`�`���ДG����,�^�r4�'Q�XܚX]�v�͖{�K�:�p
q����?O�� ���СB�""*����=����y�mJM%!ܤ�v��07yA���^Ɍ�.�D*�5w5J��{m��G����@ſ�; ��� �r��Ӓ�hs��8i�	����k�SR)�\8�!�*?�#�(t��"M4�`gri`qww�D�����J��В-M���O/��9�"�@��U
�ǌ�X����&�����+��*y�W�A�'�y��[����9$�<_�����ЫW�c�&���;ϯ ��ه(��/]�zw����KS�NAʉ���ߪ�����������8�����,WrV��NF���W�`v�ײc ����`Z��J�U)�T�$r8G#�v��w)�]@���J�V����
�,�ǻ����%�S�Q��8V{��9����d������μ�6�&���7))�su���f��f�u��I(�����Ҋt�'"nrX�<XܚX�SR�	�B��I��:@�#8h`a��	��#s],(��@�%YYZZ�L��%IV%`J�,"�p�aJ��RjY�x�(B���
�B���)�� ���!K�2�Z�dGN���A�x�W^+��	v'�J�a��bB$Y)�	pbI#�Ub��_QPEP�EA�$��:_��@� '�t<Mz���_��t�9�; ���~�#ڔ:R�4:� �m� �:�`��:!$��yŁ��U=���P������`���=�l�7�l�>I(���J��ۮ%]����&)�V�gqZ(ԙx�)�E5d�͆��k�J\�<<ګ��=ϯ ��f��g%�(P��}x�~�_��NAʉ��������� �0N���ت$(�I]�4��0��0|���D%'����,`�5�L�#p���U)��׀�׀=�fL(J&!$=w���l�M�I��!�'%�sse��(��w~����0���5��-89�1;���G0��8���#ۦ1�N�"��M76C���ޗ��۝.]�\}$���P`tLӢ`o���I�컹�UUf��f}�T>��?{��7�4���G��^��:jAYsV`k���]��	)��|`\�`6�X�6:��l�I,?UU}�����`}�|0;yA�M��:�[�M�r�jD�?{v�pwv�p����$��{��u�EJ~*�����?�96z�z]p󎸤n�+-ų�5݆z���X9�`�
�N��ջ`{\�;sֺv����c��w���P�q��'���ݒr���Ѓ�#��V����y�a�=�����{>�G=[7\����u��h%�O
������8랉�Z��y�p.���K�kK������^�8����s�ڻ:�m�M��'ku���&�!�����]��}�c��`Sh���bŪ��oLv{l�;C����l]��v��੹R@�����2'��4��w��]�%	$�Hv�� �)>pG&�n�͖�͖�&�3&���֛Q4��#q$����x��0�J""g�� v��bZt�
����U�U��I)�y��/�7�`ߧ%*2�"��iUU���f�J{__�7����������#��Gt��8�6n+�Fv-��+f�xum�j4��*R;2]A�� t�I �I���^�����XݚXܚXL��[H�'Q9%�~z�-%{j��B�D(��o��[���|����x ��>�\)��i�f�f� �`�`�`���s��� � � � ������ ؃��A� �o~��x ������� � � � �;��d�&]ݸK�.l���ll_��A�������lllo{���A�6667���x ���ϧ �`�`�`���N��%�2nl�噹���A�A�A�A��߷��A�A�A�A������ � � � ���}8 ����|�����M��*�+uў.��2.�r�T����Fî.x�M�q�u�s}���U�)�sm���� � � � ߻���� � � � ���}8 ����|������~�>A����ϴ�%��͓3w��A�A�A�A����pA�#��� �l�������lll{���8 ��~�x �F����ݜύ&4��s2��>A������� �`�`�`��{߳��A��	؅຃ �� ߼���A�666>��}8 ��;O�۲a��ݙ�n��� � ؿ��D� �{��pA�6667�������lll}��}8 ����|�����t�v����-�n�� �`�`�`�~��o �`�`�b�����pA�666?w�8 �s߾�>A�������������x��G`�9{^q�����Ň���튎T�s0ͺ��<�!���J�����666=��?�"b�`�`��~�Â�A�A�A�A�=�����lllo������lll����.ɛ���̛sg �`�`�`��~�Â�,ll}�~�8 ��~�x �}��N>A����f��6K�d��-�nn�|�������g �`�`�`�~��o �b�D�A�������lll�������lll}=���s.ܶ���rM��>A��� H*�s�������lll{��N>A������� �`�`��VA\���$�"�?8���~Ϲ�8 �\��}�0�.n�l���|������ϧ �`�`�b��X��ＱBQ�B������}׀{v��a�:��N����W�ٺ�6�N��ׯGc��>z�G��ǯ���vxn� �}��Ɍt������MT��p�:�����,�f�s&��RX�ȇR:I�$��?kw�{�ه�#�������ՀF�Z��9Q5"rX��,�M,�� �n��ݕ�P�8�n��sV`ݶ`DB������x����MA�X���A#Q/���k����f1q���%��e3�vg��75���\�k�n�\7Ƽ��ώmӓ�l��ט��0s�Z9�q�r����pg����z�R7m�	��V���:����C9�k]Ͷɜg�l(��"Ŵ��spOi
��6�縵��/�gX�L�8�ŋZK�Ժ��ƺ��-��EN��� O����-֮��s�)�l����)74ɖ�ˀ+���'Tݪ�%�K����\���쵺��]�Rp��}���ƫ�m�gM�&e�����"`n��(06���҉�R$�JG`����ٻ�~,����:�����ǲ�u9�^$�݊�����1�vȘ��ԡ�r��4Ӆ��ɥ����`�&�P`wu�Yt�F`,C�d��"`l��P`z�<�ex���Z�r=]�֍q�{��è^p�X���<���Q����$��vȘ9A���>�����`�s=5!Uj�\��uw�y�<����IB����� �7x���\�8�n�h�w&�.�?$n{���l�`sGY�`〔C��ϧ��'}�`t��P`uw+���i)	pJG`��`wri`wri`b��=�UU{Ox��(�4�,=���f�@�덧��� �esV��S���)JQN�'"q4���,�M,]�{\@nk�gۄ{R�Iʒ	�b��o���;dL�����Y����Rp�5g��;�,!D�(@�1B�InU7x`�`�X٪D:��N�$v�ݖ�m���0>P�">���Հ�S����9Q5�7�4�;�4�5w5�wvX�PZ�4����R4����y�m;�X�֭L��ܙ�}��-Z�U��e�����#tӨ�,�M,]�v�ݖ�&�4u��&�M8X}���A�u����<�ـ4���
%!"n	H�;�,�M,�M,]�vz5K�S�	Ș���~�f�����DJ!D$$�� ��C߸U�����������#��,�M,]�v�ݖ�&��0����MJC$j�^��
7��͂��ma�u�բN��!�n�Y�)��*jE! GWs]�gwe��ɧ� �l�`��g��u#��(�I�vȘyA���J7�:�$I�G%��٥��ɥ�nf� ����+eEG$tӨ����'tL�D�����0dphq��73e�gwe�����0�J��RBE%"U�P%�#a$bT�!V��ľ),��<&�����$L)���Tԃ`ȍ�!B	v^��@1�1%Q�H�h\�"Ӥ�CA:�j1�H�Q��X' |����cj� �,F$�[����$P�]X���`Pb�@��"B!M4d�,$�r��c��!?e��
�͗5)K7g���,�S�_����	�CR
�P��Hf�`P80vY� >@*D3�w�@�*�UUj��퐄�f6:ɂ��)�!��ۄ²�P�Ϸ��`�э�f��0s���i���7>7#��ϮC0�T0�'YA˚�P9���;=����p۲���\N1T�7n��0��ר�ެ��8Viƥk�A�x*�k��c�6j��g���N0��C�� q.��=�\�u��c��Y��7m��n�Ѱ>�t�t�H#n�/B�b:m�[�S�l	��[��'�Z�^8d��r(��;m��K�[��6�6vU���Ɯb6ٛs�vf-�
ݻrfk֥U��$Z�6z1�ct��W(�Ż5clU�`�pې�TbYx�l�/7mm��M�I�5�{$؉�ζ
�öK�+�!�<V��[P�@(Ѹâ��W<��܄�-�nruG n�kb*�V��I�ڥNdv��&Г!K�	��e��ZD ���x;��v\���tm�q�F�m��IƲ"�m��}��@�����vˊ{���B�6�م3\T6ヴC���}�A�5��e�\��6��.����I��^mbA+D���';_nul|��{��y�����n�B��;I�c��h��&�;d�q�n�O;.T�#��atZN�ŋ�}�	���h㗮���m��[�ɮ�^�ʮa�;W;]g�<����LLpW�\c]�q`�e��1���ʑ�tM:��=B�5Ӧ���y7#�Y�B�U`��������rv�����Y��BV	RF2�1gav�١�َ��tQ��m��V�쁪j�Xpl��/NkK�΃�����]m*�i��5�i|qw���s��jmlu��
S+pmv���6�O�2� *�Tw���rwʘt�n���&U��q
�E2Hۢ�z��5N譬`�%(�5�1���VKَ�u6'm�F1�E�l��\����h��+l��hY{[�;'M�a�C�N�r�A�6��z{m�ڽ��h���2�WV���'p�,�6��r����s�q b
��Xz��uVx�Pw�8�Q_��D�(��U�D����7
��q1C��v"4��u�������[Y�qO(�Tm�C�yR9�9Pql�N�p�ݤKh�䰚;[���Ӌ\�-�R7oWR��l�4bW���v�8�6���即�ϓ�����7\�E��N�/���̊5�7m�Y�h��
��A�����	�R�C�hn���Y�*�ˮ̦رŽ8�b��āu����	{i�l��vnf�i�s刻y��w7n��O���|`B�u�bw��U]W�|X����CvW�ŷB7?�+LPi)	q(������&��P`�&��_QYH&��jj� ~v��Q
ɼ� ��X3v_������G�:nT�N�p�5�� �:&O>��;z����]�
��2HE!`���9��`ovia��fߋ �Vk<�C�$�J����n��Dv�q��|`�w����ߟ����]�.`z(�dv��l�7m;j��a�OIp��!��&�gB՛��%w���L	�A���\��6X�<6TU*&���,�&��M"a����Y�����w�����M/�Gtu�pG&�,����=�&o(07yA�')��Օ37e��XM��tB��!D*�}xϧ���ri`o^j�2�i`�~u9Vf$����P`MΖ�=�&��o�~N�.L�v�g��q9��n�y��ź^*�x�챂9 �ͦ��%��U5f�m� ~�s����_�;vx�=���SR)RHG��y��=�o(0;s��
���1+2�Қ�f��p��x��RB�Q�D)@A�\�Q�FJ/
T(%��""�;���<����e�H����j���9D|�Q[�~�O����Ζ�=:&�2RYDRI)�F�`gri`~�������G��},�M,+Q�:lU)�PJ���a�8l��Mƭb3������O^�U�l���W��D�n`��$ӍÀyf���D���w(0&�L�V��H�7D��36_��#ٳŁ��Ł�����]������N!�,�M0��0�����}X�}x����C�$I�n�幷�����?w��0V�=:/���'$���ֻP5$qIQ8X����_|����͞,�&��Bڧ
���&bJ�lr��GM�Xe�Q��E�LKT�+n�t�&���t���`��7�4�;ܚX����n%�t9RH������m��7]�t����n_ꯩ#�ǥIN�$��u�����/zc �ȘyA��2�b�dpi��`j�k�wvXܚX�M,`�&�
BD�G`�w�r]�8��0>�X�	#_�����\�72书�ۚ\Q��5��Q���[[Q�\㓒i��K�#�i�n�䜋�Ƽ�m0���p��'g�5�[vI��ȸ�k�8n�<��x��]yf�dB�����Yf����}��q��&��J�eκc�Z�qڂ�1���r�f�L����.�c`��
L]���γ��m�M�k,�v��0�aU���b�ٷ6aw6��d7$t̞��L��v��9\71N�b���9�uH�q��N�#Hi4ܖ�M��{Y�筆�5�P��_�P`Kޘ�=�&Wv�ڀ�r��9Q8X�M/�IY�v�����ɥ��b�v�*jE!%+�0%�L`�Ӕ���++��R!Ԏ�bR8��ݖ7&����興K��}�`G�3����X�k�I����P`u�L`��;ך��n(�ҔEN���A��C���]��c�轋6�!wK�m�ש��8��dn�pn{�Ks]�s��������GY�`��$Ӎ����ט�Q����}�^ �_���l�9�X���T)	t���9��`sri`s�4�1w5�ѪZ:ߜ(NE��I�׿G����׽1�{dL��=��*I�n{�K�կ7π�zXܚX�&�TN*�8��7ۥ8;^*�K�w(V�[F nHy��Y)�QTq@T9$�J������`�Ӕ����
���+2��M�H��,nM,�&�.� �j�j9RH(�nK��K	�����QOER*T��M\B����塭�]�w���9�zl��)#��M������`j��wvXܚX��5�L�q8�]�v����{����v���Z+:�&��G`t�����H]�tnf��â;<Ӧ��y/$v�I��)حJ�)�m���&�$�`n�K`m�L`u^��+~p�9�NK�{��������9��`ewj=��*I�7)X��0O��2{{� ��r�Z�Mڀ�rHG�,?}UT����sޜ�y�;��M� C��UU���9�~V\��yH�R:M�H�wvX�ݥ`w�5X]�v��f����!<1�ۊ���Y{]����C��ۊ�(	])2͹&����0�$����5��V��Ζ��ޘ�=�&�2R�C���'r��޼�`uw5�;�,u�Ұ9��k��28!6�qX]�v���=��w�J��{�`sY��i�B��7�v����{���������]�����N!9ܒ����-���1�{dL	^���T�"�b����@��>/ӟ��m�L�4�as]����#y똥�u��Ǟ'(K��u.�v,s��;]�[{�c�N�j��\�,�4��u��l��7�`J�������֊rr�vw�d9���5v��F�s�9��n���Zk0F�Ű��Ɠ�ܿ}v��bv�q��q�ؒK%fs��4vԜj�  p-�;��[�TZ;�n�p8�;����[���]�������@?�?l�[XnΤ�œ�)�bm��5�щ�HA>���5��ճۖ)mN9�麐..ο�'������u�����6� ֶS�PI�#������A�������Vz�U���H+3���t���`�|��ұ���-�׽1�m�jj�*Iܑ�a����]~�S�7i��>�X��Q3��x�+��jP�q�M�9N��vi`~������3ޖ�Ӱ%n[5���8:�B�QZ���]N�Oe�z���.��O�O�~�v4�:�@L�Q�t7� s�����R�s�0�9����m
@��6��$�~�w�� � �2�KmV�v�g��>�JdjvN�]'"q$�:���`ff�X�����,��G�JBI��)��0:��0I�:V0$������!J9V.��|��zp�o����ViQ�ܦ騏��q��m�R)s5^�����%�'��5���q:R!Ԏ�bR8���,-ͧ`ff�X����f���$$�����t�`.�ޘ�=$O����ޡ��8�n�pNS�7w�V.��'t< �
b zp!1�HA���
jB���-HRU�Iׂ�� A�FA�@���W�2�4 ���C����!�"^7@�ÊP�i��B�㱁,@��X"�`��	�(&*A�D"B �}P��O 0S�ʷ�$	E�0%!`�RX�"��}	��H2��Ѕˀ̠6ʤ���2�1�HFI7W]���S��w�J�H��F$We �VH�!(A� &{�e�]�	��@�Z �Z������AR(��z�.U�QQ�>�������Dߐݟ��o$����9$�G[�`����rJ��UW�^o��w���8�6���������j�!nH��ݖ諭���� ���`b�k�p�9#���(Ф����36x��׎��x9�n�*�a��/nt��46��Br'NNչ���f�.��}U�g�,��G���$i�ӕX��ϵ� {���^�Y���l��ʿ;PI������쉁�+�A�uoVA+2�t�#j8��ݖ�Ӱ;ݚX~��!���`�$#@�+�S�������t�}z�a*I��9,�ݎ��_UUfz�pY�v������+���(�2���<�&�Ʈ8���ipnL�>�[�$����Pء��M��|3�Ł׽1�nȘ�"��r�H/�IUE�Y�l�]g�2�׀=���٥�ŵ��i��Q�E#���$X�݊����%�8P�#�'%��{����,]�X(J�
UM���}Ү��*WE����1%�ؠ��ޘ�7dL��w9$���+�����`m1zF��HB rP��r�U�x��o[usC\�ܔ�ר\��P�i��Kj�p[�8���r6wH��FX.Ke�ѧ9ڤ��=�t�a;����p��rT�ypL�(t�6����d�s��3�=��n�n��E�4E��R�������>��:�$�n[+��cl2��sX�� ��[lu��[s��z{�#��XN�����T��M�6�����/N���X�p6����')�l!���v��*j(
�$�p�B����; ݑ0;rE�lP`[ՐJ̤��������{]��BQ	L�k�� ���`b�k�1e�����A�,�7u�~�a�	L��Հ�� ��V�H�8�n�n'#�9ݚX�����xB������R�	���ۉ�X����͖u��`w�4�5n�D��+i)hI�Ꮂ�\�Ts,���k^4n
㫛��]�:���2�v%BWhV�x���$X�݊]�vR�5=
p�8GNK:�fs��T�wG�p|T
"��'<�8X�|��ݖ�*�e�2IˬĖ07b��zc ݑ0;rE�n%Z�@T9$#�R.� ݑ0;rE�ؠ�:�����Ie]QuSuu��w�t(P��ϕ~w��s]���q����1Jt*m�M��BZ�Nkr�7F�Ʌ�}�n��M��cf$^%2H��Q�`qnm;�٥�����;��`s�=�@rH�6���`{�ـl�]`�7x�z�g���� �|�&�m��X�|����%V"�T�$	H�"#��Ԕ)I��|� �}�����)(�(E#�wvX[�N��ri`b�k�3���N'���~��V�B�������ǀ�}�`;�,�����*1�ʍ�Di���qr�pf�\1s��n�������cKO2�-v�$����S�;ܚX����ݖ�Ӱ7q*�jP�9$#�RO�� ~�w�~��V�m�:!% �k<�C�&�ڎ;����p�o���M,]�v�XkJ��S�r������=��8ϵ��@�Q"�1	dF�j35�^����W7t*����`�k���K�B�}�x7��`qnm;�|���xt�D� �Ym4�{g���q�X����$#��zssқ���&�t〘2IHm�8���; �we�Ź������|���oͦ0RQ"P�G`��8�6��޼�`b�k���URF�����BpR1�,�|� ��\���˝}X������E:��F�Q�v�M,]�v ���t(Q	O��*�;���ɴJ��B8���1w5���ޜ�����0B��+�&"3d�TJ��-e�:�P�<��vӵ� �Qd8�\��ŷ<0s��gk���Z��]��p���q�`������q�y��V���a�#������3���;kHt�'"���YkJ�g�i���7^c�.t$���>Q�iS�:5A��[OF!#�3����8����Q4-����󦒺��y�IFv���"��[�#7�F�V�)�?|@眔�M�f�n�.q����o4t���X�ݮ*��
�4Qji)�(�R:M��x�߽,-ͪ�����%�Aξ� 󓧁M��c%7#rX[�N��ͺ�1w5��v_ﾯ�H�P�/:R2�pnS�9�ŀl�]a�;{� ���X��\��JCm�%X���{�,-ͧ`nf�X6�=i1��������� �%	z���s}� ���;�M�4�����NS�FH��Vݹc%H�S�I�����WBp��^l����vM]Wx�z�`u��6}���
�zX�J����FI �q�v���g:�C�E
X߀ z�K��+�; ��`qnm;w�V�
��H�"p�1w5�{�,�U}�]^�S�3=<XWr��Ԏ�b��; ݑ0=s�cv(0:��0�u��$L)�������v{�Ks]��K3ޖ+2o��m��6JEF�t���g�O/)ײ]mǓi�&˴P�p<Wlxo��Uu#��#)��>���~,]�v����si���u�L$�<�f!�׽1�nȘ�ұ���� ��'�&0RP�P�G`��`r�ޙȧ�D�$�"�0i�O��t��7��rI�����-OA�D��q��8�6���;f��u��(Q[�׀v��s�E:�)!q�v{�Ks]�w������vs)M�qS��I��3���=x��`詙�w9荅����́-g��wz���թB�䐎HpY�v����si���V�ܧ�@u#����uu��w�D(�2zy�w��s]�wQ�H�ƢL��Q�`qnj��v�:""&\������?yǆ�6��33ff��>Q�;��?�$�^����O߻��xAU>_��U}��~�`wG^�1�@�#h`u�L`�&�t�`n�����CEg]��=��}���ڳ6/7�n�n�.e�v��o�"r2
v+���WX�7x�z�`�|�D/�!%�-��`g����"(��M(�8�5V|�"d���9�Հ���{2�\�qIێS�9ܚX����͖�Ӱ7q*�jP�9$#�)�B�.��`�����U��J�nߋ �ͧ�D:��t�Dq�;�,�J!R^9���X����?�" TW��TTW��U��U�����*���򪊊������Ҫ ����R*!  �Qb"�1 �D�"E�1DP_�*��������򪊊�����TTW�U��TTW��QQ_�UEE�U��TTW��QQ_ʨ����(+$�k9��y >E+0
 ?��d��.;��IA@ @   �        ̀( J 8�@�T!�4��}�)@Q )B�A@E%B�@ !HQ �$��P � #�   ;u��   t$�Q��}��{������>���}��@��&�v��I$�-����� 죚��5W\z�oUT���UɮY�0` zwf�s �:}�  ���Q��@ ��Q����ҥ|}�Ϡ��=���n�p:w}��]@́���9<�m�_`��z}�  �=�{w�ࠣ���zy�!��ɞ�h)麅Z�A���}�&@0 >���}�T�h f�͒�U{����Cw�<����%R�v�۸�1�1����[���|z�|٬�8 �`�{���,�)K,�zisPl�QKX�:n
`R���(f���0:QN�t  ە�� 
�M�����J ��JQ�)@��P=��J���JPb})K��A��(���P��R���@P}��   �s����q҂\/{zá���i���@�UR�n  � x}�t���O�`8 ���[j� ��(���S�'��=�G����z���'�1�^��S �6  G��O6r���������^cs�����%w�r} M� "~��ڔ�"b B'�UJP�@��U*�~S�H  ���5IOiU)�@��T�i)H  !2��" 3S��T����������?�=�������TW����
��AS�Q_�
���Eb��
���O�j?��b\�VH�dW ��&�ǿ�[7���#/$V�5���h��!��0�
a&14t�%���ltP���Y�I��F��7&����f��6��%%/)<��eg~��=O	�Y�!�m�3�,�'P#���Y۔��4���M!�4�D��a�#Hd(i�ahAN<���l�1�^�O��2Fr�(�R ��ѭT����U�2��O��"�X#D#O�b&!�cW���7�# �\ީ�B	��i#pѠ��3F�I*֐�N�`@ F�8�a��	:�uN��&�05��F��	sxR�"��H�ٚ4��`IA�	
�M0*��#LcLjB������0�+���Cj�x��h`	
����D�m�@���n���Sr�4���2CAu#��2��cHBB��A� F��D�K7R)&��B-1)�B@�Y4�foy����I!#�)����LI	CX@����B|�ʍ H�2`d��;�>�� �6&φ\�F��-$"� P<�b�0�B�JK B5��pѶ]M��	��$���J��+��sf�B͐ٱ��$)���E��"G!b]3.\5`K�p�
C,�5KX�T�"D�X�P�"M;�+�a�	Z��A�'AC��iļ;qv�i��6l�f��l�۹�fc��
B��B�+�v$@�mat? �š��9N�4[4oD�ċh[��M�&���K����1�j�!A��X�:�tE`0.M��l0�%0��bI]!�"R�uH�����xS�Į4��9��4�jHh�KĔH�q��-
��j5ģ�c\T�@�V,�jv \4����8l�����B$ I�t�3d.�fZ��������!%2S[c�m�#)�s�FNBFa��%O�}�L,
��e��Yh��3�i�'6k��n��ַ�o��aT���6�k7���L5��*B�� �����>~H0V5!L�f�ٷ�+����L�Lp��:�g\��Q�s�����7�!Lл6�4ׁ�Ħ:�b�c�
iaV0׃Ft���i:ơ�(G�� tP��H2�e)�gH�st8�	>@�R:���:�)q��d����~�Ѐ��s|4l5��kz�/�x:�~a:�(a����\�&�ψX�L��eX�6$�@�R4�P�i(Jdjc��|�i����n%�������t�<���jH�Drtcp5�bQ��8K��|HS�D�N�P1֍�5����S5��P��$���8o��)�N%ٚv$.&�����F$�σ�D���ٵ#L4)��1J$Z.��p`WҦ̺.�Ng�*�B)�$.B�s�"��F�sDc
�F�.�
a�4���
,X������B�a�#HG������֬��8�\��B��5�,.�f�T�*c��\4cB�$�Kӄ
F%	p�E(B�)@�� }���i0��8���$M�\v�6)����r��F8k|���![f�BF�HB�I%�%P��i�Y4���bIŋ	B1#��C$��"K���M6"��|��RT�`�e�IKYV��Ȑ��!���)��+�! �YA0SCH֬#�
a�1�"?!��|�H	 A%0�
�b,(oa
D ��֝1�3�
�![�[��k5�7��G4P��)���E��M�����gxw���$�!�E0��;�J�M����Jl2��]�ώ|ne�8�l��jH��p�t������_��ϷG��F�o4KqK��).,.fFN>��.+��~tL�d	��c��.�o�n�&٘jo���97��
�o8K�a�̳e��#O����u������oY~�9rfja��\�\4I)��\5
`F�j@�h�;v|�٤�0���j7Bia�c���o�J,XLb@�)$ޘE�>H|��So�����Ęo�}�{�,���ra���ɖXkaB��|Hq�k$`W&:�5z��D�$`K��90���F�_��5�5�o4��M}��k�@� ��X��6� �!BF\��w��̿g���(��+��3��5pM�Yt@�#�#Lk��k\<H���oF�
��l�p��;N<\Ѱ�D�/�\!��i�g�IqIp�a)\!�C|~�Ml&�����Ē$t�i���!��Ņ�|�.�m�ܻ�'����o$�M��a�|l`WN�e1ӳΎ�O�[8|���(�paB@�[x#����q]ÈA`���䵕�K�/��5��xW�i~�|�R�]��N&'M�B᠄�k)�W�2��j%�kZ�up�\��0����B
&.B�*ƒ�B���gi
R�@��a��L2�Ɍ��d���!�sr��L����8JK�I��4�B�1 �`=�͔��*"��i
Ɛ�
ā �9������_vw\���k�։~���e�9C�Y���λ�=ϝ�W��՜��ۻ��:v������ާj����}�n�;�1�pN���<�><W��]��B�%��	ą	t2D��H�0`C�IGaPąI$�1P2BPŃ��4A��L�L5���D�K���3a*F�i�)�k[e3I����u�!�4]g1��H4aK!�
Ҹ��יּ�Co���V5�3{w��ޜH����%1!L
��d0ԍ*���$+��$;�#!:�t�6a w��uw�Rh�B�͜�#u.l������&D8�5�I	��u� ��h�1!\�
c�)��sF�|ȟ��ݳC�<`C�.jo�f�t���d�����!HV_��l��Xo5�v�B���`�2B0!L#pָl�Is\�K�%�RYr\!IHR<_��,�tawXBb"D��u�X4�52���r^w�F4v\ѹsD����\V����)h%�sL,��>�^�����]�.��B��p��>]�E����{V�����:���J�>�Lĺ�3u�9���kZ!���d(!d���B\T�L	s	sdi@ 4��)�.�#��$��#
�4|�)���2(W.���B)�YL+�aŗ
�$�C�����.j��%��
ka.M�6�$* �E,�s5sZ[#��hF�5J�
��
��t1��H3N�sE�)��aM�<�L4B���o���h�ٚ�&�O��-�5�m���"@#Lѽ���}�7{�4�� G���(a
�2�#����C)���K�T���ސ�D�p����!�=	8�I��Ht_����s�e��#V\�.kr�w�w�o��CZ��5�Sl�ZY/�y�t���r��׿|�i��K��X�]��䂰7�uy߻2M��L�����Е���!q0"JB�S!L�(JAH1 ��HsF'H@#W	��c�lx%�[8�m%C�g��md@�a��S5	�J��+���%�ol��6$3[e7��op���9'���Ca�c�۳��e0���ަa�[40�k`B�i`P�ޙ����2���)�i
�>C��#D��_��u�!s���'vsF�sA.|����4������	�w��F!��h�#�S4Ja3l�2�/t_�nS���$c2�)��d%ŏn9щ.,Е�|�^ЗH]no�K�,,�IJt5IT��k	s��3Y.l#�Iu��Zִ �   l[%       �  �    8         7V���l�� �'Y�$�`ͻg	(���E���m� �D�U�����ڪ�+�h�m�l2p���ྴ�,;�ͥ�� pA��m�ɦ`si6m�   ݭ�ۀd	�.
yU�j�i&�����d5�       	    l*v�G�0�5��k��]��!�S[��k���  loRޥ�xp9�M��g�����4�r�\� 6�ܛ2�U[l�9��تշa"&�
��+VtW.��UUv���l��\�����UU:��r�>��]D��w��j������'�U��i�+�����ImHN�F��f����k�6���%��]����l�u�m�l "GN�$���l�2g� $[@$ �D�6� BF�`�H�H [G�ڻm�h�8m&���k1etf͚D�  ��`�cn��{7K�҈\�G�:��u�E�8Ʈ�m�!�J�Һ�3���Z��ԁ$��:uRs����8��nmp�l��T�clհK(��F7gI�]���@���T6ݛaت��ɘ��X�b3vЪ�   m��4Y;m� �m��Mzî����p   ���v06�iKB�0Һv���`    m�> m�  :D�A,�am$ �]T���vܲlݒr)[i����m:��-n��ma�m��5U��4��n��p ��"��I$���meP6��m����& ���� $��UR��U�@t��=�5W���� 6�m�FI����w�]6p]T��UP nv�`Ņ�j׎�5��p,z����,����<�z�q��s�Z��l ��K����$�m��P!+Vҭ�U\� [dHlY4��Ͷqo$�Ëք�$ ���&�V�$���ya&� m�[y�Mf�ָ���[\[�  մ K*Ym׮��Ȕ�F��I��ؑoY ��&e�4��E�zMj�ڪ�	v&H �����m���֋��fY��˂����ڮ��d�Gee��4@�E��ռ�Z���6����9�cc�l�e�޲[` .��17�>�$�md��M�#UU��UX'�U�����.�m [[dS�ulX�v� $�m�g^  ^[���������ٗ\��QÍ� 	 #m���ڬ��p���c�ѪvV��lu�BA��� 2 "t���f�t��'I l���	��f�m�d�tl�� m���V 8m� �[&j�I�l�&�i�lHl�^��2�Hs�� �5� m&��z�H8��z��� knؖumݱ�� �a�e�류UT�Q�j�Z�{d�#��pp��ߎ�mm�m 6��[@�Ih�e�Ku��o��F{aiIj�+=5lq�Q �I��R8����SV�Im$[M��wl��� �Sm�&��:.�/�m�$�I�m�h [A�ݤٶ��H��qR��CU.���L(�$/Msl�ĥ��UJ�P��@m��um�JqU�At�[D	� i�#�ka�q+WP'5S�sT��6��	A0\�a�6�<�P$  [@mM�` � ��-饽n���ڴ�i;:Dm��I�mj��cl<kՃ�C��9l�@-���`   9):櫽(   �I�Y�:@���N�J��v�m�mu)m I:BH!�	�9��p�ݻ�i`���g; ׶ �$[ym )@��6�l��`:��mm�e�%�څ�p��UJ���Cy:��t�MfZ�l�n �l�$m� ����p94��D�Gl8 �۶��j�`'e��+��[ p 6�j@m"�9B�6�5ti���V�UZ� Ih(���  I#6�n��{5m�U�U<��p�-�m����o9� �	�B����m���'�  	�*�  �*�� 6ٶ�6��/�ɵ.Y��6�|�Լ�.�Z �!.�8օ�ck�ۮ� ��F��vN	WP �t�-p 8ׯI��� 6ٶ����ր[u�w��  m�kpH$n�F�  H$ E�
ҖҼ�q�J�]VQ���Z�����v�媠r+F�YP8
��r��Hf]���j��`���K-l	nP�iP���v�6�涐  ����f�ql�mo]��V���5[�� S�r�]ui#�5�)V����`��IQJۍ�ٶӡÜr��m�P�͖��I�k��SNJá���*g�a���uʪ���(�,����]���Qd�j��jU��OX�Nܪ����;]U��ZBF۞�#�S�uOn�8�Ӡe���k���v44�u����JȦ�u�V�d�m�Z��j���an�Wl m�m�گ;7l���-eڀ�*	��m����J�$H$�n՛/��6�q��-��(BB@'@��d ��<��A�}����	YR��v���� D�L�i-��`�Č���  �Pn��Y� �7i6@$����A����jWT\��X�l�M p�$�+E��`����j�z��h��vE ���o   -� 8   ���  6�  ��i�ۦmyYA������۶���u�m�tC  ��� 86�d�m	� h9����   [@lG��׵&��k8���bAm��l�Ŵ���m}� ޛl���۶Ŵ�gB�z���v�i(>�i{�I��Ӊ �ִ����6�f��D�4�w� �m$�Z/m��t ��������P���    ��r��p�m"�hd'@��m� r@H6� ��a��/d7ǫ�� �����ڎpX���M���VQ��Д�
�9�<kԎl�t�N���J1�ؗ�k*�uO�uh���-�\�m��]   i3G[u���,0 �m�i�Ŵ�+UKi��@j�a�WQ 3�-�Vm[Y�t�m ���h��඀ݶ)͵�v�JP� v����i~��-� �"�%�� =�l���� [�Ͷ:
�l$Hm�N��
ڀ�[�R^��� H�m�I4�-���b��UUҭ�%Z�L��-UUUa��?*�}@�O(	oH -���-�\m��6��9jjm��k��l     %�t�-��[A )V�8U���g�j�� �m�n�Izݶ[	.(  �-�6�޲Zm���� -�K,��eVy�Z�ڪ��I]�:��6*��U���V� ��>���'�&�ک�@�VqU���-ں�Ci�����\���R��J�M�&��[Rg 5u��Z,�U=�������g n�KL [���pjV%��k�E�HB�]6�:�[@�  �A�n�3�f�� �m�f�8 d kd�mtT�$-�m8�jڶ�@[I���pX6�@5��Nj�$ آ��p�UKpl:*ېq�[��UڂE���l7-'X��.�:v� v��h;�7 ��dm�f�o\��m����KY�۬�$mY@ �Y-�I3t��s�@	Lt�],��Zm$��`�����,8p[E��mj�sL����-E)���nݳ�� �m�2xl�W(����.�\4��8���jt$��uT*��zNL �)�az��ڂ�.��A�
�p�*[,�TUU@KV�e�t�;~}�|��-UUT.� ��@�n��k� .Jւ��$�zl�/R��m,͚�:B�    l:H$ś]u�I�[@H n����m���6�HXf�� -�4R�mZ�$`	z�[m���Nu}R�ְ H\����H� :K��m�H� e�J巀<�lM�]6� ԁ]Tv2�ʰ
�UP�I�  .�&[`9 )g@�� $��ٲ��L��&�GIôV�V@e���ۚ[� �HJ H8[% 	e�u^��6�q$�	 Hm�m���Ám ^έh����텴 � �	6Z q\��2�V��UPQ���t� �k��I+����'�lm�	:E����\��1#m�-�@   E�u�  6� {I5� H�N[��M�`��6�l��B�m�	 -6 m"Z ��[I�,�ۃD�6��'H6�`m[@�`�l8ݻv�mm�"tɫL	$`�"�P�5�|��Am M+ �P��]5��l�&� -r�R�S����UY�3.7J�]UURC:�g	�Y*��6��f������Su� �N�    ����w{��T���*�\��T�*�_�0_�� ��b@  /�^ �����"m��JpP:�Q�@��P6�� ?pD
���튖� ���A�	���6��*`��9�h
'P|�8�"�D*�|� ����:
�C�h��a�E��� �� � � =O'�@��
!���Ex	�E:�W�]������NU��T��E�A�&�@Tx #�� P��b�AC'����؊i��	�D���>EC�A^�h@(��T�'�(�|�<@��h��W��0P)A<=�t9h��T�C
��>�$1<���UНQkp��D*O�> �A�'P"TC���px��4(���T���'H
|��) (�%E\�'�|�h��/�D6���W�ڢ]�:z�; �ESѠ�S[@SȎq���zP6�@� ~ :�(�� ?����J|5UУ�b E ��@Uڏ�!��N�:�I%����&�Ϫ����A�� A��[U����5U�lgs��$ul-��kҌ���$�XYs��뱷��h���P��%�eV��mu�"���M�u�5�N7�8Z-���*�n.�J�֫�Q2�[��m�(Mi6�n���y��P夭��S�����n]�v�sHR(�x��/Iۧ�t��nPɠ�L9[�z�y9^���/5l!'�	��c2�n7S�N`�8��X35�l���Ӊr ;=t�h�c^�����g��Np���)����H�����4s9�v7)���+��ɹ����*5;O��G�=��$�e��:�#�������d�`g@뚇�g���0ltL�O*dձ�7k�8-p�s��ogn3fP.!�ۉ[���4�1�s��m��fԹx�<�ɢ�Q��iZ��jܳa%��ێv�TA��>ґ, �4s� 1�m�	d�s�Ð;��A�m�e���Ý����v��g�gF�p=��j��G-�6����$ܥ�u9�� ���6ݩ 9N��@���l�W�vv�8˸�C-V5.�����Eyw^�X�&� �	
���sX�P��_��զ;J ճ@,ځe÷Z�.JCd�[�%����zZ�CFN;c���h��c�;W+���:��ݫ��n�k����˴g�6��C�;L�h��x�jc��fn���6l� /D�]�-ҧ!�����l�v ��5���=�M�n�#�Xr^�5�t�������K�<ؕv�tl�7�Б'1�n�Щz�&�9��uG%t���=��X�9��^`ݝ��>�l�\"�\l
QŲ����s
rᓞ�=����JnB/^fM�rɕ�n�F�#tT.����҃�i�0r���h�/-<�Yu�l�$���aE���.'t�쵒�]t����� %9���wF�u���� Z�J��S��PT�6[M���t��:N�}��~�ʩEH#O���<����N������y�^l�q�7t�x��ve
���5����H�����t��p�q* ��<�[�ۛ2�	����Kik�s�63��\�kg��"���DJk���]�8�$�Sg�7i�����Ud���9�� ��\�ٶq6�
��u(K0���`kËl��\�U>T����zA��66�v�0a]�����r�����хՙ0؍qF���$3.f{l�*�a3��v�C<���.�d2rv�(&^�7�����ذ��`b����\��d�g�!'M��ۺ�4��uȳܮs�I^������7^ŀwkU(���e�]Yv���$xd�`�b�7\� ��QQ�[B�O�6����n�� �r,�$x��'W�iҤ���ذ�"�>RG�vK��[�-�n0�ÆWY�c��	��'=s��t�L�BScv���=�)��+��ujݬuȰ�����n�� � ��c�w`�Wm[��|��>�}@����q �`b�	�� ��s�!�*tO�_�3���rN�;�'u�Xu�*��Ӷ6�$����u�Xy)��:��<�*Ʈڻ��1
��7^ŀn�� �I���BN�ye�v�v��"�>RG�vK���,��]4��`��b���R��S��%\0�T闋��6�#1gL:�cT��o�{׀vK���,uȰ�%�+T�cn��.�ذ�"�>RG�H� �<�iS��t�'f#�Y$�s޻�1"` ��$H$b��V( .�ITf�����`��5J]%W�c�V�`�E�|�� �u�X�B��&��2��V�`)#�;%� �{��X�ʪڞ^U��CH�zy��<���[�֜ٵ�tz����N�g�΄`���K�gS�-�����u�X�`)#�;�%B���Wt]�!]��ذ�"�>RG�vK���*i��Ym�_N��6<�$x{��UU�7�� �s� �֪Q�tղ�v�����p�7^ŒQ�I�Q�%U<PhX�-
�U��D��ܹ���^Bӥj�,m��7��n�� ��<��*WN��lT��ۨq�ZC$���&�g�ӹҞ�g�'�E��)� V��U��:T�� �{�6<�$~�+���_�/*<�/]%W�c�V�`Sc�>RG�oe� �{$��I�v�vZv�����p�7^ŀuM� ;�k�wm��I]�U[��`�y`Sc�>RG�n�*�]��.���u�X������^���� �Ur�������}<n�g�-�2hշS���n�:�j��6��c����W �;�<�3��U[j����cb"m\�b�,�6��TR�^J�CJiX�ؙ�	��j/^&5�M�<j�1���N��듈^ة��sn�.Y�v�K`�v89�N�����X���qp�T�:�N��>5�a@�3�O�!ݱ-��$��,�p����I��f��XٰlJ��fflYPbp$ ���hg�Se�vK����cG"+Z[��'k@�������p�7^ŀwkU(�:j�����N��<��H���H��6<�EEGP��Z��v��`�b�:�ǀ|�� � �5��|e�tӳ �{�6<�$x�\0QQ�.���իv����)#�7��n���$�ϯӟ%�5J-��K0�d�	��^Xu�,T[<h24�z�RW��K�5���e�o�:��<{.�ذ���Z�q�b�+��oe�(�_��'�Ď��������+����,��� �I�ĨR5vӰ�LB�0ױ`Sc�>RG�oe� �a���ۺ�4���lx�H��`�b�;���o5uwu|M'o �I��UM�x�	��:�ǀJץ)V���-oj��;:,akC�uӃ<.������PxմY�P)���V��N��|��o �ˆ��,�lx�H���\-S���N�u�Y��RF�O<����7��j���)t�_��[��uM� �I��U��W*���e��'\��$�.SM�
�We�o �I��u�XT����V��vݱĕ��7��n�� ��<u�=Ǽ����9�v��vb�{]��˨���sr��ͤ0�F�%#mC�V�ױ`Sc�>RG�oe� �a����v�v���窫�UI^��7�� �{z�I**^o5uwu|M'o �����`�b�:�ǀuV�UKIӵO�6��{��r�������=��I��}������R��HA�R"� � �@�5��|}�� � �5��>+N�$��7^ŀy{}���{� ���jaw]��i�qt)�r�u�%���ږ\��^p�#w�������K���tG'����^�<n�0ױ`A�&�̩�u�����w��;�;�>����'\��	�/ ;�k�wi��B�Xݸ`�b�	�/ �9#�lv��lB�0ױ`엀}��Jn�0�"��7�6'k 'd���Xݸ`���7N�?>����T��1Y�'�Ƴ;k	z���.D�f0�"�W�#pZ%sX�p���ٺT�	r򽵫�eR�r�uG�h!rv�u?��xCƙo;k�)#L3\�3�:2�],�\6�qn���z(;&�xk�Ղ���5Έ�f��,i�+n�#\��E����%��7Iu���:��mp�Oi9�'�Bf��6��1��6e�Kv�W�����?zwN�'I��ӿ'�30��e5ֱ#�ͱٶg��a��ƛ �c�r��w\�s�� �k��K�����	�p�7^ŀ�^�Z�Tu-'N�>X���Mۆ��, �����c�Ur�5 J#��|E�tӳ ޽� 'd�?r��.��� ��� �D�R�*�+Z�k 'd���Xݸ`�b�$�.SLwJ�N�ww�}� �r�&x�	��	�/ ���v�t���w|V�ш@��V�oWk�,5cXJ�HM��\\1�(W0���S������o�� 'd�s� �y�P���n��d��SrN�;�/� H
�H	"i�5����9�����n��lM卻������^�r,W*��)�p�7�b�;�*#x髫�������X��0ױ`�K�:�R��:v���ݬwn���K�_ {}��>�E�{��O����~-Xn����G�*k��Xca���-��� c]vA�nt��m��h縞)�g�H� N�x�ȗ+��V ��TU����U|V:�n� N�y���� ��� �{$�r�n�X��N����`v�k��r�))���(B1"J0��B��A�E*�"R�@����R 2y@Є���	B U xdc ��*B�!LP%	VA4�kZҤX��`1�"���� ���d�Ċ�bC+*,���q%t�b\�.ԸP�BhH�����ʱ"���(Ju�������k�L��]�Y޲�:G�����]�
� ��T��T!$"C�K	!+qh}��S%,�ҞS_.�_�V���)��ͮ�P�-��CJ ��:yX _ �D�'�!���?��T��W`)b��=�ذI/ ;�H�):wv��Wk ��u�X;%�o*��]�q`1*5�wm�]]�!]��س� ��� ���=�ܮJ�_�$������6Ӝ���4�6�z���Y����<h��M�J�˱vS\�-���}��|��Xf�=\��y` ��x髫���-����Y�#}/�#�X��������ӧ8>�Z�o멉{���W8��g� ��\����}���ʮR]����޺�N�[��r��E���$s�=Uʪ�H&�׀}��9U�_��& ��" 5U
�5
�X�Qx�]��������@[go���b�e��h�7�?;�N������{�_��A哿���rpDos���z��K��]MX�	 A_ԗkFm[A<�p��2����}�c�����q�W#I��5]���r�#|�~XܮW7�<|�ya�r�"o�x�	���wl���SO1}�%����JG2�$�[�/�IG%� ?�hK��QZ��J-���w�ĒK{%����r��Qܷ�$�7!��%�״��n7��3 {�_< :䷉$�܇�$��e,I%��Q����|� ��]�����x��l���}��\��P�� ���ԍل&�!V�ةX����푣SG\�s��mqu�D��/+�r�k0"$�.�
1���3�&zP.�Ir�cK6�Pe�62�g����Gku:�c��^�Y?��>Bh_	aA��a&qbX�iQYlV�ݣ�5���w:%���ā�lg�b��XX-������.�v�:���+�ٜWd$�ַ�n�i���N�I��~;~v`��l���DsisH�#[j��^��=g�I�|Z6��X��L������t ��s��$��e,I$��{\�Uw�/����� �[o���iBc7�>��~�}��X�I{���W*�֒^~��I}U�oޟz���'ư���tG0�߿I�ޞ��I%��[�*���^��|��+�޿} }�)��M�K[�p��m�����I/zg��I)�X��W+��6_�$�J݆�][���{�;|�������!� }�~|� ��]�����z�4�e��E��$&�R�]�l�g�on�7�=Y�l�h�\ˌQ��%#�KI-�/�IG%�I%�r_< ���Sjm�1�,0� {�{�s��""+��������m�ٞ>�$�s)g�������TT���j��?��|� �{� {�y��ߧ��M�����$�����H�Z�GOC)q���ĒRnC�JG2�$�Rl��I#��w ��i/zĚGiq���e,I$��|�J9-�I)7!��%��P�p1�SgM	�M�����g�����"�L��e6YM��NNq\x��� �޾x ww������< ��w�������ͶK[�p��$���$��r|�[2�$�Rl�� �ޔ+�4�v��]��������=��� ��P�<�Pv��:"fe߾�\�߳��n�o��i;��V�;R�|����C�����vK�&�� �3U��)���� N�x�ʥ��_�zK�vd����~�i�6>�`�W�g���/	OYl��h�$�A����厺C�N%,�]�_+���޼n�0�L� �����H#�cR���n�0�L� ���l��H�D�j��ۡ�f�I���^ M��	�p�$j��)t�_��-�`엀d�n�0+�UT���I�`h�W)������� &�xݸ`��X;%�V��S��E���N��ݜ'�6;R \�Z�͢.��Ҳa�nt�a�a���wN��l�դ�� ����+ 'd� �%�1*5�v��v؅v`��X;%��/ ����A�6�4�ҡ	�`엀d�n�0�L��Z�F�c.�J��l��n�� �$�����w�jA�0e.1[��7v�ve`��d� �+����TW*�m����vR��ESg���"n���
mu&�-���w���ԣNCVK$^]ʐ5��kv"{W6�@�3g�^���8ڸ�p�.-�K���Qm�`-͚ɝ0��|���a�v��Z�gu����~���sazۀ��4M�Y��T�t�,������*��^kOV�Xe���@u��u������)A�@���¦��֌�h��Dp���.�hӭK�M�6�96�8̼�	�.���=��6N4��L�Ġ7#c#�5����߾O ��\0l���������yS���ⶂ�wX�`�/ ����+ �Ur�n�[M+�0l��Mۆ�I��Nˆ��V�4�v��V���/I�0��e`��d�F%F�ݫ�];lB�0�L�v\0l��Mۆ�:��4�c2�
��#F�E�Q�lݝ��y�n�;swjѸok#;.�㱆�߮ˆ M��	�p�;	2��j���tkZ4��57$�ｭ�����SU L�@ЉE"U]4�� �z`�i!�JEt�_��&oz�ܓ����v\0��H#ecR���n�0�L�=\�UR^�_� ��� ��*���]U�CN���+ ٷ �%�{�➙� ���*b��U|V�Yn� ٷ��޿���� �$��?}=���-Fַk��X���K�!8��\Ͳe�ܛ��t��t��ʱ�&�N��	�^�na&V����@�ܦ�nݴ�.��͸g���=�o�� M����\n��.��!]�a&V��2�r�9\��K�7�p�>�4nU��N� �ˆ M��͸`��Xv�R������+iـd��na&V��V�R�K�Wn��q�8�dHw]Pv�t�a��o=A�V�Ǣ�M$�WNʱ��n� �ۆ�I��oe� &�xu�*�Բ��ۦ;��ve`v�d�uȰ	���]%W�m��	�p�	�^:�Xa&V�Ln�[Miݘ6K�'^ŀve`yUUY��> �C�N:���srN����Sl�n�twx�ذo�{��I~0l��w]!IE[���Һ�]��N:d��Dם�9��n���v��s�2������ۻ.��(���ve`v�d�uȰ��ەi;�B��&�� &�x�`��X�*#k���v`�/ �r,��+ ���֤����c���:�Xa&V7n6K�;��D�YWUm���;	2�s�����$��ߵ�'��z�IN����"F�w�7"FRX�D�!�!q���a20�hB��)�IŐ ł����A�~һ��>!HP�G���d�0&!�35nLHd)
@�ciQ6�l6��M�	q��.�ʅ�IA�	e�a��
:ְ���t|I���&��q��u�I����`'����륅B! 	����X�`¤T0j���K�!u��$X� v�@��!IS���X����'���(@#��"B$�FB1�y8Y��AW��! �)J¬*A$�"@hC�����#!#A��'�#!�w01X� �!"@��|ϰ��$��2'P���������� 	������Q�Q.!�T�0�Sg�\�8��5����q��s2� j-��z��]r����:�r�=^p$\���z�uJ��v��i f�s��z��nJ���#sӚ�m)��r����m�1e�������R�Q#R�����5��],�u,̛gNN�f�v� K�ˀ��]9�͹�J�����ؑ�B�%�%�U4]�6�Ȅ�΄U���仲����E۩�|�vѝ�^3��L�qs����h[���+s>;;u�j��݆q�u�9ł�6��ķ5���90,�5�V���e�ѓ����Q�-��1�l<� '
1L�J���qY����ϔ���O*��t@�ey�&���l)��:W9%� �quE--�2�qp�[:Y������X�o���EA��낥iGb�N�F/I;U`�d�Y�rN��rXՂ$�ʧd��uT	�ʹ���C^k�(���&#�����lnFI{:v2���2���.y�r7[�v`"��glx9T��;��CXM�Ĵ�q�on�q�؎v8G��u�YP皍Ŋ�q�f�x�{U���tU�L��;ydRB�N��U[=l6[���|N�M�{j�1�6�ˑ�� �%�t6��ASvX�ݺ9�(�K����0C���&]�s=�<�0��6���e����V���w�	���fL���N�w;��`\���n0Z��X����R�p�u��l�=:Bއ��w:�\��\­��D�B<�j-�S���Q&�D�vյv�ĳB5��J̓8�64,�gQ�-��v)��ܻ�热�@5����:�����μ1��&��!�6�Ȭ�pqe
�[����nn�o��O(T�)nqX�͛fey�<�5K�C�
��-��;om�m�"�)Y�!pgC=�@knl�����ۂ;i3�T3��t�g-���e)�!�Qu���[.Q��4�n��f���t�Y��I�I~w�Ё�~@~U�� �� ��pP�� ��o�Z̶d�^�J���<���蕗3��i+���`K��^jF�X�[ve��|����6�Y�h�����M4Mt�K�cH���oo6������;7l����݋���٭�EUukH B�	wJhڶ�8�q�)8��v��sO.oiG�0t�m��Аniw��ba���#H��^y&7.��]u�ę���� BڷZ�X�,KC4��t�#Y��V��3�U�(�q�e�� ��k� ���8b	r~�0�Y���]単�]%W�m��޿� M��	�"�r�A�=����^���i�� &�y�\�+�*��?ߖ?�e`�r���/�����C`\��������� �$������_� ?{���:���\wv�˫������=� �_� �%�G"�>��Ccmʴ�ҡ	�`�p�	�^�r,��+ �l(�`�ԋ�+�bL��,2����1հ�e��HwNn���r���b��8���z{׀}� �$��\����I/�݂���YNʱ��n� �9eWr����T8���o��s�7$��צ M��ܪ�8���B�'^���[�Wk ��V��5"K��}� ������U�ۥV[��7�p�>Sc�>�b��+���O}Xg�*�	�e6�.ӻ0����ذ�ٕ�ov��o����8~��r�f�w<���2��0��t�b�m���z�ï�4�.(��%v��ذ�ٕ�ov�ꪮW%s��^�<)IQ�ݻ�춀���}�̬{��6<��,�9Uďy�P������T!;�l��lxm.W(ʪ���w�~��7I�H*#xں���+��*���X|���2�>��L�`w`��6VS��|����>ץ���UJ4��|�_���{|��|��o"�u�`��
<�Wk���Z�Kr���C���35pm��%���W�[�Wk�;	�{���/W>A�9�H�EL^�*�e�ue��wn�$w�y`�����2�ܮU$vxB�`���Wiݘ|��r,>��z��ۄ�V$�{���r��wt�:B�X�R��Xa=��n��rm@E�D?�h���?w����~��l=��\������̬ܪ�I�>�s� �r,�����ͬ��:;+6�]�v����v�Ɓ3�#�~�%�Xlm�F��'u���`G�`G"�*���WX(Oe`��G�X5uwu|Vӳ �M�?s�����l����o�~��7vឮq#�Ey����c����?y`i�+UU%$�W���tP��FU������r�v�V$��lx���|���o{��j|����F������9S�U������c������ٕ�w��EW(ℶ�lj�0Nͤ�h:՞�ɽu �nn�E)�&s[�l�My-z�J�4ƶk���y1��S�����k3qj��m�IÊ�D��[��d��ѡJ=���GD�y(4G/&mm;2�\����S$����0�,i4����I����U�|�}�}�F�\]�$jL\9uǧ�VK��Um�8Լ�:6^
�晣
�iT��:wI<�ݧ���[n��Ike*Ux;	�[D���m�v��M�
�n�.���ww�)c�M��Mmݐ/�<��X�l����Ӥ�������~�����镙s5���r,��$v�X��`)���RF�	��ۻ.�h�Xa=��n��W'+��������#5P�ۖZN�P��<��� ����>�E�}�̬H*#k���v`)���]����;	�wn��P^.���6���X�p���-��ruʯNx���L�Y4����,#��&�\��>�E�}�̬wn�Xj���/	יW�[�Wk �M�X��G��<����0^�x�ȳ�*��"F�*b��U�-ӫ-�`K�|�Ǉ���,����>�!U�CvR����6<��X�l���\�g�d@WLeuQ�3�m�9m�O����|��`)����<�Uv�1����Ny�1!66����l���a�펮%iy��~��Hǎ���v[@]���{+ �ۆ���A�?y`�"���^�I�*�����)#��� ��ٕ��${�o5uwu|Vӳ ��{�ܓ��z�iDtP���S���6K�}�t̫��|�����R�����{+ �ۆ�W+�q����O:(_���*��|��>�fV�UI3��w�y`)#�&��T�J��4Ƈ��s�:��v.�\����dY;]4r����M���R���h�3��}���G�`)#�UW�;	���_���V[�����,�9�$u{�xa=��n��?~�USd��H��P��eںi;x�߿<�6ea�UUU%$�W��ՠ��;�wWv]��v�?r�������7$�����䜾�rq1��࿑T�o��f�~���332z�'t�BwX��0������i�+ ��k�&�pT];M]v�v��(���tf�d�2U�%i�V=ql����I#e���WNm�:�������i�+�ʪ����`ڊ��OvU��ӻx�H��\�q#����$�� �M�=\��H�R��:^E_o��xa=��n���\���U�oW�~x�߿<u��LRЪ��t���=UJI�0�O<�$x�l��>�!U�bv��av�ـ|�ǀ{�����{+w�צ� &�E

R2C�wN�}�vh$�[]Kn�\�'���uݎ��e��1�h������;[Q��Bպ����6<�4O>�H9�#���\�,ܢ�e�f�A���bu��b��f�ml#���u�s����uY��N�rX�^��l���Z$$0rj�'��73���_,t��0덧v.7M=�ׁ7N:Lv�%�M١;=q�6�#u��gR��e>�t�'O~�$�x|����%U6܍.��]�@È3(,6j[�]ڗA���m����W������.����j����ٕ�n������,T����컲����}�̬�$�� ���>RG�H�*M��*�wJ�'u�n�� �=�%��y���V�%Do5t���۳ܥ�\��:��<�6e`W)I3�ݨ*<��j�X�m���|�� �]����K�}ŀ~��z���J��_-���.m�=��R�:�E�4�#�����!	�M�Uj�
�tZ*��|���{+ �ۆ�{ꯐu{�x�TT��B��k534nI��^��N+{)!����Ͽ��?y�i�+=\H���W�bv��av�ـw�y`)#��+�7�=�+ ������$[R���.����E$x�l��$�+���y`Z	~m&��v�B�x�I��z�����|��,)#�>֍�V�St�e�۳taWDh0���\V�F��lTL;��7�7n��C�$y� �m�"��3<����rr��{����]a�=�+ ���Q��lV��������{��i&V$�Y��$n�y��ժ���wk ����nI��{f�D6� � Č#�"�����B@!�!���F��aHD��aYYKH��h�Z�HL%�C
a�|:Xj�@�@�# �H�S&*<�1���A1��`I(:@ڐ$ f�]�P��V�"D$ц��t80#2�]�)�f�Dv2ʺ�Bh�X�'5J��"�c��"@�P��X@�lq�(�Ӡ��"M��J�""Em4��4��	CJ�hD�5�N�'Ƞ�P��tb�P<|b� =A:���U\�r�����X��,�]�]'J"����]�W9�.����{���:�ǀE$x�Th�-$];N�X��$�X���s_���{��X�I��N��?�7Eg���m֖��͹�$B�����܅4Z��6d��|<,��W8흤�w_��� �Ȱ��+�+�W9\�߿~��7�I"��C����t�v�	� �I2�	$��:�Ǟ�r��:�<�ؙv˵i
�`����I&V�\�W�W9M��ߞ����`:ԓm�R�'t�CwX�r���}X�O<G"����>UVW+�����}"TF�Z.���wwXT��r�޿y|a=��o{��r���Ĭ#mb��f��J�8�E��Sb��ɕ���<j�X��߾�!�ibj�X�m;�������e`I����O<����:^E_o�]��$��$�+ �#�`�Q��J���N�N� �L��lx�b�>�fV%AU�Nݣ��I6�?W*�u�y��X�l��$ٕ�wu$�jP���]4��G�`i�f��}�rN_wٹ% 0�E�w��}�۶�˱�Mi �k���:)�v��`٣��ۧ����N�Fiq�.mU=��8vA��l�u��%�\=�8Kѵ$�t��M�81�[;W;�iK�.�c��V�`l=a���;ypiʼ��<F��V'�������>-Iv�(��89\F5��uj-vkF�x�U^�Ri�v�vE����-���A�Kv�v�ݫk,�fȺ�{#�I'��y)����F��Պdɥ��릸��$�\[:��se1տ1�|��u:�0��O���I�+ �M� ��X�D&�N�X�ӡ	�`l��>Sc�${��eg�'�Ty�lV���[�wX�O<G�`i&V&̬��GKV���iݼG�`i�+ �fV���EN�E]Yc�N���2�{��W�uzy�M� �vvuɅ�F�
2�n�ջiN�����KaK��=:��)�y�y��Sԭ�1V[[�#w_�Oe`)��M� �M�X{N7n�2��M���6<��W�}UQ���tF����C9?__^<o��	$��;��E�)ݶ��t�v��� �M�X�e`)��]�q12�j�I����	�`n�� 7��?���<-��t�V'tИ�����6<�$x������lN�`6.u6g]�6Ֆ'�P�sl%�y9ˤ;�7�ɳ �������\lV���]���Ry�)#�>�ٕ�s�K�o=�h���-�v����V���7v�|�c�W)")B�*t�����Ɲ��'��ݸa���"�Q�T ��H0�J(*� 1H$D�;�s�J�]�?W�{ߞ����1K���Zl*ۺ�7v�|�c�>RG��r�jO}X�E9O����m1]��v<��:��?��I�{�Wn����Ǝ
�cEI��xM����u;b�m��6못�H�33ڛ�;x�lxջ2�ݸ~���:�W���^����˶]�I'o ��fVz���6_��O<�6< ފ�ciʱ;��M;�wn�v<=ʮ%��y��=��lԨ��b�]���fI�V����ܓ��߳rN�nDF�	"�H���r�7�'�PA)��c�����Us��=�|�~0��x��:i�]�t�땻����ۄe(��#&�ڂa��:�7 ܎�o�Ӥ<б�M�#7k����X�n�v<�6<u�4b���&�Gfx�ߏ���$��;���}�� ��ߞ�n̬�9\�$OS����:B��һ0�<�����ve`ݸ`����;v�wM'o�\�qu�y��=��ov�ꪪ�.�<�P��12�j�I��>�ٕ�~���<|T�x�lx*�t&:�J=�qr�L�ѻ���̩uhmK�=n:�ہ�d^jkI<v,R��&Va�j�We�-��b^5�WE2���=���ȑ���Z�[B� 8t�?'0��n�ã���洧ahM����;Cn��N���.
��y���S���؏W-�Hð(�]�J۝g)u�k�X	6��:6-B�A��5�Qz.�`���9$�I��$�ȾPP�=E[��G���h8K���n���I��JY�����F_󤓻����6�ȗ3R�s<�K�|�c�>Sc�>�ٕ�lԡ����1�x������$�'�����5~��m{߲���3��UW;�)��T;,|����:�<��ve`ݸ`-����TT�TYc�N���U\]�=�`e��>[��~���Wwv��}�������̶1�P�����0�v<�6<��̬�V����`�u���ԕn^i�N�tr�Ł=���'s�y��K�J�O�I��o2�*��vh{���>Sc�>�ٕ����s��O_� �����[C�n��t�v����A��?/9����ٹ'��x�>[����$�Oɉ�l�V�N�ړ�X�n�v<�6<�T�NU��4*i�`z��Sfx�:���>Sc��r�v��ՀOD���m���]���>[��)��V���>~�}<�[m��T��`���w%:)�DZ�F貉���4���adҭ����<�<���c����u{�xջ2�ݸ`-����Q�Z���xջ2�ԑ$�T�x�H��H��#T�hUue�*ۺ�$�� �nǃ�(*���H��*B)ʢ�ݪ�)c^�<jo��	8S��ڱRݶ�ف��e�,����>�ٕ�����g�}[�n�n���)���]�=�|�~0��x��{w�C\���-����p�f��,�M���'�N��=]�u�d.0CN�N��n̬{���{��*Q��*��4���3�$uI�w�y`V���6jTG���uue���>[��G�`V���7�p�>�)��P���wo��ya'ǽ�f����ܐS�P
�P��8P4"�Z޽��r�JOF�Z����ݬ�ݙX�W96g���� �=� �[i"6����N��.f�P��`�[@��ȰL�v��6�UQ�|��WhUue�*ۺ�7�p�>[��G�`V���6S�r�X�
��J��>[�����,�'����3�9��q#}[����Ɠ��w�y`V����Se��:�����⦙m�j��������'��l��v<˾��uD*^ci��N�SN� ��� �nǀ}ŀ}[�+ �p�B1 ċ0��H1$��1�E���I�Fy�(�zI��$#$`N��;�HW����BT(��_�Ӏq��|�t�!��y3I��*`�D��H2!WO
#�y���!!�k0G�T�Hm];XO��OedBЕG >l	�ך�`@��bFH0<|@������p,��R1 �_2)������lN��3ba�-�B$g�0�	� o�`C��ͦ$! �P����G��~��m�ޠ
��� ��pY��7���dH�����"I-��r�� U*���V�ӣ\ݰ+��}��ړ���]�j�T��XPy��iR�c��`�k��E��k'�d�@�[]�՘�mP�V�5vv�Qh���PV�[ګ����j�,� V� �+Wu��anՌ�C.�{J�����E1j`O#��E`K��[ܡ9���
��3�d�E��"a6,�s�n3���sC�<<��&��+4ݡ�A"����e;�
�.�۸��$�]�ԎP��r�	ך;M����ҖRyv�1�t��=]'=�u�;'i#��&�6�*�dv���nx��c�VE��z"c��1y�,F	���q����(�:J�nݱdÄ1bb�em�5�Qc� �͈`���!jƶ�-S�ۦZ�a1Y���vG5�lP��钻%uu��Y]�[[] s�@�a���GV�ۀx��9�=��4�6zOg
qs�K����V����)���cCa��l�-7j�JA�7;Q���.6��[&·S��ۍ�*6�)8�gk��Y糂�UU��]���K�v7i�,ζ��; $�Ԫ�Z�t砖θ{N�[$� *m-A�c����U�/b8�7Pv�vH=(��S؋(��sO�{:��h.l�@�3Qu�וI5����xBިWd����Wu�Ɍ �X���N&�n�N1rP�[;[3�Il�f��A�S���A.[P����wj�*��vے��c���v^K��!�m��d	u��7bz�� pf��9Vy���twj���L88�;n���!�rPvB��h6bkH�,�҇�:}�NL����7QY푹L�x��om����s�\���(e0��-M�@`l��;�d5PЭ5�4a�a��1�l��A����ӲM#uX�uE�'1AՋf�e͠6�D��q��M�u�t�����N����"�~X
�
��S�_ �DD����hD�~����</�l#ם������-7"��&5U�uA�b��Y���e�Z5�u� s0Lᰖ�r��F/N;�awJ���a�هf�#-��0q۞g���]{�� ;�n%T`��0��GiCw�n8a;Oc4"Wl&C��n��f���g� ���u]E[K@�m��bE�q��m�An��ku�)���wrxK�[3Y7R4�Zus�[��6[ �`� 亗8a�-d���������v�*�5�7�o�߾���,�ݙ^��9_ �/���J�RxP���wo �=� ��fV�ۆ�ݏ?r�W+���T~+��U�|��m{߲���0��x��X�TkT��U��h*ۺ��9ʪSfx�:���>�b��W*��R{��=��?]��@������n̬{���*��E�ݦ�㪻�v�Xy6����(:��i^�"��u��ޓ�_-c�4��wcI���O<�ݙX�n�v< �-N&7Wl�V���ܓ�{��N�� ~؊(����S���/� ����>Sc�>Z�J8���J�4���0��Xz�UIu{�xjOe`"TG��e��]Ym�0��X�H��ve`{�RL�wy�KԞ]Տ�ӻx�H�s���W�I/��ݏ �פT��WWbY�m�]��8�uD��L�V���mi�gpv�J�E���]�Ʈ�����7v�|�c�ʮUW�u��߿</Q�~�*�Wn�[wX��0��x�H��fV{���p�X��U�wm�v`^��ܓ���n<Xa�
	�D�
6"pX�P���w���`wn��q+�����v�=U��{�~x�߲�ݸ`-�����8��]��ZI]��ٕ�zI�>�O<�$x�ѵ*ժn�;V�n���WBh1V��I�N:Y���W
Fݘ��
�\4�H9�����}{ym���V�?|��{+ ��Ty��]�WV6ݘ��,�$x۳+ �ۆ~�$wy�KԞ]Տ�ۻXW��}�2��r��7�z�����:��D8��>5v��fV���{�8�^֣W� ��J���t��߽�ܓ��{)}�)��ݠ��ݸ`kذ���n̞���'߁�y�필kYB(A��+/d�b��f�8��YSa9��!�琙7��V��i+��o��,�$x۳+ �ۆ7D+%�һ�-��'k �I~�9\�;'��	%��>ױ`u	�cuv˵i%v��fV��?%����y��
�r�]�j��u�n�� �^ŀ|��˲{��'��x��WWuue���>ױ`)=��s����;���rJ���P�(H wHӧ���o��C3K��Fa7Z��9���Yz�rZ4��(�+	��oWE�C�'���}49�y���%�n1lm8
�� {Z��
�"#[���mz�sQ;f���D4�m�P�;u� �S�y:ֳًW&�es���9+6.y����r-�ؐՅW"�f�
�N�A�\5
j�V�h2�lN(�H�؍�kn(L�nA^����h���$�'��?�G���L�k���ss��F.uzA�v�U�[J�˞to���j7���xX����@��{���fV�ۇ��]a�~���B����Ԫ�>��>ݙY��U\H�/��'��{{��W�USd^��#��Uһv�ۺ�==��s�E�Xn̬k�Z5MpM$��r���<�����'v�M�
�i4��n����b�=U�r�'������|�c�;���%�t�%j�)� �%�-��IEk�Lm���Nt�ۈzWF2���wc��}�2���0�����S�t�߸>o����aa����ҩ�`ݸgܲ���W.Ʒc�>�b�?>|������Ӧ�����y]�b�#�L|��`G�`n̬{���*R�_����wk�\�s����vOe`ݸ`kذ��Q�N*�O�v��fV��9U6g���s� �=��o���x�]�3�(�n�	��� �і�D�[���hm��N��@��P�q�v�ۺ�	��`kذ�ؿW9Uʯ�vOe`�-�7n���i+� �^ŀ}ŀ}�2���3������r��ǿ�m*6�U��1s|����|�w�74t?��Q�B��h4@��o7�k�ܓ�����O�D�q���eڴ��`~�W+�]�� �/��^Ł��]��, �Q��eݖ��!ZwX�n�s�\�˞_�>�r������'��;0�l[�1Nmpcjڲ��jT�	fW��ӫ9ݸd:���[n�����mـ}�b�>�b�>�̯r�ʪ��~0�yR�,�uc����{~�Ur�;'��	��`kؼ�'w��;�=�aa�lc��[�پ�����ov�}�b�>�b�:��1JE�v텷u��W+�Sfx�;����w�rE?�M'@h x:����V���[Q�uwĝ���0��X�Us��y|d�V�ۆ*5����#ͷ/Jr��g��%�v�T`(�m���s6�&�Z���������+ ���ܮr�� ����.�v�	;�����7���rN}��ܒs�����/���w���uweۺ�wX���}ױ`�e�wfV��IJ�m�Wuue����9\�������z���+�r�����vsʗ�e�-�v���s���~�UW*�{�k�zz��{������F�*A����5�P�z�吗�g�v�\\*i�ˣ���%���N��^�T�*]s�ݫjy�^��c����{4n.��x�u�5�gS�T�v{E�I���s����v,�kIZ��.{#y��!ڢd�9]u�!zz�m��T�õ�iG�2��n���Pͯ�IF1�P�H��8܁�Q�!�%��=���Qd��[�zҭB^G��;�I߽Ӥ���M`�e-�%3��jl��7!��f�Z�ZY�7F6��֨T1�����:bwx�L�{��UUr��}=x�Q�C^�]'n�+wX�n��\���X}/�[|�������~��θ�gE�0
`�<���0��+ ��� ٩
�i4��+n���>�p�>�̬{�UW+���<�b#�be�.դ7f�ve`ݸ`u�X�n�>O��k�lZ�PL������z�ڰ�C��3�'&S�ʙ�"�M/ޓ����Xy�U�����[��	��`u�X�n�Aݞ��'��/S��uwWV[n����@�H�"�� ��s�T�'?o_�����7$��צ��wI-=������X���� �����>�̬?s��Se��;�y`[B���Uv���>�̬{�	�(!�������'��~�f_�虬�A[��7�p�?r�]۞_�K�}ݙ<�O���}�n��QjWm.s���L��F����\�͍�N7n��`�g�;���̟,���٠O?�� �m� ��2��A6_�ނ���Nt��`M�g���r��g�e`����^ŀj�
���N�j�� ��2���0��]��"����
*@��`	��$@��cM����F�|�H��B�P����@�� �ڰ
�4���1 ā!�4.<��[�����d�LS�$�$�#Ib��}���$B �@�τ�:	a� �����)��!��O�SU�����4H!AH�$	
�(�����!!��y8)�q6�@>pE:���'Pt
?��Dz��+����Xݸ`�B�9wwi[wI�u���U\���?O}��6?~X�n�ٕ�l5RR�6����]���>�ذ�ʪ�����ߎ��߲���0���M7�PC"f+2�%X5��j1].x��RZ�=qm3��[(un:5[��>��X�n�ٕ�ov��W�;�y`�
��^�-�'f�ve`ݸ`u�X�n�q#T�4���tZhwX�~0��,�����$��ڍ۫�	�i+�ܪ]۞X}5�nIϻ훓�� #A���A�3��wsrO߽,��ճ.k)[�����,����7�pگ�U�bX�wY�Sq,K�� �=����5��*;B-�4����j�+S�c�q�vZ���\f디��]�W����q�����ؖ%�bz~�ى��%�bw���iȖ%�b}�g�Mı,K���Ο�Jt�Jt��!a�U[]�l�Y�q,K���ߦӐ����,N�Y���Kı>��~�ND�,K��l��O� 2�D�?~=K�j1cˮO:~)ҝ)���oO�,K��}v��c�,2&D��혛�bX�'����ND�,K��Y�<RU���-�<:S�?���!&������r%�bX����q,K���ߦӑ,K�I�;���Sq,K��x���f_���73WiȖ%�b};혛�bX��w��6�D�,K��~�7ı,N{]��r%�bX��^��ȃ $0{��Eƺ̹�&�\�^v4��	�]Cn�� ��g��v�Թ*�c0��X��.g�Ɏ#�J#l\�X������6�%�Fz�Q	�uq�:�u/��r��KY/*�:{[\.��M��vD+4�^[��a�V��X�x],���:���덲-[��`6��qr]�g6��Ir��d�u� U�Ǎ/N�s�I1�,P�3�;��N��o�l�]C*:����g0v-u���̽�nh8�]R�3N9����u��v`�Cl��ӥ:S�:w���6��bX�'��z��Kı9�w�iȖ%�b}��7ı,O}�����\�mSΟ�Jt�Jt��֦�X�%��k��ND�,K��l���%�bw���iȟ����e:JT�m5Ε�b�ޞ)҉bw�_��ӑ,K����*n%��C"dOw��6��bX�'}��jn%�)ҝ/ϖ�|��Y�Uͥ����ĳ���;���Mı,K���M�"X�%��u��7ı,N{]��rt�Jt�K���U�ٖ�����,K���ߦӑ,K��﷟�ND�,K�����Kı>�����ҝ)ҝ??O|.��[.p�*1�N�tr�nҎ�X��h��܆+8�p�ٷ2rKY��ŏ.�<��t�Jt�Oߎ���Kı9�w�iȖ%�b};��3�2%�b{����Kİ~K>��%X�����å:S�:~{���9�v 0W�Eh �&��Ȗ'�?l��Kı?{��M�"X�%��u��7ı,O���z�e�55����r%�bX�N�f&�X�%�߻�M�"X� a�2'}��jn%�bX�~׿]�"X�%�zN��˥i�M�>V�r���g*l��iȖ%�bw��֦�X�%��w~�ND�,�P��߸bn%�bS�߰��ﺺ/;[T��ҝ)҉�u��7ı,?�H����6�D�,K�߶bn%�bX�����r%��Jt���>��)���{H�cC$��7�Ԩ���֋����Z�#=u���sV��X�%��w~�ND�,K��l��Kı;�w��T	�L�bX�������%�b_z�Og�2ʹ��<��t�Jt�O��M�Ȗ%�bw���iȖ%�b}�g�Mı,K���6�����,K�aa�*��̴���xt�Jt�O{���ND�,K��=jn%��b@i������M�"X�%���l��Kı=㴷�s2�ѧZ˚�ND�,�"���o?Z��bX�'ߵ��iȖ%�b};혛�bXȋ2'��~�ND�,K����7�B�F�:��j��Kı9�w�iȖ%�b};혛�bX�'~��6��bX�'��z��Kı<g{}0�M7a��ͻ%��2�}ay^mi�+����Ʋ[�+
i�$�'�BY��_X��:~ı,K�߶bn%�bX�����r%�bX�wY�Sq,K���]���N��~C�oqZJ�B����,K���ߦӐ��r&D�;�g�Sq,K������9ı,O�}�q?�ʙ����7p�����浖�jm9ı,N�Y���Kı9�w�iȖ?� �"dN���Sq,K��}��iȖ%�bzvYOm��:U��ͽ<:S�:S���o�9ı,O�}�q,K���ߦӑ,K�ڋ�ީ �
��G�G����~�7ı,K��e�7݋2˜�\�:~)ҝ)����bX�� G��?M��,K�ﵟ�Mı,K��}v��bX���;�Q�c[6��� �e��m��x�Z��N�0rWTu؏l��!Kf`\��̴��X��bX�'����ND�,K��=jn%�bX��w��"���^��K�����Mı,K���K��j1cˮO:~)ҝ)��㽷��Kı9���iȖ%�b};��n%�bX�����r$�$���S��d�2e��5�O�{_�ĐI����D��w~�ND�,K��=jn%�bX�gHS�3=�)��m�M�"X�%��﷉��%�bw���iȖ%�b}�g�Mı,�ȟ~���W�)�r��R�ҧ�+B,hz��Kı;�w��Kı>�֦�X�%��k��ND�,K��ot��N��N��������v�`&�+]��� 6�Pt5͆�gs���[�l�Ժ�ojN �s��`���{Kh�����r���������;��3L�
U�i]��\\��;���xـ����8�\�mձۛ���Y�7d��Mٻr䅈Ƕ@�����^��"�3Ta���r�g��y��gY�W�sV���5���t��g�x[�pm�-Wh'B�um��0�흘$ų��0�g�p2��a�t�Y�����5����XIsZ�n�8��bX�'���jn%�bX�����Kı>���Mı,K�w~�ND�,KӲ�{z̙sX]]jd�թ��%�bs��ӑ,K��w�17ı,N���m9ı,O�������2�D�/�l���b�f�u.o�?��N�����q,K���ߦӑ,�"w=����X�%���{��r%�bY��������ve���å:S��%D���M�"X�%�����Sq,K���]�"X�%���c<:S�:S��ϖ[�ߛ:Տ.�<�Ȗ%�b}��eMı,K��}v��bX�'Ӿى��%�bw���i�t�Jt�O����
���&"N-��T�]��7+�k�u��]���t��,�1*���^��Jt�Jt�����9ı,O�}���X�%�߻�M�"X�%���{*n%�bX�gHY=��SSX��]�"X�%����T�>�/�?	��9�����m9ı,N��T�Kı9�w�iȖ%�b^��i��u%��d�4T�Kı;�w��Kı;��eMı,K��}v��bX�'޾�zxt�Jt�O}�,��L��Rڧ�Ȗ%��P�O����Sq,K����]�"X�%����T�Kı;�w��Kı=�YOoY�.k��L���7ı,N{]��r%�bX""W�����,K������ND�,K��z��Kı>�=�Z:Ye*�0e��T���+ȱ+�z*����Nt�^���ïH�p�̰a����Kı>��ʛ�bX�'~��6��bX�'{�����%�bs��ӓ�:S�:_ߐ��5r�̴���<�bX�'~��6���X�L�b{��֦�X�%���{��r%�bX�z�eMı,K�;K|g35��F�Mff�ӑ,K��u��7ı,N{]��r%��P��Ah�]�EH�x� 	���"v'��T�Kı?~���ӑ,K��vx��1*���ޞ)ҝ)����iȖ%�b}��7ı,N���m9ı,N�Y�Sq,K��:G�d����73WiȖ%�b}��7ı,?�?���~��m;ı,Oߵ�֦�X�%��k��ND�,K?O���nY_ɜm��[."]�����3n�+X�����mW��q�	�9��5�:\�Sq,K���ߦӑ,K��u��7ı,N{]��~}"X�'_�*n%�bX�?OSw?L��L̚�Z�ND�,K���T�?�9"X�~׿]�"X�%����ʛ�bX�'~��6���DL��,O���O���ҵLl��å:S�:~�}�v��bX�'޾�Sq,�dL����ӑ,K�����Mı,K��m�����fvm.o�?��N�����T�Kı;�w��Kı;�g�Mı,���IR� ����_D�����9ı,K�İ���GfZ[V^�)ҝ)����=�ND�,K��z��Kı9�w�iȖ%�b}��7ı,N=ðс�KsX�����A������^�Nr��՜�ƣ��y�B��#m�"X�%���=jn%�bX�����Kı>����șı=�y���ҝ)ҝ>��~ĭb=�έMı,K��}v��bX�'޾�Sq,K���ߦӑ,K��u��7�9S"X����~�R����j�9ı,N���T�Kı;�w��Kı;�g�Mı,K��}v��bX�%�;���5�rjaIsEMı,�T��=�s��r%�bX�������%�bs��ӑ,K��;���Sq,K���z���sXk	32j�jm9ı,N�Y�Sq,K���]�"X�%����T�Kı;�w��Kı 7*D,F�3�x�X�$dIHE�B�	c$\Ga��4FD����#�l
��	F2SZ��V+\TX�֌��4���JA)���=C������N� �0�L�.B��HU�;��0�n�IB 4#	��]؛D�XRT�.={�����oA�YAƘ@p�e�L��������!'�G�h��e	��|� H�@Tڃ�U�hMa���TG)�u���$����c)�F�Y���ROq��΀�u�B��%����j )��2�Yf.U�HS`)5弭�X�t��f�3nx�"7Zp8��L�d �5��`��Nҵ��WV�E��l��V.�UE Ue��m02�g�6t���.���M��
L��`�����e�.��Y&�j06rl���5C�6� ^���D�0�n�J�۬��+2��8��+�	u��ے'l`�ƬC�H3���sUM�&8TW�2n�����v��D�T4�m+m�����N����!4�J�c��.�u�b�3��0���$�h�Mh���5eH&/#^��V��[v{q��u>]����'��$��{,2�GR����>��/��A�u��6�Rj��d�K*��)\�n�z�@ud�^���P���m�2<Х�mtO'�4]�'dH�Z�b,�\jwkr��n�<��r`��,�!�c�p���;M�:v�m���[�]]t������Z���!nfٷi���`m��NRnmׅGv�a�V�=l�=`�{
�uP� �O �T�U�U�g�K��li����T���.��	9��F�c�!�R����Ռ��z���A$%R޺�R	qH�/;S"S��������	q
�	�6�$-�6"����]��rY ��b3�B�*�UH� Y�x��8��$�t��5 5�E��8���<N(�%UӌJ���,��y��7F^G�h�����!�g7Q��NP�m�}A$��	�B�FO-�q�{6�ݵ
��v�a�bbX�W�4�K`�;2���*��[����;)�+]S�7g&-k$:���K��ve�f��i��D�.�;mȮӱu�xnT���#�;���:���M�sZ6�!sy㝓�ճ�5ק��"`�f�VڦOA�&��q�VL�f[�ֵ��>U�Dz����G����Dpl�`� ?�����r�Z��H��upV�v������z�X���/��釴	��cP��p(p���Ֆ�Q�m��[l�[�i!�;.�d#������m;�7e����8ը��X���K�@WW6�:�|�Ũ9��F��,�G�:ފ�U�`�K<���W1�tvR@����^�gf֎�t�6��X:h~����i��,Yu7��qD�o	�4af�f�Vq�n^��Nh.��N�낌���:����%*-��Үn6m��t�Jt�O�뾻ND�,K�_l���%�bw���a�^��K���Y�jn%�)ҝ/߶�}��5�ٴ��t�:X�%����T�Kı;�w��Kı;�g�Mı,K��}v���Nצ:S���,>�Qٖ�՗��X�%����ӑ,K��u��7ı,N{]��r%�bX�z�eMı,K�;K}��5��F�k.jm9ĳ�Q dO{y���Kı>��~�ND�,K�_l���%��	2'��~�ND�,K�Є��j]]�s35�Sq,K���]�"X�%����T�Kı;�w��Kı;�g�Mı,K��d��4Md3.
�ی�����qCR�0"^8�=���gs̓�Zh�e���ވ���K�SsW��Kı;���Sq,K���ߦӑ,K��u��?����,K�����Jt�Jt���l�A����/O�%�bw���i�~��C�"��'�,O��}jn%�bX�~�]�"X�%����T�O�W*de:{���}�̆�mSΟ�Jt�K����7ı,N{]��r%�bX�z�eMı,K�w~�ND�,Jt���O[Ms�\�l��å:S���}v��bX�'޾�Sq,K���ߦӑ,K�2'���jn%:S�:_}����b�9h\�:~X�%����T�Kı;�w��Kı;�g�Mı,K��}v��bX�'�(��O�3TզMkZ�:�,q�-z˴�wT��=N�ʆ�\�%�3�a�&���N��!a���p��Kj����N��N����iȖ%�bw;�ʛ�bX�'=���?�'�2%�bw�����X�t�O�},/��sqV<����ҝ)ŉ��{*n%�bX�����Kı>��ʛ�bX�'~��6��� �鎔���+�%k�]zxt�X�'ߵ��iȖ%�b{��*n%���H��"�8n&�{���iȖ%�b}��eMı,K��c�)rjc.j�9ĳ���?z��Sq,K��}��iȖ%�b{;�ʛ�bX��[�������K�)����l����f`�/O��bX�����r%�bX��粦�X�%��k��ND�,Kݾ�Sq,Jt�O�C�==��2��jgm*����f�Q��5��4%vP��]a��g�}�֗��ԙ�5n�8�D�,K����Mı,K��}v��bX�'�}���X�%�߻�M�"X�%��R˩�[2氹r虚�7ı,N{]��r���,O޿�T�Kı=�o��r%�bX��֦�eL�b_z�Og݊��ٴ��t�:S�:S��o�%鸖%�bw���iȖ?Ƞ�"dO��~�7ı,O�k߮ӑ,KĿ�!a�U��hZ����N��N;�w��Kı=�{V&�X�%��k��ND�,��A<(���"k�7ı,O��d��\��u�N��56��bX�'��j��Kı9�w�iȖ%�b{��*n%�bX�����r%�bX�wG�̙��5��X�õ6Jt����r��ѷJ�
֞x��X���!��:��m�t��N�����]�"X�%���bn%�bX�����r%�bX�w^Չ��%�b}�#�}��.MLe�]�"X�%���bn�c�2%����ӑ,K���V&�X�%��k��ND�$�צ:S���f��&f���<�bX�'����ND�,K��ڱ7��ș�����Kı;=�st��N��N�1��iw��!�T�r%�bX�w^Չ��%�bs��ӑ,K��w�17İ?
2'��~�ND�,K��e���f\�.]5�q,K���]�"X�%��H�{�ND�,K���M�"X�%��u�X��bX�$@_�;�<��hY�͊Tq�*�f&vW0$��&Ggj�tp�Ny;I[f��\�3eZ�7(�p]BC97a�nt`��p��.�sn�i�+��vB�.L�n<\�i�.w�#�	\�e�X��l�u͎�]7Oin7OW��v:�h�FMv��U.�l�	EN!Hd �SfaG7S���	�kr�G<����-v+md�mQ��g��4ݩ����{^�'��pE�����kau����n�z"9�IK��gb�evm.o�Oӥ:S�:|=���n%�bX�����r%�bX�w^Չ��%�bs��ӑ,KĿt���\�ٖ�s7O��N����瞞'"X�%��u�X��bX�'=���9ı,O�}�q,K���l���sqV1�y���N��N��Z&�X�%��w~�ND�,K��l��Kı;�w��Kı;;�%Ψ��f�<:S�:S��<��D�,K��l��Kı;�w��Kı>q,K��:C�kP�3WsWiȖ%�b};혛�bX����}��i�Kı;�~Չ��%�bs��ӑ,K������?j�\����M=l�%����ɴ��9��惎�3K�4�۰�6ևY�3Y��,K��}��iȖ%�b}�{V&�X�%��k��ND�,K�̧�Ô�R9H�k!��pi���v�SiȖ%�b}�{V&�A π8 Ƞil�Ȗ&{\��r%�bX����Mı,K�w~�ND��:S��,�I�]s��Vi�å�bX�����Kı>���Mı,K�w~�ND�,K��ڱ7�)ҝ/��|��U��ͥ����ı,O�}�q,K���ߦӑ,K�����Mı,K��}v��N��N���X_Wl�ٖ�s7O,K���ߦӑ,K�����Mı,K��}v��bX�'Ӿى��t�Jt��=��oBk.v����CJ�.�n�[�6T���EA�����[V4�N;\�U�.�<��t�Jt�Oߏ�:xqbX�'=���9ı,O�}�q,K���ߦӑ,K���!/��\�]M9���q,K���]�!�9"X����q,K��}��iȖ%�b}�{V&�X�%��t��>֡Jf�2�ӑ,K��w�17ı,N���m9��J�D"�:1A~U����D�k��Mı,K���]�"X�%��!��oC�s,�f��ҝ)Ҝs��6��bX�'�׵bn%�bX����Kı>���Mı,K�=;�_h��Ve�j涜�bX�'�׵bn%�bX����Kı>���Mı,K�ﹴ�Kı>=���c&�Ms��9N��r�n�.�)��k <]��DV�t�+�[���gZ�7ı,Nw]��r%�bX�N�f&�X�%�����r%�bX�w^i�å:S�:_�hY�{���]�K��ND�,K��l�� �I�ﴛ�H'��j�$RD��wI����zc�:_���ܻg̴���xqbX�'���m9ı,O��j��Kı9�w�iȖ%�b};혛�N��N��>Yo���֬cZ�t�:Q,�$��o��Mı,K�k߮ӑ,K��w�17İ<�聂��׷�M�"X�%��;K}�R��i���X��bX�';���9ı,O�}�q,K��{�M�"X�%��u�X��bX�'L�m�.nz�Ub=vcl�Z�OE  �ۙ��|xy�q��Ԥ�a�?��О�RYfn���t��bX�'g�l��Kı9���iȖ%�b}�{V&�X�%��뾻N)ҝ)����Y���s,�f��Kı9���iȖ%�b}�{V&�X�%��뾻ND�,K��l�������Jt�Ov��6Ѧ�SiȖ%�bw���q,K��u�]�"X�%���bn%�bX��w��Oå:S�:{��T���:�Ն[q,K��u�]�"X�%���bn%�bX��w��K��)23�}i�å:S�:_�hY�����]�l����Kı>���Mı,K���6��bX�'�׵bn%�bX����Kı<����3�\�a�<��
�b�X��d�P\��1�l@�XU��:�Ɣ�s7�$5vGjk����@�L��M�P�ŵ���wN8^,�+��-(1���:��	
a�Y���m׏7C��^
�lC�t��6�Zv�W`��n)N�!a���v26��#P��V\g�\Bx(v�ۙխ6�8]Ԗ!�q��,�
m�V���fM,Fa�wI;�I$�-<�&�vsi����4�8���l.9e�YQ�-̲��6X9v��iG3t�:S�:S��~y����%�b}�{V&�X�%��뾻�@� ����%����f&�X�%:O�[��,��c�nO:~)ҝ,O��j��Kı9�w�iȖ%�b};혛�bX�';��m9ı)���[:��m�t��N��N9�w�iȖ%�b};혛�c� ��SQ5��o�m9ı,O~���Mı,K��Lsڥ)��˚�ND�,K��l��Kı9���iȖ%�b}�{V&�X�%��뾻N)ҝ)����ق�,�9���,K��{�M�"X�%��'���j��%�bX�����iȖ%�b};혛�bX�'�z��u��E�Зsv��쇇��:y�ƦS:[��`M5],Ԣm�Y��5�j�t�:S�:S���j��Kı9�w�iȖ%�b}=혛�bX�';��m9ı,g��J����S��N�)ҝ(����3"��!��oQb���U�؞�b~���Mı,K߽��iȖ%�bw���M��L��,K���{?f[����[.j�9ı,N�߶bn%�bX��w��K� C"dO{_�bn%�bX�{^�v��bX�%��R{4�;2ҕf��ҝ)���!&:~��~�ND�,K���X��bX�';���9ı,O���q,K�����g)�̺ѧWW56��bX�'{�j��Kı9�w�iȖ%�b}=혛�bX�';��m9ı,O��ײ�YU�`18�6�����cTnZ�T�S�o3(�.u��gI;�<,+�eΩ�&e�X��bX�'�׿]�"X�%����bn%�bX��w��Kı;�{V&�X�%�~�K=L�R��\e�]�"X�%����bn%�bX��w��Kı;�{V&�X�%�ߵ�]�"~L��,K�'�S�Ia��L�щ��%�b}���6��bX�'{�j��KbSB��Cg�� H��#F��eHQ��V������B��1������l�`h�#��"A A`+֩J�#2$%���-,,%�����Y�S6l4K�x��a�.�M4����sImh���H@�@�M똥����$jD @�)��!aIA�Q3�rԠ�`W�T"�U�p�R$H�����[&���6�@4@RM� o@R Hm!A`��!R6@�`�#FVVT�Ѕ�e�Jn2��D��@�|�� r�`�����>�*m�Q" �]
�����<&�T��dO����9ı,N�{f&�X�%�잝�/�fa�̸M]jm9ı,N�^Չ��%�bw�w�iȖ%�b}=혛�bX�dO�{��ӑ,K����T�%�u1����ҝ)ҝ>~�=�ND�,K��l��Kı9���iȖ%�bw���Mı,K�E�߹�Hm4!\���X ��i���ё��盞)�bm��z��!�)��uKsW��Kı;?~ى��%�bs�ߦӑ,K��u�X�)9"X�'��~�ND�,K�ĥ���fk5s4[,��q,K�绿M�!���,O{_�bn%�bX����9ı,O���q,K����g,��c�nO:~)ҝ)���֝<:X�%�ߵ�]�"X�"�2&D��혛�bX�'߽��iȖ%�b}��\괛m�t��N����!&���߮ӑ,K���혛�bX�'=��m9İ?>���	y��ڱ7ı,K����'��Jf��5���Kı/׾�&�X�%���D
�����iؖ%�b{���bn%�bX��]��r%�bX�x�˛�]0xsq���F!�n��8�f(�֊�&^v�~};���c'=s��lO����%�b}���6��bX�'�׵bn%�bX��]��r%�bX���kq,�N���=>m/��Fc]��Oåı>p�?�+�����~���'}����0��VKT��]�`ױ`{���U�K��� �y`Ԓ����;n�$�`~�Us��������n��X�hT��i۵n�!�`M�`�l�5�-�9��f䟐C���*�������ǵ�`I���7V�˷<-5�k������g�����n����1����м�f�`�V���l[� �m����Og�$�rq���'���{m�=V2J��Þ����`K){D괷���u¯���9;v( ���i\���Q�.�x3��1�\umV��td��W�<Vѐ�g��:���k�z���r��}M>�%S�����I�ɣ��3
�S1�AaK-`�Ev���G�rs����Y�-lk���eN����էd߶�`ױ`n̯�W9ʯ�w��`�B�'m]����0�ذ�fV�ۆ�v��tșm�2˫Iݬ����>�p�ܮr���y`\��MT�S�݀��`s�]��u�� ޽� �d��"!��pm��tZ�0�Ȱ�\���s��7}��Wv�V۞x�="N3Ѷ`99s��9��&["���pQ��=3�h����f99�9.�lo^ŀw�2���?|�����$>)��� d�����r�$����aN��������ɹ'��߮��;�v�Q��;�V����ۆ�\�ܤ���n�e`+U%*v�waMZv`{��?W9\��?~X���w�2���0��T)X[wn��n��{����>�p�>�`���sv��pTGlmu�)��r̅5�!f�ł��L����L~����|��W.��N�|��V�ۆ�\��r�A5�, �B*~��wtUۺ�>�p�W+�Ď��,k�XwfV{�U��\�g�~<�'�M��tZ�0���`ױa�q���#��_�}�߷� ��`I@�d�m�t+����.˞X��V��� ��E�RHZ�Mݡ�v����ٕ�~�s��3��w_����X��+jO/��b*˨笾�ۉݩ��$����Bk��oX��%z9n��H��ʻ3�3�o�z�yi�\� �^ŀw�2�	4T(�S�;�
jӳ ��E����\�l�?~X����}�p��UĎʂ�{�m]��Sm�Xc�X{�+ �v�}�"��<C�ݱ��K��{�I��&�߿߳�N����'>�z�N(%D����`�b'Db� �Mf�w$��骜��wtS�u�}�p�>�g������k߮�A������yN���}>�k@�L�6Ve	q5s�˞�B�E�I�n��(=��������WãuΌ&��8 ��_��b �`�`�`�����b �`�`�`�����<�����׿]�<����߿]̟�S5�f[�]j�A�lll~����A�lll{�~��A�A�A�A�u��b �`�`�`��u��؃� � � � �=,���m�k&k3V˚�y�߸lA�lll}�{�؃� ؃�� ��A���v �666=�����A�A��:����gݾ��]��M���<������~�y��߮�A��������A�A�P�D 9{����A������a��¨J���;�'Rt�������b �`�`�b���^�o��؃�lll}���6 �666>���A�lll�j!  �Pm �#�E�Wܧ�fg��L˚a����{w�T��iթk���Q�n�ώ.��X�F��Xz봂���6��v�K�CF���;b���V��E)�湙��e��1�a��)�XF���f.����q�8Û�3vH���K��1upS���Α��˭�kl�v![�R�a��<V�����ĖֺPv��\�Fn�r�U4m��q=b̖c#@�f�߲t�1�]|���rmk�ڛ%:A�$�ڙ�)ى�a��ԛ�@J[�Z��i��o��w��:�������b �`�`�`�����<������~� ?��A �`�`��k���A�lllo��2�5s2fMM�5���A�A�A�A�}���A����׿]�<��������b �`�`�`���{�؃� � � � �I==L�2��5���ѱ�A�A�A�A�u��b �`�`�`��u��؃� � � � ��^�v �666=�p؃� � � � �'�����a�&���]�<��������b �`�`�`���{�؃� � � � ����b �`�`�`���߮�A����[�~����2��Wb �`�`�`���{�؃� � � � ����b �`�`�`���߮�A��������A�A�A�A����sYF8{�V��yǆE�Z��P"�1�ͅ�hKtRAI\ٞR�`� ә`�w���A������yw^�v �666?w_�]�<����ߵ��b �`�`�`�������5sZֳ4e�fh؃� � � � ������Q�i�y~����A�������؃� � � � ����b )�$�A��������eѭkRY����A�A�Al�ߖ�9�w�2��ذ�EB�x˷v�m�k �=� �ve`ݸ`~���߼�v6��ll���������7�p�>�`G�`�+�^�>9�>�c5�1�6F��,ە�X�zX�N�p�A�]��v�l������*v�l��r,��/���u`j!��8���եv`u�`f���>�2���0	�HJ�A*v���sWrN{;�'�w�7<*�`{vl�+yUʡۗ�}�b��KTI;�;n���w�2���0��X�'��C�����I�Ȫ��R���ۆ�Wv����X{�+ �����b�.�3,�ےq��)��,�������6t�\��Umħf�\� �=� �ve`ݸ`mh�S�v��M��`G�`�̬{��z�����b��,��;��n�e`ݸ`uȰ�ذ@�UK��E;�Tӳ ޽� �\�rN{;�? `1��  D`��@@��o��ߦ�<��o��*�+ZWf޹�{�ˆ�ۆڄ�p�Ƌ�M�5�l-+1��r�t˲-kVFR�,T��B�($hL�VQN[|���-���{p��=\���� l@�E䓵t�HN��ˆ�ۆ޹�{�P�'���n�
��7�p�;�"�>�b�;�p�$�P���un�)[N��r,��,��{��Z*��]��Sm�X��X{.�nz�X�����p�QHA�FH@	8@��AI0�T%8��4Čc�#dJ,i) &�FQVU`bU#2Ru<��J@C0HF^�� E�	#���8mK���T���0!����5�����"A���؊p$j2�H�qN, Pu2aCL �DIaL#�n�i��D�S�g��n���_��߰  ��ޠ 4j�6�y�'nۙ33Ki}��BAИ�cT�T�8��n�GU��������[��l���RL�5�s.��Rtݭg$��x��Z�z�R�gdJN�s�NI���Vެe���M�"��J�nK!��5hi��������AW#�}p��H���JI}���n�ܝaP;mjzVנL�Oo)6VT�!��ɑ�2�e4�*B4<+���� t1� V�U�O�2���v��)(�S
���_<y�g�tF�Χn�B��i�U2�Q��n@!�7�#�3�Ow��h�ơ� C=\s���.ک�\�͖��]n��t$crgMtpcnv蛖�t�mc�!ە����k�V�,��g�]b����p�&F�88���Ob�N��Z��&�y�e���vsn�jUs�uv�v��\l�e�¥p�ܔx��-�^s�RZ�R�ݡ�pl���VJ��eڴZ� A�t�;-F���7��_'�R�T�.5�6Fd�q�s��xQ�ʧp�����=%lڰ3���__}�����ݘCgt��j&�آ�l1*C���*gn���͔�[vv��DI!�mO �TU�N͑^m��=��B��Uu��%�q�i�p�-�!��<j�r�N̸@ҭ��F9[Z=K "����K�ڹz����:��CN�!����L�1��-��X��Q�f�vn���m�:$�eg��ѝ̻-UQ��W+G�6����,Z�uq:"qGm������l�m�52�r[+F`�pZ�溶4.��MacW)P�� Ҙ�FȜڣ8��e^@Ce�ª��hK�Ĳ�^��Y��m*������y�%���� v��:�h����4�Ac��[��v��J�Fk��6{�g��-��9�؞�N�A���lb�i�Ɨ�� ��AAl9�m%,�r�ܘ�j� յW�	�C�P��j@J�n��t���H���Lf�ˇ	c�����l�#qnRͪ����׺b�]*m��;Pu�8�tSH�J���8�(�<
|!A�	�����ө�/�� ��l��lw�hu��&��/l�!Y�)��N\i���b�s�7k ��Ç6�e1�&oaҚ�of�v7=.�KЯf��j�۝�m#(��+�q��l��.J(�Kv�֥�\=��&:2���{N.�<����n	��@&��Ͷ�����:�'�	ާ˃^!0�2��'��o8"����B�aZ��{�|�o</���0+Q#f6H���_Fm�6^�!|xy��.�q�k��J�E�-�����;���\0��0�Ȱ�ذ@�UK��E;�Tӳ ��� �\� �=� �e�?r��q"#�o��J���V�ـn�y`G�a������&��M��� �;t�eЮ��{�ˆ�ۆ޹�t
���v���i	��;�p�=�W*l����}ŀw]#jZV�y�n#���zz��#s����=�y��杷\3��X5�H�ȮvbR�ym��צ޹�{�ˆ&����F�Z��˚��}�{��`����j���_�\��5�?<ޗ��7�p�;��IN<eۻE6۵�|�ǀw��ov�w�E��Q[i�j��n��~�9U���q�������`�`~��]~�x �U릨E;�Tӳ ޽� �\� �M� �e� �R��z�fZ�bSl���D6��ɮ����u�k�\�Qf�l��{&�����H�����\=_�\�:��{��?{�!+U�J��I��Wk �M�?RF���<�r,��-Q&�vݥnk7$��k�rN߻���!�UN�`�� �Z�q˂�1"�)����?r�I���ٹ'ol�V���wV�+��9��g����|�ǀw��I����b��v�7o �\� �\��Uu�y������ܶ�=���)Uj�fAv��I¸������W��7qsxN8d?�{�������n��n��uzy��`ݸ`�`u"��6�v��cwo �e�?r�"l����� hj�t��wJ�v`ݸ`�a���%���n��`�je&DU���һ0?r����� ����;�p��W*��8��@�T~O� ������~�����%N�$�t+��|�ǀ~�W7}�>l�z�Xu���Z�t��������a�WUO@t�:�x�sN���R����Z���t�I'o �e� ��� �\� �M� �i*#���ݷtЅv`ݸg��W)#u�� ����;�p��\H���/<V+�waJ�v`��X�lx~Kw�� �/���Q��[wh��v�����\0��0�Ȱ��DuM2��ݼ��{��r,�6<��q�s����R� ���"N���5��l�.4i��ヰ��vǎZ324��K�g���K�"�V��1tk�9�vݝ6V4��Eu���8.%7:t�g�3�7։�u�j�5����1Ӥ�tW5q�lsYLv{���]qЧK���y�#��7fG���1n0�pӉ���i��fF,f�r�
�up�ت��8��-�}��a�Mg����uFa�A��`{�;���~~]���y�ԫ�aF;'Br�
��Y;s�ɱM7��[=�g?s�6�N�U�wJ�v|�K�0�Ȱ����\0QV�RdE_��+� �\�?��I^�x���ۆ{��P*��5N�&ںJ��^�x{.�nWdxuА�D��t�I'o �e� ��� ��ܮr���<�	J�?+Wwv��Bـov�uvG�|�ǀw��}[[b�����ثg��˷\�Q�����]�G�;�"nA�5f]�6�f#H":��������û�ˆ�ۆ��Q��+wh�i�x�ly|��r�����Z7}~0��`]��u"�uM;U|����w��ov��W9�RZ��xW�� hK��8��SN�{���<�6<��TU���IU���һ0���u�y����ۆ�=�V�MZژ�B���x�wD�/\�=�q���<=�7X�,��
��;x�lx�\0��0����BB���N۴�v��`ݸ`�E�|�ǀ}֒�\V����˭M�;�u�'{��ܨ�� W���#��΀��n��܆͸`h�(�]��]�+iـn���.�nw��)L�+v_.�X�lxd�`ݸ`�E�oy��Y�t>�ݫt*WVXI���l�<!�Ӟ�q�ڱg����k���A��F*�cwo �{�uȰ����:p)���4��7�p�7^ŀ|�ǀ}%� �CU18���Zui]��ذ�����`ݸ`ڂ�C�6�ݫ�X������~���rN��znMED�b�TNԭ���.����I��-���]k.��i$��Ip�7�p�7\� �{���d�����JDU�Dۛ�-֡{NK��f��\Mtㅭ�[[C��<i������π�/���X�lxd�`h�(�;I5v��f��X�lxd�`ݸg���H�ȩ/2��ݗL�N����vK��ۆ��X�J*N��ӵW��xd�`ݸ`�E�����C��SG����n�`)����m:�r����D��2�w@�f�Q���/>F�#Iٺ��L�2�Rq�m���ֶ�e��ŧ88H�p�m�s�qF�` �����].��uʝ�-.����LC[�)���j��v\s��h]�Kk.��]�b�bS,���p�2kSɴO���;d�ؤ����U�n�D�ѿ�>̑��v���oOm���>�yyB��6{��?{t���c˭c,%�i�y*�낪���pǕ��(n��[YϜ��N�Ut�N�+��$~��>Sc�;%� ��� ��Y-&;hm+�V�`)����ov�n��t$-R��t;v�N��.�n�`)��u���]��wMWf�UW9Jl���X�lx�r�����Iy<v�j����f��X�_���o�~0��0��ֺls�֜��.��W��gSm�lqմaL�TlV-�y����:��e�#�Wf��~{P>ݽ0���;׺����\m;T�cwo �\��B���sj���f_Lz�X�lx�8��v��f�ۆ��X��xd�`�j�'Ut�N�+� �r, �l��\0��0�
�+;��wjݬ �l����{<|�~0�"�?g�o��풘*�F��0hL7XT��s!u������)	qV��.
�%����;%� ��� �r, �l�� ��wwn�
��7�p�7\� >�/ ��*�=�*K��[waI���$~�������)��K�(�BIYH�##0���H�	�FU!E��YRP��FB6�8	r��|'D�1b�H`�@��>�.��y�oKc:D @ wGh�~&D�8��b���%b�� �Zȇ�ʤ 4l��Ic�JI1	��R��3&����0��z�zq#۞jЏj�~|��@D��g�E���
�0 �[S폇"� B��:gbvK`Yg �
�"E�H$H����T"1`C�ی�m�w�'u߀��CD�����h�RN!ǡDmB�!����@<�DX �Ap!�x��<��y8��1T������znI�{^��}Ӵ�̬e��ueڻX��Iw�׀w޿�n�R����*u�ӵO�ӻ��\0��&���?y`�e����/k6c5�1��v)rrϣW	�ݞ�N�J{xy��@�Pcu�m���ɼ�;0��0�"����\��7޿G����%WL��һ0�"����;%� ���=UU\��UUM����?�fFZ�V���������x�n�ذ�T�JJ�hI��Ip�7�p�7^Ł���U��)1�e`@I$"��V�Q%x�T�R�H��^��w�ߋ�����P����q�lB�0��0��s�\������.�r���F:�S@�|���w���m�@ʹ�#+�--�k��@�iΔ���v+n�)6��#�X�����`�p�;���mV2�캲�]� �Iy��\����� �_�u�X�J��Rձڧ�i���.��0ױ`�K�:�:EN:�mN�wn�ذ�%�{��U.��� ��xb~��Zujݬu�X�����`�b�*�ʪ�U����yתy9ǯDI����rR�Ys;S�7U�sǁ�=s۱��xv��sl۱�S��xW�2s;j��C���W@m�/c#�>��L��1k6�Bbѷ�%�P+Îm��k�#�g��r�]Y�ㅚz2�q{g�� �"�X؍+�p�m�#N֍��+aX�õeHPmWc�`m�_���|��Uza؜��0�kV-�WM�5��U��Ó���˚�L���v��\`���t�����l����1^V�s��iC˰**}m���z����u�X�ذ�T�SE��-�BWw�}%�?����$s� ��, �IxzЁl.ݻc�lB�0ױ`�b����}%� �H*I�Wi�waM'k �{ }$��.�UqIs� �QR�j���e՗j�`)#�>��n�� �{+^�u(�#4]j�0�%�]��wNn@L,XǇ����C��������-}��.�ذױ`�K�:�:z�����L���'{���^�Q(��r�z����y`}�^��QN	U�-:�n���, �Ix�\0ױ`�Y,wm�
һ�n� }$��\0ױ`�E�wt�����Y]�ܶ�w�o-�O�I.y|��X�H��ۤ{�j�77�lх�!R�(��K+
��3��3�tγM��3P�Qk��:mJ-�����r�u�X�H���`II6e�v��SI��7^ŀ|�� �K����?��$�gH}�9��k����{�nI�{^���4���bD#Pg��s���9˹'���� �QS�]�Z���x�\0�ذ������@jdE:��N�z�,�UU����K��>����>[������gc�6Ytrfٿ���{����M�k��^���g�:�urb;9�t�]"ӫV�`]��)#�;�p�7^ŀn�Ud��n�J�m��>Sc�;�p�7�b�:�#�U$lt
�����m�I]�w�� �{���<�ĨR5j������u�XWdx�H�Nr��Q�U*V�P ��FM��6;�k�rO�bBM�vݷv�v�����UU_���~�����n�� ���.RWB�(�vqdH�%��e�]���͍-�\s�������84b:�決��[|;����u�_��s���x�*�^.حS卻x{.��0������USg��*��U��f�z�Wdx~�K����7}~0QQ)t�]"ӫJ��:�#�>RG�w���UW�<�	
����wM�Wcn��<�W+w���$s� ��� �Ӥ��N>�v�]��݊��ma,��k��5�e�4�r)�d���$k��zlƵ2���u���&y^�sA��\/]�<�u��B+W��ZKl�����.:���i���D�Ϟ�=p���7N�V@�b��UwU�;K���Y���hkl�)�ˌ���d��e����QOoO2���yu���9�S�5PZf�5Yv�t�:I�|�y;���lk4�n�)��+u�e6�N�S���X+�����2Mbᕰ,�wE�i%v��~0ױ`]��s��O���r��p�|�.[�7^ŀuvG�|�� �e�?��U$w��BM�-�n�)��`��x�H��\0ױ`��J6�lv]X���)#�;�p�7^ŀuvG�uh�*u�+T�cn��ˆ��,��<�$x��yv��|We�n��z��NZ���W5�
41�81�~�3�:Au�CUwE>]��'g�H��6<�$��+� ���E�^T�뤪����j�I��}��Ո?j>��yʫ�XZ�� ��u�X�eK�wI�WcN��<{.%#�X�O<��H�):���m�I]�{.�ذ���)#�7ZJ���V��v��v`�b�:�ǀ|�� �ˆ�ڗ2��:�J�;�8x��Q��tk��7)����!�]:N��Z�A��ں��N��6<��X�\0ױ`��J6�j�wWV1;x�Ȱ�`�b�:�ǀuh���]�Z��v��`�b�UU��\uʯ,���w�y`@j�tS��t�'f��,�lx�Ȱ?UUqM�x�"������Zujݬ�lx�Ȱ�`�b�=U^em(?�2����ط^�"!]�ļ�*��݊5�g�x6y7ź�p�Y� ��`�b�:�ǀw]	�]�E�i
�`�p�r��$H���� �9��T��Z�wC��+� �{�6<=\�R]���7�� �d���Ym݅4��r�UKs��f�~�߮����ܕ 61Q� D�	�4 ���z�I�����]���N��r,{.�ذ�"�7���/���I�V�]n�0�l,u�nz7\��tT�r�qqD.�����Z��v��p�7^ŀn���U��a���� �?%��W˴�RN�u�Y���8�#����y���j��1K����Z�k �r,�$xd�`�b�7H.\�Z�t;J�ջX�H��p�7^ŀn��t$k�v[�6�$���.�G�߿_���~��n����?�TW��TW��@U��
��@U��TW����J�������
��@Q����+����+��TW�+TQ^����Q_�E� *���@U��TW��
��
�������)����w�/�8,����������0m�>�'c�� *vTض��,�R��q�̫W���6 @$AI  ��B@
� P����� ��=� 48�����c�OF�a�2���;�۸A��v�'�k݅�X(2t���p1{��	zc�'x�D 2��sIW�m�gZ�H��M\��2�Hz�5KF����9����TѮ���lz�U�W��U����ѯA�{�L�@�7F|��;c�BtUa��9:5��Pᮆ��^��[�X>�½�hkA�=n�94�ֆ�}�UG� �`U�۸Ѧ�kG׸W���� :º93��+���]�sv�i��6o�   ��    ����{��h
 V�A���vқ`���+�N�
b�(d����C�ttӓY4V:͏j��  i��IR�h�    ���R�F4�  &10`��T��E �    ��5RaJ�@ h    �J@��)�Dj��h`������� �  � ��_�?l~�?���71�~�d~�PCe,?�+�*��*�*?p61�<���cc6����t����2D#Q8�TE7����61Y�������l6R�Lj�ԅ��~E~�񚿓���հA�A>�Mo��ϲ�\F:@ڻSh1�� B�qЌ
2�<+r�UXk��!�d��p!�!�
F0/5�rC\���/s*t@���B0�� ����ǐ�BX��̳���^�%g]������.������\Cs˫셗V�˶��a�ĀRF��%r��x�$��ea��J�*�BHPbDe����fYʴ&�,U�X&l�l�t[$ܖ��(R�U#G҆;�c�	M��Q&�u氳�].�	�!z���L�Kd��xx��m0�����A�פ)F�\
�g�ʂ쒴� Ȑ�"YXʹKze�� �X����Xw����xPB[�`�h,0H4��`1J�-��nS��-�Mk|D瞽�j�����[U�i�F����@B�HH��1�4Pr�R����y��S%�����\� ��"Q�N�[5fQW>�+*1�2�m��_��
j�ɫQq��$�m�#�KzB���;�7s��Ǩ��Z!�i���w�q��#�zs,q�q�[�ŴT����F�sq�1�K
B4Y��cfˣĉ@k���u�m&��8ْ�,���s9ך����si�;9�8M!�$q�V���	ޞ:�9�-8��8ĆX
H�j2Ͱ��q �h����p���xl�'.�4��/�x��@���H��1h-"��.rxW��͜�N�:���B�,ǀA����,
B4��U�kTJ�TJ���%Y���n�
���%�{,����l�ѭ�|z$���ʶ4c! ��ɚ�3R��w�Z5�e��޷�έƜ[��n;�Ǝn�x�:��vp%xbjYG���/_��BlNZ�%^0e5����*̅�<4�D�	�-pѩ^j�\�k	��1`�ӈ��,1�Ai��H!z�Z`j^�ʳ$V��U�R��/F�!%�-|��v�q	'�g�2ۘF���F%���)�In[���V�.-d��:�=o-�Sy���N�
#E!C������s���޷ֲ΋8%��=s��rsw�Q\�9XW�48p���R<8<�N��Qq��5a)�kR�L��a���˒Hƍ,Vh�4����)�57*H��NԄ���$$Is7	������*��s�s�<�q8�Ֆ���<{�N$�[�(���Y��㤅\��)�Bt 2�Fơ�8�M0�z�(�k��,aA]nU�k�K��փ�񔗛�k~J!���Iwm�˖\��T$�a���{�D׌$a�C
��xӎ�v�㥸�9��60��R��%Y���H����m� =���y�t9qt�I����C�'��K�p��x�ixXRʭ�i��(�<I@�\E�ͭ��#�qf���m�v!���m8���5�8jbE��i4
LM&�%6��!���Q���JT"��H�I����4i�g�
l1	� E�"Qnkg8�8@�.ԅ^_��\�lx�pM��4��4o|NJӳ��Ξ>5�:<��x���ٺ�z!0�%���#/f�Q��E�C�fYݦ�o��՜Κ�ۆ�B�����8��0m:��@���)m3{<ŷ�addn���s�j����mԞbst�M���E�`�4���7Om��xm��9����M�wo19ׇ�C�w���a��"PXbE ֻ��04�h�`�,�;�J1ѵ ��f�J�5�f*B�`Qdi�4m�Y���`ġ�ѽ�
l�[�@�����k
Q�݁��4�6F�5�y*��]»s���l�j8�z��;���ϲ����u�77��월�`��(&BJH�-��M����Y��*�vn�YE�1eݖ��k1�7&eVN^�B�ε9�Ή�t�\i�Օ4-��D�<%�a&l%$8K��B��\С[�HUd�ה	���f���<���D�� �h儍����A2������2h�Y�q}*4�y�@�!�Ka;�p�[��e�%���^^5���F��r�v��*�y���� ����R=�R0�b`ILR]��Y�/~Y�r��f�A>�!x������"M�%� (�kSXב�p���8f���{dP�B��Æ�̔u���$(Q!9�tT���~s�? ��h�>��S�w����������?��   H�m� �    7m� m�    4�5ն9r����S��y��;bW�A4�JF���ȩ�s��N�Yv���g	�!1��^Xv�9�m��l�v�R��ݎ�ms2�\U��h�n��W3����)	��ùtX6��%��_�@y�@�\2��T���B�d�Kv��Y���v%'���q����[R�<�G,���]U uð�K�ffTJ��ʴ�WX��=�/'W��N���t�&�;q�H�mu�@ M���� ���� hF�<m�k�+�6sJ�!�D��ٵ����`l���[=��@w5�}�]`�)W(�Nյ���*)�pj�Vn
k�Kֺ�ە� ��F�k�Mzl�h�`|��}8Iͦ�b�6۷"@  ��[\�m�   V�H$�n&ײt�I�   	   H-���� ����Z	  ]6�  :�   ��&����� m�     p    �  �  -�@   ��  ۶m  ��[@ ���l 	e  m���m�ͳm�����,KT�UR��@   6� $6Z��    h $�6��n9�lH�u�� 	�   ��z�C�  H�g��	m$�i�m�	)@ �ḿm "��^^v&GmԵS����i8#X��F��I���Ŵ$H m�!&���u�6݀�[�۶l -�6�&�t$ida��#����m�["ݤ��6��m�L 	lu�M�	  �^r��ɰh�n�� ��m� ��4��l�2�T����UT�-mA ��ѷM:,� �|����6tی�/���  p$�mq$����n[3LH���m��6�z��JQ��������y�]��`H  @  sv�Hl�ɰs���»P]=�WK���aۋ�g���T�j����I��P�;���,�0Ԁ$I�M�c �%k��q6Z�i].�q�M�m�\� i�V�m� s 	��`UG�AնY��j�6F���d_/P|7��� �  ֱh��;��	m �I3�:�d�䍺���mQl�ԉ]�ۀt�m�[k[p�[B@[� �@ku�8�D�v�Y�̀]g�i�L� I��Lۆ� k���MQ�$� -�l�4��[dr�b{w��,ބ��n�-�m���l���e $6�6� Mm�6��` ��K�8Ýo[i&t�`%��r��j��xMɶv���ʰ�5�8 a����V��`8   p [Khp� ۶�m�v��:Xm��JQ�n�l�:  ڶu��GO7$�K�����v���� N�lm��Kn� 6�p m8m�� .� �$ XI� ��@sm��g�����JN�̪�5�9k�6�ַ$�  ��9o[d�m�`� �	A�˦l�  �` 2ܭR�٪�MXW�S<V�UUҪ�@@S�'@n��^��i�u�g�4W � 	 m��ŴCm�� $�z�!ŽD����`H$�lN�c�YZ�d�l��m�D�bm�     -�@� ��p��Ύ`-$-٤Νz]6Z8E�b��� n��t��I���r���t��l$ t��m���;e��ʾ+��Uڨ6�ہ�l�n�DX��k=��d��:�m������۲NH(�.�l�\l�}���m�  [xY����m��� k<�nm� �L���<h�8q���ɐht	ݻ`����ܑ#��� ' 5��X �  Hh����N1Vݶ����� h�  �$���`�h����86�	6�h�j�N�]R��<���`�� ��� �ZͶ   HN��i ��pk�v��m#^]  �Ā m�I 	:@�-�kl��Ā�`R�k�$]V�����c@�j��.��3��mǛ��9��v�8�j��,�U+̫ 5   �vm��n��V�4�l$āq�   �`�m8���6�m�-�@ �(�[@q -�lz���-������!Ŵq�mU*�R�1T q[Ŷ� q�� ���ݰ�e�N88�6�m��l�h�!V�pz� ݬƓ -�[&�} �VK@p�d�{�k�c��n� �@�$n�  ��'].��K�wJ�Q�N��۟X��P��h⭕j��
]6[Amm��l $ m�i��z�6�m 6� ��	mp�nͻ� mz�+i�  l�i�Z�m�[d"�!oWm��a�@lӷ`-��uT����UUJ�����Z�%�B���ﾀ   m��*�֠#�����V����  � -�  l  ��v �\�  ���� Gm��8-6v�� im��$�W�@۞�,�����?w��
}�|�DT�T����
z"���y�b�����@$
����_�B���� ��D�Ae/4�#��W��2��M	�� ��x��T<��@6p� �(i�@6�)tCA��+Cm&`�ؽ��O 4)۷c�n���l
�:�<@ +�bq���m�L�}8�z��I"^*�����<])�w�g��>�}����@ׁ��"C����Q�y�#���u`����0�
<�%��8��R&���h���ݔ�)�E�Z�ŵ/�A�*<T8���b����Z/���h<4�����3�:8����,���H�|�Ah8��^�M�`p4y�#����})kR>���ETt�#��b��8����^<�#�u��H��a�X�B,�M��%�������X�Rx�_�����$��B��H�"AX�u�>��Ywr�f ͤ�B'-�fɻZ�0�h���hf���ۡ�ۉ���9�W��N�h��[n�z��]Y;XQ*��E8m)tn6���,]��mn�6�p;Mk�)D��-��^�����:o�y��ŒFp��A��'$��*v�]�9JPi�U(3�����Ŵ�"�r�<M�[g�i�"���C�����MC�=]����F�c�X���&�6x��9v	xhw\yTؕ�ם�n�5��ݜ��f��s*t�F];�^�ɚ��u��鰖����j��4�u�U���Ȓ8�:A�ݬoN7a��`hwXUp���m	JC2�.�P�i�����uj�I��a��K�=���F��q<�����Hʢ��9�=��Y��v���6w]��%3�Ӎ�����9�=���M���, ,]e˚xsS�{!�����K��x��˔x�u� �U]�l�QJ��bt\+��ی]����b��Hs��k*$5���T���d��b����=�]�m���mn��PT�+;g�V�n�d����.�y����F�yYM��d�&C.T���j��z�� �^��
}:�:�|4'�AG`��ț���e��e�.$�Y�P��5�K]Wh�Y�(�$�Kl�#v�=Rڥ�\�C)�;t������E�Sjη,��tqVEk��Y�kh�kgst�+]�<pD���4���CR�V�jP�[�˴M��ⴉ�p殮��J��������L��;������q�r��p@�c��E�t�rr�t;�:""�!��+�������}�eb��CM�~����Ka�����i�z���pXi%��1��mj�'}��nt.����6�YU(�n����,l�4�g����������h���%&c}�舑!���w��0�nX�5�l���c[M��-��H���"�����,�n7�$����!��w�E{�q�z�V���I��q{�a�z�֨��S��m0�>1��mj��C�puL̰��pfad7	v㭺�n1˞7��F�4�nLv�X����f�lh-��n�樬�l�ޮ#NGxXi%܆!�R�Q=�)SS̳Z�ݞQU~T)'CO�fbZ���Z$�m	I���2�C�CM�[��b2Ԥɗ"G�N�HJX�YF2�պ�)C��D4����C�f7q
�'C.QiKq[�a���֨��S��m0�>1��� " =|�����\�l���v���{`u���H��TTث` xD(�� �f=�a%2[	���<���=��<���]�k��$څ�˗Q�3�ɹӔ��k�۵ү�u6cw���"ezH��>1��mj����h���%&cwP��u6aV���^�N��o�+u����*���E�-�n���n�Z�� �B4�V7a��zm�8+3��#���j�uŜF�@�9��"����sÂ��gg<Gៅ����9�B��k�4I�M�a���=Xԝ%hӰ�m6vW��:��w�:՛7IUp������$�Nu99�z꩛��2n����؅�&ݚ�.�}�Nfe)I�i��>8c3��P�P��Z�l�����+�6a���Jd����y6cwx�n$��P�f7q�Q^�tϓ2%'CO�e�Z��t�N�v��l�X����2���s72Ҙ�V�Y�����y�Q]��d��Oͭ�n���z/���c���l� ��:_�����̇(�����2��CkTm�)�d6�N�v�=�C��Wrw+C�-��}�tDDz��{��6�t�!�:�q���<ݻsN.6��Tm�����w:��=� m���Aa��^��>������'���!Wy��Ps|�4Z�`��5���a��%&c��2�En���*ӳ�k�CM��r����f6�FwJ�#]��ҙ��00q�,]-$*ˁJ:5�����g����Q���V�m��i��� ��آ������9��mɎ�C2�Wrh�~��Jd�����CM�I� XQ(���9Y��8��I�]]��{�ns����n?~��|����,+BlM\��rݞ+<�Cw%r�%<p���e����P��P8�BRf7چe���4хZN���)�ڢ���6�ZN�.Pi���P&6��Q���V�m��/f>��1��+� @n�g���r�V(���a������$��q��X���l�w7RPӭ��z��C���.�76�x��ܛ}@��g��V�[�k���c�Nr���h1��CM���`��(�z���=]���Yy�S
��P!�� p�J�2��m�"s���ƺ�zI(�3!6%4�jKe��/1�Q]�+f�ޒS%������ٍ�H�4`%��Q��+&=z�ި�\��M%'Q�1��m��A풁��-�o��\��w:��OT��V�^�5�.C�AY�cJl�s�;��o�����+�Q]?��U�+��A�-��*� �:0E
���Qט�WCm��3f2�#��/u�KCR[-1�jx��TV�7�$�a��QY��~��>�;w�[M.�4�p��y�nt��M�i��v۝��+&:��Q�#|�$�:x�g���܃�%��%�c}�e���8F��J�(SBB�eYV��8���l'�R�sm�;â��)�rU��F�Z>�(֒Z��F�[�4ӝJ�o1�so�y����t�D��X�����H�M��k��9ܳ��N�u��79�$l��Ql �uB�@!�̱؅�[,ȶ"mz�lB�ߍ�!����K�FM�?�QE��R��R~� ��4|(�Z,�|�"� ���g�bӾb�j��ٹ�ކ�?2%�cDDGw�/u
?�"��*��e�A�-��!�.|c�����;��e�̄l��nt6��p[MJ!	E	O�D����m�NǏ��:�@��|���	l�ُ��� �<������ ؑw��-��n����- ���g(�q����6�ps�3g�=�_�ْ�Ċ�]!�q�q}@���>JG���<c/������BlE����gn'S.�U0e��MWj�W'��߰�yEw!G�*?t��D��v�����7qZJ�Ԡۖ�P��7q�Q���V�m��a�x�ި��.�-Il����C/=�(����{9�e��`�K+����W6�q�<<�[���v2��ѱ]����T]���$��۷#�Nuf-�� �tl��۸U��q�>�n�u��gC$ݰ��d촤,�l۞$h��V��87)�s�#�?c�~��A�qu:B�mhb��{��%lS%�ޏ���q~܆(����yF���ԥ܃8cw��^;>m�mW<c����A�k��%���>#�����+�"��;>?'��i����8�}ށQ�>��W�%��m���e!#���WHm�ۮ�g\�-.͆R��_r��<{��w� G_��WCm��\�4>��1����C��G������-�1�|�}�!��>��ş�Ut�Ĕ�l7C��oڅ"���n8x�R��3�
>7vr�X�;O���.3�CSc,I�-(A�n���ʹJ��eߧ~_���gＢ����İu6���}��A�����x¡���?"'�UX>��+u����4�E� uQ֦F�w�l�]�ݘԷ��Y��N	�K$�sd��z����a5D�O}'ޔI���L�sd��9�{�g��mcM<-���SX4��3lnCd5�mfO��J$��g虿�l���`&�Nq%2[E�{y� L���I��L���Iے8x�I*�L��l��� 9$��{9��$ޑӭ		6�}<W�$�҉=�������|"<�_�'�rOɴ%�k��?�Q%�g�� &o��NO����޻�;4���=u��� �Jї�S �s�4�!zRYn|I����f�[$��9L�=�D��é�H6��'�s��D��҉."'�,��͒z�K��{��O��$�D���=��&���*I��/��-�4I=Ҽ"d�<�&��>���s��K`���'b~ߩ�o��'�I=��s�������\ŗ����S$Нz[+��Ž�dY�MԈᆠ��"�e4f��P	�[�o	j�Y6��61��K�P]5ɯl�ģ^526�-�v썫c����e���[�t+EuX��{�|�ҏ%���3b��38ܛ�)!2HM�MI(�I,$�sd���K$���O_?@�$ޑӭ		6�}<W�$�҉=�����6I�����%�h���K$�<�&���T����p�f��-��L����7����3��D�ޔM�&���r��ܷD��l��'{� �ˀ����Ӿ���fnh�H[0;K���Τ�u��d.�g�Y��<��I-<��>���� M�S$��k�R[,&h�{ez"�B�#jq
lJD([pnl�Ãw;������d���>&rt�Mڜ���-���DOoS$ߵ���3������$�7Xi%^�&N}�d��(�����{9�I� ���Tݒ}<Q'��K; D	���d����&��|�������fd&"�s4�☀�m!���9:��}P<����$��D�cG�4�$L�6I���&�[$��Q$�J$��I	�-�&�[$�������O{�$��R�Ö�n�9<Q$�J$��d��l���hjKe��N�N^6I���7:Q$٭��MjZ��.��V�a58��,�Q� d�|�@��� {��uI�������~����ި^�y��tw� w��{���}P:��7�frh�wer�Mn�Nd`}��1�(�����D�sd���$� ^�Q'w��wpto��1MZ0��n��%���WJ`���K,X�����~����ި���ox�������p��@��T�kD���	�$��D��l�[��nt�MR��K`���'����o��&�'��ޔI;rGXi%D��l��G��Ԓ|�\���fI,�|��U!��֙(�O �+	� �=���o����f��[h�9W8ӆN.m2��okX;@0×HA�CUH�.��&	n��kP&���U��� �py���lR��Vڪ���u���V擉�\;��S\�f�ME��kI�ѥ�{nǈ]s���[8K�^���zU��)t{���go9�tmi��4��j���*��j\Ck��j��mH������^�-���,F8��[%n�.�S.�	��X��@�u6x��g���F�dXG%�$ֽ*մ/([R�l�$49�lv�c�Q�U�(�T�	"��n�.^���v{e��Ȃ�݋��l2m�c��Єr��v��主a�Ĳ�V�Z�.\6-��9vY� �Di�xcr�b�C�TV��u88�됶k��6�pق姒��rt�$��3���q[�ϓ����	�TZ�ŋv���-"��aE��L�1o1�#*��h/]�n<�a��aXҰ���SXi\e��Y�Y��o*ǇM������%N*6�M<F��U&F�T���V��9kE�W&�9�f�t�j��n|%�����̫j������6�&Mi���f��`�mέK<�]���ʐ#lJ�0:S���um,*�hjLܨm��E��Lt�7Z	5��	مv������0��WTU��2�]\������@P�(���.!H�V�������REk�V�h �i�iEo脓�Hsru������^9SkC��[���ZA�a���!�i���t̘�� \
I�0��\R]FWh��YjQ���h� n�b�˞���؝ ���p�t��/u]t�&�$I�ΪEc��͚\	ܓ�������۶�%A�b6眜X0�����œU���n�B9v��� ̔I��� T�}͒o�AaN�!��Ol�: H�<�';�$��Z"&M`��B{DL�6I��l�^�fx �O�OzQ&��9H�r�����9:Q$�J'�OgS$�y�K���j�9<Q'�5�}��_|�}��yv�
m��N�^n�}z��<-����%�e͒Ot�N^6I���@ Rߌ���>��pހ�ϗI&��$��ڪ{�'ǚ���d�u�'��}C��O 1�n�����r�{0��@�����B9v���ـ���zM�S$�x��KY�h�ӥ~�z��}͒nx�M��̙R[s&&2��"!gL��Q
�wi�!?��"Zf�=��&���7<D�����~�>�5z��(��	;��;z�@�?{Z����	�$��Q$�J48D	����$�sd��<$�[(&h������J$ﵲM}�d��/��n���[�\�'�"N�
�:��� �������mm5�a`ۍ`�-�s����[}���(Π1�o�w����>���q��͒vrO#a�ҢI�J�$�҉=|�&���&M��a%���4I=҉9x��	��l���]��'�"e���߭�s��M��#� A�B t:�en�'�R�ԷD����=�@>��>���ݡ��b��R0�4j�����K�.~�])J���j�>�(�s%z��h��l���p�岂f�d��_ @���kd����7?�&Mڜ�r�sD�ߔ��Oyow� }���>��c�TO���I�҉'�Q>���d����H�i�����~ z>vh���l�_(�������(9�ˋ�VЭ��xه��y��Prǒ�Cd��C�[��Чj3d�[�62g�]��'.�kf���-;rF1+k��8g��)��ѝvl��XԠ��MvcWb�$�m�2�nB��ߤ��&��M�	��&�r҆�elgCl[�W�.�v�&���=҉9X�&��EI9<Q&�s�!=�&[�$��6I�y�M�I;��&���S5���|�~���6/��(x��2l&����Nd�N޶O	��d�{�p�[fBf�'�Q'�}�$����~�����gV�B�an�on��ێ�d�uڃ���$ﵲM{͒nt��D���I���Ia��o��$@�S�OzQ'���@ hH��H���iQ'g�'2Q����d��l�]��%/2L�?Dt��Q'}��k�'�@��(�~?��"e��O���&��z�����p��{����ļ�j@��M	XF6f�l�t��lV[�Nw6I��D��<��͒{<��U�����r��ˀ�����}���S�I���f�'�Q'/2#�#�4Ff��d�O�$�)����\�>?oԁ��T����������;mD��l�ыK$���O_6I�9�NT�q�	(if�LE!��A�n��ʮ���x�۠;����o_RM�6I��%����i�$��] C	g�$�sd��+��F�>��D�sd��~l�^�g�� L��(�{҉.��F��m�tO�"D�u2NN�d��K]���<�"7��'��zm�r~(��$�Nި{����y�z>Pf�4-恨�)ZFm�kn����䓜��������I��D��l�_|�  
�rx�Of��A�E�{��D&�[$��D��+�D��i$��J�>���7>(�� p��e~�͒znO�H�4�TMF���(�k҉=|�&��$��%ɕ�D��N�O�Uo��M�I�@ |#/�+薃�Z�)4��]t�1�&�+&���P��g����F�㝔�Le������v�ٚ/8��.m���<V!WWC��9�qƢ�T�kpj�,�30���ܥ�٣��l�R`B[�x�/]u���η��7��c*B]�͆i�%���ruf����-�����6I�y�I�2~�$���M���I����~�=���#@���?�(^53�6�	�$���I̔~����7ܠ~�� �\��{%�}p~�@��?��}7������%F�o@y��W��&�J$��D��@����%�(9e��x0���>fq�7:U�3TT��IA��}��&��N����l�oO#a��TI��D0`D!���b"��IݔI��l�_|�&�	.M�N�=��;�ڟ�������9��9�P��L�~�d��(��=�D��'���r�o��Ob��'�p~�@����f�f�7qi8;I�i�����~��;�p��I�I9��=\�"���l���|	-1)��$��53���ou�Mϊ���I'�"��ؕ����מ)�_��h%$�H���9W�x,9w� ��"M,�F�S��Lp`��Q�LVG0-#y���i\��m��wn74M��A.[qj�gyG-�6�m�ŴŚ�ZAu�F�w*{F9ǭ%���$���AW�h�8"m N��0
�����&��N�T�I�����>��ˬ�$�v�I0��IA��� D��2NN�I=��=|�$׎�#��m*$��D��K��P:�� ���o�M�*��V�2vҙ�au��99���z̓���\�P:���O�� ���Q2&�>�Ҝ��9�O�~l�^�d��(�w%|"	�W��SH��n�9��''�� H���9�͒~�3?ۄ��'W�O�(�]͓b���I�x�����h�wez"��?}��������-ţ����KWۓy�@��|��;:5���(y����F��� Q��IA�J�7��''�N�Mn��$ޞ*F�	�����Nd���6|�}�����9:�$��������k�$��Q%���S�Q
S�$���O�?�$��(�~�D��6����ܩq��{W:���
ڄtD�J�Z1p�u+� Z'Y�)��;^���1zv�{ �b(�����ݠ)��[	�$�Ŝ�ۛ�
��:��je��n܃��2fq���Y�=q3�5v�홚{�:� u�����Մ��<$��;fݍ��N�[8f�"��x�w|0��^��{޶�<���_M�-��u�[��s0������IݔI���5��;���7���߾�y�����pyg��hݷ@~����=��:�� �����[�X�a[�<>���[�fÞӞ�a�Mc�e۠<�����}P:����RaU���+RI���C�OX��L	��[$�y�I�J$���&}D)Nl��͒k�l��?l�I�J$�'�RR�D���>�D��(�l�8%�S$�)��Ŧ�7D�OI9��5��&�T����ۦ�
m��9cc��3�im�;"��2l�{�k1�Mw<�Z%OI�+����$�sd���$��D��+�C�	Gdw�%)*$���NO�0b [fL���f��s�*��+Dɿ[p���f|�~��������˷@y~0}�[��� 	��d�͒X3��)3D��(��"��M�6I��3u|U���*�ݮ}91EU��]m��g�6N�&�����(y⁓��舁�l�;(��������-�$��7�&IݔH�L>�:�)���MǷTfH�_rܢ��p$�̧46'�Ӟyf{�R#�0��@})�84������8@ \_�Q���}�|οo����0�l���3"�ls.h8�M�}�Ns��0r���Q���uC�Ҥd0�J7ھ
�(�i�ϖgϗ� ��~T�	U�A��;�b�F��j��>��"G�kϟ,ߞ[�,� ��u�jz_�t˖�_r�g�nL=�6#�F&B�倡��v��\l���K��9�5�su��xK��)���yK�=R=5<�`R�im���1�X��f�DD[�ۣ9�}�l`��4a�3����0f,lp7d6�4q�������ma�,�zP�E�ˍn�)��5$�B�nL����{����Zl&�3�fL>�ꋻ;���2�����>�Q�����oϞ_�U+���@�h���A�(��Ɋ�����z= ���{o���Q�|�n��'r�&ҏ���u���s���s.JdG��t�c�u�V6�Ke@�7� ��NI�fm�e<�釘��_�� �����|�6�QS��ߓW
 B��ƣ��nO�V��<��ķC;�{<��aiL�e��lt=��ޘ}�xD]�T{�=����E�n�<���Cb'A����.e�b����٬X�h].����J�S�t��A�(����H� ��B�WA�Qޘ]��ZGyȐ�m(���  ��6�� L,#%��@P�������yo��I�%y�)��0��rD��+/Ͱ��1|����g�(���8M2�2�&MHb�#u
�(�6-mR�e�t/uE��7&+u�Jga��M�n���zb��}�.��Jnd'Q�1Y�=���Q��@�������A`��� i�������=�A�T/�G@"3��1]�m��nQ�����l�"C�۶hnu
�3ۘ�D6�Ha6�f�Ɋ�A��d���' �u��>���_�(��] �k��l=�)�o� �� ��Gzb���N"˖�_r���nH�M�!�iL�6�	�������Q�� G�hm1 `<��H,$iǘ��8�4u�-�MdLE�����K6BYia+R�P��6���A��b�4��I���,�����&͉Ϧ�m�K	#���/,['G�{]6��V*�U��uY���n4А�cj��-酺Y�Lkb�܏�p�.In�v�b����;&39���Y�!@�;m�Q��%�k��ꆪ�r�4��9���4���Ӭ�Ho ��l�i-0�2��[R	1�KJ�e����Ub���LW

%.�v�m^��댚��v%qF%��!sHS=b��0Ⲇ1��`�1�P�ʝ�-H��$�+����)�x_+��z�OZ#��f觌�N�X��#��wk��;ր���5�&λKʯ^�R:u0ց�V��� 5��^c�c�)�\@��n`-�W�g(Ư/4�:VH���n(�	k�F���;�[yBuu1�JS�%b��coGim��@)��*�	^;N����<���i䫎�{v�v)uoh҂��:���k;We[�V4���1�*ŷ	���1"�N�P��#Z�!�H�+�E�kh!�كhۥ�"쭤e���e�&��v^�k�]��ؐ���5�`aW�	v���C�8s�UF�U�e �x6�Ū��	X���Se�˱^�-U�P�B�UR���@�/.�%��Q��U�.Z����lH��"t<� �`p���W��� 2s��۫���%�&�2��)5�1Q�f�\���Ĺ��.�i�G��5f�Cd�������$s�'6��T�Ii�j��`��Ӟ'3�h|-H�5��6������W\����3u�p��?NNM�N�GZ�Pf�7y�3Z��R*�k7!����*=@7L�'��Le��t_rfs�-�.c��;���r~�� .�H�H!���QY�d�ި~#p�!��A� �9ܢ�1݈x��nd���NA��;f31����mJ�Z%&�Q?�5�Lc�E��f]�*[�
���EHo�i�p�9�߿ �?ߔnLS:4)˙3浭����(}��^ޠ���-��~}��?ZJg���M�n�̑�����v{�%'$'Q�1��=�8 �!vg8��-"�;܇���Fw(��ۮ���G����)ځ���ܚ�)�$L&ĳ2 ��B��⽪+'� !�@C�Fqx�!��n>�VLn�o_���L� ��=���xM�F�,�ۏ{Px-~i��r���}�����	�%,�n���/wT?LWv�t}�74a7t#5�`R�Q�6�.N�d��%{����Y1[�=�q��te2Bu��_��vs��B��a%�[E�f���w(�L6vGa �*��3ڢ�~/���B1 h�=�)��G��_�d0�m��E�b��}|�����m�i����7jSL��;iL�0�[��Xҗu��{�y�b�����Z��/��9��_�"#�{�b�����2E3��,JYr��s��QY1[�mZS���AKq��+&�WgT{�=��)��͘��޸��
 ��'9��$��75�k�۔�Z���%�.��X���#�+AS0K�-ֹ�B7m��-�k�Lr�E��cf����[(�L[q�ٌS8�t�4�����
ф�hV���&���Fb���p�ع�v��V,iNs�眝Ns�C�:�h�e|y�e���:�KlTK��y��h��������͘�=#� ��B����=���1]�� �����fC	��o�(�����+s\Vi"|��LtA͘��޸��_�e��1��>��g�=��+&(Wt�(�]��;�f�{]l�.���%�
�K3*�o���TVO@�Gg!W=<��aKq��EDC�B��ޠ����@��?|	2�)�F�0�_�7u�9���m#�D7܅fy�w!@��N��BR�{�q�" o8�LW�i�R�7��R�V����E[�2g=���es��\�^�n����� ��vs�ç��\șN�6~"��+��gr���&�y~���9N_~�K3������R�+H�`C�
�S`o5��5N�{엒��)�� ���z���+$}��Or�p����> ��g ����ykDփ�XX��lTJ��D$�I��`����͘��6�p /��=�K@�����.�E��$U�>�BR����Q]1[���L�awwg���mߔ�~�}T��R�Ȏ�vl�+̉��3f8�1��+����*�lUK%�˅���͌M]e@�*ۛ�(�z����{/weG����+ҥ�ӡ���(��׫�">p��[!�R�}�(�����ި���	)9)� ��2��_!�C,�x��-��;܇> x�F}��^�>HТ�.���\�]K�ʫ�����gdƱ�-��1�x �3� �J� �p���f���.l�x�(,609�������)	bc���#n#[D]<J��1i-7	�EœE2�]��˚�U�͝��ˎ��Nn{99�����6�a��eґ�n�#�ֻX8�MS��l&�ws���7+g����w��,$���_   E�b������:Ͼ��+Y)�{�+1�Q{�=�Kr�S���x����\@��Gx��R˖�w�E��m����"q�㦜�{�
6�"��mt2&J�%>Qn�@�aKq��+$
�Gw�w����]�B�G;I�ǆ�4�W�Bj��r��_� �?x��-��{��C� N}��:��BeP�r��!GH�@�D��(�#�s$��J3�����!��<"6��\�e�s$J���9�S�ݚ�TS~�g!RITșO#~���>��^�E��ܿC��=ܾ�>�(ϾQ]2 ��3�d6z;�ۿ<�h3��t	�c�z[]E�b�ޞ+��c��}�Lz�� Ea�Cpx�]�$�ŰJ����ik[͏�m�:��u�5���4�,���l��P�G`$yF	0�$=��m��[,6��r^u&M�\hIg��������mm)6ֈ�i �+"
�%�(�v�6���
��C4��Ѐ6�< �iK�S~n�5S���Jj[ 	߾Q�1_|���;�����͘���vr��B�����,`��`{8��0�{=Z����w
e��ZE�f�x��h ���CNH!2�o�E�V�V��7�,"���A�1[�n�Y��I^dL�B�@�����m�����Dvr{hX�k��/�����!��/�
��7��Ԕ#���rne�z ��tM0
�$���,��n~��+�
�A����A�Է��1[�m�� @e������1W�u��B���Y-���r�Q}�T@<a���$�ÙT7ڢ��Q��� 4I''�>�{:�]���j,�.�j���;���8HB�N6�X�c��6l�Y��%{$hm�n6�C;��q�%�r68�ݜqS,=xG��i0��%{v\�7i4Ֆ���D[X��;'l�F匶ې�C!w��Φ����rs�܈_צ��fA%Cl�P�6�v�0��V���*��|���/�
�Q�86H+̉��{d
�B�T^�F/��~����VbAϾC:@��s8fC`�C" �Q~��n��I�S �e7��D�������t�%��]�`��綁��3,(&
)�Jnd'C� U���Hs�l�%{�%d�f`s�oo/K�����=�6����I%�2�n�E瓀́[�(x�2XJR}܇�@��;�G���(ϙ[�� t/<�v.~����w�pl��Y�/Y�f�X�6e�4m����o�r=qVO��̵���1� ]�2����#�y��W l\��2��q��2�&F�"	l̞�g{���|$��d'C���@^y�C���|�a��Y-7&3��q��uHu�bE��e9B��J�0��WP��]	�>���H�MI%�2�wj��!� �A�����s%��(���" >�������v��:�r��W�� ��(��+���2��c�|�e���*"����6P���z /��kS�Q�v-����f�8b�t{��f��0���6�<
WE�-���JH2SS �i�Df�6b�>�>��=�?|	)������7mE��� /��d)JLo�!u1_|��o�}9$�ʡＢ��i�:"b&��X��\�iJQ��a���� #��D���E����^ã����('Z�kv��Y�#nP����uȒ�p�1�-��u2�q'���d��]4�7�˂��@*Ǯ�N8M�!���7l1dMZ^��AH�-ܷkkn^O^�����Dx�^�͎	ƷiE,1�/�1�3L�-���C����h�������r����ڐ)�j2NCe��Q~���=������
*������=��T�]�wZ��;����	�ܐ*��Q��t�HO��x�p,�m�m�d�qs�s�t�`:�a�b�m��/-E�!� 7�vrI,9�Cw��+�4^�����tvw�*�uj3u���7܇u��8:J3�C��vHx���+E��m�lw!�j/�Oz�t�y�ɋ�ᄼ%���G��5�Ьtť�V�h<S=O}����F+u
'u"SM8��0ъ�Cv� ��;����	�ӆ*�}�Ìj��� ]���^���W9	Y&[rc;������0��ՒIa̪����i���؛+R3)JE��e�Rڐ%�j �c�D=���m��I(��0ي�CkTz������� 	��C��_r� �	|�ئ���eb���6�
gӢA�l�CsT_��wM�0WA@(Uw�l�N��E^)n3u��P�����	���$�dc�`�9�P�v�N�y2�$�̄�o�
�CkT�/u���
d���=��_�_rl�cgVI%�2�nj��!��V�����I����܇W(��%�!�t4��^!�v���yH4�4�;HU�d��VJ@��;�� A]��,FJ	A+�������(�)�4�D��)��e$h%Xʱ"��LF��!F��!:7�s����9k5�l��PƯRB�B�͖����*$-`ĥ&K�Q+���!5�
M���5��,���shk��!L(�TNƢ=ՔGĢ����%wM��඀ݯk[7c�mC�l;K���g��1n\m>����w���vw��`l;u���v­l;���{t��a:1����D�ڢV���[].^��2���oٶ��H쐶���q�l��S���k�$&�YnV�[M�ht���v�n��lK�B�֎��arӅ!\\l^�H��;Lf�^���s�ġ4��cg�����+[b���X�v�G�e��q�l��AD����'McF��q��B<�v�Ө4���8�i,���`ڱ�����͚���A���e2d�^ѸNE:��6��P�%͸��WmU���f��]��![2l��+&v�J��QP��rQV"p@'F�E�s�*���xמ�v6�`ĂS�^��޺VU�@�#����W8L�K��2n��a���4�#�;6��۫��c��N��m�Ȑl�)z��i�I\�E�H%A��K�v^v�1�	F���h� ���
�;rq�΅�x�d�	��K�d�s�"�O�"s�<P\�;I!蜩@�|�<�+m�+.]��Z9���WE��,�u8�,����c0�v�P�4v�	2���umKog�}A���)jX�hMmL(N@��mU)OG`�:�,o��$�9?_{������6�si-�7fd�Q��X4��$r�Ҏع��&^�����q��$�'/&��9=-�w�O���t�#j�+�\�g��UV�<V�t[Fv�k	�s��z�g8�ͶCf�h�RrrHNu'�O�:w��ˊ�����N�<5sY��[d\�X���\\���t��/����񌾙� v)��>Q~�l�n����ܦA�Է�C���6�E՝�Im�	��@��!��>@���3&{)��,�B�^�r�������]���7S"u�:GMe��K��$���@mߧ�}���,�t�mא�$ʬ.���{k�hp��r\�����!N��C� U�|��Pz,/ͷ�i����eb��C��]l�����(�yEl�n��u���d��nmÊ\6��:�0�L5J(O��d�MKq�|��b�����Q���[fBu�x�ި����r�{��i1��/1� @(C��5_7nj��eOy$�eU�zw8�j��> ��(�#�K�a)J3�CɊ�Cw;���R��`�IpĠ/����l�ko3�$1�RB�P�����^!�j/u
�h�m?C��=ܿ>�(ϾQ�?��$]t���l�C��/�_��_rR{��2�M8��T뽷[0
TP��=��:��HL�2�옫�7mE���3%�,�n�,#]�A��Il4Ԓ��Y-'3��娽�4ц���&L2��w�_�Hs����u��&��}�2\�	JQ��0ъ�Cv�z�N�	/BM�ӆ*��C� D s���m=��1�C2�_rh�����^	��iAj�+.�`g�<f��kd�y��J*47�k,��P�lbu�����>��''���,�]l�T�l��h�(�b��vϮ͂��vz��z'�f�,���줅\q�����$Τt�\;�$��v��
��CVi@U��h<S?������0�F+u
�;;$L&�f�q���7m|F^�Am����x�u���.��d0�rc7P�����0�ٝ�Ia̪�Po<ƚ1[�p�9�NT�a�IA��u� Q�.&mm�.Hl��R�{�4b��1��U��B��e�h���a�� ,3�!���B�Z?&ߡ6�{��Q}�i�
�gB!���(�y4b�P����A��i�n���V���عݔd�,J{c�9�̛��|�5��a;��[fCv4ኼCv�^�fw2i�1��^Z��CMll��$��W��������;6�H�䜍�(��IrĤ�f�l�n���*��3&W���i� ��6�E�U72���-Ig��=u0��CC�3sd�R	��	�n�&�7�����6�x΄NCe������nLV�� �I��$�aKq��2�+��QugV�6����w�,�~ٰ�+�P m_�g�I� �a�\ǽ�]��Q[1�K*Z�f7x���P{]n� �!6%ɒ�$��T7ڢ��+g���QZGx��I(�����ިw홙2��Q�1Y�m��A�~M��I9�w!��/�
 �
�΄NCe:�Q~�ي�C��Б.T��S)�����Ec 7��ۥ1]��rʶW���h�d�n�m�'�C3��.�Ӯ8��(��[Iۀ w㔹�=�u�jM�=���ю9�b:����Ƙ+�#�t䮼�d�w{�N�w$(/Y3p8M�Ֆ�<5�z��t�I�4��.6+�>�U���D@�c��fa��Il��Ft�f!��/u�;�4����.� �r�����$��C�� |~q���ܡ���K�%$�7TVLV�z�r����m#�K��j�Ƭ�I��ҕ32e8-��ي�CoT^�w.����wyO��x�jx�>�UB �ڢ�VO��D�K.[���/�[b �zb��b���e5-���|��1]�wb���[6XN��b�����޿nۣ��B6[m��`�c(�1&qu-�_�Fz�.m�}��E�(ۘlN�$��*����6�+uEx��K�%$�7Te� @K.���@%�ԉ����%d(�WN�6H�R;b��Ф���+Z>q��-�|z[s�ǻz��M�B�ۅ�,��l�kV������cm��rQH5���bt�T�U��~��Ї�1
��n��
�>Ѐ��4�)���mSśp�D�̳Z��ߟ*�J�e:��CkP��Wa*T���q��eb��Cnc� ]\�$�2�)�L�aKN��h�u� ��q"�e�-��r���럈��,\��d��M�w!�1[�mj� �w;+a�N���f.��grS=��m�>�>��2�����8���g0�Pr��Q��oP����}se|��RR,L�Ԥ]l�uٖ�\��{����Ae�I(��2�+u�P��3$ϙS��+��մ9�ڏ�|�]��j9�r]r�,���{j<�-_���ڏ��[ײ��ʪɕ�����|�^w����^�j:5S���]��`/;�Q��]��]�]�`YJ�>}���eR���=�\v��n�VBăY�d˪��\vw㤍�s\��]��Cv�!�'r��:�Ê��:�z-�g�9ct8�:�2A[vsv�i#=\p$�o5�#�OD5,E�AFU�{y$�$�s����,ˢ��Ea�X�0n�m�$�r�8A6��t�Y� Gժ�H��}�n��$�a��y�7\�]�����.a<��I,ʻҏy��<�}R#�(~�`��=�&L*��C��<���|���mG�{`��;URyyD��(��A�(ߞ[:�}� GVNKL�@��d�$�'����'Qj�Ș�FGj�/(���{j<�,}톐����f�s�Tf3J=�lv�Q�=@4	����׾Z��T�ە%�]��n�u�ڏu���]�r^ay����
C����~k���@����J6�#7T@��@D^�N{���u�A����Q��ڑs�3�����Yt�g�J��@e]�G�=�]��Q�t�����u�;�L�U��/;��*�9@���Q�^ڞ1\�EWk(�y�{@��,_�!$��h��l^�j9��u�̲��C�'��j>o�߾ڏ��]vk��U��ҏy�ߞZ�n@���#��0����4�)( &%�=V�hI�y]�=޻Z�tU�]��ﶣ��.���{��.���w&I���{��7疣���]��Ԁ�W�I,�3&�ﶣ�r��#�}�y@���{�̫�x|��y�mG��%�T1�����!��d®��y�ڏ7A[� F�"*�|�4T�KfA8BWZ�q��u�z���w{ܮ���VQ.�j=�뜵�v���u��uʼ�e�/;�Q�7`��mG��]vk�_%цfiG���w�/�D}���mGF�{�*�/3yﶣ�PDV��";���3̲[a:��(>��ߞZ����wﶣԊb.
)��`���[=ｾ������`K�m�`�ɑ�ZD�j�R�q�K��AC��Q��m5�<��a�m��Q�	-b-���N�y�-��� ��7;)�������!�~ye�2�1(qe͊"�Vf��ٙ���N\���
��{��v��u����\��I���IA��`DW� i�� "3�81S��.�N�If]�ҏ��`�疣�P.��S"��r&uv���y��{j=��7�����]�{��9j=��}�뻒�yd��^w���n�w�ڏu@���s.S=p�nI�/�ְn����i$��-	L�6� F��(�REn��RwIE��m���D @�7H7ﶃﻱ:Ey�{W~�2��z���e2�L�S)��}�)��e2�L�S)��e2�L�S)��e2�L�S=�}y�)��e2�L�S)��egl��e2�L�S)��e2�����L�S)��e2�L�S)��e2�L�S)��e2�����L�S)��e2�L�S)��e2�L�S)��e2���y��W^<���L�S)��e2�L�S)��e2�L�S)��e2�L�����S)��e2�L�S)��e2�L�S)��e2�L�|��猦S)��e2�L�S)��e2�L�S)��e2�L���猦S)��e2�L�S)��e2�L�P�iɔ�e2�L��޲�L�S)��e2�L�S)��e2�L�S)��e3ߵ�ϧ�����l�S)��e2�L�S)��e2�L�S)��e2�L�����S)��e2�L�S)��e2�L�S)��e2�L�|����S)��e2�L�S)��e2�L�S)��e2�L�~{�YL�S)��e2�L�S)��e2�L�S)��e2�����L�S)��e2�L�S)��e2�L�P�	 �	 �	�E}���o*��k���6\�71�.&mm	���Au���	��' N)��e2�L�S)��e2�L�S)��e3����L�S)��e2�L�S)��e2�L�S)��e2���e2�L�S)��e2�L�S)��e2�L�S)�Ăo���$A$ �A}��"�����YD����(P=�H$��S)��e2�L�S)��e2�����L�S)��e2�L�S)��e2�L�S)��e2�����L�S)��e2�L�S)��e2�L�S)��e2�����L�S)��e2�L�S)��e2�L�S)��$�H&��ʯ.�ɗ�A$A$e2�L�S)��e2�L�S)��e2�L�}~~y�)��e2�L�S)��e2�L�S)��e2�L�S>��y�)��e2�L�S)��eg��<~o��=̦S)��e2L�S)���<��e2�&S)��e2�L�S$�e2�L�S)��g��u��e2�L�S)��2�L�S)��e2�&S)��g��.}s���<��=�e2�L�I��e2�L�S)��2�L�S)��e2������S)��e2�L�S$�e2�L�S)��d�L�S)�>����e2�&S)��e2�L�S$�e2�L�S)��g�κ�e2�L�S)��d�L�S)��e2�阜�&S)��g���<e2�L�I��e2�L�S)��2�L�S)��e2�����>��w�x��e2�L�S)��d�L�S)��e2�L�)��e3����L�S)�e2�L�S)��e2L�S)��ec��&S)�]u��e2�L�S)��2�L�S)��e2�&S)��g���<e2�L�B	 �	!>o���ϗr��aY�Z�f���e�f�%0R��e�b]D�H��mj"�T@����J6�#7T@��@D^�{��'����.��G���Z�w@��l^C��Ʌ]݂�n�u��&��P ��AНHl}�������]�{�뜵֠"/uDf�oSH��R�����fz�:��s僄� �K=2����\�]���=���k���ᙙ�y��9�ڏ��]{���K�^e�y���mG��]w��6�w{+Ye��u#} De����{j;�WN�32`/|��\�]w����.LU�4��R��"�w�Z��y��X�C��y���ip�:��$wl��n0�j�b���]u,L��/��X��e�F",`�c��ݕ��Y�5*�Z��j�O]�y��e��K���3��ru�x�)UAV���V��4�2�mk�F�������j�a�c�v�uc���p�hHH����zSӝH�\�xktM�iED4�.�LF`٦�%�Bƛ`ݪ���&H)�k�h[x� �v���\��ݼ�q ���4�!$���t�`/E�e�I�� p��Ks̼Q��Hް�c|yo����e6�n6�UK��6]���ۨM#����%v�̫,��*�U�.37]ozF������7qZ�b��t���Q�[�|�fTt��6m�*'��WlyCˤ�ۅ܂b�4�[e[�l�lݱ�v�v�;n3r�@7V�t����)�iIn���m�Ѷk0�`.D���j-0�P�_!^y�ĂBcwh�-[���E`U:��n��m��ɐ��w0q����%�垛V1�pص�P#�٥�[W.jȣm�N�.�j���k���Ŕ�}���#�jwCx��*rM+Q�pU�;���&A�G��HkiZ����&�&�v�E����`�5�<컗�6�J6���B0�����Ӊ&y�m��GS��^UP�65���Z�u���!�Re߯�4�*>��@��AsJ!ĥ v"��Ťp�$�=��;��f�Ŧ#�氛b��ĝ�å�������[����g�.�����>
ض��g�=�ɰg(r&�9���x�9wX�WQ
�����:j��( �!�X���H@�ffL�I��埭�֝m��.y=�W�ӱm�fल��R:rļ��а��-�	fYwꏽ��u�-G�p����w��0���]���ɸ���{�ڟDAb����YD��(�;y�Z����u�ڎwr���y�V^@_{��]� F� D*;%N"n�njA��{j>�@_w퇱S[��n�^V
�,��mb1h��c�v$�n+\�l�s���s����9�ﶣ�v�w��;�̺�f�{<�mT]a�a�N^�G�v�u�-OR su^�\��32�/���w�X.���{7s'������(���]s�Q��D���=�]��	�
��߾ڏ&�.ި�Z��ۼ)ks(��2	-J(��><�ܦ�â7�إ2v"�]�{<���-G���M���a+���@��~Q2�]� F��������\3���}���{j�T�@"��,Ԉ� �-p�ϔ@�Op*q6�M�}� F���mG���]�_\ˬfiG�ȃ�m)�w���mG�n��f]�/&���r8인���u�t�0Hm��Ph̰�r@��j�u���P�f�.d�t�^a����yj=����l^C��Ʌ]݂ｵM�^ﶣ�v�s͝��ɔK�Ї�C���<�u��^�v���%�/��Y32��-G����mG�pIק�)W�/	n�f�pM���Ѻ�o*��k���99�~�^yj=����mGZ�ޒ^^]��ｰ>
P�r��mu�׵��̺p]>1���_(��.�xb3,6ܘ�rX��P�f>�
	���QY�4��{�'�}$濾�����ֹL�d�P�ҡQΦbCIf:�;(�v�g��D��R��#G����e��� ����$6�3Y��
�<䫶mf�����1_����f���\,R��3*!�)�����u�(�v;HԼ���&a�6	 �s(��,�)%��a�_�mj��"|��Rt4���!��+�l]���{DKL���X���6aV��)NCM����!��� @�=��ܞ�Bi��q}�a�z�֨��x�a4�a2D��)�L�+4`�\�lI�S-�SN���.��Q[�]L�����rc}��D 0 ?f���8ن�68l7CsTVyt~���}�W�\�)%��a�z�֨~��<�h�>1��y��Q]�ud�̔
nN1��a������]���Rr�/�N��i���2�Ew|�0�J����t;9E{�i�z�T��Qi�w�ｳ�p֒��=�1L7�{gv(���^��.���6�En�u3���mɍ��u�+u6b���vK@�F�`r�$5�u���Ҁ��S,0Pa���QY�4ٍ�Q^#p��I(��0ٍ�Cv�?X:W�N��1��nڊ�B��_$�DKL�� ��!�b���(D؈�Xb��J��Ô�wyE{�i�z�{PX�i��$����<`jr]�ٶm�8{-6��4�M���0э�Cv�U�̭���]8b�ݵ��d�%�ۓ��e���4ч�6����CM����w�.X�)E�!��m���Nr}�/�&1o���n��J[-cl��S"��Q�k�ֈ�J�\$�4,�\$z�<e�X�'8�$��.Pۨ���/]ѷ
G+�J2��n��-��2�-�5�"���g[6��`-i(�5������7޻�-�s��n�������u�3�$�,��A$�|t�^!�־"����W�=�%�c��P���Fi�I��:�P��4э�B�N�Rm&��"��<l�v!���:et4��q����{�K�rv��`�K��@�:Q���:�n1˞7����2[-�1��fZ��<Y��X�PA���+�<��1{��zGx�R�_rh�v!�j+��4�	'CN��7mC�B��_%��1��fZ�܆�0�k���X��g*��e�c6��� �(m��������枚1��UI�*CM�ۊ�C��7mC�ٕ�Ӗ��^b0`^��P+��Н���.K�@���R��eC��=Bq-M!ť ��F�R0xBI��Mabh��-���F!�v(x�,�4Swr���%�[$~�o�����-m������< F Ia�4@5���bq)�M*�j��I� �7�<�]ݛܯS26䏢w!^�܆�O�Ul�Pa���P��i������r�R���"J��5RgٺɹӔ��76r��J+u8cw8 ���i�N�1��=�up��L����4����������;)$rN��~���6�W!DP"I����T4� +~��5���%̻˗�+��w{�8e���R�a2J���e��m�[)�_p7eL�9`��� ��+��<<&Ke�����{�+�����J6�{�y�wW��9be%��d���=����̄��� fbuC�S}�'��|r��w�]�kU���`������]�����.S�[�/$��#2nO_6��8�]��e9B:��pC���bz�[���\�1y�Z�!�B��h�Dg՞�i둷��>��ꐡ�b嶀�V�d�NI�d�����;MU*h��=k��	s�\�	�"T�e�s%L�⪤MS�����!� *�u)G!��^��!�n�RthE��M�n��n�uC�ٕ�ۖ��Le�uEn�TgF	��mɍ���V�pǬ��4�̄�-I�$L�B��p�e2.6��Tm�0�N��y�4፽Q^#pe�)(�����Wgx��}�Y�r���h/&d$�:c/{�+u�J���R&���b��CNT4jR�CMн��!�m�DU��M�d�rY$(3-��b�<���*���嬹�&Ԧ�;�Æ:�����el6��i�x��Q[��jL��2[-�1��b<�"+�� $H(�僫�q|a���J6�~��CN���'pXr���C�� ���r��÷�m��B��]���2�T؋�LB�4�g%�g�����w�֨���*g�UH�Tc����܆�0�hԒ7CsTW���1��UIѨ�y�w�ｳ�q��f�dUCাߝ���~���||c/�����׍zP]���k�l��)�F&�lV	te��ӟ{�����_}�1�Ul��Pa���QY�4ٍ�\���Aa��grl� ��:�C�(�3!��oN��y�Q]�=�Q�ު�-Q��C+>�4لl� {��ڶ8��y�, 7/p�=;:�����ʻqJ�É.�d�� �ϵ=�ˀ-x�%-��͠I�eer��m�ZD��݌�F喽z5{tg]b�b:�cm�+=�� �׃f�uv����dg\�ߏ�R�6a/	n�k��CX�Ҙv���E�I�����C����*��ЋI�-�n���n�Z��gQmʂ�i�CkTV�Ft`2-�1��2�En���?T��Xa���QY�4ٍ�CnM�Ԫ�z����\WZ9��V��%�I9��&(4���C������Q[���2N��#�z"�O!��������J�T�I���2�Ew!��*5�!��nj����f7q
�'Cs(�����0ٍ�CkT~��h2�M&nm�8=@�ny�p]�Г�2rԤCmʂ�v���W({�]р�l�X�C+V�r�M������^�#߀��Bː/�!&�d}���I(���oP���6BKĄ����2��Q[�|_��I�(��ȶP���fV2��t�dR�RK�4ꐔ�w�eb���6�CF��2n�樯y�oP��t72�����C.@��6�E]��!���i��,�e��JG�G�& �P,����x�ܘ��!��+u6b���=��%�q��uu��Hms����-�ج`�X�O{�s���f��E!�=�����e�ۿ}�Dx��C��=��^$$�>1��mj��A풿O�R�1��eb��CM�U��Ic!��nj���c�@��?� ���� ��5)Sa������'�� ����͡Q4r������u倫���癝�m���Vm���QPXE <�(��E ��1�Ű3b��5�O���/����l?�u̮��Y���OB���r]�������i����~,4c����FQ�?ڜ�~w���������t�661���l���[����/_Ǐ�B�����}�$�(
p������H��@P�އ�?���q�i?��7��~;L��}���ԁ���ӄO���>O��M��AAF�?�D\.�
 ��S�Cg�W��,�1���ѣ�?��†��ڇ$�}g���� w�>W����?3?�������?R ���������'�������W-S�>���/�������zz������(!�~�W��/�Bc������y�H?��A� QA������������4�H�ꢇ�����,�J0���e/�3�DPB�Bݐ&ܹ���-2�!A��W�(�@PC������������� c��O��_���Ϩ�g�O�)��mQ?����_��%���p�@PC�����>����ϸ���<?�����P�;O�F��G����S������{����h37��(
}��/�>����|��~a��Oפ'5��:���A���6��g�)���?��y�8Qg��Pk;7K�k�1>��?R��� >u��.�p�!��0