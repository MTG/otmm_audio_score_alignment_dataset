BZh91AY&SYy�x��_�px����0����a{�      �W�*�z�	 P  ��*   J'�P!  �   �@.|    e@�� P��I(�IHJ(�(% T��UP�A@@�%PH )"!@( P 
�    � ($	 P
��� S�*Y�l�6v������
=�x�m�O6{g��ڋ�
N�:���� �Լ��7}p����;�.3��V�j��]Z�s4)W�P4sT)��==8���Z�j���iJ �< B�]4A"�l.���y��z�ξ��͕w��ױ���
4���r�[[��z�k�;�{�唫�OG��d��y��> /�ǺW���W�� ԦO�ޛ�u��mGɮ[�} /g�_W6��͗����j��ZW���@ �*��)E�����]�ﲮ-W[�N�n��\�}����+�����]<�u���U}�K�Jͽk����   �G}���x�K��|�eҽnm}z�}�z��yy]���wS��| {�[�]+se��ŕ�}��z��� (J� �`��)VO}������}�ź���z鯼 m��/q���sj�n^m��yt����=޶�6���^Y<  Yso[{��wMk� ^*�z���y�U�'S͸�]��� n���g�R�Ԫͻl���W��< D�R ��c` {ԫ�_[my�_.^g�Z�ܵ�� ꞹ���v�m�ͺַ��R��!@<�+���վ ������yk�j�(��+�}j]�uﻯ�*���uw��w�R��i}���W��/�sj�| @          z���J�J4  4    ���6U*JF` 10L�4"x�T�H� # �dщ�  ��U*)䚓P h414ш ��E<ԥJ�     0B��I hb5��C��d'���S�	�����?����?�o}�u���܂�������DEOހ��W
P��*
��,�T]G�%?�B�
����~m ?� 	@�*�T�*��A�����)@o��B����r�'p"=H��(�)� �@�� �҇ҁ��"?H��}?B�҈�(J�� }
B#�(B)��J#�
�B�}
"?J � 	� }
?H�҂�@��
��
?B҈�
�+��} �?BJ�H@��'����m��D��N�N��EC�O��O�~�>��>��AO�G��� �>��G�S�>�O�C�C�~��C��O�O�]ț�7&��>�@�@��}��L��>���@�!�*}R��?J}	���½����@������~��W�W�S�p�7��O����>�>��>��{��O�~�rЧ���)�'��пB?J� P�K�+�B} �B�Bw@�>��<�5*}@?H��5&�O�~�>�MA�'��?C�����BQ����+����>���C�S�{��S�O�!~�� ܟJ}}B�'�?H�H�НK��
߰�S���)�S���)���O�>��@�Oa~��GR�M!�H�@}
Џ�P�H���?@?BHrS�O�>��G�O�N��O���9/ПJ����@��5 r9���G�C����_�O�>�������>�_��_�~�~���C��~����~�������T���>��Q���O�����C�O�>�>��_�>�~��S��O���~�~��G���>��S���~��W���@��]�����B}B�ҟK��?K�}��?J}��'ң����>�>�~����C!~��>�>�>�~�S������~��<��:�O����,��q~Si۠� �h���yka�4����٣i�ެA���Nl�[�C�owן�^~��u�Ϲ�s��>�H�ȓ�iT��IT����=)ɶK�Q�Ƞ�h4;�sa����K�|6���G��a�X�0�vZo�}�Z�v�%�!��цb	BP��d��{�{�g���]wᳫ�I���Y�3��&���h'x�%����&i1U��kT�YHfX�ó��x�c��-z*Oa���4���=[�i8%Z��i�B�A�HQ�v���t��C�kQ�;r�{5���"��\��p���:+Z�zx[����o|׼�F��F�tu���Kmn��R����8�o������lI�8H�3͙T��Ǒ��x��Lw�� 7��v�%��M('�D֕!����k�՚0u/�G`e���-�B�A5/���8�5�~EZ���y��"��%&&bq2!(J�������u���J6�R�$N����r�5�a��N��^w�4d�5�(��i�"c�����Sȉ�"���v���ϡ��0��ttj0��k2����(+5�|L�\C'B�iu�2{�0���# �ӥ+9K���:���9*�'(,#(����^w�:7׭��^nۡ��8������z�N8����q�(_i���%h4�ԝ{;�I��m~���iE	BS�9���[޻μ�;-��:��u�c�tfN.�������n4e�oW:zczp;�9�]�5�7 ǷXh��6Xh=�{p�a��m�{pѥ@7lJ���Č#F�@$��fb	F�3NX �I�Y:Ƨ
���� �<�hl�[ks��{���^I�d%	BX�A�@a:\�4���94�4X�BP�LL��D�q%�{�-A���X悵�X�	��]��U�������!wv���v�sH�{�DN��UQ&R��UQ��v��fÃ�m.�6:���ѽ�4j7:I��A�5�p֡��tFf�4n�(��(7�eNN��FBR���]!A�rM)���;�4� ���1�;�xUO�r4�.VA��{A���A{��ԟ5�'`¢�O;��Pv��9�lh���kV���Jh�^�����O7�HI�ңR��ERഇ4M*)�y0�F���:-��dD	C�z�Ѳ�{6Z6��%	�`���(��#1���r�����|y��=6��J5C��N�����NXl�utt6� �5&1�㬷�xtkGL��+i�=���;��$ѣ���Ph����S����|��0|���{F����q�A8�`IP��/5������7&<5`i*wAGg ;9dC�Gr�'lBP2���íl�	5h�Lki'VҢ�<y�<���Yߜ3�e��N�h�Ј�`Lda��=<���i�J�����2N'0J���8z�[<��UI�e���(�y�qs��ƳZŎ��n0N���;���9��u	I�e�fNc�y���P�	���2�,��s�9�%�Ɍ���o�;3xT��f�Ed8h�����SQ�O5��z������7	N�G��C(s�ӑ��jq��[�l7	@p�0#!(J��,f��&O�Rq��;��-o�a���:MY���w��M(��~z�k���(��Ǐ�ټL*˛	��0��K�5�k�����}��i���[��bz�"��M]�M6���@�C�cb�f��ɽ[�(�PR#Jb�,�#-I�Ԛ'�sQ��o#�2�2�X�X�<0�]q-h'f5 ��ٵ��yq&�P�����H+I�բ[HM���]*�q*�%&i��섻��Û�=&��AѢtf�1!�M#�޹�۵�4҈彭���O��XAFS9TG\2��
t'y�h��`k���������ʍi���I	X��u�C��]�������Y��c�4��1,��(0�{���[��x��[g�z��q#"�l��Ġ�]Z��ֳI�5&&M�w͞A$cZ]��цFjـpٯj��xtq=r�N���	Xd%	Btf:\��)�JA���ýf��`��C6%�b�4��Z�)��fi���,X�� �C ��d����d�]F����Jl��ia�BX0u&;s�r�F�[�JLL�]j�Bs0t���-.��k��8�FvsY� �"�qu	BVF��2LLY�[C��(45'zf�]Fh2��MK�Z���A	�O�G�`�%� �g��< �K|:����&�X�]�\�F�+��#�21�1���r\���`�JF`d�h�m54�二�-������5�n���.��Z�{M2x���iÛ��S��%9%����MF�Y�k��y��f]_ ��]g]���θ�N���:޻��7�Z�<H)�8����θ���8�WJ6�Ѫޔ�3�75'g&�߅á��$���Ot�&I�Y�5�<�2��~�ֽ\Z���fѨ��Ǩ�����/'y������Զ�����<9�w����:��������A�f�j���}Պ�)�sj5���DݫB�E�b��*�,���*�U��]"�5����sJ�P��QDM��l�ٰ�Z��A�8����{d�&�P;�ݸo}��k����l-����TNA:E��9��^�ѓ^7}�o!���&�\H������P�{�����"�Aj��s}�ٯ#8�3K�0� �r7.ZA�5���	N����J��Q�ӵ����ʹ(�*~�|��w�+w.h�������Be�7	������N�����";:��.�w�XVl�<���)'����=N�����	Cߎf%6A����a�9�ى��δf���dk2e�9.9��d�Fa.Bj�VTs�T�^���\�~�4'�!wv��HU�-���Ån6ͮZ
�������Vٳ5�l+ ��C�٭O�r{ӣ2p�2����Es1ΰ7��k���塐M���kvhA��uFA"��5�J���c�Z��H�آ�zQH�z�;lU�کM(�B��uP���QS\ڼ[[�|bک�Ҩ&)��5�W �+ ��%	BP�%)A��vx��Ñ���r1u�6�Z��a���%)BP�%	BP�%	BR�%	BP�%	BP�2����P2��(J��)'�s]�k}��|��c��J��(J��0J���8.��# �Jz\���0J��� 7	BP��`�c��%	I�6���Y���p3DjŰtX�L���쌂���%36Fp�u�Ӯ!�JR��%��� �C3��)�� �f78��%��	G�i�h�Q��~��:����j��_���q~J�m]j/?uu~�\]�(��3���ԙf!��G��CS$��%M1'��BZqy�u4�Bu�()|� �L 2LL�5bj�Doi��XB	N$d�-@{����U�/Z�}nћ��ۼ|gZ�\���2�2p����f�7q�7h$����i�a�5��a�����u	�`�%y�`	BP���Ն�0���=�����P�dh �J�!(J�N���I�J����$޵�;}<��f4���${�RLQ�BQKS�NԱPI���ֵ��睝]`�%	F!�&l9&K�;�0p2������%	I��]�$��ԙ�Ș㖣�7ߛԇVu�6w�
B;�4���o:p4�:3��!)�[������6r�5��	F&�uÇA��ow�u:6��t��I�\�;kX9�^!�Z�u=.G	,��O3 і!�bf�����3DZ��*��ph���z�޳������h�GO-!��+�8E֡9j ٩��	�f����0�t���ѬSq�#F�q�s�i���%?k{w��M��o����?-MJ��~W��\5Pnﻼ�'Gf�?��Tvj�������s���k�xÙӼ�V�a��d��	X�c����&�s�i}(���2�UVF�0�h���P�f�:�m�gM���hߺMΗ$;�0�&2L�jέk4�-�Idc ē�ߵ�$�!��xqn�\��˞:�Q�5b	`vA�i�!(Jl<7 �Nj6�+X�E�A��;�a�J�m�Q�%a���Î�N�g�:��'f��\��A�)UU��'4(Թ�]1����sg-WP�d��̼]I�a�����7��f��]�$�;#��9u�9�m�޶�-�koDv��3F�ݢ4֬t:�u:�ntj�b(�On�<.���ap:w	BVQ��9��s�g:5�����,��<3Nh���h�X4d��k��l��9�[3g=��8���u4Ejh�]��n���b:�VsŻR���\��]�8ݔ܆9�k+���왱*PlH�<��{f�g[��Lq�sT=��K;��We�x��� x��sj�r���p�x�;t�f|㳰�`���q���^��.;���݉T}�9]�˷l��Q�l��_߷1^�\�_��r�ڨ8�d � p��� )R�� �@
\ Am�A�������� 8�� #�@
P`8 p�Ȱ� ������� ā��  �� r�   �-� �� ��8�p � (@
Pf@
P`8 p �� ��2 R���� )@A��: d �G � (  n� �[)�         �           @        mۃ   ��  0 m��s @���)�\�2 R���� |�� �p �@
S (R�A�I!�UԪ1�J�V�)-UU@N�j�s�U�J�.b�5�m�m۰K�EYZ�z�vj�s�5�k&8��@ ��#��[@&���m�d�9m-��NK�K���[m���I�m� �   ll ��k�m�m���Mm+ʭ*�lU@P-_���l�6�!��8��5��Z� &��HZ7 
C��j�b�r��`��N
(j�k<GL����m�q�׭	6ۀH�E�ɱ&�I7[�d��#m'�m!� ����i�5^aɑu����&w�I�cm�;b�l;���pF�8t��mUP*�cV�;�3��:�G��l�=bv)��l�c<�ζ����G�W>�J�a3�8�c�����-[EtqZ���
v���T��eLh��VǪ���3�&b���[t�#k�����)YT����Bڒ�==ף��Y��k�㴊M-%�m�M�m�� ���)AL�힂��hҎ�����gvv�(�&��YP��ғ���<��61�Ĭ�=i��ݫs��G�u�n�n^7!�D��ad�7�Kn� |}o�K����Hi  R� 	ֱ���V���6ض�@^���ZlH�kV�r�sm���&�`�M�n�H�<��UIҶ�1�H�Ѯ��m�mm�l� P���l�G����7m[=��	�jj{m��M��/Y�\j�r����pT�+�K#��*��j���-h��ٺ5� -�d��="�3�Z�&��=��4 5�ا]�Nv��a�����Wi瘲�	*i���Yx�/N�[p�V�˳u@@Gm�LT�[Sf6đ5l�`�کZ7Eo`\�uN� nu���6٭h��J�VՌe&܎��mM� �bkt�$k���՚��:w0tk��d��\�X[cm�����jtnN���qŝ{v����d���ˀ7e+I�$;m����O���z:�@!*͍W.���Z%kb��jpH8-�l-�-�����v��[��u[J�i�٥�z�;��25U@�kXI�� ���h HM�	!�Mշ���6H�Z��ִ� �8  PT�mc*�[�`ۮ�U����BuR�\��Hk7�lm�P���vь��.�Wf<
��hg!�gm��G��6�nq�<�k��6��Z�I�mo^/ZOH�}�.��ں�B��W�u�e�cm��c\wcW��7n�m�(�.�R��[V�yz���N�%��4���#m��L�:�R����j�d&UQ�N�L��UU��` -��6�̃��c���~���g�[@6� E�M��z+�����Q% .  �[�ٻ6�[�hm�v�k�����u�M��� ����m�HH�Ac���r�1i�;m/K�B�psn٢�kZ��Ͱ 6ؑ��Z���U*��mp�t��,�Cm$� �`�p���m����װD�7`ݳ�$��YGꯪtI�6�7mS6����%�oRG�$���l�J�@[)�V疪��k6��:CE���H��u˶�#�)��z�6�q�ln�M36�F����lI� �e�h   �|    h��۵l       I#m��ڴ40 H�5�� m�  	iІ�I;IV��   �.���շl�n�  6���m��mn�!$���  p[�4  s�$B�m:7l�A�c Ԧ� ��A�3Q�|m m�6��v�yS�5!5n�y�v]Ut���d�M���V�p ��z\	muUV��M5���*˵N���A� �v�E�9��/n�UGP�%�"]V�rީ8�m�$   ���loP�J�$ !�ڶ�d��i`�H� +c`  -+6����%�M�;^�+vd ���؀n{���>y�p�S�5��-���@���V� �fͶ��� 6�     �  �n�� 	vY0m��[p     �m�    �m�K-��KmݵI�1a��8�`
^Zy
��oK����6m�6�#��۶�j�X)W��P.�]֢� �� [G   �       �� d ��ͩ����BUmH%l�<��Ӕ����5J98�yZ�B�(*���y�H�-T��1-�9&�M��]Ei �&����K+�*�jˇj���6��K�PU;;mFyķIW\k�2DQ!�C\�aQ�mc�S�UJ��.А޹bb��1#��jp m'a�6�e  ���Ar��-E�J�;7��	��E 7R�P��/UN�T&]� [@�j5���` :F��   �6� �[,s�����m�m��*�#sl�U��\�y�[���9W�����@@)���� 8E�F�ۇ8m�`�on��-6i��m�����lr@6��Xm'D���5���H	 -��l6� �g��:�۝��m8�m� fײ�/��O��ds�          Դ&��9����[x�����a�����.��� ��@�
 �
�Z�Am7m��� 6�� �knqa��m� �6�d �i�6���m� e�   � �r4�����۱��V� Td�i��5 �4�6�jBBBBڐ�� smض�Y\H�9l�,��I�l ����6�   6��nHI����ͭ�-Ԑ$ �fL�M���-�6��n�6��6��#�^��;7
�!;Qg����ۮ��t@�4P�L�I  8�` Ӧʱ���p���U]A�[��i6 6�1Xwa��ڕj�G] [,��U�Ć��GEjj����s8�63��jy�KT���U`�^xk�8 �"�|pUuP'Jz%�����iV
Z�UZ���]kv�n��6�r��$A���A�n�m���2 �۶�'�2|$ �Sv�n��<dZ�wE�W*U*Ɉ�I;�[�:^�&�Y��[�m�I� ��Ҷ$pm�6c_WaK&����  W.�$6�m�Kh���>���o�   �   ��݁��O�m�l-��i4P m��a�  �k)oP��mm���i6�I�˒ޠG$84P��[p�e��R�m6� 	  =m���� �	:��lJp4�nXs=*� ���n���v�-뽷a'�m�Al�m� *���6����er`�U�\��FB�+jڢ$v�m����       � H 'K8��@�U�UV��m5 x*U����j�@j� 6U-�Q{j�U�UT�bD� h��}��m�!� Nt�/[��   ���M���m��   -���VvU�
 6��@UT�6ۀ	�  m�m�����  ܴ       m�ͰH�M���S[�m$-6Ԁ ��a�@ 8   N��I:��-��tVi���a$���6���k�l�p�f�p$���   ��    6�[d.�I � �I��c���   p5��H��lԀj�6��m�ړ^i���-i�� 4IV�0 v�H�m�� �b��  �a�Gi�޲c��`&�ղP۶�A�Z���*�`S?U@ECkl��I�d HI�m����_�   mr@�׭��W�~���u� ��&���hh�l[��` YA �� ���oIdA�����  ڶ�-� ���`A�m"@�����c -� ��`$�#mm�[m�!č�ݖ�    �mĒlpmm�m�$qí�    � @ Mَ�` ݴ�im	�l(@J�+*�V�*��   p:E� ���[- A$�8��`  � � H-���_���(���߀�� u���h���D��H                        UUQETR�UUUU_����?��O��=��Xa!`�J�1"8D0DC1�A �JPL-�z��_n����	�����r�9�(�(����r�Q�9G(���r�Q��(���r�Q�9G(���r�Q�9G(���p�8�8G�(#�&GL�0�&	��`p�&Adg�����n��g�܂8��(����u��ow��ϻ����~!�QM!�T`�����C���e	 ��9�r2@H��N(���T9�����+�} :	A<}=T1wЪ�:A�΄o1Uw����9'���A�A�E�M�t��� M�f�=@�T�1�d��CSե�<U�ԏ�E��N�zq�G�_'H�t��y0�z�;�Qe�@�҇�R��F �6>��ǠW���t"��zt v/�!��6��~��>/%f!	}P bTЀl�;;DO`v�*�
�U8�@��UN �4�v'`��h�HP�P|;Px햂V"daB&Bx���P*�@�D�4ʙt��s�U� x��<D�VE�](����< I��Q��P��2v����<q�Dt�	�� � F�8� CH�ϊ�8J��J!�:Px���4�z����8
�����i �R)IbRAi�R�Hs����=�����&(HH�@ = �G�T��U�OEb)Dd���0��(�b���df*�bJ�%�=O6@*��U��(���M��
s�D��z�zE�*��Cv����?�AU�������_����k�#���?��o{� �(�EUW���;�������{��b��T�(9� �`�)QRhLR���� ��V�u�������F��ckq��4�F��Fj6u��^�<�}��H�.��R�A�� ����}��[@s��-��p �$ �p� m�L    ��g mS[n0R�0l"�b��mʶ���f
�H�ev���VA�
���1�%�Ży�\H����k�֖�Ʃ{vQ��e{�����4�K[ʼ:�^y[��(��5c\kͺY\��[Y�G��*���6�q�M�d�*1˥U 9Np]v���j�z=/*BR�=M�N@"\l=ғ�vd��T�ԁA�P���9Ѥ����ղɥ$ �����㪔�Zک��l����T�ɹ�o:�L�gv�!����u\�n֣R���t��իq=�y�Ͱͅ6lֲ�uMZS��6���KtȲ��nJ����0%\U^�8�ȼY6�9��$��C��2�����G	4�T�UU*�'�J��G9U�8If%�N*�j����l��\S�KP�9kR�Z̈́ɺ��b;Q�l�&5�p$ͥȋ��z�d�z��u�d&� �`���D.e�\V;Xݘ�
�Z���x�^A�#���vM�l�r���١�8ե�gkp���4cN{�:\����S<+��S�^���s�l��u�GHu�gsjv��:��uԮ�n�UUR��Ƹ5�e��m;2�HJZ�e�U�nͬ��nD�#���HL��&�qƇt�9yj�UV�`.[mJNN	�ꡐȱ�6B3�@�MF:���=�D�x
�S�-�Ά�|s��HMOY8��ԫM�UuMA���63qg�
����G���ӱ#�Z	И[N�Ͷn�ok�j:�5��2�f�����J��um�j+� /H�P��Y۔�/
�n;5s\6qC6���(%�+cl�����g�Xc��[���bt�<a�'M��V͵H@1�U]���v�/bNM���N"�f��mTE��uֻz�������Z�f�7���g _}TC���v����>`v�N�Q�)���A���z�"��]��g���}V���処�.���^���Q��8�E��ޞ�b�q0竜
c��:7'&��]��5�e��UmF��uT�ǂ��/@i���a獊����"�+���{i4�j�N��P+���V�.7B�1�n1λ1�]c-9��sq�lo��9�{s7Y�L釖�h���m�\n��iձ՗<�Xz�Gd��{:�m<�q&�WH���3feg5��6��W�������¼��ɍ�6y;��7�Mϰ�����c����� �{���}���`(a��$���9����-6���Ͼɰ9�_�:����0�Ү�����r��r� ��^�x�V�Gթ�n�4��;�6u�e<� ��^ r�xܪ�b��n
��*n� �\� =�V�@U����U�1~�_Lu:�u���-�JR2^�3.N3t�zv10:�.L��D�8�\L��΀w'x˕��JU�};�;��R�;j�T�n����wσ�T�s����Δ;$��`�����H�%AE���[%���6};�5��&���]�{=�`s��<��d),rK6*�8��S��^��U�(�萕 UO�UWU���x��������|��w�Bk�VIaB
8�q������ᶻ=;�J6$;%.]Ňn��g7:�ME7u3 \U��ܹ_ؽ�#�������y�ju�Dժ�n�����=��=w����߽�HY���暕
����Y���|�=窚FD�};]y�w���g��L*&n���"�ູ���Y���u���׺��߻�J�CVZ���\�y+��u,���x����#��`���*���':��ء:��fs�M�ljp5�nZ+g¯r�{��.��NGV�f�����.�S�{ܳ����w�E*����ʺ����)�.>��]�y����^����eD�]TŐUU\���Y�y+���_����?t^�A�ch
��޺�{�\��=�����
��`�����<�$E35�8u���{7k-en������YS�~��,�����Sn�&�ms�;d]��uX��q��r�������]3BәT�|����nn�]��+����'?w��>�%n"#�5�y��K��踙�.*.�f�~�{�i)_ؼ���<��or��4��P:�ڇ{�[���Ͼz�������9�X�����mO5��3��r����,�D
9��zuUS3E�u5UyS�~qܞ�.n���Y�}���$�^��׻�[-��*��r����bzsp��r=�m34�5�؇v9ѥ�ոS8l�ImsPY������Y�2���s3�9�v�&��U��mjs�`]�u!��F��[��m���`��K�^*��B��u��9Cn��ͩ�1vS�9y�E�,�Y���%���.�uc��[aː ]�Y���F������O��7����P�Od�2ֶeІ"��H�5Z0�;����o@���e�h����G�k���Pt�+;�����r+(�MР����s���Gy+��dw*W2FF�
h�eYSqWW�w%��5�y�9��ܲ7�ʦ����������{�G��}�>K��	~�=[R�';Tv�^���}�yr���g��L����d�������ܳ�_ؽ�>JyO��"��GS4��M���N��j4�����\p��ݲc<>ʡ�Z�Q�h�CNZ��,��g����Y	O)G�b�'�jq,
���*h��{ַ�����/���T]p �X�,X��Ȅ��}=����ʌ�gX�@b�uU34YWSUW�ܧ?w��>K����d{���`@d�bIi���z�N����S�F�
�(�WS0\]���r� ^K!)�6Go�dytһ>�.�j�v�/���	�uD��]p1��l\%3K�m���R�Ƣ���+�[���kޞS�o�g�r��yp��*����n���!)�8���\�}���ؽ�>�
%T�E��[4n����]��O|�`��A�Q{�%�����<>�����ԵIj�����\��^��yO��r�ùD�*�&詢�뺫��4�Y�)�:}�>����r��פ����v���s�Y둸y۵�$Ilu'�5�uV��������U�dZ���O)���Y˕��Y��A37��M�\���,��+����<��lzh�&]��uy�i�ؼ�G)�?w��=�����6Z��S�Չ���=�=�]�߾��  q��@׻~���׽�"M�XF�n�}���~����_۫�G�TҊ���.������1���$g{u�ぽ��p<sJn١�0V�v6QTY^�s���{�}u�{���<����e�Wqww%��ܹ_��JmwϾz�����w�OѷR��][%��K#�򟼻�gܹ_��UUS3E�tMU�r�S����\��ԖB��AA�a5Us����G�i���O#��z~/Ϡ?8�Gm�J��A�Z��oXI��:tnt̳n����կ�;�/����i{Wn�I׎lm{/g6�J^�&� �y(�e�H�tH��AN��ͤ�nV��\X�݉%8a���1ّX�6�u�x�_6��h�=k�N��^��ckJLg��D���v���9��-%�y����M8�t
ֶ���;>5&n�S�mb�<�F���b�K��CB t�ε�oq��ݼ�[��;�']�k��, ��$����j�z5٣P�P[K4*G�uVi�e��u�{���T���Y��J�*���
.n*�����#ܩ\��%�rJ��	%5_pE�S7au{�)������>�9'W���Ͻ�L������ູ�����W��dyO)���_����-@�z��z�s�ﶹ��=~�������J��������M�[�mr�7%˵m`7;46�gmw=���k��Okj���N�8K�\�S�����Ͼz�����kZK��s,<���s-��
�`�]����.v��85�=�����޺�<�t^��q7�d����$�[���q��^��<�퍎%EI%R����늺�����ڹ^G��}�#|<���.�jB*ˊ����d>t��ry�y+�������d&���9�NEe�lrWy^��@�wr����rQ<�����x�V^�7h�*f�.j�9�s�o�g���j�Y��!M7UCATUW���}�֒Im�w2��{=��Ͼx�B��y�CR[e�r�K���{����D1�f���̨����˛����#��ڸ�,K�.i}���Rʿm��K�@�`d�]�a��$f�[�����a�)�]�|^MQ8G�ܽ2};p:z�)�ںq�8;l�6#�hHh�"���:�I����&����BP�|�64��I�K@a��Va͌AX�2`NITa�FBT<NNJUц��������%�I���&ll�"��MQZ3
J�Ih�V����;��Ǉ��WDg���4x3X�Če�0�#T=�z�(vt�>��UY&5�ð��PRSj(�� �:!�w�5�]��B�~���S��<��W�+����Q?^���E��b��� t)�� ���@�1��J�U<T6�~�yлG?1�	��YQ"B߷](�!Py��r�Ԅp�V�n��	$\��6��IJy���┥'�y���JPK��]�H5�\�;��$��TK7�����pz��<���qJR�D}��~��)J^�����)C�w�}��R��KE���%nF��]��"��;^����N�	{#���,���n��v��{��ݾ{��Vgֵf�qJR���~��ԥ){�o�k1J��︟�0�)J��_��H5�]]X|��W���]��JR��~� ��������R���o��'������ %�=�_�a��ckv�Y��R�=�=�D �_<�*!BY��ҋ"kH�}�ih5�X���M�:�v�޷s�ԥ�Hy�����L�������JR��~��$?B~�òB�L�JbSH�	�$��bkB.�%]�)�
�"����~�=@Ҟy����Y�[3*٭�f��)JO{��R�f!�	B�n��D}������v!G�}��:����n���$7g9�mI֢ٺ�9����Fq�9LOkﾾ>��᪮؆���)J^���┥_y��_��(5��┥'�y���)KϏ��[6kV�m��{��7�=}��pz��<���)JO|�߸=JR��{���)K\����$m¢Y�n����i~�:�B�LB\��ҋ��F7/��!�~n�Y�!<pH9��"jE��f��)O|�߸=JR��{���*��(�!B�㪈A���g$�k취�n���z��/O=�|���U���?8=�R�~}��)JR{����R��	��U��0�v����w���]Ul��f�ol��ƖE�����6�C�VM���nᱲ={7��%�ζH�ݮڮ��ܛ�n����d�F�In�A�� H�`�l�f���� ��qt��q��}�{&���Z��	��&��U���Rn%lg,ը6�hh��@��66nI\����K��l<c�̺�n0�mnƷ�3�u��M�3v�����iԚ�o{�j�{���Ѽ�3��p�R0��RM3����=:K8���;^�7n>��Ws�����y!�~�����(��TB�!Q�β�D ���@җ�{���)I���}�i��3z���s[��JS����)JO{�߸�JR��{���)B��������)N��\�6R���ZA� ������?bC%/���|R�����^ҋ"D/k� ��RB�3%�g�d�o{��Vo5�R����)JP������R���w��)O{�߸=��R��q���f�j�ݛ��|R����=��ԥ���矟k�┥'�z��Y�GHS��ڈA���9����s��,��&�ý�uj�k�����`ssP�랻������v�u���3�_s�ԥ)����D�'�����?#%/���|��@0@MJP����mk���Z]ϗ�#@=�PrJ��"R�����Q�	��T��8 $��F�_j!B��D �_>g��?J�)��������Q����1ٽ�|�)K�~���(z�Ͼ��"�k߳�R����pz��;�`&�Y+�c�v��H4��Z�w3k\4��k߳�R����pz��K�=��ZA� ���̒$J�d�f��ָ)Jw���8�)C�{��JR��~�D.L� Qo��E�"�Q�׳�=�t����,�گ7F�',3ѧ�[f����ݬ�3�͸�
^ӧ.���L~�)>�߿8=JR��{���)C��:IY�!|�����!{ْ�3ޚѽ�{���k|�)K�=�|R��-��QdB�|��B�
3��J,� ֑��br��R�V�m޴�Z@=}��pz��;�^�����	���B������u�ߜ��)Q�}��i��K�W��rIp��n[�pz��=�ﹻ�R����pz���g���D Qo�ҋ!P�H��K�XU��n�Y��R����=��ԥ){�o�R���}��JS�����)?@h�~}�h�6�7���N�9�uEnO����h���A���.�a���g7�U	&��`���+ůƴ�ZF{>��R�=}��pz��;���qJ��;���i��t!��	��V8�m޴R�=}��pz�JS�����)=��ҋ"D#<�j!BMco��G:Ff�7�\�9��R���w��(O}�t��	A�o��!�~n�Y��i�nDXXHR��7� ִ^��ҋ"D#<�j!T�B_6���JП��X�3 �t'Gb�> ��]~\O!�JO�7���6f������y��z��/|���JR�:��<��;���qJR��<��R����
����G$Cj���Yb,�kc5�Nm6۷Pd�3��l�Dc�^�g���{��}�w�Z�kn�����)C����ǒ��~��n)JRy矟q�R������5�_�*��c�F�Q,ܳuk���O>�\�YQL����?8=JR���~o�R�=}��B�)�~��^�®kXn�Y�����>��ԥ)�����B!�����ǒ�����7� ֐i{����z��.ָ)@�}�)JP�y{�ג�~��mqL��d��=����)I�}�O�$S�Z�n!�v��Z@��3�y)@�w���)I�~}��JP�}�ih5�_�K�I/�������Q��*ٲ�i �n�8�4km� \]��WMv�L��F�w�D�;6�㢇F^8�7=	m�i
6��7�2n-V�H얍=�?$�k��^	2YY�:WN�u�c��9w5p�ګ�݂�ÝsY4�W��xf��$BA%�7Y���ت���IA����TW%��[�;��+k�s�	�E؜]���Wj�K*t
��M}����ҫ[o��ٹf�ہv�e���\r�y�b�5��u�Dд�E��u�{���WٻpF���9��R������JRyߟ}��R�����|O�T�J�>���R�;�s*�I �ѷi�iZ.�����?������J��Ͽ6<�q�kK��|mk@��K���V�mIj��o[��)J^y��┥ }��JR�w���)I�}��R��������V��y��R�*K�������)ߟo�R��y����/1V��KA� ����W�7
�f���Jw�}���)I�}��JR��߷�)J���%)N��u���S ��X����ZS���#��r�#$鷕��:���zo��p�6�v��:۲��R��y��pz��o<���JR����j�R�����\R������ZӬ>��N�o[��)J^��}��	���&*:��Tx��A�qaWB����f����ߜ�c�JS���u�iJO<�����x�%)��j�Zѯ�xn�E�o|R������R�R�k�}��@"��t�Ȅm��D �A	�۞r�fl��Xo|��lz��E>�>�\R����>��ԥ)}�o�R�=feZ٭ ֑�y�'aT�
����E)I�~}��������}��)JP����ǒ���~��)JRw�����J/=�z̴�8�v�4]�m9�m�v8�Ͷ}����"�{4}�����g������������߷�9��_}�ǒ���~��"Ҕ�w��pz��/�3+4*�P�VYn����g��l_��)}��o�R��������R�����]�$�/���y\rB8TK7���cԥ)}��o�R��vy���?BhP?GH��@8!L0=�!�(�K����y)~�\���)C���v<��<�����s5�국�R�'�����ԥ)}�o�R���:QdBK�}��!g���n�����T��Z� ֑�^˽i��_}��)zw�┥'�y�mk���Z^}2a�Kk�ء�#�P���um��۔^�^�넷׵v���l<�?{�#h�	ۭV�U�w� ֐kIs3(�R����w�iJO<���ԥ*3�˽i��K{0�A�� ջ7��z��/����R��<��R���j!B�������d�xU$�K$�zҭ�H4���mk���Z#��|R�� �{�����R���2�ZA� ����M�mU�P2�w�u)B����)Cמ���){߾�П�4�hG�֞�� ~��9͏ҽ�l!0�����U�ܜ���ԥ)w�?>-l0�Z5f��z������~��R�/|���JR�����R������)JR��kK��(�wV�l���Z6���/^�tpzB��箣FÂ����h}��ݽ���Qlܳv�\5��3��z�����(�!Bc�%�!�x���)O=�����\�a��k{┥'����^�@R��~��(z�߶<��/{���@�)=���Z�h�7��;5�o�ԥ)}�o�R�>w�}����d�C����┞Òf_�k\5�����)�XQE\�jR�)
��~lyJ}���┥'�����JŁ�����JR��^ϾPn��5n��wZ� ֖w.fqJ��H�=����)J_����)JP���ly)Jl���}�9�sZ��ִ�]����$V�j����4�X��'�͹�Ɣ?6&�ﳀ�����-��0� �CjHt����:;�қx�U�y�B�tlN؂\ECb�a!�fB�Gx[:���(C�2LA��F2�ĺ�DI�fۣ3N���ATK>@�Jt>���D�9�"{���j||�i�	�蹛5�UI�adٙt����z���
R�3e���8������28�`ݹk�lq� )\�� �J-h u� (��  ���6Y5Ͳp �Sj���e�4<��B����$*��ԛ�N]I�:���XqOn;6����0@��O\N��u<v��	j�FwX�<�R���n-��r���r	��ՁӮS&��23W�m���9�H�v��cb$6|۱O=���59�ɺhU �t��i9�+���Ջ/e�Ꞧ�us�ݫ�3��Zc(��lմmU��I�轋���s.ak" ԑO�*˚nH�
���Fv卂���۳��m��H���Se�s�#6ѝn1*[��^d��gSj��.��q©�bHm��:�a����{j�`֭��6K��K�ƻP��E���,S�;a.]�B�<kn8� 5��m�� �Քې]��f�I-�uK�2��#�gk���fltL����vq��2 ͊�$��u����G:s��$M+ڗ�m��Hm���z�  �j��:6�wj��U�l��a�` *��t8� n���R�bj��U2 )kP���v�� d�I�� ���b:%%GhWv@<յ�h��m�H�lőge���3��*U��p�3MUT�p#��:�e5��3�@�LT�&Ir��ZT�ke�l�Diy�8`����٩RX�˸�]�"�V�G7L۵Uw���Y���)�C�=r[mp��l��d��l��I@�ԑ�[�U[�'ir@�J�jM 	�Y�3�w�eRy	�Z�]��\�]�.�3`�2�U-U�.�ylƓ��g!u�����-'[nS��	 �*�USu�8��퉽���ر��/Nݬ
 n���*�Ŗ�+J�<�R�:7�VΐR!������g�M@3v��
�W�������L�%�apN"ř$�
�W<�ðWU[��s[Ֆo3Y���Z���#ҧ�@�*�������
���t������(3�+��U;D<�?Bv��;�۷��{ֶf�+:��:��@:Ē7���Ş�c��Rk�f�P��M��ڔ/h]�-�v^����5�֑��A��ݱ�@�Ý1��2�[(\��jx1�`��HI��8=.��[:��
;7ZK�۞N.����GC�2Q�ў�=��9 ���$v� ��53ͮAV�4�ƌ�Z&D�C��%�r�أ��tX�Z5V���%��B�G6�4(�����;W<���(qo-{���,�힯��=��
��Uh۴�Zi�s����JR��~��)~���{�)��|mk��4�����ڶ�]U.�t�������h�;������3Q�Ы"���v̀s=�`g���"b��n݀n���+1yW��ͭ%,���ZY�\6{�� |��}�G�3�;�9t���@mƨ�$�����s�$����\ ֝��рzn.�.�$��7b����$�t�`K]�<&Te5n�l����rRYĒ�-�Mm��z�Yw����Zw�/+FD}{��<�"��"��
(������Kz]޵�kZMh0q��E��1N�����rO%�7@N���*���.����3/@|� w��� i;�y;�H�t\UPvL�ـw����� [��В��L�F�ի�����ٸ�	.�t�� ��������� ������=������]�V�TW�8�h�::�s��;I��/:�^�U����Ok��s}��
�(;�,�`�g����_��g?����3�??,X�~rB8TK6�e��� ���ސ�x����}�(�f!��4�j�RJlw�}�}�o���'�C��P:DN���u�A��\6�u!��gζ��R���Z҅3��i }�{@g��(<��k��!Lb�eMQE\�`#����y��`>M�I��ӛ�f�d&���g�k�v�sծ�\��B��MGK��M�/a�͌��<P��r �Eq5o�w�gr��;��7@l� ��֝��J���⪀��fn����4��}.� ��_�����ح�U�P5\��Bw�ۼ">�;�рws{�A�-//{
�HU�A�Ye��ѭ-$�ۻ� ~|e�{]�~P�-jb�)�����D�/�#�~���W��x~do������7xw.��ִ��}��l�3��ܻ�;x�npƮ^�b��3؆�w5���9�q8&���7M�s�[֒��C�l���IM񳽹���� ���D`�р/r"��"�[i�e� 3�˿�I�����=3�ݮ��^n�1S�q�xTY5w�Ӽ������w�S�ɻ��$&���񙗤Nـw�����ɐ֝���D��*�v��M����� �Ii?�ϯ?<����|��w�ʿBiL	DRʀB���D�نETD�F�����k��W)l�J��+�g-�-��ӣp�]!�y�֓\rvW[s�Unrc����vퟥ@Ys��9���^0�Q@#���Щ\N�9=���j��g/E歔6�;q̙^��K��6�n� � T��ݮ�K��\p��+OQZ���t�r��gEM���u�=)�[�\��m2Wm��ڂGB���2��^g��)A�4�kK[]�]���g�;s@-&�Ri-kSI$]�ʤҁW��0�g�X�PGOK��3�i��<�LQ�)j�E]U,�����v ��^��F���@$�n ���������i�(�+f �~���������p��nY��=�\6{��#�<Ӽ3�����gܠ�Dh[j5D'	M�KG?w3�� ��˰��i��}��F��T�AN&T�Wy۰�q������۽�3޸l߽�s��&���Z�vHYn�3�����=:ܓ�y]=���p�U�:�W������m�EES�݀w�e����`~�oc� �R� p�e�ՐM�]�&����+�(_�$�����~�v��_�@����DBR��3���z�T݄�v`����4���7xv����a�ajة]U)/8*}�{@۽�=������y���,��u&ՄQ�R�v�ٗ`~�\��s��t�;��U4�"�v�<Y�6-�Z��3Y���'K9�y�k�C�L$��$I�^��"�[WnHG
�f�wx%6��M�y���n�r���ж�j�RJl߽��|���ZZ���� g�{D���w
Q���9��n#�6���^s�LC�e�f]��J~�,��w& Hv���������r��<��p�1�H���a)���������� {�s
ﱻ����Q>׽�Y���\�p,B-�{�����o��KQ�M�y�x�n�$?Du6��nffKG=�X�Ӭ�t!�F˓���V
$v"Kv�<ۚ��p]r�Ea[�#1�݀����=�}I%@f{)P��y"��ة]Te� Fg��kH������R�����""T�,ժn��dQ�R�v�����}��?~��� f{.�����+�HG
�f�wxx�P�� oh?(Si(P�J��@�Q���ߝo��ʾ����&�
&*����� �/�t�� 9�]����k`$���	��]��dq��P�W�hٝκ2�u�u��t���峆+�dz���A�UK/��}�]�w;�`%�# �&�� ���SPS����鸫�� �����F�P��i�~�kI��}����y�� ���k �&�@T� ����'�����*�欚����'9��xϲ�{�������R+b�uPe�� M;�LW�r呀w&�@�#���֖�-i��.C�����V���:���Ǜ�-n�%�y�r����u`8��5��t�oN������c�X�+��fI����O&��J����1�۱q;�^ێgi�;I�&��v�T��U��-G�yT�b�.3��Ch��s����H�Ib]��`���j�n.�f���/,L�{�}� ��KA̵x��c�s����&	v ��o+�7�[$>@���(��F�]�f�+�ŎsM�.��e��)ͦ�v��nYl����^�z�5ݎ��^���m�?�ڼ�,��t4� �P��D��������O# �� M;��6w�˾ii�~�F#68T)m[~�n�&���Qxй\`P�5qA�UGo8��]���_]��w�[��}���}�t��mvu]�� GЎj���r�06��lϳخ��kA�k�KK���S	T�]D7��Eg�5qˑΐy+Tӧ�y&��6�}2�gm����g�?3��k`~�fs��e�Z@~}�M�s��n�	��3V�r��������i���8�:�;�2��E�x)�����*�>����kZH�煉ڤR�J��L��� ǉ���|�l(B���"ƽ�[@w���p���u!�����h"�<�dɜ�R�>x���!#w�l�:	�������'.������"<�y�	�x�y��#�]7���MMԷSbv�-�qhݜn�;,^�e���nT/����/����K��ɾÎGC�{�@{^��<}�=/�Ȅ�},����ly{�նH��l�E�� Ǐ��~���e*A�����D�JMߛ�r3�m�=:���?��`w����kjs�o7��{܄�I�Kk��m�H������>�i�O})��Vo�7��R-�<��u�f#��pi&� �1HS��P	�ٱ�m�a�kN�5�,"p���ӘB�Z�jǭh:å;N b����T��Ob����@�"�/!
1 ��M7��:N�C�4"$ >t�ڪ� ق'ʃ�l��b(,'�/b� pS^|�b'@�b���\ Cc��j��*�f�뿹�����{2�]A�nnp�����9��@N��j� 7�=VE\��U�;��� �KF4� ��`	r��?����QU3_�������103���#��=Ͷ	;$)k�s���"�{4~}��?_o�x9��=l}��׽�=/��3�J�(@y�w`]��!�����v^w�`{�����x��1��D$���y������w��A��,k*��5������~�{&���Cpl��MPV���B���x������3��*F"ȩ�@7���Õ{�襤�E�Q6j����e��ֵ�:�0�d`d�r����_�_��˻�.x��㍷�0�v�ЦPtr�u/���t�Yh�5�9���[�$Sn�a�۰1�F �,��4�"#@N/ rn������.�2�����9��@3=�`u�}6%�9��7UR@��J���Ot���"�ʰ�d`���jX�n*�y���ֵ���{�{Y2L�>P3�J���was>^�L�"�iTwV�n����M��ZѬ�g��n�����J?Fʄo ��\�jY�ζ����ruC`�ԻmZ�m��:�E6^NV��,�g�-<����26v�#��V���g��p��b��\NF5�7s+Ʌ#��֢�!���n��v����BTY���1������x��G�NjR8�6t�t�p�^��1������8�5r�T��G7�ִi�f�c���	d�J���������ZIyij�Ii�<q��L]�6����xA:�:P�[46sͷN�\��TN��:�~������r:��e�V�˿�呀sr��i� ������$�fی����lً3��m;�;����S�#" P�LUU��������`��=��!(L������ �ct�)��\z*�[�;����� �m�6�x8�ݱB�]����ɘ��33| �̽�I������甭��Z��`1�g�wj�G�3����[�۫R�<��f�m,huU"��I-�`~��� 33.���5�o޾��;�M��kz7Y����j���͟��<O�e*� !%qW1���vh�nMo�fg8?.�R��;�\�`w��	RS�y��@��� ��t�s"�p��Mݾ�D�c�~��� =�J���{�x�m��m���]�`|�w`����ɠ39�4�MD/����:�ڣ�ݶ ���s�ɫv̹�EYɜ���`*.��C.�8﯎�^j�d�໼��߿^�MN �%8�fs�{1�$S����n���3�`%IN����m�@97wQE͒��w���f�o���M���ľ�)E���AB�N�@�]�}W�]��˷��?{�h�uU"��I-����� m��;�� ��)�{͙mGK[��r^p32����Q�%IN�����yN�**	�����'k4�G�:<�L��J�rAN�V���^���M�v"�9F�Hj�(�r���6g3&�����(�K�ջ�����uȡ*#D���3&c��H���@n��h�<��f��&�f��]��h��ͷv ��h"!D{ϘPޞ��^^^�H�F6j����Z��	N��h��(����$�TkI%�KZ����M�}w�߼ڲ5>vZEV�v��r�؃ZKZ���6F�ffs��˰=��;�%M��(	�Z�g�'�H���.��[:���ny{l!&�U��ųu�����g X�2lٙ��fe����a�}p�s�x۪�U�s��y@}����p7w{H�w�Xd���6�V��ܗ� �̻�Z0)*���ot��ʛ���**n,.j� �V�.eJJ�i��>ִ����}v�՘�W�"�p��G����s^����٠;������>LG���S�кSHq�z�{�[�����U-��4P�oXI��:F�z�I:��ܭ�����u�ڭ����n:����f�@l�8�6�\<MQ��)g`輶�%A���j�ӣ���O��k�
\<QA�c��l�5ڧ�����n�,n�X��J���7mn,�h
�*�v�* yx�\cXkn�<nCV�-��8)�hJ�9�v��Qrf�du�3�ܚMچ�����Z֥�F�JJ8��B�H��E-����Cq;���m�ø�ZzZ�5��8��Ld&��������;���t7X��`~����W��rI�&�T[y�3&d��;�`[td�~M�����suvT�]������`7�d�{�2����L���͜�����JJ}��T�'��x۪�U�9m|w��s�}������`{S�(g3&��׍��\�=,u�
<���i˓mv��h	y.&����L����mث���Dڍ[c��r^p��4<�
��s2uDBW!��۰��^�ỡ����r����|o�$�]ֺ�$��{͹�7�ͻ����y\rjB�f��=�1��=���i��g�`w�l~��ۄf܍�P�����7�t��jрG*Jpu{�$r)�M����{&c��~x�:np��� �E|Dâ,�+b��C#�of!�]���aK���mŇ�D����V��ZG���{�z���i���p	�s5�͓_�sW�h	�s�y��@���<�Z6 ?{�~m�T�*���`w=��{���9~��C�/$�$� H (FBT�P������Q�����{<c��V���A�/8#�%0���@{_Y@{9�4�� ��y��"��*9^���=�-���Oy�xݫ����]�Gg�c|������V�溭�g=��̣Iڜ�;��җ�@��jmȤ�TG#����1��ot�����0ld�F]5S<��I�f���wz���7f������������N8�_D3U�pd�4�;��R�H���u���v����LvZG���{�I���g3&������K�PDB^�����#Z��ZY�7���_{0���2�Wo(�1�
!%��1�>y��_�}]N�ݑXȅ\�F�).p�l�9a��4V�c&�Ŧ��<�JG0]D�T\��5ws�sM78��G�Z��]�����g�yP�j�T�݁���~P%��P�����|�s͙��(�U����`r��#胚n�@N�' IРq1Ȥ�TG#�������������ɘ�I������M�͹5B�W84��	��y�D`ʒ��?��R_���o{��!#�H�ݔ��d�Mk[���[So��tt��BhM�@�ή���A*:FB9�
\Z08lWd��,	aI���t�t�)��,!2Ē�L��@H�H�Q�Q6M�B���p脍�q�J �f�� ��iR0�B	7%MEUS�#7γ$@�H`&�6ʐ@D�A�4M�P�+�d/� �S�1<��B:":0Ȩ�af�e��ӵ�X"��#M���a7�m��1k̆�%C^� R��U��@)\[Cn�v�  1'$ �� m�\ 2    V1�6Y%1� ��N���jQH{����3�h�,��u����P ���b��Ñ��f�!7�:z�`Su��Cc`�u�9���s�6�WIĺ���1�!��o=��3[m���km0��Y�zg/hMnu�V�+,t�����T�뤻�hp�
�	��/8.6Fx*%�ʛ�n�і�4�[n,�÷��-�-��E�gldֱ��l��
R0��ƥA4h�[���+!��5vQ��#����nN��V�:�����݄h�)�v'5�̪��@����\�]�<��W^�S\��>��6�a��Ϋ6���xvm�a�E֋B�����Q�U��8Ӝ���mU�,��]� �X �nӍ�ܙexkv��$�歝 k5���_\.���m���yK�]��۶iDme������[9�uUt6�)9gW<��� ��F �w�kcg��Ve�f�#i��f ٶ�iG!5�ɬ���Ѹ���o��JR�i���/(L ���X붶�l
�=�ce��\\W3*�V:��M+�z(�'��		�p�ˤ,l]{ �:�0����k����+eK-���R�vٶ86���6��%`�	�bu+P�8���at
��h��ܝ��F�˭/X����ck�϶"����;�+��͙#���k����7RZ5:e��`0�/j��4���cv7KnM�H܆�E�ݻl�2]״�:�I��6� ۱(C��ɝ�*,hg1�P-]��iu� E�5�V����].r�q�9����Q��Jv�  �K*�i��� P[���*��<�˰J4�5v�Tp�碩^T�����Ss�U8&՝�1�F䒫-v�ӂU��j��	ej�����K�#7f��p?�����FDa�a�a�VfVXqB	������PO��T��\^���	����~���4
��Q]�tآv@+�x~�>�ZJ�ֵ�i�K���V�Gh9#i���/j���k��mӗ����q�M'�k&�4]Iry4�t�q��ƭY]N�J�1 J�*�b�n�"��j �ݗ3@�m���^��=�ӎwc\m۞�Y�hD�m-�]���S�L94�Y䙲�sW%v�T]C�I#%J���ݭ%�����0]q�2�M��X���瞬��T���t\K�K�n�R�ӻ^�m��?g�z�'l��+���'79��fw:�fvôt��pr�yd��{�ӮrF�{j�۾���>����6};��N��a������[���WY�����jрt�)퐖���U�����fa\�h����͜{&c�9��@N��ɼdh8NJ��ӕTڴr��I#��,� �Lǰ?g��������=�3��"i�ն8�&j�t�9�+Fʒ�4�8�2�(�drD1֠�u��g:ڑ13��pt�ӗI�e���P8E7��ǻ�����I�R�W�>�\6z�������3�05���:�yLv)#U�Sz5˪�}�\�/�e�=eC`*�*G�[v�f� �;�y�W9Μ��5B�)�=���ܙ�a��kKF{���b�}|lwǦU+�FV3U���~������Y@{��(!$�$gٙ���j�I��ʓ��^��{�[!%g3&�1�����s@_��;r�rc#��v��W�r�mcv^ձM�2 �(�F��,��h}�ךk�ߍ��|nhm7vg�V�BP�F�e* ��22����բ�װ��ٙ��--Dȷx�hmҠ>�fM%	$���D5��ۗ�ޙ�������
�C�K�K}����nh�[��//�3�m���Y�����+�*��(���R��7�5�v y���'���c�I���v�?fM�kZֵ���H��ݐiE�.V�������ͱ#�s�ң�9��V�.F��'p࿡����}��#n���TB��g�}�8T��+U1}�`
y*�7�3*����TKy�3�1��I$�}��{�&�����>M���Ղ��mn��{<��s��jC3�9�(��K׻��O�{5��E��WR�˷�1<o�?7v�75�'���������T�00D�քA�3�������^�9�'��J�mZ9l� _˛��np���O%Y ~���Z��H���H)��T��+��*g�SI�l\�6Ц���Q7!#���k������5��ܻ�u��}��3��{y�ޛ���pZ���&�2�Ȥ�T�����V�0�$s��z�n���٠8ή��c�HB�6M���&�M7�}}�5M� �Z0��@**fr����&��{�5M� �Z0��^~������q��3U�p��+F ���4������_��$e��GR��!k_���\�*ٲ�vY �o�ӳ;��kH��#O�4���ݖ���^��Y��Q��Y�cN�c6U�M-����Y�p&(v��!rv�۳���۱vrܛ+�i]Þ���S;�EU�k�,vQ�)�m/ch�ZAVb;��3�:�mX꽣�ӭۇP@�e��/r�ݍ�<&��y��a�e��S�Z�ҕ��cTv�5�}��%�KI~_���MZ[\-��BA��VY��G(0ru�ܫ�iΊ�n�K-a��N�9RwqT�@|��(���� f�s_�$�
�n�vh�ר�c��:��{tX[|��"s��kn����@?gp�a(HL;�FUS�Tڴ��6|g�s�c��}��T���� i �(��&�fk0��� I�f�[u�8�,�p@uwɼWCRE����w����R��4���s�y'������.��'v{<��i���;uӍ��MTY0�݅��@�mYm���pA�39@7�݀��J�7Y@y����rx�� Gy�P����B��BV��o7f�/��*����~��6r\q���3U�p��|�����G==�6sٜ��mR5#�<�N����V�JJ�i���� ?f��B��Ym���2lZ�s��@n���,��B�:"��U��Eg��vn]/j��3����=n֡����,� Z�cU��)-�p}�}�92���eDB�Nfr���f��,R��ܼ��1���߳6���(��9�ԦDH6������.O;9���n�������%؄�I4�!D\$�BI5�M~��]���~٠��^m52ȣn�.� KIkfL�ot���Y�QS3���Ћ,�u�2�8~oZI,ɛ{;�ml?{�`g�HL-���@YI�͙X�!��*9Nk�ѩo#�lgAa�[6��F�J�u��C5Q-�0�3���������7�kI��g8��jGx���vy٠�e*ԡDɒ�� �۰3&c��Z5�i0�_}�̴����x�?�~�4��	�s�>K# =�O���-Be��ٰIh��y���3&�~̥A�ZI$�/D(��?}r���|M7K���y�=�1��D�Q��c�2[�Pf�w`c�>uqqJ�Μ�n���M�:=�n��Z�H+�I��i��Nۤ$m؊8�vCRE�Y+��{# �IV �';��i �Ss�����"�Ȫ+d�\�3&��{3���K�s@?fR�����$�0L��9�w���۰1��)P��������+�Eb��o8��f=���J���g(6�/^��ݙ����㩚vW+��{kb��HצfJ={�`c�s@~M&�BP�D�JH���� 8 b~�Z�ލ����޶ml��Y���g'Nn��tLb.Z2��rՌ��l���q�M��4ƣ�X���g�E��;b۔��3��n�@j��#Ý[���+��ƻ-��c\=���v�ٰKTۜ���k�퇵Ι��u�p�� ;-��S!e��Ra��ۀ�[��ힶ���G2닐�Yñh:��M6�4���`�����"5Ӯ7��W�֖�崴U��6MGʆ�8:gsԐb�ݨ�A���V''-�3u˰�f���+kԲ�%�h��K-�������@�ov N��l���0�zN�DMń�%%�́��g9���ٟO�{�fml���6���]�Geܼ���.d|�F���4��P�xCRE�Y+��{k`u�ޛ���pd�{���<�Im¢�K���n� M7�t�����9���	IG$C-R*"2Uj��@܏5��n͎ITOOf�z�|㩍��/f��]]{d��@N���%��)�U�~���n2�5Q-� �z�{�S��1CN�)~'a�C�<���8����`{=��/�i&����>�R��f��5s��7`Ғ��M7;5�fJ�5j �R�o ��ɴ<n�_L�㩤

w�@��a%�Ie�`{�fs�|��׾�|��ٛ[�wޛ�~3שׁ@e���&��$囡4�H�%na�b��F�t�m3d;2'6��w�o�؉�C�J���o7f�~̥@z}��\��׻v ���Tڎ
IR�W�3���Š:w����ύ�lDB��b�5��9�I��vd�iX^�(�����:JDQ�����}��0|��M�U^U�~}�PaQ�f`�d��?<K��8`�cX������A�/�:������0|:%H�m�����ț��Q��1$�fl�X��Xa.�$M� ���d�4���q8H%�#|B�V)���q�I8�IfL��M�p���� ����8p���h	$ �hq�\Z�1�$�L�th�]']l�{X�;Ѣ$)�&(�H��I����b���;c4�0�f���:c4ƓA�l4%����i�=�Ԕ֢�132a� �Hl��dm�	� ����2˕%.e�T$�L4�I��`AL�9��#$��z]�·D8hꤒH`�� `!�Z�"p�Y��5k6��9���n�t��i`�,a�#5`�9����8����'��G���#�� �0�00��04_��F�G��:�'M�Q��-�m4˻Z�UQ��#6F0#0���`�dp#������01	��j%�V��v�zi�1�鉌x�fe~��P܀~�?p�~�]2~Ȣ�ۂ�+�(?��v ��	�~��(>�	DG�*����^�3f���Q@}�@gL�T�MY����otu� �,���Ӿ�`~����q�ʢl�D����sAS���q�����@f�w`���ARJ�t�۪հ��,�9�g�[�%�n�[�ԛ�jt�I�+�,�9R�x���˙%��l�U�&�ߴt����d�1:V�R�y����d�	��4t�����¨������.ʺ��4����+Gl�K�6g��Ni�X�\+���4�����;���g(?-�J��B\DJTц,�1z � oK�_��8��6�Tڎ
IR�W�3����(S>�;���ڰ<���DB��v?���z.6�ȅ�6�ټ�a+Js]V��p��盲�n�t�{e�J>�/]t��/]��I��9�V .cy�s�� |���?m�8���;f��{3�_��G��>�`��V�
*f���TL�\w�2���a ���4�
����"���N��{��?�3�����@f���!/>74��!�u�F��jYe��~̛�-%�{�~7��@?{)P���䄒�
&!Q���%�!-k���)k����!�j���6L�k�i�eѫ�t�gY {�+`��!^��z��I998{�x��ӁF�FVӑ�
�ں�9ǝ�7]������U���G�a6p|$f[N�m.�#HU:I��%K�N�Z�;6�{��jů<v�a8�V�7�X5ø�JH[kk��A�cr6V�2$t{
�3f�K��Iz\�H��%-kK��sSKIS���[l�آ5���ۅ��k��冥h�W<�Ai��D�a����Z��ٸ�UI(&ZK-�s��?�p��9����E�d�|�7q�!ș��¹���3����[��ޛ���s�����ر��Sj8)%J�vh*w1ڡ}̜�D$�^������uuS$��El�k�m/4�`	�{�s��ܲ0rS$�M��)�ٰ=��� �%��-/}~٤�N���g(I/�N!K����u�9A@5in�x�h��t#s���MKQ�����Z9�4ԍ�d-Q4���ɘ�3#�e*���l%r^�����Ns�ϔ����w������i	I$D(x�Pw�s>���*���9�O�1��f:�h�j�,��p)����t�j���%��G_�����閒�f��O>Ͼ���ߧ |�F��WZik�.���;<���b�ni�(��ڰ��@{�fs�/fS[drD2��-�D�ΚT���.1�N���lGK�n�Sy)����jK�9^�ٝ����}�G�ٜ���ή��d�!����p)��$�H���o#$�{�G)�9j��Y����+��LR�{��9��ͭ�?w��(܋�iPv�g�c�3ٔ��e*��u��`f��Ns�O� ������ms�>�fs��}�}��&c�--~���]KT���v�ΟVKKuFܨP�p&��m��R��@p>��r��B���e�����������ns&E�d`{�RUa]�UWi�����d`	%��i6}�`}4:X�\+��� ��}���{m�`�{�	B�E\L�Lp�9��<���2���J��z�~���=d��G�zBCX�k�_��������3�����H�TV��VmҠ1�w`7����J��Z֒�\"o4�T(����D+(92=nv�tu7d�j.������s�z:~E�n\�/#o��W�o���ՠ�s@���@ffR��|Q����U	���3�~̥@ffR�1�wy�!(��p�)����A�@�ٛ[w��P;�}�}��I��tFf�
�V���k�ffd`	��@n���Y��������J�����fSOw@iܹ�%�ȯ}����-���f0����g�!�I6�&�n%��ק�DA��ʅ�$�vV q��F�j�.��u/a�g���r(@�����=��-O��IM�cö�ݼ��n8m�vl�-�Q��/'��k����:�X9��)燣p�u='m̶��í��7Y�HC���/ld�:]���MJt8�UݡfQ�d��W�.�:z3!�6��8�L�հ�&Gg�=���ww?:�#�3��k��D���!$mB4���u؇�1ۍpnx9@��@�M���%k@����rY@$�F�s��/7���j˪I^��<�g����x��	�75�	D�}��vy�J�;2s����](�a(P�{���3�3k`~���୻"�SB��T"$�u��`n�vh�e*33k`~�6�:6j�������,�;���M�����Ϯ˸u'n{.8��kO��P`N��v�j�dJt�Ѷq�),DmX)�U'Ke8�Ǒ��z���fW��t�����l�j��K-�\�����W�I%�њZV��ݫ����@?fR�쩿{'��DܬL�$���=��� �e�g�KZ���&ml/fml��1��+�rO{v	D��i@��b���3�n7� {�ͬ�&�jˢ�M�������J���=�9�f舄�TLK��9硍��bK�ãt�[tpz�S���ȴ��V���#v�Tܐ!����p4�`	��@9�f �,�$��fr�����*���{�sv̀%�`u�ޛ�|G�m�u��P�� ��o�_y��p��î8��*pqB%��~ �GK�������ik����f����לٍ�#���3e�Y��|����� _�{�w2�]y�c�WtP�jYm��~�X�7�:c0�g���_L�Ja��\�$2:��u�j��7q͹ض܌S��x9a�ɛ��k�ی�5U� �ot�ـ>K#&z�d ��y.�]�¹���W�3������6�{3����X�Ҧ�jˢ欌�o(��%X���7l�uuS-�)����p<̛7v7�R�J>��.BBQj�q~[��m�m���C�l4{<��	�f���:RU�?t*��fF�E�Ѽw9'd�#\&-t4��t�mӪ��أWe�ˋkc���]��~ M�0�Y\�t�� ֛���&Ek�UN��� K;�U�<��V �okd57�Щ�C�˛�&�*,����h
Zu�i��8v�����9�xh���bd���6i<�>߬�� ��J�aB����P��_���B�W#��ٗ�3����������?���@��Z����������"�H��I$$�=$����j����)F�HA�k��������$#{T{P;!I�Cr���Y�a4�d�%$Д%!�� �t�]\���(`$��GD������A�;h�`���H�E<cE)�����m�b#��T�Kݷ���U����Mbk\�y�z��@lǼo�`F�%N�l��j4�Tx��Ѓѯ�� (�.��^�����Q@q=є��`�4�zP�q���.�7���k s�6˦a\l�88�s����������D�p �۰�n�      ��ZI6\� �-�ص�W�&�B�x´*+�pQ�&b� P#�FiM��4c��P������,GQ˵���H%�.�Y�#�v�����n�Ywj9v:�Wp�;9����@y��cn��[�n��W�ͥg FF�dܛ��(q��X�U�s\�����a����EJ�4�[��OY�	$�vQJm�S�m���x�	��Gm�9��sǱ[q�Ө�!ni��WaŮvӤ�`,�H�q�kgeC �{n�g:ӱ�1p�>�9�6:{v\����oK�SI'k\Y����-�(\v��gN�q��P����_A�1�������M=��c�].匀�Nɳ�Tu�m�l�l  �Z����󱙪�*����nŻUꀕh��r��!w3�5��:�f�`r8�9��]���7nfԊ�I(bm&lurj��gI BGm� zKw/D��gh\Ǥ��
������V���Ŭ@%q�ܲ[��4�g��㊊()gC;���HmҮ��1kJU*ʹ��:[��`��Z�6�]U�����34s&��]��ZR�U�޶��6v�)mć��Xإ-�L�l����P�����A���[GR�S�<n#*�%]�z��h'���UK&�������i�T��Yڃ����d�m��oC����{cQV��K�9����!5*�Ғ�1U[�'6՞9�)�ȭ��p�������U8�<� ���U����]Xݻa1�m�I(B�j�=�i<]7kjy+�'�cm������[��Y&�ν7]`�wh��@ Sb#M�U��g���en�v�Ufp$m<���!��USÆ���c�Ed�K�k�vٍ�i%��P��fV�A��t�=�*�p�Z��Mk�CBz Α:|�'=ENb/�z�������D(��h�� ࠑ�Dt����>]�w���{�9�U�d�׉ �d�㈮�����k;3��e��Z�N+t9���t Nl�j�a.6[jC� �%;K��u�� tv�m�U�Չ�z����V�W���"6��ۇ�ծT����Lڒ6�hu�'\���>A���3R�,k&�5q�v�����d�n��flqPj��(0�㰏h�I�쑺�����.��L7VSd,v9b)t���R��U@�Nt[M#��X����պE�j�Q�.n{u�i��;9F�El���!	%ӮS���ͭ�Ғ�4���@&�� �u6T��72]�h
[u�2�o�nـg}�h=�V�R6݊ID!�6i���v��YO���=�&˩��n������v��YO��Z���g8|b��
�r��t��0�daS?�Tۭs$�_�ozA;�`f}��	�0v("3VY 2�.����=8��l��zq�]ql<��v:�ϻ�M�}�wE+E%�յ�}���fs�{2��Zֵ�{ml�f6UI(&J�o7�r+��~���D$QC1��IG�BQȰ��‿���Nfr���3=�ɦ���Io8��`g|�0��`@�ot�P��7U�UU�75f �,��%X�N�@��Z�e�`Z�;���#�Ճ�j=�%��R��v���J�2�/v�+jG"4GZj��P��X�:����qΝ%�]i�'f����������w�?|d����� �j� M7�nـ>K#�Z���d��F(���j�[�	�dn�T��s�GJ�X�Ot���|b�ȭuʣi��M����l3�}�.�'�r݃����4�I-?f�Ӷ`a���,��ʻ�]/����{�bo���BI��/��;�<MUT��d���6��o�nف�,f�ȥ�X�!4�� �O�ڛu�s:�[k�X�al"�����i���^Ŝ�ߎ����[|�"]�B��6 M�2 �K(��%_��~Ͼ��3U��]:�M�u~�el%���m�f�۰1񌨈P�/y�aA��#��w��y�d��ۿ}:�&^�t�=�����3�&fn����	��y~�	�f@]l��A��	��^���V��e��?\T��`]l�:RU�s�������MdrV+��m��rũ'qͣg�[�0�܇Ym������13q��Z�nZ1:[)�?w���3&��W�9���.��ƣ�)Z)-��X-�V�DGy���۰�t���f�$���TNJ	��JK6;���9�f�l�:y*��_L��A2���|������:��M�9߳9����,��!	%ӮS`}��(��7���۰<�Y@oRQZBִ/�z�Z]�ɋ�J[m�T�b���ް��I#p�w��$�hݙ��W�U�z5�S�	n�Y#����1\`㳵�d�=�ٹ�6x!��6�߾������w���..�Ş�8=�16I��<�'	5��o$�Zֺ�n.ƃj�V,�gTl�$N	��n:�������]����^pk�4�n�EkY�-�x0���kZ�mv���0�a�Q�u�[f���z���rF9f�X��E�t��;'I:�2�ۆ0�ے��8{������	.bn�"k0`��Xzg�9��9��i ~�f��Fz���$�B%]v�z�w�7l�#�������>I�������G���� ��\6�[0�:y*�7�{�$;M�\]���$M�uf������y������;�f8�V�Kd��2q�Q�?c�v �}e�yҠ5$�|�O�츀�kn0�7dV�0cZ�^e�D�,����MlB�G��զ��<��\wWZ��߷@��ysϰ��M����4�vA2�-� �e�s�*f�|��o������w�G ��d��9�=��
�M9%Ӯ��˞F<�`Dͽ�9�f@�q�P��Ӱ�r�p?fM��m���0S=\�0��*l����j��	��y��sv̀y;��}�9�a�j�l��Em��+(��{]��c3���lۧ]�=:���ܲ/M�8��s7EO�7{�sv��O# ��������x�)�U��F'Ke6�ОF��V����7l�<�n8�r���/ ^kٓ`s�fs��(|�D��ӤJP��4 ┢-z/����{���J�G�/bQI(&J���lBG?}���2��w��`���.��.����� o# �����褕`L�����fC��L�G$BvM��ܵ�=��͡����k�ܱ�^{papr)��G�}���h���nn�y<��%X��� {36��9��o(ڭ;
).� �}��y��t��ή�B�31u�ԖD6䠉,������3k`~����~��8���L�n�=U�a�!D���ڠ=紨Nfr��(Q��(b�-��u�p��uW�^�&Z�nU[N�ڶ��ͭ���zl~��p�f���i%����g֚���+S��8�ܗYxcKԜs#��l3ԇC��(�^�v��'AM�8�V�Ye��<��E�ۻͧKaBJ�=紨��ّ5��2TKe�s�ٜ��ͭ�?~�ml���i3�^x�,u�2�W{�2so# =�L�#���}��1�,��)$wN�V�}�>�7�FN7����ϦR�N�R �^NZ���T��EVa�)M��m��v�0߽p����ʫ]��h�$n�����(,t鎥�k�j���Ξ�))QcnM�CWV-���G2[;&汻J^��"hl�-�6E�8�ˬ�ʑ�kP
��뒷l��]�s�C��&vڄ��g�M͍sӞ�4
gHI���q�ݬ��Z�Y�2���r�>�Sk�,!��^w!�p1D�O���vެ��f)�Pr3�9�v���]Ѭ^�m{��{�4��_��:#Ԏ<��f��M�\��ȚbQ4�=WUo��n���x�K�2��t<�<?߶�6�P|���@u�ޛ _���<�o�oUGn�s3# }�# �� ^m�wqvܴbt���w���_}��-ikOJ_�v���T�mO'�;(���oa�fe�-� ����y�y��>�y
���%D��n����� �7��>瑀t�U�sc�*i�]���#�,v�\p9����c����k�s��� � ��⮸X났���y��'y >瑀t�U�/6�@r�8&���kY���{�_y��9���(����%@��� �0�"B]��R.�7�H���� ����Z֛ؼ��D�ڑ;
Rݮl~�y /6�@9�x�y�2*��چܔ-�����}�8�Ϯ���6ͅi��������x7Sz�Sw� sn���� ^�W�/6�`����Z+KkRѠ��L�F�U��v��nW��lU��)��Bp��������J����n����l���=�F�@=�����jk�˘,���� �'x�n�@=�� ��FG���Oi���PL��n����� ?w�v������������E$�I$�I?��z?�'������{H`Z!�����a�<E�Ԉ��&�E���IJT�Vd��NbtI�d���&���t,�fHA$! D�#� ET�0������T�@fk4�tnt���2� �]�Z�)�2�4��@PRTAxDY!fTFI�Q�L�9V5eI9D��a <��^4�RSALM4[�Q�h41UT���C$IT�$�L�Ԛ�p�Ȏ$����4LG�t�����"��	"`��$$����"1��'#�RÈ��
��]s���=|�="qT�"y�G�h �5�@��&�� b�+ ��yߜ9A��.��ؼ��vMVFX���� ��}��������Pɹ�������.j� }�# 7�^ ��s������O5-����R�j�e�˓B6͵�ǝ�m�]�/�h#�9�͚˂���n�.��#@=�� ���;�Ƹ����[w1V̤�nJ;���ד��ls�ǽ�7�t��̻@~���j6���U��{���� ��� \���VE:��&��E=]�;�A�w��P�y����wZ?	$�	4*�RM����65�,��8�EU����ͭ���%	�Y;��/b}Ҁ<�G�fs~����z9lծ���ڬ���w�v��t�xA���$�3p6�yk��mUq��y�w+f�?w籠{���>�,x�cvj�2�-��������Ҡ=��P��vjI%I�ƴ�9�)!.��6˿f��\��ml�$�y��p/e�� �W���;
ff]Ɓ�o# M'�u!��Y��i��rH�(J�[��g8�1֖��7J���)P"x��	(4�Z�#I�#��[B�k*�Y(3��d[���2��Yj����b��TTK*g�趹2��9��.�"��.ۚ0��9֎�v��Ʌڃ�G���>>���Z.�۴�-�\u��.7Gn���E;��P�f0���u+m����N0-�������n|u컵��Х��`y��v��ݝ�.�s�%�:p�J�]���Eah:�B-X�u-kZ��[Z�nF�	Gm������y-۝�2�Ů����K�k�r2�+��]�j۫=���7Sz����3�������Yi=�<�dS�.�j�&������=�+# M'��l�<�pT����7W5W��y���&��r�l��n ]��=*��L�r�����v�:e���W,��X�JHݚ����y�=�\6~�ml\�0�=�9"���E|v]̄�=���Hspiv��!�ՏW��Z���/g(ڮUK#�h�������sk`s���~x��}&ν�(�R�x������Gv� ��ͭ�Z�	!	!4�"D�`�]*���}Ϻ��ـo��0��'�A7T�M�w�Ot�ـj瑀j呄z��A�x7Sz�;y��-$�ٿ����T粕~�w`|��]8��ٹ�������� ��# ��# ֓����`{��h��N�b��8�9̤�ݘ��%�:p���`n�{# 1&Wu]�n���&��n�4�o# ֓�%l�%��{� ����TRZ'*%T�c��P�"&F�t�=��T7����֒M�}����XFY%���t��-{Ε�)��%+�n����`y��Y*�8�AG)��kO�����o# ��=���`�%�`�&j��ɩ��ɼ���Ot��E�`{�ͭ��I�]�	����V�@�.2����t\��]�v*�2�ٮ��q��:�����!��Nڳ�Ͼ��3.��ml+���-��˩�yF��ު����Y[�L�3j(ۥ@^kw{�-6,��'>�W\�6��Jl��ڠ3�T8�������(�,l8w�3О�N����K[�j�=ݻ���|�A:�cS��$�0JJ@!����D������yw�B�)-�9U�ͻ�6�i��;��2���_��@!��ڧ�-�z�C7��V�uã�5���l<��1k6���b#>�������l�9$�4M��T6����3%Q���(�6�w6�Idd���nـ�ȗP\5K���ÕE���T��ٰ��{�Ҁ��~6�&���lB��p�����7˰1������PjQ9�ڠk�m�7Sz���w2�>^����;�Ҡ/[w`?Fĥ
!
"`J"6"'mw�܀��Y�3:��@,������-�y��}C6ő��ݐ��эtk\�@�/6�T�+o�ګ�KŘ��շ�2�ܑ��(	4��e.V����Bv���t\�	j�v��]Uv��敭F�5+��8u۶�QY�p)����<��m��ԝ�P��W�v��3g��E�e�{GmbR��ٶ2i'��vn=�91BD\]�ՠ���={��}�{q�;�gu�Ulf�&Ҝsh���䔰q��<�F�÷WA�A���[��!�*[M�߻���>�e*��n�%H��P���i�n��t��8}�������n�ڰ37�ɠ=�u� �_f!uqs�M\5W���	�s�wu������^O$u�MXFY%��Ɏp�f���7���)M�UF�r��J�{ۆ��}��fg8rf=�1k��Ps{հOOrAƝN�ɶ�fs,��N�I��ݎnE6䮭�8{������nE\t������6=����)��;ۆ���mzͱ
z�󪀼m���"b"�#����>���`w���9������o��7���t�_� ]��"�,�Soc@�e52+]����M�<�ۆ���{k �����`a	����&�,��4M�`�{�rv�ަ� ���Of:�m�����`�C��u�˕�Z�I��M9�jq�yu��w��;��u�E�WUU��~_�{@���MN��~猪g�`�]dՄe�[��?w�X��p�<�ϛ�"">��sq-�8�S`w��^���{kg��i.�iS�w�pA�e�`���"���M�9�;3$ro# ���@������$�����=�f&�ō�
�5q�{�7�'l�=�jp鞤�0��"�Ym�5-����KmaTnhٝg\��#�s�͒�s���� X�O�]���0ޖ�l�+Y y��pa�S&�vJ�i�d���L�آ"}��T��݁�}elB�=��;$�L���]��N�����7�*f���������EQ9U�RJ�"P}珗`{Y@}�M�P��
9舅��{ڵ@{�̝�9ޗ�������� ]��prY�ٙ� ���q�-���;&�VЖ]aWH�2+�g������G����Sof��Ix�wW5pMY�?u��ܖF ����-p�. �|�Dʘ�U֣{� ��F /4�@���`Pp���R��*������\6�_G��`�0�Q ��e�qR}pU���1)�0�h�#ܖF\ȟ7���Qc���-Ӷ�M����;��0���9;f�z;�_�ww33쐑�$�I$�KzBh��Z"&9�@��áz��e�с'����H��mS�kLHc�W������`�x�y��.t<C����^��CH��5p͌�fǇO2�6�e��m ���qG���⁰5�`H��!!,��$�07�����Dx�?t��]�z!�(��:8�x0G)��N��%��06���T$�&�H��#�J���d��iQYj)��-6�.����WOi�"�Y3:��v se������J8�2 �,�9��m��JD� )@9�m�L      ,1  l�M� ��iu�itic� m!�K�q�!%\�@0W4�f��C#�����v"Zx�,Q�+�q��Z�5g����MWn�s�c+yd�k��g�����q��[��;g[���}:z�2��2��i�m��Ļ;�-a6f&ٻ ���Nx�lTgv�/8�.�y4��r�Nwq>����m����
��b.��<=��e+^���.j�� }�`ݳ��+��f.��r���:vݱe���zL�,�k^�n�4���-�t����ŗ��9{:s�;j�[ZTB�g6�J0�\��!ja�Ӂu\WذYغ��s*	�>�]=;��l�f� m���I�f9�%�������-�q9H�8��f���rKYI�D�%�m�Q^j��9A�v��6�3I0�K��	-�qү[u �Ŵ�zJ6��j�8��x"SL�` �H5Ӧ�6�l���L86�K4t��d�Xx)&�����n���M���S��u���ɷMϟ7����ډv��g[m��n]��^յZ�s�hM�UUJ�*�v�X��6�d6e:dpR�ʫ؁���yJ�h:yv@�RuˁcEP���qA�o���'2*��)�\����%�ka�j��,i0v2�:؝�om���Z+k�d�n-'FE�7l�-a�Ą�m��p��d�ݲ�$�Y�5݇pڔyM=� ���}�\U���\�`0�H-�'K*��'4�����2�c$�t�u�pAŢU���I��I��Y7HM��h�:^�� n����۬u�T���*h�z�+vQ��dXm����(j��V�e�#$6�*SWv�ۆ��GN��W�४#��-�uq��2�[U��A9������׼�(Ӥ�`~ ��X]�i�?���M"?�%���qh�ߊz��rBÇ{�n����[33L�b彦I�[:7�:���YG������>
OU�Ǫx�6㜻#n�X�C���`A^,�m�zKVnp�۬[��l�'y�ku[(klGn �s�.q���ڥU��Ե����+�	���u��h�����2�ۧ&�^��,#8��t��;�������']�M8�Xʵ�n��<j$��������՞��@�͒�K����y��v�s�8zRwV���8t������"���6��-��w�g��IVD�]�sW�h	~���'����6w���zw�
�������l�{�rv���`�2>��	��KK� Ym���\6go���5���6���}�m��مQ��+��5f �֌ܖF@	4�@�>���s���KTc�WZ��8 �6�COtNف}h�+
��_^a�I�;k!5�,�s����,:��Z�Aۇ��(j��#-�B"�H!HR;\��c��n���0�р.�S��oB��n�U]���\6����-hIk�J)!y)J�@�ݢ��t����}��cϏ��"��j ��Jl��� =�^	~OtNـ&	ˢJ�J��E��n����a(�{��׷`w�p���6 �Ӿ�UE%TuZ]��	4�@���-�J�I��f��I�%c�B8ƪ�DanT�>6���a��Fx9@ݳ@=Xҵ�]P]]����0�р�>��=��� ��a,i�[er������+TDD)��7�&g���ԦA$������Ln�֠�E�g�]����~뫴�*A*D�"�8 �(n~���\���߷*�����!E+��-�-��s�w�p�u� =�^�R:�	����.�W�C�`���3@97x���gfe����%M؝R�F��u���.K���dS�iq0ІP[3��,��|���]�$M��Y�5֌��V �OtNـs7DQQd�]�sW�h8�+R��۱=��w
��^���j)*���m����p�o�p�-$g�o���>��`g�^XݒZ]Y��{۰�ǵ��:���g(������=��x�rcv]6�,�Tr�WZ0*c���\�`	�otNِs3%Q9�m�M5\��VG-�Q6��Wh1�f�ۑ����7U�'9@�����"��4��`	��@��� ~Jr0�@����	]��l�W�����DD��Ҁ��*���R����!��ٞO�;�݁��\(���Z�D7י�`f|}�8 �E��%'m�U�I``��`	��@I�0�}�����:V�廜�3&�5��m��3Y@9��*���J�Q-i|���/�}��m��BF�#��d�כ���޳l����]p힝sș��f7%b�3�ٶ6}=s=�e�F��ϗ��m1db��+�pa�s��\3�G�旕c��v+666G%[T��zRL�Q�Wh�0�6 ���Ƕ�G\���~��|�Y�8^�n|��i��3a�ulUԭۜp����˫����ћj{�]�����n=��u�x>�˗;�3�6K��8��ڬ�ٶ��#>�%n�����g$&o,����Ue������� ��ᰯ'��:��M����2I$�VB����bX��J �;-�P����3��� 4��مu6�l�Tr�fr��s3�L��۰��@�x��T��lkc�����`s33��ˆ�kZ�w�˰y��d�c���[ot���� ��� ��d��%vZՈE��V��r�&vֵ̤t����\��F�t]�˹�7�^6��{��w�$�������`�{�wT�(�nJN�%6��ܼ� :ie`�{�&�f��EE�^�f^�JV�����(v� �{�`�;�*�J�uTY^����HGS�`@wr�gܫ k�H�Y$���Em������I'���Ͼɰ9�fs��fJ����h�;u�M�T�`��k��!�Վ�k]�״��^�S�����e�J��Sm��{�`r~�r��w�$����(�,d�\�3E�La5w�zy:�5��@�r�l��]��%� fh�[ @��	;�P��vهYE+��l$�Z�"!Hb�� �h��4��{���*�<��l/˺�cP>n8�E�� ��\6�����g)���>������l𫙪��&���y��6}ʰ>ox���?k�y��	J�rF7e��c6�����Sƞr*f��sӇ�`$��ΧQsQV_׳�q�G���ϛ������{�]�.�{ E%U��\�(=>�uw��"d�>�@����}>������0Y�n�� +e���}p� ����N׹V��i���˚���%�J��Sa����$���.�_�}�`}�c�@֑\T�D+w��@庞D��[ݕڸ��e��s���V� ���Ǻ��]LUMՇ�p��[pݓ��;4�t��HUk����\�8�ܖ��6Żd�ev�6�糜~�0SW�{�`
=�3SQ7{�G�[1L����6}ʰsOt���	[��[T��=��:��֫ �sOtr�d���LTY3D�׹W9z������ܭ����e����UE%U��\�`~��{��g�� 55xϹV�_D}���S`��Ғ�6a�w{�_��{��n���1[T�[Ām�s��E�I�v�Ω��	�m��M��Y3\�u������F{�`1�ԁ˜p]I��ô���,�3�X��Y3�,sS	��]�nm��J��Wi.�;��.v��b�p�c�&G��S.L��������$eq�l<��랂���mHWRK���܋�
NLH�h���v���a���xw@��{�{��绿~�ﯿ?��@%���S�,���š8�`%�vm��nl�W6x{=�-�k[�GQX�-����� ���.����O䵮0�Y�8}�ϊ�le�J������x���`�i��V�9�׼�"��Z-�m��?vɰG&���l�M^ %
�QS\��UwX����{�l�M^�䴟{^d����b��pz�����l�M^��U����D�cێ���gu�Ez��Hq͉���d�ې�$��h��3�L�j�/;�u�6�l� �U`dﺰ>Y�o�рy{�G���s{���n�kX�����K��P��������x������/wkKZ�f5�YH��)*��J��u~�Hr�`���r��!�K���U�[����m s��8�w�`���g8��a]M��-�� jj�ޮN�_���#ܭ� �߮v?uʧ>zjK[/<3n3Y���n�qGps8ۖ���ܴ��������w�wz��� \�� �'�@�ߝ� f!���t�[6���� ���x�^��U�tzHJ��O�	�y���˰���?O�/���m�r�*���{���{����x�bL�j�	ʳ,��30����ul�����\F�ͣl�������W�5��j��`zD�N>�k%	��Aؐa1(� �p�
�G�BV�	4H����NZӽz����+����!gf�A��d�ĆG��JDx�BP�`��о��S �	}�I�A:�_A��0S���A8�q�3��=M�>�:x�ꤪ<CHz >.����QAQv�*8�*��}�9������^�:,p#�i�U�݇��w��ﳔ{[.�R�S>ǽ�=����WI�.��ʼ����2��� �'x �g��cK������i4(�B�A��'X���Nt�euQ�k�&�(Zs*���pZxUU-+uR�g ��3� ��e[ ��;�BQrǛ����$�&z��"份��� ��:&}<���=��ﰮ���ʁ�-� ���6|�`�{����a(u_I�$�de]���n��Ǻܝ�(��O�apc�]�h�E��EB�?:�uQw�}�~޵�Y6U��U� ������y'x ����������j�l�q5��I�Sэ�Grqmm�5�F�	��Αf�W6q`w,��M4�(dz��-� ?{�v ���ԕ�荐k���1����r��Gm�~Y�ZZH8��M��<w`f>��S'�A=Ӈ�y<;;y��zK� \��	��N�����t�B��i[���6~$����}���y�� ?<� �!+�{9@6��5���
�Ym� ?{�v�3�z�?{9AS�x��.��B�(BI�D-���{����;�-j�[�1�hԺ��`u�$niI�+E�	�v�
��$`�[q׆��^̋�����r�_L�H�RB��;J��Wi���:XF9�ku�V�+e�X���<�g@�X�͂N�v�h�Б��6^:��k�A�\s�,�vplPfW0���)wd�2��p<�e�x�y����d��v�܉9�1P@�au��Q*����U�7C	�<N�����w��{��}�✩4�&�˸�I�]4V�o:�&�u8��nLg�Ȧ����૛��	�n� k��L�=ʰ��=���]��GՌy�m1�WZݶ��s*" 3��\�ُ�<�~���b��RȜ��Ɯ���_g���{/ ��z�N��Q ��T�a7{�I�`�W�F�r��>��s�s�~��'��U��Q�v���`oW)�ܞh�'x���]���݇m��&W<m֬u�B�0ZzP�,ۦf���4�vꓞ�ͯ7����`<��w'�@I���� !{�D*���v�v݁����E�$�kA؇��+���*�W�����˽��}v~�f���5b�����y'kde��ʯ ]����a]M�e-��`;�v��׀.��@9'x�J��~�r(��쌫�� �n�ﾈ�]��$� 3��v�I.�6�i楲�S�%+M,�W\����d�t�.h9Â7㷗�����u,���l�[����� ｗ`�˰���`u~^L<�,�=PNR�nd9'x �W��^ ���>�#��x�H�:�
���gs�.�����:1CB	�*�t�B���f݀c����:�\�ӕe�W�w��M� ��� ��Ϲ��`/z�M
��� ��ﳜ>�N��7x�+�5�E4��^�I���b'n�ŘM�k/�
4u��������,n��VIy��� 7x����=�=<�q717wupIwx ���I^ ��� ;�eސ������-��ɻ�r{�	@���� 5G|yK"�����`{��s����<���^�}���γ.����b��Bj�r�p��]�L�Q��ڈ_ nl�h�7v������V�ՠ������]qn,`K]N�q�ث;1�ZY�fy�Z���`�.*n�z@��e��W�.��t!;�;��jR"KX������f]���� ���� !.�_qqt�A�v�w���`��q��ִ��o�t̻��fv7QX�$��l�u� n-���3���y�~�:���6��[*YM��;�v�fv��{��yfu��"�Ĉ\K����{��{�w�z�+��Vºnp��IAc�F�f�].��l^��i�r��7=m�"91�܎�.������X:�zI@nvc�M&��q�B�F��A�uF
�P=tM�˺x�n�M��6Sv��T�7��+�6�B�Ęn8��u	�U�nCub����/5�s �ӷ)��ڜ��z��ڇB���=)]����i��v+6	���O$f��ٚ���b�#��`	�;l�����U=���8��h�k��-�k��b�t�^{<5]����s���ﻱ^��s��l�_h��݀{3��
!+�7>��ٯh͕ȤRY	,���� 䭘 ���� �B�����&��@�Hf >n��������g����L�DѴ��e7�� {��w'�%l�2&��U�TՓ{�yz����=�9+�`�˰>�\&���ܒj��*s3��ݫ�^ͷsϨ�ۂ��q��xᲄ���I��UZ�J嗀g��s�����`�˰w޻;�`�K
�
��$����-�_S�((^��
#�P��	�/^̷��2{�~��қ"��f&����0�w�l�U�.��`�����?b{S@�$�]n[o ��� ]���[0�;���𢶪*��*��{�� 9+f y{.���6��֗��7>%�[�x���K}z�έ;\Ӣ�Jѥ�b�7M���st*�U n�T����/��?{�p�T�w�or{�&8��Eݓ1!u7V`�w�l�U�or{�ro$�9�se5u�y��zSu�o��pt�`a�*� i��=��˰����f{$�EUZ�)7u�o���$� =���ﾈ�RY6��?�	aShUE\r��� �ܝ��L�*�7ܞ�������):/K$N��-k�z�"6��-�sm�G/=;��������pt�Kv�*�ܝ�A�ܫ ��=� �N�t���v�]n�o ������ZҌ����o���;�5G@(�����ʺ�*���M�y'x~�#艑5�����76 ���a� >��r^p>Q3����7�Ͻ�����ARHIi4�Ĵ��K���w��m�Cv�1!qSwx �W�l�*�7ܝn�{�˰9����	J���KaJ�m�'V����E�z�v��>��W;Y�ͨ��&.��2�JN�����w��K\`{=�����&����R�K6���@=�� r�x;^�Y�&O�����
�
��������w�˰==ʰ���	Rwsq3WquW%����s��O'X;����trw��:��F�p�[����c}~�́��7���΀}ﳴ������� ���(�IU����"��t����(�0���޹��v*� �B�(��!�D0�T� TQ�TB��UIQM�� % H*2� �+"�����*���Ѐ��NJ�$��`JT9"�b�L�
�Ȋ *#���̪�ʪA ȴJ(
�B(�(� R"����("��PԪ�@ h��EG���߯� (* G�~��������%������/�a��� ��:_�H#����?��.�_��](/��4��]�)�����D��?w�r�           ��������������������P]�)�����x !0������'��;�������_���������AU���W���������*���?J �� �+�_�{�{�dhO�H��Q�������G� ��!�`����!������������PU�������_��������N�O�����s���O:�"�������1�
"�R�I
$
J�2�H @)$(��� �
$B�P�@)J�"�J��A
$� ��������B)*$#
$!
$����%  2
�0
A �!
$�*$
�)(0
@�B�(2�B*$� � �����@
A ��
L��B
HH)!*$*$
��*ʉ�*$ ��#
$@)J�$(��)2�@B�B�,��H)�R�D(�
K �0
C"$"� �
�*$� J� �B���H�����	�,�@�@�B��@B$��� 2���J2�@J�	"�$��J�K!����22HL�!HA HBK! �H�) !!"
�@$	*�H��$�JH���!"�!
�	H@�B@�B@	!	!!+ @�B@$�
$
����!	+(B@L����0$��A L%(P��H4#HD�B0BH
,$@���0
����(@H�����"�H+!��J	+!(B�	 H�@(�*�� ��� �@��!"�(J�(J) �"0��B�@��
�������d!$ȅ I J�$��$�0� �*��B��*J�$BJ
-I@JH��J��	,�@�+�$	�$�,!J 4� L$�)Ȱ��,
��"	(ʣȠB
°�"��H� C)0,H�2���JBL�$�2�L���"��(�(�
��0���0�  ����H���� 2� 0,#"2��*�,�((A�( Ȅ�����2!"�� 
B�H��� �@$
J2@��!"$�H+*)*�@��#H ����������O��UZQ�����A�~���M`���?��������"������ֽ���?�gi���Á֏����"
������� �W�~��������W� �*��?�=��EPU�����&���T_ס�y���s�zL�����ʀ?���O�k��ǣ��Z��u�v����F���������*��?�ڪ�A������?���
���{��*
��?������ѭ�f���H��;�����.��?/��\����y �*�+�+?����	�:?]Tv@�=��3�������k���APUxC���*9����W���v�����?�O��(+$�k0~=��ھ�0
 ?��d��0S�� �@��5�  	"%@P   T  gs(��� ��F��
�������)J��J$�P � � 

M IBF�u�@��PPP�))N̢�EP/      �{���  �C�@w�{��|O�o}��j�n�m}�Ҩ�Zk[�E�|�W��z�si9o�T����%���`�g�� ��uq��ހu�*�:qi��c���{����kq֫��9�v�g6U��vvގ:|��� �h�PS��e�﷔�y� ���M70 h��P `[h}�@��s6P ��u��4 ;��0   Z�(l  7Yr��l��; :{�ҁ̀�Zq�
w1�/w � iE,�R�s�4 ��B� ����RS����0�w7����\�����71�=w����w��}z|}{��:���  3��m�7T�wT=����͸ s��Ӽ��w7��� {�R���U�<�s�v���|{ �T� M4��;oI>�}���0�oCY�һt���xг>^���y{{<C��
�w@ͯ3�^l<�` �6S��;�=���v}�K�wc��x���,)@� �m�����Ӌ�8 � �@ϸ  < rπ����
̓����qovyJ�lr����t�=�۞Þ�� �rs�S��P�å��3��;�;��e;�Cl��vy{�=��=7`     D�M�)*D� �O��*0   D�*�EOy�ShF�`�������U4��5O�j�6�U(2 h��"B�� �➢}����_������R}����k���_����AU�(�*��AU�`AW�(*�DQO���?�
�(R�VP��]�m4�FI!�" D���F��fi��H$�	-�zx�Ѱ�sa��.��$B$"B����T�H]��O�m=`@� �&ݜ��Ǹ:xE�!$����Q��B�# ���C�C�i��L/<���I!0"B5outz�(�_WwSn�c�J�QIЅ�(J@�)�)-���3rsO�f��4�#�sTD��D`��t�����
��p#L��ZO7�l��<�M���!8Ł)�+
��n��Ja�y�s��|�F�$�K! D�H��^��A8B��������\eevp�$��M�g�,)#������t�$�����.ׂ@��,!���	��H�+yODy���H�ܜqbM$c��)�%/-�MA<��1a�/���8��$eaX�P��IHV�S2]j\�.B��(��f���S��e�;���L�Z��i��G��s��n�^�_��Ffl!��Ȑ"�r��e9|�-�79/<�5���nc�[���!3$,ּ�D�h�a���|y���5���m��3ї5R6
�I:y��O�5��q�o�uBe�>��7�xA~CߜS���I���#��k����RX��4��`vD�B��jJ)���R�2��8R��!�t���FF#�vGHH\�@��'�?����Xi)4��o�R߹����_>�)�^���O 7��t|z�~[����&s��9-�'5f��熹��=&x�!u��By�9����!�(�/7�5�,s���:I�����덐��͇���dH���e�����$,hB�i���t��$B��A��\��SI0	���� �Dh8���v�b$P�HHP�p) �$Vdl
)��Al�:��i)��J@��yLr���Ȯ�^p�N��Y���m^��k��,d��5��f������.�:)#>����o;�[�P�;����y�ߛ%�����ۚ�W�"b�Cy\#t�)�R�`�I	$L�-r+b��(h�ZJB�����1$k��S)8sy�g2���NW79�K���].�(m�$bP,"B�M���6R!~��}����g��v]_?��w�w��TQ9�@<tĐ��z�c�^?��;����a��§��&���sz̜_o/6ۢ��8*)q_���zn��)g3���rg>�~�]�[���뭥�e���v��-�|����ϖ�_NC��絖g{�U�����k�Mg�X1�
�bS����`�I]y�a��3�����ק��ߩ��S�����*��������
��Ŗ�yzi�T���ow������9�ҩP����]�Map�H��g$�7假��	<�>�|�/�֡�ѵ��
��J���b¬h�(B�(�

��
�H᠍X1�$#@@
b`���) B�
�`��F$[$K�(�b`m P����¡�J*�"D��a=��Y��=�<Rf�<757�{s\�)RC�I|��p�Ns$��s[�@���������)�V��O|��yL����$�Gp) �H	��r�<"�@Y�zz.�p2L����ɓ��>b�z����9�h����Jbݛ1�HZᬙ$&�ᐸ��. `�8;��&���f�l�57�y������p�]��Bȑ##��E�(D�R�+R��
R4
珱)��{�s�7�r� B�"���H��4a���_\�M�y���$��Ny�m
��� ͻ�v���3�U��;�2���T��T�ܕ���]��J��8R^0����)��$H1�K��ߑ���$H���%�qU4�_ww���v_ݡm���nK'��_{I!���.���v.�R�U!��;��n�߹߬�_�J�8U�H�e	Mp����S�s�z]�8{�n�h� ��L�_Z��|N'���H��_<�=��33Yy��S~_<���*w��J���/�0|3���_{���umfw�����ܫy_>}t_ՔR�t|�����o�$�3;��g�B��W��AYK�����U:X�&�mb8�߹L�<"F$c�<5�f����77,���~6B����FI$�JI�.L!`D��bB @�I*��$@"�`	@�� � �0(�(8�A$Y�	$��ņc�Ә����̆��I�1��V\UO2�T�~�]����E���ƌ]��HԜ�k��$��$6m(L�f}�"�p< ,	�<�L���I	�����|��e!NaM���@�()�-�\H��O�I��XH�@H$}�4�p�k�O���Z��H��+8�A���kF:�d��J� Le2IB�H��@��@�!c�A��܎�S�!%��`Jy�!sl��/	a���������lƳR���7S�׾S�m5���t�.2�&_ap$jk&u��̼��]0��n���������Z��x�L7�0
�j�"�`JI ��D���w�Ӆ*�u����k��\J��b/��.gm����߮�֯�[����mٟupY}���ky�߻\�I������ٛ�&C*GP������a�X�2���d�	&h�#@!�@�P�Xj�S$"��qSo�)w�vϯ���W�N�T��*��]T;w.>jut˗����s��
�E�#�(}����Kvx@%�<�.]��o�.�\�����<�=05�� �F��\,�]:�Mxo~6��ϼ�CbK=�*�3Fofi�!g7�޼XV\����4!r�D�H�ԁK��D����T�d�W�1 �p��p%XЈ@�4F�H$!��`aR,�Q�Ƅk(c�)"��!���"�1b�r2@�ł�`�ȬXE��	0��ҙ�!$��cR6H�Ӛ�i�H@�'�!�RC�h��d
11�
�R,
�J�RbS�l)��~o3^捤Mf�9��K�	������e�˽R��FXҘP�)�6ߕs�CP����e�&��-�ݳ�s�y����I	8p�Y���9�Þ�SG�xa�i/5��ādߪB��ގa�y��aS�d�8��B�o{��|=7wy�e8R���z]|�;�ܛ�w��ܮ������'�Uc�N�jy����s�N_~Y�_X��g�Ӭ|�S%��P��47$H�3�F�K�V�՚h�[��P�V�eZ�v���Y��Ia�ީ��F1�q�ƅ�l�bl4�54Y)5$a�0aG5jS<4���"�B0"���ZDJ�  ������'�3�	|��<p4m�!F�B�-��
�:�|�A��xT�n�KĂ�sLk+�d�i۳����b1 A"����=H�y��N��O�E��Y,HX)BZ��|l> �6���,c!$dB�����|`D��r�

��Y�X���,T8'�8Bs^N���$Í�l�oz=�\ɳЬB9�)��ON`i�vd��0�Cn���6����7gƍ����<���f���2_8s'>�Jg�)�y���D�.�B� X�H�Q���$crHP1�����+���~�f���8s�.�S��6gm]K��o��Uu����=y����yE���9��K?��3���9NR_,����++��� ���!R WjJa��D�F!t�
8�ji^3n{'�o�}����������G��{ͬ�OW����@;�����Ӣ��w��D���K;_(�K�v�(N��N%2���\��s/y�8�e��f�#�j�h!e���Ox{�򏇥l���ʢ���_Uw+x0��)�T���O�$�����x
��Ea�aj�¬��J�$���|N9:� �&p<><<!�C̻rM+++>�џ^gw�J�w±�	�!��ݛ�4�B:1�.���hB�ZF� l`��`�rS!��H�H�B4�B»e�l�ċѹ#B,X��@q#B$`"�� ��pH1�AX$HذH�%X�R11�R.�BYxa�c�5�-JT�sY޸��y������zs�s���<-�����޴�(�Aii�N>=B$�o�>{���G�&�E�*a˷�"}
��Yݬu�����R|'�U����4��!o�+�wکCda D�A�������T��x&�!����V��s{d�p!L`@NH�HE��$ѳ$���K��7<�ngqt�! D,da A�I LD�a��4®&�i@*�E���~O�  �   �                               m �   �p �   �         � ��   e�      �sn�mv�(J�2����"��@�Z�,F��nP�?�l����h^ݰ�m������u뜃d����S̮˺��[�r	鄖��RP$ �gj��l�m���U]�V�7c���T
5�\�
�Z�c��XbJ��ro�@����}�c|���AU[@-�-uʹ"ʕ�jn���Tڝ����m^k]kW��
ܐ'.c��ޠ�s��\g �|khr9���Xű½�����LcS9�^i0�n�u�� �f��2D�6[xvݭ��h�	F�m����z�oi7e����6�ꪕ�U���  ��j���Bj��6�s� :�m���Rl ���@ %�% ����f�i>|85��ە5�$��ö�[N-�۰6Ѭ��mm9�Ą�C잎t)�8@�(��5�M&On�XV��n8^&��v��6��6�96�U�z8�emmK���m��偫jX���n�ai��9����}��T�egz�fvZ��^}>�kX�ɏ6F��u�m��+�mu��H�6�)�ru�b��Z`l�WGWT|�9���Q�[Z�vDIe��7V,	�*���;������\�z�1v�	��4[mҞTz���h�nAݻ����UuR��^��ȔJs�-']R�:I���d����.[4����EU�6 e���t�5�� �AJZ��,�V�t�b�8v�L�=v��ݟ��r�A��UJ���v^	ꖥ�lnٯk(ݻ`p�N�ԩt��� �Uڪ�t��$AUT�N�t��6�m�M�ڧEs	�+H>+��I�iҲ-ZL�T�jUU:W���Gf?}�}�/o���춎�Cv�d��\�@Uʀ�E)����6�v�iی�\<�jڪU���U�Q��%���� �6Kd����]��\:\ʷ]��c��x��$��2k���Dνg/H�UPR��0� zKeS��v�D��ݶ۶  �|S�cu�����-�mϤ ����Z���Ⱥti�ʼ��T� ^X�#�m�����m�T���bv;��l���Pͫ���7��m�)���s��K��In���:E���8r�e�8���C�&�r�½�1l�ι՘H��mjI-�5[K�ʇ!�^�Jd�,ù$i��jI�,����7��F3*�ic�]m��Ԁ� �KQٸ�n�ݢi2���jm�E��B�ҙ8L�j�"dv�.��'0\i��%^���;����춝�z�ŵV�`z�4�Nv�*�']p��bu�pY��ro^�ۭ�ە�U�uI��;U�L.X�˱��v3ųK�C����:+�/˴ݛ=�����0bL�Sg�����e���*�<�n�"6rF��]����۵YU��N�Ûl	D�+t��bY����m� ��@,����!@l� kj�շOS�d�M+ʠ mmd,�D�-n�n�[��&�  ۷��w�w��v�m�.�-�F�d6[[�GV(�c�ջj���l�� �ce�B�Z��ݦ98�UvZ�ګm�[@� �� ,�n�%��<I�yl�,�1e�sm�YD�����Ѻf ]$�7���m��m�-��`8�x���-� Zl�   $ m��  ���aiU��8$ ��]t��I۸��I��pf���:���m��H�h8@6ͱm h� [M�l 6ӛY��-�f�`,�����8� �m [e�       �H2I�m�[@����U��e�#��K��m��mB��2�-����K����9mH  UUmOcp�	�@@�- m�h�m�8[@	�d�M� 	��mm m�-� m��m� ��ݶ[d�  ӤΊY4Z�m�!m  m�H�8�{D�� Ѷ�$�į����B�� � ��٢�m�m�� �P����\���`x�` $m����    �[@ p�j�|l 6ZA�$��
ݞiUT
���(i�[[l��v 	m�i�e�8�8 �`�`��m ��[kY�[f�eT�W ���� � 	�  �m��m�k���n$�֖�=.�ܴ��m�#m��	�i,K�T�z����А 	 �   km�6�m   U�k �UP)�@ee���d�i�l�%��	$ٵ�m��iؖ\ [�   �h�m�[l� l�P  H 6�  h � �m � | �m�������e�]�����`4U�m�@M�hm��h)=2�ɸr9#6ؑ�,�� ��       M����n׶��Pq��kY6����f�K��m-�    hH     m��`pk��d��Z��˦�,븶�# � m��DFF���G���Lݮ��c��-�   
UK9u��ו�n���Q�N�p�`4vn�ڶN/��V���Y�v�X����!��*�k��k\n�q5��u���R�ӆ����J���&���^Wʹ���I��n1��J��W��{�r�&؎�]*m��a��RqK��i�cxv��^�)]���`*��m���̭V1<[�������WJ�ԫ�@]S��/�j��^���^AV�
�j˰�H��]��z�[m&X6�۵l�p6Z	�mzu�4������l*դ~��W����z��ۦ�n	$���ܐ^���.@��pm-k+t%���� ��Y���]�^�j��V�F��� �^�Y׈d�[
�%^vݬ
����Mp�r{p�l�⫆�+�9by��ڢ������{��yV2�.��9��W�uR�{�Z�Ę$:�,�H6�oI��/1bD�7��j������C˹n}��[�mq=rCt/]Z��n7F�9l�����)|f�ƀ��ǈQ��Z��3���5��<(r�X�6ċ��#v�ì�*+bvܕ�[���;v➄��nd�nvc�������w]���E�]���ݫ��K3lL��.m�q�c� ���3��+�tC�u�� ���Y�ٴ�t�J���Z��Ě�� Ui1
�t�⦎Ll��	-rIpn��Y�$K�e1F6�V�ca��Ss�l�.�v� $�m��k�E�*�
�1�P��`9%�k����a�  6�ېI��l{��p5��� Z��� �/��n��l�e�0$��MI�a�pA�"ہ�:u_OK]�% ������� �[l� q�5Q�6+e�+�s�f�D�rK��v��͖WL��8Ë��
��'��C����pu�G>n`ڪ��kx�[M�  m��`p6ʹ�hh��]�ꪩ]��cV�l��nl�� ��~�| l m� � ְ8һ0�l�iV���`��p�/nJ��am �^�&�i�M���[\�Y@�Nr�;m ��|����kX
Pll-�VU
� �/R���)l���"���) 8������I�ky��k��`6ʹ�m�a�i7H��  4��۷6m�8��[���m"�.���f�(�DH��6�[@&�8�Ͷ �����hԒ �@Zl�(m�����#m�m�G��KBT
�����@�)m���` �	 �g;m��6�$  �m�f�%��h�:C6U[�$q�m��ܻK�kd�d4!e��MUuR�����PR�G9a�N����mz�� UK�r�+HW+u8�(\BL�JKA�2�UuJ�lml\-�h��M�q��>���&t޴$�(�U]U 5Ul�Uv�i�UaŴ��[n�]$J���f׭Ʃ�j��P�V��J��P d $�e�fI��[N��l�-�Z�[DUUAUYÓ�'	hHLg)<�UmC��Z��d�:h��-z��ʬ$ q�T��[P2�v5V]�m�/C$	;+R�QU�ԙ�U]k��	{K��,7m��mm�  �u��ڶ��Z �g-�K������;4RV�啒@�z�qJ�lɝ����8h8[�  �Ͷ����E��g -�� ��6ݶ�$۴��ݶ ��l�cJ�q�Hi`��U�Z��/Zs��� �]mNu� [m��l�� 9$����ݣ�Πn�2��*�Qe�R�XL����vH[C$��w,4�r� �>4�d��X�v� &�+
�8-��� ��b��`  6��j����mí����d��PZ��kb�h  ���ReW���>�U^���!õ�l$� �n�P �T���b	0˶iegH��8HH  -M%$8Hh���km���m�khI�Ć@�a�r�����6���{���{��{�͢?�N1|Tj@�+E��)�(� �@	6cHB�!����X ��N�TW$xma6b�@؋�,����)�!  ���*�~Q��Q*��ئ��� <P4&���>Gg&�v��`�4	h@�� FT��"H ���
"A��c�v�����|O<@� �|@LQ��h/�q:S�'���_^���(�H�"( ���:D�A����	�ɛb	�R`�@)� �A$����6 <C[E���a��==C�~j���LA�£���P���k �a�����<(|EW��aGN��B��⃤O=��{d6�����=��� ������&���Db���1B1 ��F)�>U��"*� ���h��� `�����~�����抉�H؉`0T�N>���Q�TOb�"+觀pT��ILEb/��� S�S�Z1h�>�bz �TB����Gd< ��"�H���P�Ab(�6�5 � Hx�C�t&�| OQ��>Y�,$E�W���%
�X��!i|�}S�P�8>��A]�i]������� 6���|�!-%��UI(J�)JB1,���Vح)(�JDI,�X@�BYb�- ��R$!`(�#BY)K)�!H B��QP�),I=!=G��|4;���$�c	B!$H�Fm�C�a��8��B F���S�0��|BA�#��$��6�%hUt�l@�dZ����i0M#�G^O�Ux���4�& Q�0`�@����21
 ��
@2�T �!I
��y���      �I�.Q�� 	 �h7d4�J-�ZJ4sG��L\6X�M�)v*f�W�P�;��{��u�u���ձ��"�n�sm�c�2�젯4���Ej:O2��=�7'C�����W�m�J�mܥ�h�����^{��͈<,U��)�`h2�7���	�)�(���5����Ws�@r%�P{#WR�m�l�Ƕ�ŷ����*�2K��n�Z]���L�N��M�밼#+L&m&�KR�<	kl��:�њYP�͸_l��s��'a��q,��;�쾮#��fi����e�1#[C��b��]�]F���<+�mRch�>-��,��]��;F�[��&�f��ƶ.^S��m�� %H.�mJ�ܜ����]��%�+872�YI3VVv^�NȬ��\�x���o]�Ӱ#�Pe���X�^:U]�uէ�p.ŶZX� �I@+[�n�:���N8�UX)]����&�d�u�gE(v�x;16$a���@2.� �9ҸԭU@UR�e��k�k��Y���X���
�	��2q���8:����ۋ���;f.Ӎ�1���Q�#���Zʀ��e3܎�܀�8�A��6�Mlrݵ��l �}Z1�{�,��n,�%۷:�9���y�������Rױm��-���m�;a�1�ح�
;1h�5�������T�[� �F�<�nQY{(*S�:l�L�1z��J�YՀ�V�s�lᐴU��K�B<�L�uu@T����]eZU��٠c��[j�ݝ����]S �k
b0�d��Wj�	�o\�<v�뇤e&Pc`��B��qmѱ��Y�%p[��+	p�,k0[*�٥6tl�y�t&���q��=`}r��U�k;=vq�*���g"۠��J�t���i��`���Ks���V��,А���b�l\��݅�Tg�ڲ�V�)��e�s-�v��[kDn��΅����0P� ~Q�"��� h�
�O� ��0A� ��)���A� |E�6=��y���s�3�ԅ��a)X��;m4�cFP�.��slT��+��Y9��h��K�kt\E���=h��I���upa�����,��g''i�mz�tt��d���hN{: �Mڴ�z�@��<0S��:Yq1DX�L�;��Dp�|v��t���ܽ�NЛ�0�7n���iVܜ��%]e֝ (r�ȍ/��;��Ͻ����/"�n� ���e�&��p�=�ݑ۞�0��st��N�U�)#����߻z��;�<�ǧ�M�:MZh(������=��`�X]���+n��n!PƮ� �ۆ�{v< ���젫�$SN��eݘ��X]��]��	ݸ`Z=�F4��]�Zn�`wc��e��p�>ױ`�r�{T~c��Z�����byy/a�T�j��g5��۴���e9��|`ɇ��m��e���ZI���z�	ݸ`kذ�#�;��v�[wjՍ�WorO��_M��6\B�ՂJ�]9ʜ�r���B��� ��ǀn��:��B�v�-��eݘ��,.�x{�uI�{e��5t�I��V��c�'v����-��	ݸ`{��.y`��BuwV�V�
-]��7n�I�+ĒQ�G��%�{����{^ܚ�=7#�>+BX��D�c:X��i�*E�n�n&]	a�Hhe��I/I�>�$�{�I(�#����$��e>cE4�v]���$kدIG��$�\��I%7r}�q��P�o��6X1�������o} ���ٻx�Q"s���0TL�3'����$u�W�$������*Ʃ���|�]rc1$)����Z�[Ē]������۽�j;(��af� ���I%�e�I%d|�]Re<I%�~��k��[�A�9L�iA�E���Øш6�ۇi�����ե��[����En����$�췉$���K�L��$w��������فQ�rS+�߳�~�s�
�fY�{�[���~�g9m����x �~�,vŲ��} K�]�I)��}��)�����$���?�I)���2��I��$��܇�%l�>��v�~�=�9�i�ǁ�H�T(��_ �?w��uŘͥ��� G"�I%�����$���I|����I}!���4�r�6���Z���NX�6�|�����Q��u/c��g�x���Z�F��@�~��� �z� ��{���9޴���+Ē[R�Ճ�ĩ�j���{�� �߻��wz� ��z�����ͫ���| :�G��$����s���޿�I!{�w����ݥ���h9���NI6~���$���_�$����$�^���$�k����չ0e| �����Ϡ�߾�� �W����䳛����a�t���f56�<�5�r:���T�l�B���c:*f��#���Io'j2�{6���v�o0�cvb����Xl38��-�v����J�dwF��m#kH<��<r�Z�x��:�uV��]��p�w���kh��H�J�LKH��x�f���\��S����a�9�{b���{\���1+V�$��X\�������{�����䵛�%k���Э6�Cih�����)^ubըЅdBR�PL[����g�����} �]�I%�%��IH2�P�P&�I7n�$������r�i)�]��K}�_�$�?w�� ~����������@*��I%�%��I%�]�I-{#�����n�6Xhֆs�s������}|�I{޻ĒZ�G��$)#�I��S��Sh,���I
H�I-�/>I!I�I%�%��%��9U��#�S&��aԗjp��r�Fh5�Oj�Oi���@��E�=��3t�RQQ������HRGx�IvI~��Wz�I{�_ ݭ�ԣlW/��S��k<��k�5C��nHlt��/<M���k-��y�r�o�޻� ���}��rm��{}0���Ƀ9� ?}�Ͼ���� ?~�_} �{�� �/��]�1lnW�@�s�������I$����HRGx�Ivw���w�β�n�$��S� ��K����I.�/�IIr�$����B��E3MUI�a����Ֆ`!�˱g&؅m���{<�n؄L� ���{�(�����޽������zP��Vn�fխ�����$�.�$�����$���I{��{<�wX�6-fVy���S��{�پ\�0�D�����u<�>�> ��}���Ϳv9�n\�ئU�$�����I)%�$��I�}�I.����ݥr�M�U}� ?w��I/��W�$�%��$���|�Dt�V^ee��+)yF٨��3��=��n�7���GM&N̸��p7R�f�6+�I}$���$�.�$�����$�O�����{�Gb�3�@/z��y���z��$�{�W�$��}_|�RL��wbL�!�/I.����$� w��} ���� ���Z.r]M�����ｏ��~������[��C����c�؂m�UWs=���9m��h��[�e�V�� w��} �����ޗ�$�����v;Ē]ۡ*TDۉQx��][Ti���B��[��aT3hF�iA,�#*[]f\GY�Y��} ����bI%��|�B��x�K�������F-ˑ�\.� ����} ����$��d���$�ɌĒ]�͂.��l�w��S�{� w��} ;��� ���w��~����g-��q��$��fC�II2�I%׻�$���| ��.ݶ8��}� �{�bI/Um��ޤ���;Ē_l�}�Ij��YbH0��	 �`��r�UK���l�j���lΰ�1P����̺�u�o]��2�[m#\�iGJݞ!��M	t3:�,��ZQ���l2�A�t�tlՃ)]&�kڊV����l�-�Rx]�H�jwd�T����͐tj�IQ� JbR/�79�8]������6s�s����p%N���jp�b�IgR���OlV�&ݧ5`�!F��+����������ӓ�I�<�?���m�X��:[i�`p(��1�mM��]������lu����[t���[��[�����﷾�S��| >ِ��RL�I-�ȋ.��c�P{�;�������@��7��~��������,ڵ9�}�!��$��fܤ�I����(���,e��Eӻ� �&Vջ M���\0���n���v�U��wXV�x6K�>�p�6I��n�wY��E�.�͡bl�4L���/m��O����Fi䳰��%�.�lj�=0����$��d�^�+���5I��>��e��]��fi�^��^����A�A�`@|X��P E؆ &�BO��6nI��߳rI��K����Um+M�0�e`[���/ �e� �l��+�j��j����I/ �e� �&V o6Kj��v�'V�+��d��I2����r�l�ׇE����F�\r����vԡj]k��9�CtkuƱd�2ɇF;mvY�cn����|`�2����we�"P)�e�l��t���>�2����{��/�����9�~�}���U#����������=�[��S�xsBCA�e^�L=�7�� ��0o�m82x>��@�ăPĔf��C���=ñ����=6��N�8B�%1�|0���K`�x�x�[�*��I<s3�s[�ZDC�p�J\���$���$�0a�ۄ0�����zˣd�kh���|��dH���5~{<�qǐ��֎yb2x<9�s[���n�K�چ�g�dd�|u��㨐�J���ww�[2kZX,�O�oɼ'.�^p��5瀌��9���P0�8��0�ks�7u������D!�f��a�;!�ӯ������V\�ɰP���!�߁| �BO�7�0aV%����on���.����F*���`+��)�a���� ����T�@4 xz�ZD�D�M�8���H� �6*@��6�U��:Pk�������L��3`��IZ�i�m]�vL��n̬s�����ߞ���I����ݎ��m]��ˆ�W==��5I�M�+ �ʪ��'���wI�N��s�X�n���Y��앋tۄ�ݗ�T�9q�Z?r�KBfr�V�'vt	����v<vL�ܮ~�s�7߯�l�R�F���(T]�`[��ĉ=�����;��s���'�6����2�إъ��x���V�ˆ�q-��V��^�������,ٱ5Y��<����vnI�����<�=��L> i*ᠫD�B#F	��8�B�R k��	���?{������wX]%l�;�wfݓ+ ��r��_���{���۫�>�N���v��m;��Ά��1� ��TMl���G�;p۝J(<N��9�2�˛���}߾���2���{������6�wV�v�6����7d��r�;�_�g���o���~�O�l}�7�]�.�S37j��o����;$���IH�'������*�V��N���R�{�V#�X�X���{<`��FvZ�wX�ذܪ�+�s߿~�t����2��ݮ�
TQ��ݖ��71�3h�@����hhX�4���:��h4���N�
�M��<�ۮƼ�Ѯ��Y���n�ۛ�F�az�j�Į�b�PJ��;j�v��/<�@ld<9`�^�y�V/e�zԧR�ugM�3�ߏw��|��G�E�t6S�N-JT}lu��@6���=rM
3
U�����51�>9twE��պ��K�jճ.h�h�;�����T�0E��hc�Y��f��I�O�����J�v�W�rnJ�5������EEإє*߀o�~��>��l�+��|�G<�V�ǂ�M��n�X;��>���'��G<��eg�UID
���;J�M���ـI�e`�b����_������' �����?�&�YQ�e͎֬�z��Is� ������`z���=�}X�1��Ʒ5�h��������~�9��߾�t~��+ �{��A��-��8�Pk������S�n�<On(�㎶0�k����{�{��ԳY��;����� �&V��/ܮr�s�U]a�߿e`�!?ȫiZh8�ـl���zqB����j�5�WZ����n��X�\3�+���U\l������;T6+wX���l�+߫�o}���~���[�۲�m�I�ҡ]�UqO{�V���l�+��-�=x��ߴu�e�6!�p�z���������'��L��9�U-��Z4Y-�pr����\���c�ݺ�x����l>0d����ukn�e�p���΁�߿e`[��$��*����Γ}�ѫ�bm�����w>�䤉�{+ ����7d��W)#i��]�۵i�V�����x�.��j��f���Z�ִL�k>E>��k����){{���5I�wi�	�-�wc�v��������O{�XV�x�W��� 7�=�;.��t�
N��6I��{��9�O?�'���>�p�?s�P�ݦ,ˣHME��m.�[���gA��[�¢S�A�s��lΩ5�cq?I䑡3��N�	���@����d��}���Ur�� ����T�c���N��%v�d�����Wꪮr�7߯�{���XO߻��I�r���}�\e�$@���_�d�X{��)/G�, ��� ��Z�VR��.�ݘ�����`�;۹$�����<_�Ch�A�dW�cDB���:Gj;T����f�����h�j��X�Wu�Mr,�\�Sޯ_�yOy�d��?y�?&�X��c��5bux_a�g��bm�6x��ڷ7$�a�s \@j�h�Ӓrk8^RqJ������������	�e{����=��	�r��*��m;�hi�����Us��U\��������� 'eK�s��A؃�T��I]&��ݼ�=��Mr,?W9���q���~x�����=�'��
�3gCi\�P/~�{w$�{��nI���r~TOȆo�~�`��E'��ƊN����ݩx�s�_��W���Ϡl��+ �dxW�y�Kd�y���U[�nd��h��m��E�5d�p��q�'S��O���6�7$�YRL{��u�7nDz���T���b��t����qP3�o3@^U�HEkK�_b|Q�;N�wd�պ[ b1�r2��M+�F�[�֨�u�t�P	Ǝl���\�!ӪtnΤ��Stk�<6��vz#lݷ%gg��lFr�H�y�v�����s�Ir��wt����=��?�����1X��F�aHC Th�5qn��N��)X�Xml �b�4�O��+旈��n�7j�$��y~���d��"������+׀y
��YJ�Sh�N��vL�����r�?/~��OW��oO����s������ʤnnZ�<����ڗ���ļ���ｕ�|�����We.Юw����O<۽�_� �����>�X�+���=�IO�_�;k��k���{��>��|�����{� ;�K�>��7MYc�R5jj���m�x���ې��ϗ�7.]!�Z����I�s���JM�b�����=��E�< ��K�*�U_ ���6=F;���I_��-�����=%a#%1���<B\d5dad�hD����03q� X
h�P��.)��$&x�A���� ro�Ou�'�{� ��eg���W	R!�6:But�N� l�� �dxz�UUIw}��{� ����V�Ui'Wx�*����ｕ�E$x�9\�%$^�Ȕ���vE�wo ��e`���9��~�߿>�{�_� �H��J�6��q'�v\v���"N�Db4�a}��1� h�MPG��I����;#�uI�]��y{�x��^���\�>A���pe>��}R�)v����޼����S2~��~��=��훒}~���UKgҟ�^�;�VӺv�ڻ�<��<�f�W����@��F�(l#30X�-@��=� y���9� �߷��~_`vY��e�#�p>��|���'o{�ܒy��nN�%�w�x½��L���%t�;�)#�=U\➋��^��7fV�^�D�p�I�j���7\�ܫ�r:Jݱ�-*qX�W-��	�E�7e��fL,�h�7k�	�xRG�Mٕ�U|��~��7x��$��v��m]�I~Ȏd���ٹ'����ܒ{���o��������
mIݼ}=��H�Y?(��2~���[�~��~��8ߏ~5�]\�AY�I�rC<�߾���$���ٹ6kA"�1�D����@�N�ٽ���5�n��``�WH�J�N�������H�^��v&���	5K�=�s��y���=��H�X��%����C��^�v�CT�э�s���.x�,���L���]��$�#��Jy��32S5w�^��6L�G"�9UU�W�	�/^ MR�Ԙ�AV��6L7�EQ�w����'���$���پ�2r��>��0b�fym���ǀ"������R^^����e`��6�liK�.�7��y����O&�~���~���d���U�s�r���g�� ���?�V�Ai����� �_��r���~�tߟ�� 6E/ �S��UQU6�
���	��o�B���Qߞyb��C���˰�	B6#�,I#B�#a) Kd�Bu�̮d�e���F\���y�T��X�#��utHq	fY�`�'5�! M`���$�$&�����`�!�t5J@��Y�b}�%ڦ ��dU�BR��H��0dB	��<�">���$�Ie%��$e�Cp$�&�$ B�O|�糜���y���TUUUT   m&��i6  [@��q�N�k�Z��Ny�]�L�r��<=uַ���zZ��U�Ǧ# �p�1Í��Hm�F��{"1��Ar���Λ=25����L�niҝ�g���Ȏ��z=,�<��\�ۀZz���l-���'=W���(L��;�Nս��$c�ۖ�'6ѻ�ݞY�]���zG-�����|k�T9:�"Nvi:]�u8�������:�pA�%�=%������>�{$f��|���DQ�u�XlP�۔�|�嬦*��[t�(dH�JLB�gD�ԗivƖHHâ�E��]+���"M�e�<e���U�r���g� ��X.s����_	�E69��/l[p�`Z��!�<��P�ɩ�a���̪9S|}���J�啕S!���u�wk���@�X'DFPaבctmS�6v�)�k�VH�H�UYh�K��9��ڣ\h��WTr�IO�(ܐv��O+J6E��u���\��^)V��4�j�VV��Q�'n�x�dͰ�SI�ݢ�Bj�3l�R)e�P���ҵnKb�n�������HEg>��η=�����3��Ť�Ɓ�W/����6��\�G���5��%��ܩ��gHkq�l�S��{cf�]7�˚�F9%���s`gR�d$4���)�l�V�$�pd��O@l�(�͏
�v���V%��8*%�e�A)Zkv�l;� ��J�ˢ�keV.Zrs����P�J��P�����g�cBuN7!m/l�mn�'��( o��T� �����hΥ�K<�׮����5Y�'�����1s��"�q�������y��� jè�ۚAV6�<���[+$@�]��`�upr5��	*���7۵[���'[M��R��HZvm��)-v��sv
Й3v#��PX@���B!MHAB:�+-�&�j�T��y��~��~M��\R��j�L�\q8.�{�SJ�WB���*`�P�"�v�DO� ب��R���>��E<E�Cࠔ�<39�kX[&�լf���ͮ��;��ŋ�f5�/
1%����1T���/�s8-7%�]j2�^:�-�v8�t�M�7u3Xù�Y�e�e��@���ha���UV�3`�\�*����6�����#7Q�r��,�ٞ;ob��GW�嵴��WP��G%�@��{b�ƴ\��ٌ�ޣV۞Nx.K\ s�.l�dw���]f��q?
���[d�Vg3	������T�-;���M4V �5�b,���l�aI$�3q<�j2���}���X�E�"��W9U_ ����>�rs};�v���6he�r{y�^B�{���9�1L��,K����[ND�,K�~��6��bX�'��xm9'$�!y�^O�_�K7�Zm-�r%�bX����bX�'s��m9�Q�,O{���r%�bX���>�r{y�^B�}�{)��fIs.���K��;��siȖ%�b}�{�iȖ%�bw��fӑ,KRĿ}��m9ı,K���N��h�t\��k6��bX�'��xm9ı,C��{v��bX�%����iȖ%�bw;��ӑ,K��l��.W�u�=�q\ŞD���m�Y웳&���O�'�[����$�>��˨�.��h�r%�bX�w���r%�bX�߻{��"X�%��w�͇� '�2%�bw���6��bX�%���3?��Yp�f\��r%�bX�߻{��!�I�М~AJ0���Őȉ"���R0bI��I��N���lC�FD�%����fӑ,K�����ӑ,K����fӑ?A2&D�=���~����D��˭m9ı,N��߳iȖ%�b}���ӑ,lK��}�ND�,K��ou��Kı>Ϭ��;��֤.Y�浛ND�,U,O����r%�bX�w���r%�bX����[ND�,�G"w_�~ͧ"X��������;Eɐl�<�����b}��iȖ%�`~�{5��Kı>�����Kı>����Ky�^N����,8�0Ƃ�iu�˫0�0��*mY]��@ǚ�WZ�&T��I$bs�7���C�����^B����}_�,K��;��ӑ,K���w����<��,K��o��r%�b��G�O�s��fd��|�����b}��si�bX�'���6��bX�'��xm9ı,K�{٭�"~��"X��ײ��4d�.Yf��ND�,K�~��iȖ%�b}���ӑ,j����M�D�K��ɭ�"X�%��w�ͧ"X�%���I�=���t��9=���/�I AL��߿xm9ı,K�߿Mm9ı,O���m9İ"[���y8y y�;;���)X�j���H����I�$�>߾�6��bX�'����r%�bX�w���Kı����K.�� �Ķ��e����-��f䇸a�u�7X�vs]��������yv��njkiȖ%�b}��siȖ%�b}߻ͧ"X�%�~�{��r%�bX����[ND�,K���>3���R,�sZͧ"X�%����6��%�b_���iȖ%�b_{��m9ı,O���m9�,Kק�30�W5n��5��r%�bX�����r%�bX����[ND�[��;��ӑ,K���w�ND�,K�'O��5��Դ�Zֶ��bY�X!�3�w��ӑ,K��?~��ND�,K���m9İ?/T"�*��
8
����p@=BD�o�����B����~��S��2���q���r%�bX��{��r%�bX~ /߻��i�Kı/{�����bX�'����iȖ%�b}�ݙtff��d��4�ј��!3GB���0����yyur�Ǭ���n<��y��gX0ű˼���,K���ND�,K��{��"X�%���vp�"X�%��w�ͧ'!y�^O�������� �y���bX�%���[NC� ș����8m9ı,O���ٴ�Kı=����ı,K���v�5�]-��kiȖ%�b}�ݜ6��bX�'���6��b6%��~��"X�%�~�{��"X�%��]7���Y�]ԚѣiȖ%��'���6��bX�'���6��bX�%���bX!b}�ݜ6��bX�'���|\�GY!r�5��r%�bX�����r%�bX~U"��߿ki�Kı=����"X�%��w�ͧ"X�%��H0d�	K(��(����kY�ə��`u�M��q��;�8��{�0���ۧ�9�g+��b�u��	(�u���3&2���۸0�egd�5$�t�J0�e-�2&.S1�N
��>յ���5�se�n�HId3�!{n׊qt�V��{q�����&���^�q5��g8��h"9�R�2��)5�D�p��!Oprm���ykB��KE�C���m�l�jf��5����1_G�Sɛ��&��<�Yj�b���7�� A`Uxn�n��dxC��Ԣ�'��כ��^�-̔m9ı,K����ӑ,K������Kı>����9ı,O~��6��bX�'�N�KL:kS3R[&kZ�r%�bX�}ޜ6��bX�'���6��bX�'�}�ND�,K���>r{g8^B���c���S+�̆kF��"X�%��w�ͧ"X�%���w�ӑ,�,K�{�m9ı,O>�NND�,K��|ޘfi�.Yf��ND�,Q�=����r%�bX�����r%�bX�}ޜ6��bX�b}��siȖ%�by�t�%�jK5�IB�4m9ı,K�{�m9ı,?��@{����%�bX��߿fӑ,K����iȖ%�b}����X3n��ÝY���}o�v�C���/e�ZOido:ؖj9��'��4�HnQ��ki�Kı=����"X�%��w�ͧ"X�%���w��9ı,K�{�m9ı,N�jF��[��K�a&jh�r%�bX�g{��r��#ii��4�Zș��w�ӑ,KĽ�{��"X�%�����iȟ���L�bw;I��]c�!.d�sZͧ"X�%��{��ӑ,KĿw��ӑ,Vı<���ND�,K���r{y�^B�~�����.L�f�]h�r%�g��3��~�ӑ,K����8m9ı,O���m9İ?�ȟw��6��bX�'�C��i��M\�I,�k[ND�,KϾ���Kı>�����Kı=����r%�bX�����r%�bX��ϻ2�]��	�vV=��ۂ�q����[n�=.Wg�lar�~����Z��nc��6��bX�'���6��bX�'�}�ND�,K���[P9ı,O>���ӑ,KĽ���rL�7E�&�Zͧ"X�%���w�Ӑ�	"dK�����r%�bX�����"X�%��w�ͧ *6%�by�t�)�P�RA����^B����|��Ȗ%�by�ݜ6��c�CL`�����"*0X��*�,$P������O8Ъ�DQ5��y�ND�,K�~��"X�%�~>��Y�.2��m�k[ND�,Ͼ���Kı>�����Kı=����r%�`~`�D����[ND�,K�ƤoB�2a.�����iȖ%�b}��siȖ%�`>��xm9ı,K���bX�'�}��iȖ%�Jy?y��{��~¶֡�V[��p�V�)�(����w������a��g�N�����Eֵ�O"X�%��{��ӑ,KĿ}��iȖ%�by�ݜ6��bX�'��{�ND�,K�>>��TR�3��r{y�^B�~����'���bX�}�g�"X�%����fӑ,K����iȟ�RdL�bw	�v��~���Ԑ�ֳiȖ%�b{���6��bX�'�w}�ND�,K߾��"X�%��}��ӑ,K����)�εT��6k<������y=����r%�bX���xm9ı,Os��6��bX
m��*�A��6Ȟ��O�"X�%�{�>;2䙚n��L�jm9ı,O~��6��bX�'��{�ND�,KϾ���Kı=����r%�bX��}�r~���z��=N�NW�8ظ�H���k�Vv�odh�:nI��+��%lbSy%s�Hlͧ�,K��;��m9ı,O>���ӑ,K����kȖ%�b{������^B���:v��]�1�ͧ"X�%���vp�r�bX����m9ı,K߾�bX�'�߻�ND�"�"dK��܎g�]fL&�Y�MND�,K�~���Kı/}�u��K�2&D�?w�m9ı,O���p�r%�bX�g��;��H[�4f����K��/{�u��Kı=����r%�bX��{8m9ı,O���6��bX�'�t���55��Ԛ�L�ֶ��bX�'�߻�ND�,K����ӑ,K����iȖ%�b_��u��Kı1�M����������mN�`;N(����m�����f�Ԇ,�F/;���}��k��mv�,�;\��y��|�d�+��}{[t�K�g��fO:=:���7��R���K@�o:6�2��HZ�)������N�9�q���M�*��T�,�ܩ�ѥ�y�no/����\Tr�F��B:ۛ׮�7U�\!\b�<��K����� OD����˗`�^���T�6��R��6
�m�b����Z��[�QJ�ٿHr奜R�d	�vӑ,K�����6��bX�'��}�ND�,K�߻��Ȗ%�b{����'�����/'���S�C1�u4m9ı,O���6��%�b_��u��Kı=����r%�bX�w��6���ʙĿ�N���nf���3Z�ND�,K��kiȖ%�b{�����K ,K����ӑ,K����iȖ%�by�:t�����eusZ�ӑ,K ,Os�w6��bX�'��g�"X�%����fӑ,K�ș�����"X�%�~;{?fY�.2��eֵ�ND�,K����ӑ,K�C�{�ͧ"X�%�~���ӑ,K��;�siȖ%�b~��W���݆鵁:,{f�A7 6������-�E�U�:�����瞋����<���jh�yı,N���ӑ,KĿw��iȖ%�b{����P9ı,O���ND�,K�����r:�s&�ֵ6��bX�%��w[NCé��P>0��@�6P�`F�Q#31�"��s.�p��@�Uؾ�"dK�o�fӑ,K����ӆӑ,K����i��Nr���������٪9��]����bX�'���6��bX�'��g�"X�TF
)�2'{��ӑ,KĽ����r%�bX�a:}KL�K���!��fӑ,K������Kı>����r%�bX����m9İ ���[ND�,K��_�2��Թ�R�jh�r%�bX�����r%�bX ���m9ı,K߻�m9ı,O���ND�,K������Р�%��򕡨��۳a��e:����u�P��qO}��G������Ƭ����r%�bX����m9ı,K߻�m9ı,O�����&D�,O߿o��r%�bX����˚ѫsYer浭�"X�%�{��[ND�,K����ӑ,K��{�ͧ"X�%�~���ӑ?# șĽ;{?���Ith�35��"X�%��߿NND�,K���6��c �wda5:ec	�0�}L�� ��^@�g���;Y;~%o���It�!cF��oz���a���vE$�"Ǟ2� ��InG o�I��d52]z."����s�a��4��Ⱦ��Ғ����<�����p���4�K�m!��O�ᯯ�:	Mx���9��~���+
E��A�;]��	aP��l֖ Fc�aBHB�cq�n��&<˚�|oW7D��y�qs � 4�b�zJJL����u��燆��i�׭�͚�a�>1��1X�_T�`iy�!QLWO��(��|�����& ��x���'��^����4�: ��A*�9��(��]��x�z&D�s��iȖ%�b_���iȖ%�by�M��N˫�Z�֦��"X�!bw��fӑ,KĿ}�u��Kı/{��iȖ%�by߻8m9�B���֝��kl�o���B%�b_����r%�bX���6��bX�'����ӑ,K���}۴�ay�^O�?}�z�Zl��31�:�]×[���׀�����̜aP�Й}�%���kĎ�����䧒�Jy=߿~�ND�,K����iȖ%�b}����~R�2%�b^���m9ı,O����S�jꙚ�L��m9ı,O{�g�"X�%�����iȖ%�b_��u��Kı<�����,K^O�~�e����1�E����B�,O��ݻND�,K��{��"X���DȞ��߳iȖ%�b_�w��ӑ��/!y?|�ϩ�vcs�T�ږ%��b_��u��Kı<�����Kı/���[ND�,���`$X0 0)�(dN����r%�bX����\֍\�eˎ[��ӑ,K��;��ӑ,K�F�߻5��Kı>�_v�9ı,K���bX�'��]�g�[���I�٘�v�d&9:H�t��j㥢�Ջ�ly �iW�NrO#�jJD6����%�bX��߿�r%�bX�g�w6��bX�%���[yı,O3��m9ı,O>���Yp�֩e��r%�bX�g�w6��bX�%���[ND�,K��{�ND�,K����ӐBı,O������u��MZ�m9ı,K��w[ND�,K��{�ND�Rı/��Mm9ı,O�ﻛND�,KקKzrk&�r��f�Z�r%�g�)�=��߳iȖ%�b_~�kiȖ%�b}�}��r%�bX�߾�bX�'�N�R֮��Ԓff�iȖ%�b_>�Mm9ı,����ӑ,Kľ��u��Kı<�����Kı=���>��� Oߋ���ja�NXļu�\���e��z� 񎛌��zs\>��6-�g����ݍ�raC�]��S�,��(a�[�8��3���7�������Vs�]�lN��J[&i�`��(�ŵTFǱРtb:ۤ �'J]7t�:�6�okx��n�����
Zt4���c��ѻ��9���%��Qkt2�@,�ѣ�MFX`��
7CX���D�V9f���?Ns�I���^*����\�t���@V8v8��]l�xӚ9t��;�(I��y��K�	��cB�����!y
�'s���ӑ,Kľ��u��Kı<�����Kı/�w����b[�^O�3��1�ՂZ��r{y�bX�߾�X�%��w�ͧ"X�%�|���m9ı,O�ﻛN@m�/!y;�}>�
�l���/���Kı<�����Kı/�}٭�"X�`"w;�ٴ�Kı/������^B����~]�)�0r�6��bX�%��5��Kı;�w�iȖ%�b_~�u��K�,N�]��r%�bX�w��s;�2aI�R˭Mm9ı,N����r%�bX�߻�m9ı,N�]��r%�bX�߻�[ND�,K�h��$�gn�����c[�� �IU�K�j��h�k��͖5�.a[�j������/!y�߻�m9ı,N�]��r%�bX�߻�[D�,K���6��bX�'�N���[���u&��Ѵ�Kı;�w�i�P<��XXx�#%#�+��OT�D�,K��zkiȖ%�by���m9ı,O~�xm9ı,O0�=�Z�Ԓۭm9ı,K��魧"X�%��{�ͧ"X�b{����Kı>�{ͧ#�^B�~���S�l5Zf039=�bY �X�w��n	 ���vlI�=�ﴛ�H��|���m9ı,���w�v��X%�[�'�����"{����Kı>�{ͧ"X�%�|���m9ı,O����r%�bS��I����Z�p�-fmB�U�J��jk�)cF1��s���.N1�Y�y��y������35sF�ؖ%�b~�?��r%�bX�Ͼ��ӑ,K�����Ȗ%�b{����Kı==�{�fJK�L�E�fkiȖ%�b_>��[ND�,K���6��bX�'�}�ND�,K����rbX�'�ݵ����Y�R˭Mm9ı,N���6��bX�'�}�ND���h���$ 
)�>]�W��	"w5�fӑ,Kľ{��m9ı,N�|o��1`mY��r{y�^B�~����Kı;����r%�bX�Ͼ��ӑ,K,N���6��bX�'�N��'%��f:�Z�Ѵ�Kı;����r%�bX�|��5��Kı;����r%�bX�߾�bX��~���6k,s����lf6�۞�ix�c6\^e��m� U�.M$�7]�G��c�RK��ͧ"X�%�|��5��Kı;����r%�bX�߾�Ŋ>DȖ%��>���r%�bX�?�e�H\�Թ�E��[ND�,K���ͧ �bX�%�ﻭ�"X�%�����ӑ,Kľ}ޚ�r%�bX������ٳ�%�-���^B������9ı,O���v��`�X�%����ӑ,K���o�iȖ%�b}�}<�WU�t�67+�'�����r�pȝ����ND�,K��ߍm9ı,O���6��bX� �灴0wș��u��Kı>>���e�V���fkWiȖ%�b_~�Mm9ı,C���ͧ"X�%�~���ӑ,K�����iȖ%�b^���ᄙr<tbގf�F6FK��uú��W$=�f��F��y1x@)T�39=��%�b}߷ٴ�Kı/�w��r%�bX�w_v�?*O"dKĿ~���ӑ,K���\�dչ��2h�kSiȖ%�b_��u��?@ș���w��r%�bX��߿�r%�bX�w��m9��ș���~��NK���u2ۭk[ND�,K����iȖ%�b_{ޚ�r%�bX�w��m9ı,K���bX�'�N�Y��f�kRMf����K�ȑ2&}���[ND�,K����iȖ%�b_��u��K����ȝ����ND�,K�����Ң�1������/!y����ͧ"X�%��9������,K��~���r%�bX�������bX�'�mS�	x�	"��9l���=<�|��[��kJ��Av�a���]m�&%���"�ѷ�c�1���`-�5kN��>9���n�o+A��Z�I{�03tsj4�S�T��N�k�'X����N�A��1Pȩ��sR���w<`ٜ�	;xn��zG�E��;g;��ZN�;e�&˵���u���O>eP����GB.�V�c�V�'�f3%v��XM��О}�r��6��a3����w;n��;Wc r���asɫ��=dm�����˳3F�aud�֦ӑ,Kľ���m9ı,O��w6��bX�%��魧"X�%��~�fӑ,K��Ӧ��Y�WM���r{y�^B�w}߷����,K��zkiȖ%�b}߷ٴ�Kı/�w��r%�bX��k���Jj��E.kY��Kı/�w����bX�'��}�ND�,K��{��"X�%��w��ӑ,K��㻶�fv��fj�\ѭ�"X�%��~�fӑ,Kľ���iȖ%�b{��۴�K��"�"g����ӑ,K�N�Z|o�2m�LVeo���B���}���ӑ,K���w�iȖ%�b_~�Mm9ı,O~��6��bX��|������L�:��˂���V���<Q�.���؋�!�|eQq��#�L�Y�kiȖ%�b{��۴�Kı/�w����bX�'�w}��(�"dKĿw��m9ı,N�?=��#[b��'�����/!��}9=�"q�������"X�&���6��bX�%���bX�'�k��NA�,K��R�'Ki��K�4[�5��Kı=����r%�bX�߻�m9��C"dO��߮ӑ,KĿw��[ND�,K���rfL��53�����r%�g�>����r%�bX�w_�]�"X�%�}��5��K��̉�s��r%�bX���y�R���l�h����B������۴�Kİ��G>��ƶ�D�,K�����Kı/�w��r%�b�����	�!�5xU��eM����� ��T2��3I�/C��̝��C���?ˀ:�E��ӑ,Kľ�ޚ�r%�bX�����9ı,K���bX�'�k��ND�,Kώ��Y�v�e��YsF���bX�'��{�ND,Kľ���iȖ%�b{��۴�Kı/�w����X�%��ڗ�552��r�7Z�m9ı,K���bX�'�k��ND��l"�H�����" ���P����6X��{���m9ı,Os���ӑ,K����zgsV�RMf���"X�~��;���v��bX�%����r%�bX��{��r%�bX�߾�bX�'�N�[�`�.��S�Oo!y�^C��}8r%�bX�w�ͧ"X�%�}���iȖ%�b}��۴�Kı;���%m�lv2a�0�Gmn#9y�e������]�h-�/���s�bw�Ea��m9ı,Os��m9ı,K��w[ND�,K��݇��L�bX����kiȖ%�b~�G��3$4f\�Y
k5��r%�bX�߾���"X��~�ND�,K��ߍm9ı,Os��m9�eL�bw���U�t�!e���^B������r%�bX�ϻ�[ND�� 0ș����m9ı,K�{�[ND�-�/'g^���!�ai��Oo!y 6%����ӑ,K��;��ӑ,Kľ��u��K���Ty,p���"3�|}@{"w���i������~����b�$)����Kı=�����Kİ�$������,K��u���r%�bX��~�>r{y�^B�߾��h0e�2`J��.����c����!����Hm��6ɞ%ژ�k�mL%���Oo!y�T���u��Kı>�]��r%�bX�ϻ�[yı,Os��m9ı,O^���p�5�E��k3Z�r%�bX�}���9ȱC"dK��ߍm9ı,O���ٴ�Kı/�}�m=���rk�^N�?ܺo�r���ؖ%�b_{��"X�%��w�ͧ"X�b_~���r%�bX�}����B��������~�#��`f>'"X�~�~��6��bX�%�����"X�%����nӑ,Kľ}ޚ�r%�bX��G{��u&e�5����fӑ,Kľ��u��Kı=�]��r%�bX�ϻ�[ND�,K���ͧ"X�%���|�0�˷T�|t��5��O<<��#BHBxl5����	:y��m���``}��n�� �{5�3{ѭ�w�v�~}=�/%#1O�Q=g��i�z�g��|=�6���HW��n'�dFMp9��.�@6��G���ؐ)���1�@"ajF1 �J%!9�������*�*�����   	 � 88�{Y�����=sg%rF�.9Оce� �&F�S��F�gl�]���Y��y�X��.�p����谭�X�� Dn�p96ȸc�d��N.w��nXw�������fT�v�u9&��'i�NyȐ<�R�֭��'�82͇D��`l1B�lZ�kR�9k�۠�:ӶX
`udXn�8� �v���r���%�i���T֘0M�m�X:���!=kjt��);k�L��l���s� 3�5	5Mv�є4&�X3���kV�.4�l[��H��(j��8T��s��<X�@�A��W���(�Dz��F꺠�#N׬�½��%O ���U ,n^������-�>nd�%���eꖳ�P&xy�S	��Sm��m� %V	V�9v�Yvw]�(�F�: �hG�Y���j�F��s�\A s
.mIFfe�YP��R���1��*����=H�r����*�*�U]Rv�ؼ5��ٺލ#l6N�v����U��V�,���
e���Z�T�!kD���wnN�
�.ܣqَ��pF,�5������V�ehb6l�ni�c��X���%���c�>�k:�I��e�nx�6Z(�p:��1�����M�ql��g��`�7\E0L��@qc��ٴR���c��Xn7e�M���q&�����Uvt9�A��S�$�*چ籝[mu��F�
PΜ���K@T�f��Jz J��laB�7hi�v�@`��d75�m6�Ґ��k��M���؜s�g\�F�oN:�L2\��X⧗�x&����m���n�S�F4l��U�vh �����Vۉ׶de�`�J�V�9�Ԃ�u��P!V�U-�W,��*��k��g��@Y�m��m�ƺZh,l��f�����Z���ѓlڢ��;t�-J�����k6d4��ѫ��F�)TWH��|��&�4!t	��V�_�G�	�8�å_����_� ������J���s��M�������6T3�h6�]g��ss��dú9��M]@�"X$
�y����D-`�1�L�E�aSfu���gh�*� � -�)�����m��@]u�k�r��1(�%[v��r1(�)@i���n��Qz�ɝ7<`�.�Q���2�v��Fc����Ǝ��Wk�[A7��4t�,��:twGXv*��Ѕ���̳���Ӝ���I�'��˪9���:�bY�/#	�wc��f�\�Bc5�E�%ص���#<�D`�m��2���y�^B�w��r{ı,K��魧"X�%��}����"dKĿw����Kı>�?7���F�<�������}ޚ�r%�bX����m9ı,K��w[ND�,Kߵ�ݧ"~���ߧ���cn���|�����b}���6��bX�%�ﻭ�"X�%����nӑ,Kľ}ޚ�r%�o!y;֝7�MM��u�]�'�����}���iȖ%�b{��۴�Kı/�w����bX���}��ӑ,K����zp�sYtY�&�5��"X�%����nӑ,K��G=��ƶ�D�,K���ٴ�Kı/�}�m9y�^B�}��|cF��%s� �.���l!�X�Ƿ=�g�	���. (��M�䯇��<p�(�r�r{y�^B����y��H���'��W+���l~��6�j}�҄va�c����O<��$�ܪ�q�~�Us\��y�� >�*��${]{�'J���[)S���'� ���\H������X��\�V��ۤݵV'w���Ke�� ;=���X�\�%�z���B�i�V�ut�;X��W�{�����/�6O^�r,��~�δ�r�1*��i�k�w�sፉ=��\^��*�R�<��>y�PV�sd� � wv^�r/ܮW?W*�����x����S���V�n�`we��W*�I���ޫ�;�E���#y��^����X����� �l��͆���z�U<�8Ur��_o\�`���7�N�m�[�Mr������������	���������-��,ki���IU�t���xuȰ�T�O_�l~��>�%,�a��ţ.X�)�Q�E'm��!�ӄ������&�8��ReW�q�ݬ ����X���|�c���g��s�e�l���=����?y)�|�~��O?ߖ wv^��jJX�@[*�v���K ��U��M���x���`ږ�D�(i��	�,���-��, �=xuȰ'��UW��~���6�Z0Q4Eh��Q�4*qE=��~��&w�,ߘ��R���MHj�`{%��"�;�%,��X�I�I�އ��֛)+ͱĶ�{���'WTf�#%��_ű��@4v�Be��4cm]"��w��� �\���`we�֧�m]�ڷ�wk �\����r����� 6O^�r,��b�!%E����N�`�"����;�E�}�JX]*(�J�i*�R�wk�Il��c����)`�"�7��zꡗM�lK��|�w��}��_z��l~�����9��Tn�Wwwz���-ď=;��0	=N����v�l�\A9����f�-2�]X�T���ȑ�8�OV�sP�g��z�l��s���:�n����v}��8]-An��n5��������l�:�Pdl����Y�5�jx爑ࣵO�%�-A�E��-n6Q�.�N)ܦ��ָ�x�Y��d�gg6nr�Ǜ7n}PY2�,HZѳj��a=��g	9$��4/�`g!V���v[�\n�+zԘ���(S�Vy�=X���Mj�.ipJ�Z)�쥀w\� ;�/ �ݩh�(�;T����;�E��s�I���6?y`k��z���D�D~�i���.�����׀w\��ĵIJ���i�t��@�m��ՀMrR�;�E�ݗ�oZ�7�]�ڴ����>�%,��X������%��DR�ji���t���;p� m�\��
W9�n&��ziل�9�DlMͻI�,��X����{�\���oߥ��I���J�[c�fV��}�[TX8�)�4Um�{��䥀w\�?UW+�*��ҿU���Ю�v�ZN� ���� �9)`�E��/ �k5$�!�ʺT'k�W9U���{�?~��O����/ �r,����$�c�LM�,�Ȱs�RO_�H��}����9]ٔ;@�4 ��D0V�qsF�r�7�d���͊��F��-ۚ�cMƑDMq��|$���E�}��W*�A�~��7��%�ʷv��C[��7\�?r�;��R�7��X�%竟�\��F�RO�-Sf�#��;�~�/ ������vyj-���m),*�bƀ)�W*�9h��^�9�w�j���ջ���X�U\[��� I�^�dx��?}-�?Y��4p�*yhn�x�r���y��{���"�;=f�k-�12��o
-�'�`��j�tѵ�s�I����p��c�㌺ė�7\���S�xT����_�ʯ�{׀mFD��!�Zj��$��d�y��U$o���Oz�RG��ܪ���_� ��M1Z��wW�{���`엀j�< 쒯 ���b-��MHj�`{�I�^���U��r��@�R�0
_TW�����`�+�7v��!����RG�~�9���s���}ߟ�� 7d�����͎!�X'�������#���\����,�T����Y�D�6�Պ!���;$��69 n�~��"����񨼁$[��wI;��69 n�x�#��*��r�����+��n�I*�R�wk =�߯ �$x�%^������N�XUfٶ6���<�<~�߿< ��~��69��9�JOz��/]ۡ
�n�Rn� vIW�{���=��߯�I�����=�}�nI�� ��H!��K���ֵ�L%�P�V����h����:�P8�Չ,)k[,2	�1X�sm�㍨	Eq2r�n��Y�n��҉Kӱ��ҍ��pؓ:�S[M����"/j�0��qy�v���M�Z$^M8�y�����*�8��8�5
�G\{z9�A�}�����.��j�8�8����U6gQ5�v�]�.�*������g�]x��!r��\E|UĀ���y,%��0ն����37r�B鸖��wXk�d�ܖiu�%9�79�+�$�b�M���'����/ �$�U�}�U���M��6�M5aM]� ݒ�RG��U��>��}/���#s�+巧�}��vIW�lr, ݒ��QF�+�ݴ�o ;$��69 n�x���v��E�!Qn���$� ��X�%��� ��Kx�$�o2���ktX�k��4��kg1�P�m݅�$\�0j�lm�5�#�G��P���Y�_ I�^�H��䷀lr,{Q�nP�d"
�m�w��^s���̈́��P�!	LnCl,$! B3H҄�h��8n������~���/?s�IJ󻻢����T���w}~��lr,?W$�� ����>��R��i��,wv��E��^�H�?W*�US���ְ߾�m�.���U� ������UUG�y�w��X�E�{��W+�q���qk3�pe����ݦ��.�Y�56�D�aCv8p�������vX�q��n������}�r�#�~�>@I���>��~�T*�˶v���:���ʤ�y�� 6{׀E�<��1G���r�e�������òO|�_C�!��I-�<�π� �[A�R�^��<ZY�<4����yHܗa33%)mH�`!.��fe�:YL2h���`�3\�2��}%������B[�U�a$��K���D���3	�B`�Ws�y��kT$Ij\8]�%	FH�kV��b��!�HE�`bD�1 F$�vL�W��`�O�p��PG�!#e&fݡ�&s1��s�@��n2��5J:p @"��IXE��sI�	t��?a�EwT���L4�_�M\i�����ї.H"`BK��.�x|dO y���B �X1��/L0L̗	rM��CL��<@#w�2��_��=Et|�qB+���� ��S��U��S��Ϗ84U�D[uu��rO=�_j�I����6]:i*�&]�����z�G�,���X�"�7��K�v5wt۴��wx�"�=Uݙ�_����/ ��l��L�ZJ���vm�����͑�l:̈��s��̝��C��ek]��ҡ;_ݗ�X�"�엀Mr,�]�ēLV�c���Mr,�ʪ�A�޼��� ��r�5ꦜ�m��j���`vK�&��v��w{x��uݗf�e0�r�k�`wnZ�&����I�QʨI�F�(5*�$0�#�rO$�I4�c޿ߚ�{����7cv���-`\� ;�^5ȼ���'۷���a�!qL&L��W ۄ�;���c{se���8\�e����8��wV��v��?ߖ wd�k�`�=z���	���5�:�U� ��y�$z?y`�~��Mr,{NT[�ec�lJ� ﻽���[��K��� 6{׀v��4�$�j�P����vg�`��Xݒ�=Uʪ�Ro�y������߉m��L��\� ��-�������v�UW"&��TH�� F��[�3UT�&�lt�^�����Ō ���e0ESGehbz��.�sc]Fkj�P�3�-pZ��5��hC�K�pO/kQH:4[��cb�(��Œ@�}��ʹ�O] çE�@�eDɹ��)�Z�3��&]4[B��@l��bۜa����*�8�f��*��W#�帊y^�ψ,���(��3!�(��ɔ,-&f����ɬ6D$�j��
)1��{t��^��X���拍�x��^��&x�߸��~򨈗d)|��^5Ȱ��-~�9�r�A���mz���n��wHe����\� ��r�5Ȱ�%�����5���j۴[�����l����Mr,?r�č�߯ ��������w]��Uv�p=U������߿^#ذ��-`�����Um'v��vK�?s�W���ˠl����E6<���
��v<u��ɞ��sٌ솀�ܽ�Wb���E���vP:�E��,U�%W�w�ެ�����@l�� ��D~���d�IsWrNy����b0JBV�4 HEj��KKXG�B��0a~�p�ɶPVC �T*�k�	́B1!��$�3n!}DyU��||��x7޼G�`v�t$�Lb��.�����K��I{�y`�z����Nq��M5t2��ꤷ���^�x��[���/?O<k�5�1;LwHe�����ǀ~�Us������ vIx�GN�UnM��l.K[��n�}K`x�n�\Y�Ō��q���i��&mr˳��-���u�)��f��"���dm���i���"� vl�.����w�ut	�t����N������ܓ���f�P�F�X�"�9UH�s����e��x���v��劶�U��;��>_}���}����O^)z�6�I˥I�xV��=�Uy����z��#�=����c����"�56���x��7��vi���vөx�pn|�\簻��J���<���͗�E�ջ.��]6�14�i����f��"� �ݗx[�窹č�Pח���!���w�yo����w�E� vl�kQFYv;-;�-�n�ջ.��c�͗�*��R�P`UR�H[)*`�2�&��I0+LM\B��V�X��R���^s��9��� �v����U�������nǀ�/ ��<�v]����Om,���L����R%:|�i���v��xчU&M�(8x�-q� ݻ o�� ��<�v]���Ry��o�깶�.]b*�ߝ����"ݏ ;6^J��+���R�ip	7`j��x����x�dx{P�)���2�]��nǀ�/ ��<�v]���7)���mXRWk ;6^�H���w����}w$��	\ T�P��	�d�O�{;�UGSy��Z��g�Ga��svgmΝ�b���p�&�,U�鍽P�=�����ғ���0�b���lT�����Q��t6�Ѷ�7BЛX풹5��+2X���Dg��KM�
��^��b�'kd8֩����KZk`�;.��)hBN�6,N� [/������ٷ��ۗ��\!�[���'^9t�6�CUn�X��`�؉�=����z�񅣴f��m�@Ĳ��N�Ztn�[r��s�����@4v�Be�*%uqs�I[��"�<�v]�� ;=��=�����L��;gp��z��"�͗�j�<�9�$mJg�T}�f*��^߻�������I<�E=�m)<�U�"�j�SIU��wk�ʮs��g�xS�xinǀw����f���V\��U��{׀v��xV�x��x�v�-&ލQY�.6�)� �t��$3c�f�3���0�J��V�XL	��<����xV�x��x��X{P�������|���ϞIɤ�<���\���T�m����Xinǀv=tܱ���mXQwo ;ݗ�}�E����K���x�<��hkPڜ�i7wx��y`����:�c��=��?�k��l]Zܰrl��/�ջ w�/ �\� �W8�)O[����� ��Mf(���nD�[�����qsiY;,;f^�½�Iu6�[�O< �v^���.��U�"R��T�Um"۷����>�"�>��ջ�NBݻb��N��� �\� ��ذ9Ï����R�B	`�Mb�d����"�h��4`@�7�z�Z��UJ���� =���K�B6���[.�
�`~�)�s� �'� }6^�r,�R�	�&�&��V�`Sc�=���US���}�����=� ���h�o�Gm������DŃ���tR�z��`��A��来希�.��m`�e��"�7��/r����X�P�E'�7t�E�]��r,��6���7�y`�e竕�$wZ��ՖݫN�um��&ӞXT����URG}=x��,��ꦘD[WV��;��uM� >�/ ޹UھUQG+��b:TG1S����ܓ���.�4�[H����e��"�7��,�lx�t���N�5M�V�ǍDqD�V��nN��O~j��s�z�q�X�XL�U�.,uW�����ߓ{��:�����}=x��y���al�@��{Ob�:�ǀM��o\�<��W�P�<�hb���ݬW�� }6^��Jk��6���7G������M�7o�T�}=x��,{NE��UR���z�������豫��7�E�oiȰ���f��.����r
D��`&��h�=�'������>�Ҧ�޾�ɚ��x���"/8fqi�T}�Awx˅�	sW5��oE�y�q�3^���r^s��
_g��0ϼx��C�c(2#��H�X�Zg�sZ�[��`JȠ�)��-8C�"o���oz��� �=�"[�xy���,�^2�h�H�3���M��YM?:)�|!l���0 ���9��-�q��o�G%%�KO��AW��b�"�����.�<u�j�"<Ÿ���5�S�bf�g��T�����yA��� �!XM��}�o�,�8\ѭ��{��؄���)�r���g�c�
���'�Y#�3����99�|���}��ʪ���   �Z6�`�8� �J3���msڲ��:����r�qEs����������p'����4\(��jm�[Ar"�����="0$&ͭ�y!!ȧ)�����9���J���;�#n����\�Ь��K��b��0��"����2��l*))pJ1���u��a��2�7;0"��n]��]���T��b7"m�ӷS��9����qN^�!Tp�Q���;lN����=!�����u���$�&�
U�ѩ���l�k��!�]���a�N���M���y���n�.&��L9\���
ɗ2�[5����{ld��jwf��] �OK�cl�&y^�:�M����2��D�%��@I��t5u��I#�*�k�@Y�d�����JV�T�s�9��)V�=��E� %�����#��;^( ���"��d&�j�Լnr%���s�kGYCͤր,3ij[�X�sR�c��l���$�	��ut��\��U),��3-��g�Ռ��`q���l-���͗\ h�9wH��l��εU��x[f�x�.j���{pY�F�ڭ-r=�dGs�M���1�3C�Sbg�#�tQ�]K��7cc�c�������V�֞�->�s���q�ݥ������ƪ�타�ι�}����b�פ<g8���)kc9{�N�լm��7rD�� ��!ֆ[�UiVs�iT�+֡�+'f�ڲ]�.�1qPPض��mS�P
1��H#�OV�k�{-<�2��[5J��J�E�eZ�1�[=�s����C!����.D�<�=����+�\qu��\�5�n�VC\���\�UK�WZ�-�ŝ������q*��d8]F��mX�N��i�A�6x�۶đ:�,h�Wj���]�eZB.���h�A�#p��\k�@��di��`*BiPm��U�m�����]�9���-mt��Iu��C�Ǫ�N �N�"��b'�6�z ; S�P��J*(A&�)�q�Q�=�D<@"���S�'�<�������!6h��t�WG��A�Fl�1�m�\2�5Y�r\<2�ր��a��^�����gf�rZ��`K�Ԫ���b�Z�uci�������I����nd�m�V�yL,�(��4���FŻYˎZD2�׬{//R�.��e�+˛I tNR�un�񮵰�����p8��7:3s�ɷ]�C��e�s�j)M�t��?s�I<|G0�a��J�D���D�&�� vV�V�4�n��1���K<(�1TU�n��X�9�6< ��~���,v��7l���XT���e��"�7��X](��N�J��[v��e��"��Ħ��|���w ��]2�Vl���^�6��M~^xT��?s�OO^)mD��-*���v��<�+��~� OO^�r,ܮW){`��,{r�X�M�$�1�����ny�V��lE�tnq6�3߾��z�>�T�#��_�m�~x�K�7�E��UU_ ����	?ZV&�,(n� l��r�����h�3s����=�>�Y�'��?UURG�P��'�7t�E�]�5�� �\������/ ��j���v���۵�j�S�:�ǀ$�Ur�����MA��T��Z�%wO ����S�����,T�������j�\���`�Fm��X阷1�
0+�Y�)���p�y�'��O۵��H�i*��m���~�x�ȰRJ��rrz[���o-����l휳eԎWw�o\� ղS�:�ǀ�^~�T�^���o���Zd��ӿ}7�O/����x*pcŐ#��I"e��$!� ��V���X˟K�${��'ȝ7Lv��N��~�r��O< �{׀o\��W9����5/ZVLl���x�%��"�ͅ�Sc�>��k�Y��`Y��p�rj���B.'v��C�o[;���p�SK���f�/�7�ن-kWw�_���axT��U|��޼�����`�ټ ��z<�%s�I�<�Oz��g�Uq#v��4�	v5aj�W�� n�x~�S_��}<^J%��iU��n� n�x�Ȱ�ax�s��s�䜼��9���/}��������nȳe«j���`f�������=��w�i�.tϖ�sF����W�s��741�P���Ɂ$).}pu;�^u����[���"�'k���xT��vK��s�_�����'�'I�v�����7\�?�ĂOz���� vl/=����y�:_�P���	V���ߞ󻽼?y$�F�x�G�,�(9��AcWw�v9 vl/ �r,ܤ��� ��}��`�ټ ��z<�*K���{׀v9u�{��*�$�$������ӳo�Wkp-h+���8-�C0JYbUC�:6ݱ�n�j3�H!#՟#T44-�Pn���uj�5�,�@�h �dv��y�&mi���=���kfy��<��M폖���Z�p&:�%Q�lon�7f3�K5�q{��B�ǁxؗ�]lڴMږ�D"	c-i�٤�r��59��:mҭ)ӱ3�׮�A�cu�f�ɢ�nP-٠��'�s��+�����.)�3�8]h�y�pj�Z�1����$A��Ŏ�e�F\û.�%vƕ�Ӳ�����/ �r/�U|��O�yh��WM%V�j�� n�xc�`f���"��r�$��?8�s3\��¾[}����ax~�%�� I�^��"m�-�iZ�t�����5M� 7d�s�z��s�I>?14�j�N�T��vK�6=� ;6�~�r�w�|�8�tZ�5X��*�M�cv��,�p���a���a��g��/����ݿ�7�׀l{ ov��U�_����P?�����&������Y�1H���HbB���"�P���#�-�,	��o9U�l/ � vl�h�N�Z����x��z<��{�~����'�~�߽�u�P�)�m���Ӳ�Sc�͗�lۆ ov�E�#��ݪm*���v��e��������Sc�>뭍�v������렣cko�'�7A�l:|g��՝l���S,Vd���r�{�Ӏ݅��ǀ�/ �����iZ��;0{���"������6�w�����حSiݗ�j��nI<�ߵ�����qd8�Ȅ � a�FRY���Үr���u�?�X��^�ֺN"Ʃ1���ݼ�Io�� �s� 7��5M� �pS��4���b����Sc�͗�|�q	�6`�vd�c�><�`��:�O1ۋb��,f׍댜
 �}%o��1�.��= �<^�lxٲ��b�7Z�Ʃ;��V�N��5M�;^�q���'����Ӱ5|��We��V���� zl�cذ{��T������0Y��J�^�$���o����ܒw���ܓ���f���)�P�����5�ܡ4�E�Н� ��/ �6< ��xǱ`��=��X��g�3�IttNԛ�Ӕ�`^# 7uN�4MA�C���s�߽�ޣ�W�5��m�_���f��6=��9Uϐg��$qS~E�Rt6XZ����/ ��, ��/ 'd���H� ?P����wx��X��^ N�xٲ�������1���x����� {}��͗����� ���ۻv��Zv^ N�xٲ�	�b�~{���I���)��9��X��0�s
�^.	@��Q�m�.O���g�[,Gnm>�kv�P�لv�ZKp!��kFn0I�*��JOW];1u=��uYQ�;[�M��\Q�҂�M�
)5KXg��XJo&m�b�t`�R�e�s���%�GZ-K�:��1�۵mh���7��r�Rb��v�̷S���:v�f�4qj���K~?l�`��w��{��{y����Y��)��\^ϟp[�1���m͖��gvt���������������^ŀ݅�W�9�����=����ˌ�\X�^�w�� ��/ 'd� ��y���q#�'<�~�4�*wt'k &���^�r��9M���^��ߖ��]D������6��x;%�f��&�� 7��7^�n"����ww��/ �*�^�<� �<^dx�I�p��tyŶ��+��t�T��Ӥ��֍��b� t6�m� ���{ ov�E� vl��9Wj��-óx��z<��4œ�#$�F� !D��*�Q�AQ#> ����'n��nI<�z�	�b���$H? o�Wv���-;/ ��y�f���z9�g��:[���8�"�-�I�O������߯ ���� 7��"� �l�w�.29qb9x}����{�����f��?Us���G�&۫@]۶����gp�:�ɝV��Xl�q�	����&띧���$�x�!uYL��� >����]��͗�uwc�;�K���6�ҦջW�|�#��/ ��ǀ�+�s�I�����Rt�V;���׀uwc��y�U@r��J��ATD��d_�� �P���P4p�|��}����s�I�}����~$_x�ۮGp�q����Y�%�/% ,�u]4�Ye�rp?��.�� ӎ��.Ye= ���aB���&]ᴡu	�3SSPL�L��,Յeu�\ @�	"A��3��!8 ���O��_=�'�~!���5���j�Mie3d��L���d	�W4���2�"�O4L2� ��F �!"B*GI�	"ؔ.�)�#!�*1�ɪQ�CR�4S2n.�0�0�KHa����qEt��
��P��8qw�ȏȂD@��SB zb���>���P� ���U� �<����5vG�l pU9t�aan� ��ǀ�+�>]��z�)���6��]��-Ϋ���x�7�� ٲ������N�wn��ٙ�ػq���a�ĞT�;M�loY e��xS-���:�G-x�7�� ����)���9��]`{߿+�5@����wn�V1
ݬ ٲ��q#��� $����������s�.ծ\X�^�{�����Ħ���׀j�Rr����S��x�Ĥ���\��~��nN���b�H� �"� �M� 9�s]��>{�����s.h�b�j��ذW*����~�����< ��k�>{����<l#n�l��z�8t���]�t:��mcD�PrCff�#��vӵ�6^� nȯ ޽� � �6�r������~�q ����;���/=UUʮRG����1v��[�����~���a�W*�7����y`���2[V۶�]���~]��� o���;ױ`��x�M(���iXĕ�X�%���۞_�y��`��q�
䑀A���he���ךЂ��%M�s�;\����Н�� vNq�V�V�8�Sk�7E#��u�Y�Cxa��e�]q �H�c�V�/R��܏`�s�[Vt��R͎�Pq&ـ��bb�k(U��h}�+�W7�3�#e3Ae"�mM@�6��]	�rα���sx��h��&�l\F�pa�R��˃:��6�՛�>�,�R,Y�l�]�c.����$��ŗyp�f�$mi	H�!��%�hk)��z6Y��3\|ܙ�=nh#S+�n�r��r��w߫ յ#�;�"����� ��y~��j���0[R<�{ vIx�ۆ�#��RlM�t�����>�ذ�K��we��	+޼u�M�j��馬)�k���K}�^ݗ� �n�x�{��K��S�M������u�^�s� >ݗ�~���3l���p�D��1�Z�Z��SC�`�!���"�����@<��jU*xWv���Q�u�X���U�|��/� ��?ZV۶�Z���>��wx�ˬ@�ћP~nI���nI�k�~{:���������1J�����nz��"l�^��ٳq��f�,G/�O��~�~8�z�^�{ }6^���Ԝ��j���0{�/ �^ŀM��}�p���Mht��y���hZ�U�.�m�e�r�q�mh��{Cn�ѹ�� Ϲ,]��#R�i�]�kذ���n����^�����ST�vӵ�}6��+�Ď�~0l�^���=�RG| ���.�l.��0�~0{�/r�	6XHOPPPus��o ���ӀO���fgk����N�W9UIM���;�y`M�`wn��hT��v�WWx�{�ۆ�v�ݩx���Y<5v[�E�/-���g��X�dz3#�Kv����lav�6c�L:���G'����`�"��Լ��, �؝�WE�v�b�Wf��z��	��x�|ym����>�{���|�ɛr�*�	��x�����0��`qi%SM&���wWx�9Ĥ����ٹ'>Ͼ���8K����1A�D4
�	H(M*'ɡ֮�7��<�=�Ϧ�0��݀���M�`G"��Լ ��x���w��ntr[�j]��0,�\�2�Rڮ��D��wD�s�p�M�n����mշf�� ov��we�����>O���)���ƺ�� {ݩxݒ���0�`�[LT�E������%�M�a�r����ez�P���wi�c�����0�"�5wj<r�-����y;��.�i6.5v`�"�=\�{+��	=��>�p�>Ӕp�U�W�}�M>�䙒n3o�����DWF���n�n�l�#���یu��=������7l۳���9|<���+ݺ���dd�+�����Rʡ�6�mX�[b�q�m@Ug���v�3��B��;V�t��[[���p�A��3���J7�L�)�k�"9�����&Rc)]�m� ��ˌ܇V��K�%��%��=���ୄN����k��E.s4������Լ�x��M�#�.�w_�m���ۭ:��S��Ѵ"��j��k6�"�unӰwv;��~^�_� �{�ۇ�+��|��w���M;t4��ױg���_�z���, ��K�;��D�'I����]����X�ڗ�n�� � 9Bn�.��][v`G"��Լu�X�.�g�kG�S����Ytմݬ ��K�7^ŀ}6�}� �ݑV�������'���rU26��4�T��+��"/W&BG��dv�� �r,��Ƚ_ &���x;M~��u��j��wק=��А�j��UÕUU�����/ �r,���A��n����$�SWf�~���Լ��X�n��*%n��v��v�<��^�c�X�n���y`⇽Ɠm�an����6\0��0	�E�ݩx����{�s���+��&�c���loU�v�+&4�g:��V5��w�l��)ڠ˅�������k�`�j_k�8X@)6�r�6�����������7e� >�/?r�������w`;e�M[Iـez�	%�	�r���ʃ��$���)������9%� �q�ISr������	%� >�/ �\0?s�ʯ�����~���z�?7n�ZV1RWf }6^#�`�j^$�`뭍�v���#t
�W�j�9U�-�Nw=r���%z'�1���$M�r�d[n��^����ߛR�	��M��n�QQ+�V�;wc�X�ڗ���H�����z�	�E����#�P���m��-�Ӻ��==~0��	�E�ݩxz8�R�lN�ʴӳ�U%�O^�?yd�{��ܛ6~h,ND�U>@xU�;~��{�ԛu�[��X[��$r, �v��K� }�/ �uD'�H`�vH-pewC����\(�n$�;s�jNw�6@���|鹬�;D�� �v��K� }�/��W�������M�jY��;g\���^���;'� �����ڗ�j����v�+�+� >ݗ�H�X~H����~�x��z�X��m���;�ެ ��K�	$� �l�����+�cV�bv�{�/ $����I����rNG�s��t��kج��"ITᨡ��t�PۿtX�@��6q�k?y��8�>O9�S�B��������] ����\5����N)E"/ ����H1|֍hq�>�X�.���/�P�}w�B���ξ|���e�����˜�S~�Ӹ�.k{�Q,a��~�Џ���.����o�I�O u�~����7�� F���|5�K�hA"y��y�y���1'���z�߇>|���w����V1F2%��{�J3^ku�$f�<��E��H�0�ys[%�Qjt�� ��B�<<��^sz����7�� �!(H��:#�d��>��wZ׀ͤ�̅�5K�%��g���y��=���9�_w���H�Q�A/ލ�xNa�9�o��-��h�l��/�9G��ٿ&*���Zֵmր     ��m&�pր#Xt%k��JN�]nMؖ�l�T8v(RcV�@6�y3ԛ���~K۾�؝��̹����Թ+-d�;�6�� ��+��KAl�Z}��]�võ�v�s
�om�jSm�{\m|}��}xx��>��iyby6�z]�ѭ�8��l>M�q�7m����yog4���<�W��5X^�;:�n|h+�`:��)L�Sۤ�a�{M���h����"v�	Z�1���e�����g@p���;���Am�3q|}��v�����W�S*ۑ�XCy��)f�)S�f��u�9���ݷ6�qƼ�m��9��e����ҥ�ST��� M�vgB�Z�j��+���x �Bj��Ö���9p#�@$X���C��jP�BX(����VJ������
c�,��\��cYiu.�]�jv�*��jxd��V�j�UZݓ����I@��>ivybe�eܢ�*ڇU� (1��ʁ��˩�m�W`���UU�Z�L�<6��J83�p�ۊ�͛(�o^gK@ ��M��n�����"l̳$�&�B���"���VHF�p���Ll��w1�8Xe݄����kt��n;��ܷ�e㵛=�o'gح>ed�$��m�rt�۝��8Şܮ�zq��ֵ����zw��k������[6��^�f�������v�&��v�+�阥�%S"�U]��Ӂp��
*I�ѕ�v�u���v�����}�r��iv3ۨ��ʼ	Si�8���X*��eLr�J��l�L�k���i�E�'cJ�h�N]��fJRoc`��qX�%y��RB���^�t!=�};� �dCN�a�M���]uƸ���@��jW�8���A��R���Q�V�xȕ�j-�.9�Q<���!���S�n"�oV�ˇY!0�A�L��%٩�Kc@�Xh�V�ۗ6�#��&�Y0 ���a]���fkk�&����(!D^�U6��p `m�� ��T��uC�W�桤��	�"PM#�� �=} ����3�kZֱ�f��azH"�2Qa��sv�7;��[�ok�@�򗣷A�v��7�zxfv���e�9ݱ��q���4����(`Τ��S��H�B�rݫR�Ms�+9��R����x8㜋VR���=�g�q3��xջ�oV��B�1s��+��%��3��S5��U�V�]Nn���Yf2������oQiQvrI#'�&=�֊gf�1Ԗ���;el\��Oh1X�΄�k�T�|Ť�i��31M��Cl���~����/ �Ȱ�ڗ�w� )WCi:M�bn� >ݗ�H�X��K�	$�� �&�N[��X[��$r, �v�����=�z��z��Jwc�7i4+I�X��K�	$� �v^�/z��H?&���J�v���I/ >ݗ�H�X��K�&�R]��Eq�γ7�q�5i�O�A T���d�i�ʑ�tr�'f\R���h��,�����G"��j^ I%�we��uj�ur�������C�xy ��C=OA]8�CC�~7���]� ��޼ �v^~�9I!h(�Sv��N� ���ݗ�n��>��}Ť��6�v�j��ܪ����~� �{��Ip��UIvJ�����i	��:e��� �v^�� ��K�ݗ�wZHI��k��9�v���1��s��,�zw�֌�E��e�M�Ϛͨ ����ӀnԼwn�9��z�ׇ�S���I�ZN�`۵/=U��)#ޗ� ;'� ��Y��9T�#�b?U�I�L���=�~0��x{y��Q�r�\�U�\�r���, ���5@��j�ڴ�Վ�v`~K�z�y�, �v���N |��ثZ��A������%z�ޗ� >ݗ�|�"Z{[uM]��6+�9�(8�E�a��!k�n���D�
�5#0/����-�	s��
�|�+׀I� �v^#ذ��d�!4۰lWWx�p��e�ŀnԼ�ԥ�ұ:N�i�f }�/ ��,=ʪH�+׀OK�} %��s�Sh,-��ŒIkrO~�_M��BT�(�j�S8�9��krO&}����n�hV��X�ڗ�{�^�� w�׀H�, �V˺)��wn��cN�����'�����{��o�!d���q�;�V���Z���$ۆ }6^&�0��x���+�v��i	;0M�����=�~0-���m�?r�����j�kVۨ#��w�߷�uvJx~��K�~��I��>�-	8��Ɲ�k �l��}� $�x�ذ��d�!4۰l���>�E�~�8����	��"�>�s���s�@����������������G2��V��u�]��8�rrS�� C
�+F�0e�m�K+@@f�L��J쑖o	�Lj�l��%�D95ƕ�sb�y8�9e9<v�ˬO!�5*�n�0�Z�oN{���e�fp�IQ"��}n���cg���6�vP�֦���mqmAfH9��Ç����Ν����b�"]F��T��u��\L�Xb.aF�;�O�M��\�3�	&f���Zjh�%���"�����h��(��@�JƉ%$1��&�3�me��o��￞�������` KT���X[��7^ş��s���~��o����	6^~��Og�}�6b��.3��>�~����X7e��c�7\t�T��v��o �9 I��[��{�'�7���ۀ~�?R��9εjir� I��]���ǀ}ŀI�C�\�9�E�cu]��i7	\``OOOBg^���}��:��õ�B�J�mi��[<��ǀ}ŀl����P���b�lWo �lx��WyU\�W*�w I%����qV�HBi�i'L� �=� $�x��x�p�7Fj%�c����Zn�`�/ �ݏ �^ŀ}ŀ}���Nq�m���Wv<��\�����X��vLV�un�N�V�����T��6�[	��;k�C�;CDl��:	A��l˘�������{x�w�� �v_�U��y�?:hC���v�*���>�b��e����kذ�j����ڱ�wk >ݗ�j�f��fͥ�l¹��&?�q�w���rNw;�܁�[8��cN�M���ױ`G�`G�`{�UUJ=�xd.����cT���>�b�>ױ`���-�����V;\V�'v��ld�V��2��I�<��D��n�{&�l�>��p�n�N���>ױ`���-��ʮz[���ǖߧq����j�S�n��y��*���'��9�o^ŀ}���Nq�m�N���{�{��<����ڻ��������UU\�����Ms� ����OP��/ȏ�'��|�G���b���ʵv��ذ]��)���b�=�g�5wE�[N�`d''1��۴,`�&E�C����]�)h���r%�� ��b-�����,z�, n�6����v�����,Wv<Wdy�W;�].	:�!�V�wx��,Wv<Wdx��xx��)�)�݃��v�]��]���e�{�T�.y`�Ԧ�H����v���"� �.�z�|���I>7H���F �$�J�)��� H�,U ���0�'$/,�?>N�*�Xq�%v�G�=�5[9(��v�>�����bj�6WKi*�VٝJ0�4TV鄚�0���;��pn����PP���ˣk��v�l�3�0(��M��E+�lݕ�v��ڐݹl�)u�r�s�B7$͡w1`�����ɦ�=�1ؼ�9�X.�w���,]��@�lW>yv��P9v��o����ę���H���P6�����ɚ4SZ��5���������I��#vy.�l�k76Ns�p�M��m�ͨ-�����w ���o �ݏ�W>A�� ڃ��ݫ�nݻbt���;ŀj�ǀj� �vG�N���m;i�j�`]��]��.��Ǳ`]5	�J�&'jĚ�xQ�������,W9ů{�p�����WU��3Wp�����XWv<Wdx��'��6x�2e̫q����4W��U���c�6��km0��b�_t���Uw�>��X/�� ��V/�^�(m"P��3fY��ܓ��f�Q$ hEv�R������3rO/�}��y�~���rN@�O�ٷЪ�]\e�[b�y�.��	�b��e�@	V��eZ��]�v��dxױ`{��=ʮR��y�P~�[��ڷn؝;v�	�b�=Ż=���>]��ޝ骑�Z6�X��*���15E�iU��"Tm!3�4*��q�bՃ��i��[��X�� w�/ ��<����A���H���cv�M���"� �M� ��, �� �[*��Z���V�ڻx��xױa��̮p����k�5R+vz�o���Cz2	�	��h	�������㘞�h�x�<&x�D{׹	4g3A�゠��V����F F��W4M�p%����1�������R�\��LK�௠��p��8� �'��U'���7��[�pַ��i�C9a$`�TV1����|Z@�<6��~:=}�4O��rfSA7ǚuv�iD�N{�Q!L<�
a 5�8� D��3m$�ͼ)"��h��{�@�Л��>�5w}�#��
�ҞE �%�s7�nf�3Z�t���"A&�D�r%-�S��߃��ـ� ��"��jh�T$n��D|(z���h�}��@|�\Aj�O�t����HAG��c�T�O��Q��{�k^�rO/����s�e����S�J�Hww��U/K�X6z��#��+�w�׀o�^j�ct���n�`�e�vG�M��v_ ?��:�39�6�6̱Mf4,HD���@Gh�-f`�U��#��w�l����%͌����"� >�/ &�Ur���w��xϰ�Ժϩ6����ݒ��e�{��]��T�����;5�s�����{��Ϟ�������x뎚ܥm;i�ww�|����#�:���z�r�s��Up#4F�G��!!5� !��&H�US�
Y���l]<���cv�!;��I/ ��ǀ�/ ��E�z��n���;VՀn�.�ˑ�b�]�-ˌz�]�]=>3��D�j6eq���+�-nW�o��~� n����}�^���'G�ڥi�J���2��ʤ���� w����س��$N(J�T��v����~�����w�b�7ve`Q��t�]X3T�O-�NN��|�m��w� �ٕ�}�"�>�(�&�YV�����n�̬� }$�$���T�C�$�צgu�k	b(�ˍ�;h���5���6�g�� SF0"�W��Fzܺu��밗V9Ҋ�$N�]��NɘqN.m�������6Qe��]�`*ڨ�/�t�<��њM�ص=C��dr���et��[���@��]yux�#�a�W[*Yut�3fvBL�<:�=��x��^�������y��Nywmv.�D�\�����fe�Y�d�֨��G�E7�]�g-���vH:��\q�s�7��x"�Y�;1ٙ�o\m �9���s3�b �,L}���߲��Ȱ�%����<���Ml�[n�e]���� }$���,��+=\��H�O!?;n��ݫHN�`g�xu�Xu�X��X��Ƭk��Z	��/�{��vŀ}�"��K�>�.���J�&��n��{�� }�^�ݏ �}�S�r�YteT��7g��J:�����7�M�Kaw�m���v_gRx�V��wk ��E�l��uwc�;�b�6�[M�Rv�Һe��� }�^es�q!,"z6�)"����E>P> ��M�9˹'�g�]�9�{��J(�&�YV�����v<��, >�/ �#�S��ڶ���5v��ذ��X��x���q�B���m2�v���X��x�v<��,�\ﮗ�wGڻ���SCn6�ˢ�={���eˣ���(�t��d��QvJ��v��Q�2��o�~����xu�X��, �[*��[���V��wx����,�{ }�^��t��JV�Ɓ���{��=��gN��T�U(#J�	肣��� .Y�7�n���y�j5Bi�N�n��X��, �d� �v^�{+Z�nRV���-7v���s�O?������ �IRT����YV1�l���7b�ܻ��5l��G^��R5* ��i�2��mUՍSh,��-�����{ }ݗ�w��Mڻ-�wln��x�ۆ��� >���>[���M�n"�v��f��� >���>[��wn��I9v�[�.�hN�`��x�v<���ꪴ�Us(��"	��_ Om�k�$�y�˖��Љ����{��'�=�x��<�����9�s��J�WGj���������vQTz�eL��1+56�4f!H��<"��C�̠$�%˽��~��}�b����ʯ�v9�NG<��t��ݗv`kذ��z�,�������9����f�B�F-�6S ;�׀o^Ň���%ݗ� ���>�(�U*Ʃ���=�6�ݗ� �M� >���;���]��;�7C�X�ۆ��� >���>ױd�π�H�҄' �T � bB�+(&(0�$#L�fgڪ��x����7>�f)L�\G8R!���+�:(�i^dwR�@آ���Ƅc�b��tA-���FҬa��t�ŐK]��e��;�-�zt��ۙvJV��q]��T*��n�b�묙C����J�Ѱ�KG\EhB��(�h�
+m"X%7Q	�O5E�w�|v����nn�훮	�1@����K�+NNrO�s��s����������Y�-��6�f��bk���3���;�N�'�s۔�m*A���3�
SˌV�N�c����� }ݗ�|�c�>�N��{-�]�T��\���=�|�c�>��0��X	���Wv�-Z
����ݏ ��p��%�� wg� �CK���-%k��ݼ��� �^ŀwe�-���EA6���컳 �^ŀwe�-�����U]���H���AiU��T!��-�6&U����dŗ��0�%�,�4���wWc-7v� ��^�ݏ ��p�>ױ`mm���cT�w{�r��پ�:g����	�0�H�B@߁�Cq�	�hB'�'����`u�, ��/ �#���v];v�n��x�ۆ��� >���>[���T��*�c��N�ـ}�b������x�ۆ���NZ�v6;Bwk >���>[��wn��,���e�WI���;*�Xĕ+,�m+����L�a0��~�1��G�s�֍a�M杫MX��j��<��� �^ŀwe�hit��B������v�}�b������x�v�A6���컳 �^ŀwe�9�*��B�Y	E��к���f���ק ��_fݗ\U[Q�[������x�ۆ��� �h�Qc%1�m�����v�}�b�����{�+wBb�[m%i;�H�2��4�b��"�K�H}�����ns�H���V���MW�޿N�����we�-����PB�Zc��N�ـ}�b�$���:���>��0]6[��F��ir� |�� ?��� ��p�>ױ`&�+w�Nզ��ww��R]�׀we��>ױ`\��S��АʘUP�<Pݾ��nI�j����p`�� ��p�>ױ`��x����SaMR�	;uN�RWuAƚ�@6�/��5Z���گ`���l��sPՍ�SN��eݟ�� }ݗ�n��s��~0T����wN��Mݬ ��/ >ݗ�}ݸ`kس��GjP���bT�I;x6z�	ݸ`G�`wc�;��v�ZwnՍ�]�s��/l�|�v<Wv<��(!J�i��Iڻ0�ذ�r�{<����߻z`��Uʮs���AW�*����`AV�*��AU�*
���_�"
(�P��AP��AP�#B
$��T"T"EP�	B(0T"	B 0T �B�P�0T B*T"��B 0T �,B+BBB!B!BBB)BB)B#B!BB+B#BB!BB!B#B
AP��P��P�B AP�BB	B@T"�P��T  �P���P� AP�B"�P�P�AP�AbEP�	B@T$U�B)B)B(AP�EB �B*#B )B)P�+B"�T �UBBT @T#B)B0�AP�� �P��B*0�!B,B$1T"�P�P�B	B$B0T AP�BT @T#BP��P��T ��@T"+B @T AP�EBAP�	B0	P�UD�	E�P�BB0��P�$B�T"*@T"DT")B @T"�T!P�T! T$0$U��� �
���_� ��AU��
�W�*��AU� �
��PU� ����_  UO�U���
�2��Z��������9�>�!|2B"�!"�$�E*�D(@*%AP�%D �)$%AP�i$��  $���(
�����@��P
�H��@B�R�ATJ �T�*���U*T�*�APR��)�       �@  9�}�]ﯸ�gw�-W{>��y�מ�f��s��;������hX z8_3��� 
�l��h&@{o���Ը��i͟+��oUp ��{�m��3�y�]�ݼ�uo&��*/  p     >��Š��T��Y�=.}�vΧ��y��� 6�U����wWx��Ū�n{u*��ޕ�=��>��8  �������ڽ��窭�����㳶W,�e݊����1���^C����.�k^� � I    q |C;逸)n�0i@�}(��悔�h��(��� R�ܥ)C t�JR��OGJ  ��`�
bh��=5��R��e)Fvt�Q͂�(͔��  Kw�(��P��
14� �`    u P\0 ����
x��.��O,��uzx��� tX�.������}�W�CK��+����*��� ��a���> z�<>����<n���ɫ�\�=U�x ���������t���� | �  �� � �ƆO��q�׻@��OA�����T����<or���n }u�®/.}�s^4����۽���}n�}������=����7mŨ��C����!��w=� �x   4�3�T�   �РIT�Ǫ�SQ����Ob�Rl�� �S�BS=J�� ��jTS��0G�u(_��O���#�~����Jc��"���DB����������PU?�QQW�����aQQV�������)mC�S�1���E���cR@��D�W�)/?ן��f�^H|d�o�.�0��gh�|�]ǫ��Z���s��"���bj)^I��ぅԔ�y��%��Jf[pq�����2s{�3��Zni�,BqA8�!Zl5���7��]���<��wK�O�L����{��Vw��\UF)��W4��̳��#k����T�Qa�UC6����6f�_~����o3[�xO`�3C�2y]�2�g��ўS��Ń�B+`��������g=��w}�oWZ.��ь"���v��8(��t]1L�\]�5Yu���O�N��
5��a�j�ںX,���&�^[�pւcF@�@�8ek��g.��j���C�B3���5�gSJ��l�)�-!���|Hr����V�*��)  R1c CL�h�K��kB �
$�EH�k�!�
�HB!R1N�Y#�A�!��5��|
�!�k)Ij}��L����\��Sۛ��8��}��w�]�~[�+�nߪ4-Bh{{�RL��I۸o������3���jCs��v\�O6��97*3z[����SF\�̱��zcF"T(@�dL�S
�#YF-0&G�u٤����ޅ�t���	<�HMEP��e��7�z�pQN�)�sC�9+����==L�2W�`Ǧ��� �c�p8B��R�P��5��XѮ���{ҜMvY�n*9z��Mw|�xI�ӛ�:W����D���X��3��\޷w�����i.{�Ǒ�;��h%<nHg��Nk��H�Sa��.�,%&:�,17}��],#����)�f��o^Д��4�8m8��
`E���$O�za��
]�$r�Y���k�k�]#,�ﵮw�s�x��6�a�3*�Z\�g`�9�DDuf�uV0�!p��5��bC5.i @�������s�D���׃�y�0®��!w8��B�-,Τ	C�(D�RA�I`�-�`�,dd������F"$�c���&�߰��1�*B��P�4�cq`�F�S�o|ZM�TS8�n҉1�!�I]&�7�ۺjh��k� ��B<Ņ�$5p��NS�ɗ�p�ܸh�!�	�W�\S{� H&G\�-�]HC�5��i�{��E�J��L5y�$I$���V4���c�yt�ǂ���{�ػ�qlH3z�ف"��akL2�(C1Ke���7��F���4���8'1V��sh��V���F`���S�{|���5º��_dć��ֺ^ni�W�t
�k{֖�vo���r`�J�×3�H̘ĸn��i�7�o�l�g����'� ����EL�Za��&�
峜��h�A.0J#�i
��&�٩��F�5��zwL׶��W�n�w��搢Bdޓ{�%��;�&�پbX��s9���Si�Qe�2eIWJ�^�֎��dֳBMJ�k�����q� �v@��o(���7���ZV��n�=����搤ҫbռo������D�o6n��a._hCc)��(��a*1�0��V��V����$�7�z�z<�n�jd����(�]BFV��	D45V�[N-�ڂ�b��w�i��S�F\ѹsCY��f�0���#F6H!\�YI��%ā��"P��	�H$��#D2�B!��I�`ň��I
��LJH�:HA�R�q�h�a�&�a����b���G��3�G{��h�x�y�0�vr3��kc	{��f�F��ѩ�2��a���3n MM{}��r�>�b���P���B48��B��W��Č�GZ!rp�T���	XT��Old&��f�i *D�B����h4k>;{����i�M]�S�<�G��H$���&)
�K���jIsR�f"���um>�mq!HʭQ*��I40�Ѥ��;y!���������U�.�$tJ�և�0����W�d�BB# @F
Rp�w��&�j�v����w9�=��|(أ���[�!������gw�8�䲷��W��\� �%�so�*8T�X�CI�>bb@$Q[y�n���c��Z�O����`�U�+F[���j*�з�b�[�[�f�F�W��m �*}P���G3�Nw����g<��f���xr�,ki�cq.�����=}#��{Ϸ�(�^�[H�\�i����7�@c��F��8lL7�s�n)�Fyb�B��BO!I!|Hā�����s8ɧ��!L���F���������V5�F���,[C�6�ڸ�(c�hѷyqq.+缌��}8o] x@b�xE�z�]}�Hɭsk#	v�c�X#����s��!��$h�$��c+���*0H� @l�l�a�MH�`8Lh�D���j�0�S.h��3�a�'��<��p�6�
¶�[4d�y=yu�\֊��#	���CȰMA�n�7�1㲙���B�����ǒA��.y�:�]An*(��6���eVĪ�%Sh��#p{��S�������i���%nU]쯒��Y�nu{�jp�O{]��g�M�1��ĳ����T��+�|O3��h�ui���ב�s�zA[�N)uw�{���\���o���A�!(�����P�4����aqBJ����	"��	SȰ�@�R�Z�FHU�.��I����;��!r�WP�SB�M]8��5��J��tF�WfLɾM��F��0����ZF4,�d�N\��q��ohNnb�iSKHje�h����v��4D�[��"���hM�]iJ�B��TZIU�����GR��5�����I2X�0�vB��rI+(h��
D�VR���S��!"K�$i/$��졣�院U��a�7	L!|�{�7|�J�jf��x-gWf��ɔhT�HBƷ��8�n#��D�u���k҂�w�|�[.�f�P��FcXa�)�3^��e!]nH%3D.k��߆8h�K���S	��FM�jI$�%#I ؖ͒��
q"@ �[������"Q"@!� Q�%uā"C���A�"��a��&ͻ����B\L��$���#RFR`汁K�� bA�8j �40��0��5"\�I�=c�3$��! P#M��9���]�q��˛�$�rЁ��@�0�ND����g��߫���k0!=�B͛7��fq��U1���Hin��S{�ޗ��a������Г�K�a�W���H6<vX����8l�#�rI����O�i���4}na��a���f�m8p$�0��h˓Xdߙi��=#X�$�+��� ��	J��y�ơ�H��ѐqa@���B�t�`f�r����޶�H�J�ǉ�Y��|�ٜH��R��2x�.;�q���
`F���l�!�C6B膶0!
�1`@��,ш@	��ط�h������E�Di4�3Ft[��{p��0|[&.\��o\]H�kY��@H�U:�qZAZ�[z��/u���v�����]].�5��PB�9;����ZHMEu�}OXU-o��>w;����|KBI��v$�M
]�0���[
����h��t՚����3�Z�&���#BC&$�}�eZ�����q�OZZ��j
`��H��F��Z�s,�Z�vBg9sE1&�CQ"Fa��<t�]�*�xMk\Mɂ�����(�mw{}��[Shr��\FM.�nim!�\�ETWc��	�9wA�R؜W5^��ʪ��\�˭�f<�f�2�1j0���(c� ��HO�;���khN3Hgx�qY�$>�oQǪ��ŴR���4�E�`���
d�ג�M�6�l!��X[��Jo������a���1wP5{����IJ������tHF'�Y�$eB����	sF�ܚ�R}�a�k���#�$�b�H��2���f�Y!I���<��HSh0ɟkeaP#Hۚ2� ���)������Aa���ZA�.�sUhq"�%Bh�``�L�fw �&��z[�"q�	�Ņ\u��| ��J$	eB��5�i��פ�g1Cp��� ��4S��j;YX��.kэ)2D"�H�1�xE�f�,���i ��0%%��u��!�4���ap��N�k�0�I�]�)�!EkcZ��ZQ.YR9�{��{��׵4
a�'���͙�C6i��9�w˷�^�;u�s1��(�ζ�[�`��3*i��7�t74b�����Ꞟ��7���ͫ��r�H��~�҄���9;�9��mq�0\�Bi�B�.�,������!*������s\�ɤ*����\pEK�;��Y��!v���o��5̽HO"�M]��"j�0��v�$��a @I���ֵ�^��������V��C�;���g%RwK�ŵ�׆	9�.q�S�k�����e���s��s.��-3[��3G�rs<�\0�z{7i�B�1��K\E�\i��mbFUųU�i٦�: ���+bmqk���Bn���ߌ�2��h`T��
��D� 	$i
� �,B����c��$�  �aXT��00��C%$H�#��`"�@�Ç��浬9�zs�
Ô��i��@(�$B��������ow��4gQ8�:�Fjk������ޕ�/����[@h       -�� 8 ;9g88Z�L�6��Luc�2F�[Y��2�����}�A!��,� �pM�H�J�MkN��U:H�Q�V�q�Kv�г.Im�{*��,�bgҍ�z����v��cx����w<ZS�SeD�Z��(�:qSՔ�t��
���IV��`�����y/\x���c�nM��P$�{(�Ӛ��c��G;������A�Ôr�s�pj��MmU�/�C��A*�oiU�V8.VPێy�l�vwl��-��v�$�gK��1�J� V��?s�XX��v���Í��1J�,R�V��	V��mό��u�vvW�;U6��r�k��n�Y����5vc+��nm��m�7h��0�7�%:y�ƎNu���kͤ�K�rB�ZF����v�1:�<�m�+U*�V�%����v��}��CW+�:�����85�tF���YW p9#i��gj����UZ�G)�!�iem��Ø
p�8�{[l��w�U�[G�hh�[Z�[@-��j����]��nf��Y����A����)3��d�zٺ�;m�- ��r%UUT@�5ԫWb˻t]P/l ���t����/L�
��F�V�Kkk�sT���O�@W�S��HS��Y�UQ�N�� A����$9�����F��o��k�j�iI`�CT���9w]h�h����4�:�L��*�Z'DҪi5���E�d�ӄ+��V���L�N����G��pZ^�öVCr9��u�S��:�VA�@���������X����~U�æ2 �^��Q�+̓��]�x8���p���'e�.���cj�è�Z�L�aD�޲�����`w6��Fx�'�zڥ=E9l<��*������qUU,$ z��Z�	��Z����X
�y�lj�Q@���G@)���fH���Ŵ �B�V��^ �`/F5�R�gN�Ͷ��u�+2u��`-��m��n�ݧU՜��/HHp�;-<�+t�<�L�����l�M���Z�p2��[h
�����:�؞#!�S���i�g��w����UU�ʴ��� ��ր �m�&�WH`s'K��\�erK)i��0sl�i6 j���m��$H
��W<g�'���¶�Y��[@ K,����K�4kn�M���$镭�p5K��(6-Q���k`*��i[d��ɴR��z�R��(��q��amm$gX��Ac�=H�S�(�C�P��p*��3ِWz�	&۵;G@�B�Yv[�Vv��kt��Lm���g�X#]�:��+����$�s����p-��/E�4�iQ����\;mvN�K�m��E܍Ŷ�vUjt�u�MLb� �\8�KĽ�׋Ý{�g���`(�t�댼��mL�O��l��'>�n���:m��WX�t�H�ڐ۵�$����N8���v�<�f�9�m�[�[[U��.5�ܼu<�qݓ*[W���gW=����ac�	웷Kq*�<�'��/p�� ��r��N6��:�'5��������iv`���*@�C�&��*����r�$`�* �l9j�6�
T�r��&4�]�W>@��Z @��4�ZRN��n�g�:r�r���	i1���Mu�)�i��5K�8��]]�6n�	��l�F�N���[t�;��*��&�䖕h��7�Smݡ:�L�{�u��l���'@�b��	-۝�$�f�pY-������U�U۴ gW q��ut�n�t9��NB
v��(���MV�tӸ�햮z�B�k��l��n4Q�O5�N����R�B[T�`���nhn̻-\��%�*���aiV���u��B��t���K���g6^X�ڭ�^@�جq��')��� � K�$u��L�l�� H��p�n�ln٪�U����}�l�]V�t�Uq���2�l���$X` ��9Ėյ	��N'j��U�e^��;.�[*��!V��T��X`�4�u��m�$�J�K� -��u� �Im 	m����m��kh� �[pr@[@    -�  $H l ���  z�:D�f�1`h]�����9�iW��q���Nn�]���NnR����ɀ�N�� [�m�]/[z�` 	$�kSS�mI��[�H	-�� ��[%�@N� �n�  �H"I [@   �J � ��G8�d���R*֞�Z�ڠ *5��-��� ��[Koc��ސ jӦ[%,]&�l޶�� ���k���2�[� )V�с9��Y`�ڥp��5[�� m  �[s[�}�� 0 �m��  lhp$d��}��$6� �@ ��@-�&�K$.��M�g8�`��l���z9��V�%�m�@   6ڀ���]�����-0M/j�(����i!t��n�l*+P�U�ӻ'F���Mp�b@qk@[@+5  �It� �m�I��e��@ H�Āj�P��-�Z�ꩶ�I��L� �Y��   �l � 6� m�ZN��	i�8le��bAm�7e���m���9� *vߏ���m��b2�4nY,�gE�Z]d�� �ã����U�M�]T ڤ��F$���f�p-��,1SY��mJ�{n�V�1����݌��p�ջp  5�؋,;)��{eUz�U=�#[U����m��%�]��� �I��&e��K�j� �m��[6��� ����+���1�Bڠyey��<�8�0&�����.7FO-�h�F��8�lq�z�Z�@K�A�ۮ����F�ʄĻ��e�ؖK� n���P�Tq��&�@��6����f8�M�i"�:kj��[]cp���L�u��>���[]J�Ĵ�	���ev������Y:v6�m&R�8K+�u�i75I�D�Ƹ m�l�U@mm,9De�n��ck��ݷi5�N�  � &��յ� �I-��h�%/`M� �;j��E��I6� 4���n�a��ph � � �� k$��   6�0�m���m��o��'fBϩ��U�RZ��e��Z0���)-U��*���]�c���K��[Mk��Hp    ��  �4R��UUl&��4�k�[��J[�biV�jV��P�p1��85�!�v�i:GU��	G]�h ��*ҭUBO�٪^q��i���a'j��7 �P,���t��	 �h
���ӫ���ꜙGؖU�j��*ZӍ\2��J�yz�MT쫵/<�c�a�-��E` *s��ܻH�mt��V���p�p	V�;;`��m��4�ݷ�m�u�����( �UUW�����檩^v6��-�4�I��BGA�۳V�Y;^�ڃb���j��r�V�Ɇ(�YyP����kָ�˰ -����d�9��Zڪ�� I"Qz�� p � ۉ�&9��$m&̂mr�r� ����݋�4&�UP"�mPp�lh�P�V��@utK�ݷLm�-vl�@d�n΂D�<qd����O�﫫m��i4����6��#���tv78��1%�[M�	��j�v�f�rdP麔u!-Ut�5W�m����� ҪRZ�������!��   � �Bi�����ie��s��	zI�h)Ζ�uM�T8��y,�۶�9v݀u*�m@U�\��mr���]��Ҩ�����$�-��m��l��6�c�r�PT����Ҹ�@  ���knm�  �v����+��UP ղ����N #]� m:l�hD�Bl��[oV �knZY�� �a  �ݭ����6͈ �5�@I $��dm�	���Mpm�s' ��>}�Ȑ��@S�����l���^�f�{X�E�;C�BE�085�+*�[��8���+\q��J��Ʀ�
���0�p�]��UU��5����8:�:�  �h�S�d�#�B�l�:t�kͮ�ڊ i6�wk�v[�� ��PQmn����d��6G�,���:-�E�S�tݯ` �i ���:m�jrܛ�6#�m��9:��ֻi0 P��l�@UWmu�`�Qy��@�'m��+��U��v� �lhŅ��*����Uy�P]���!����,�̭K̭U�ښN���A��tga�WURv�4�ķJ�U�f6���6��E�p �SU[O'�A� m��i[j�@6ضC`ංC��g�m�-6�d����6�Z�-�mfvn�(����0���t�B���[Uܤ�m�լ 9�ٶ�c�BmsD�vn� ݲֶ��/>_��iY%�20@4��m��>[F���\��m�m�	��m��a���m�i �2�ZE-��h�H&�m"���/6$:����٫����]u5�[�5�p���d�\@6��$�8�F��U����*Om��]Pyb[X�<	m���+SOllM؞�h	HM��3ʴ�\}}���5J���N���b*�왦�9Mn  ��n�&�����u�����J����0�A�v [�g}i�m��6��$$�Xf� 5�&f�5�� ��mCB?�M	 P؂C�_�?�  '��1�d�H0VwV$!�
����Rǂ�#T�����&����Lh&,P< H
�� P��A(|�h<@*���N ,US�b�a, �c�����È���M���B	"�b)(�*�j)�|�I$!  CJ���&�b�`'6� @��~cQeh ٷi�	�S�k�E"�U=��A�� Wj�(��C�R��臿+Ǌc!V!T5�@�~X������ �H*HA���Qt��.���<W��Pc�~ �-����Q_ �� �,X�h�s�[Q���� <@t1">/� � �H��"0] ����_�z���T���� 0_� �(�߀*4M*�D�`���	D������A]��O^(_CRE�!D�~J� q=D�Q4�/�8\�hP=>�"f�OD �P�GX��<R!V��
���� * UB �<Tv+��>
���mC@ ��������P�! �`B#Hd�$&!�
P	�J�W�@B`�⯀�"���d���`�6*:6�O~T�H�*�| }G�RD"�	m-ZE���!m$)��eIiaZ����#O�OP=�!!"� �		"��F2C�]K#F1H�ER�@U0 ���!�d	$�|�TW]�� ��4(% �>q�}!��EE_�'��A��H�e!,���x�x�g���V��S%��z��n9}p��q��ms/s'mu�����p�v�Ff����/mK�g�vP��KGK�ˣ�f�⇶{i	p=MFA��El�^�vz�Ȧ/]i{\�ˊ�pp���w��̲��@��+���lQ��t�R���j|���-���9��畒-M*Ke�:��.w<횎6��狇V+���G��rl�grcJ�z|�S�e��n�ZɷV5��jZ�$3�G%�ݎ��3�u�Ƈ\���n�"��;\�<�����g,�z��nz3��(,�ݱmv�81��]���m��v��F�g���s�.�s؞�/gC�:�l�n���_Gc���V���g;���:��ڱ����gO�
�tڜ���';jÅ��u�CS��nL�a�&I]�kI�5[�u�:ڭ�cs�=v�Aiq�[aV����J�gi��kj�#�lnO;<�#(:$2��&�zUZڔ���{J�s�m��ӱ:,�ܨt�v�ɸ��*�I@���ڠ�qgYN۱���r3m���qĄ-���gZ��Q\�c# ��YeU���u�8�LP������m�lU<�`8�m��P۶Uxր�v媉W�ێ�ɸ���VS*D�{s/�_O\<�Ss���{;[&U�v��aV��,�5����Ĝp�UI�mEN��K�s�yd��O/K��Á[7:��l���m�
���u�g�L�l�pk
n7:�=g˯N8V�B :�Qk9&r=�2o:�ch�^;f��r,\�Э��en�}gcR ��Vvӥv�.Zl�-s�pr��ڻ$����֖�4�4�MT�V�����1���b[��\��[��6Sk��<�ç�r�kv8��$����f��ٵ:�7.6]m�[kۄ'�h&�gt<A��[�֐ꥍ�[���T�= 5]<��m�̭�Q�Gf�*�Rs�V�k�]�vp��7hn�'-�R���9�X+�R�֦k%�j殳3QC��6�T��C�i\EO��<�x���(	�?���_�*
��1�|Ȅ��m�[\�r�%�l�ol�z�k�㰀躽���c� >�n�{v��.�l�8�.F���.����9NP�f�9��t5,�q�R�sᛓ��vm�M���.��l�JYmcY���<p�F�rĮ*�Pp7"ц�Đ�Ǡł�e�z{rcq�jn�e�{s@<�C͹ك"%/�c�6#s��[�8`�����ǻ޻�����vp��&0nr��Lrs��W���(�n�ϓ�m�˘�P�"E�˔7�����k�����{ﴴ:�{�,�:KA�9&�w��@������� ���WJM8�l��'&��k�����y�4�h8$e* ,��4����/;w4�٠��@����
��!�6,Q'3@/-� ��x��:�ŀj��V�S+�t�A����y�m����g%�E��p�y��{u#\�9�S�%\J��`�����U�^[�����U{��-ev�n��gW����;�o2��Y4)���	�.jk��f䓞}����]ΝW���U���U^�|�ŀ��2o^�����;=]�BH	�ғ� ��h�l�/_r�~���}�.��(��C�h�l�/_r��s@/-��=�P��ve)kh+r[���;�7%��ʚ��me|Och�z������y�%��dWp���=]�-�s@/-�y�4��R�T@Y1���ȴ��� |n������5%�ɲ�4�h��:�@wﮀ=�����E��lRTajBF ��).�TD,�Y�����9�Nݪ�%I1)��&�^v����@�����f��U{�	1�D��/{
���� ��h׶h.w�������ln���r�����K*���e��8�oG"��q��O���j�����74�٠^٠[n��Ws���T���T]Z�ۼ�	BS!�{x��hh�n���]qDH�`���>��o�Je��, �ݼ���T�q��C�rhۡ�w���rI��}��Ӡu�t�,=1��bKx���@G�4��(:G$p4�s@-�h׶hۡ�yp��\��6M���Bs�#�LJk*iF�d4��z�)q����8��gv���V�SL�UZ���^ q�� �x���{s@�y�Ǥ����rh/l�-�C@�-��m�֪�cj@�G&�m�yn������4���y��,��GP��45BI)}��`���]����U��E 7���&h��ٟ��^��n��`�x�i!"G�ڸ�%Xƽ�`�ל%n��`����cN3V4�,w,TP��C<-���R�Jp'&B3m��u 㗷�7g��̀[<[��u\���\�롐�E�e��Y�aG,q�`Mծ���~�d���9,bM�AS��khpwjX�vh�H�.���;�su�2U�ˠ�B���]��]ד�N63X1㓳�lS��fNƼ�n���F7@��-]9������ǻ��w��y:��z���Ŷ�8�z˓�P��3H�u,�Gn��g�^u\��DY�4�$�����m�yn�[l�;�:v���m48G&����o�(�^������]��K�LP�ۙ�w���m�@>��@���4�)FUX�hH�s4=�
gwv�����u� �:�`J���Ȇ���S#nM ����k��;μX �w�j�I)����73%UU^S�MI�Ż��:���*hш�Ԁ�����BH�x8�x`②�I����4� 6�ꄗ�5�����w5�[]vYeZ����ĸ�H�`����$�*E���3t�HHFCI�!��P�kD,$�mo@�K1f�I,K�on�7�}t��|h
��tȞLo)1
L��f�^����)�^[��w�5�dQET�Ww��!DL�{x5��>7� /-�qgN��&�I�Ȝ�תـlow~_ k{x ��x:�2��� �N���v�z[��r�F9X�Mvz/�EA�hv�k�S��<F맶yy
�`�۹���@;�٠v�JhaJ2��ƛBFF�h�l�g�ؐ[}4꧍�۹�^��
��R<J+-�@�}t}�|h��\A�H�H]���P�A}������9�.�Z�x`�q<qI4z�4�n�^��@�}t:���V��[lu��4׷s@/{f�w��@���8����M��a�5��7g۰�Lv��q<,;M)5��&����8�y����n���7}����v���S@���h�u�D��!94���H��x�9��� ������/�X�N4�C�94꧍�۹���@;�٠GDy?&UTȤQ�M�w�Z �{��$����ܑS��J�p�K�k3&���h4p�:�Q��"��X ��x�)}{ ���|�w4���cx�X�0MF9�6C&�t�F�q	����m�z?߭|�~�����5��{NӑH�)��'���@�)�}{w4��m���as��@�l�BS'5�, �{x�u�Ϊp9�'�d�5#����s@9�٠�l�;��hu�1�17����4������,����s@�1�l��� 	!94��xYM��, �z� �a
G�	LA	!��������d8t��Ɨ�,��Ɲ�\ܝ��ZiHW�굝�� ���@	v��Fs�w=n�
u��ڔ��&:��g�.����U����u���*��v�]�Kul1fۥ�Ì��JR�n�@����O�^���nw�kanuc`�Ƭm���q�0-jvy|�n�w]Q���d���N�r�m���
Ր]��<���Glvk��&j�s5�[��kR��W�P�M<��s���ՁZ�l�\m(�R�;D��!v�<]v�t������wN��$�P�NN���4������ �{f�}�t�\d��7��4������ �{f��S@�
S"�cČ���w�h{�4ԗxKW�$���RIs�:�Wm�G�L�I>�$��l��K�%��K��ǩ$�;�>�$�����0R9�cȤ�RIw���m��fv}���m��{뽶�$��m��\�@'�`�hm��,k���k��9Ƴ�j��E�t��='6�����7���s��{m�>�Ji���{뽶�$��33܍�t�|������R�9n7j��m�{���	����) ����L�)|���s7�f�^��}�Iqv�=I%xdK�F�����|�\o��I%����%�۸�$��{g�$��L�Y��&�hd�7�$��Z��$��w��\�l���}��m��g�����	[^��|}���m��w�{m�I�I��|�}罶�ؒ_�h�����z�g�6�n���E{l^x�n���7V�.���u�k<rv�n{:��#�L##s�$�{}>�$��kz�K�%��K��q�I.t�\M�8���ܓ�K������]�=���%�}��$��;g�{3�6���C�RLo&28ޤ�ޗ���|������7��e�ʗ���ĩ	��N}�9��m���³�@�k�%3B�
��������E�F@�,d�sWA��<����3ώi#%��FE�F\.D�_�����]��,�=���Hx��>�ISR���l�f|����7և����0�k}�DM�͇�!���F0�&�%�d� ��A�WV��ks�sCj�c4b��@��.1�	A�:��ך�%�lDbH0����n�~r�����X�p�!�7�|��V�;�2��S`hv�O�j>����\ܸ{��H����6!2'���P8�|��na���y��B*XIF@b]��	����!�"�no~�g�v�;�ˣZ]ňH{Ǻ�Ki-�u��+��\��4'�l�o�|�O�W�(c��/��*!�*����������) �B;A��>�0Ch��@(�;�P|�]}���-���f�c�U���eR��pv�����)��o����|���M��1Iޚ�罶�}~OB���D���t�m����o����$��Z��$�v�MI%���v��rvF��Ga�;��1�GkX��؀�y�K.��������v�n�N֭�k�c}~�M�����{m���T�ŹK���|�^��<���q�C"�z�K�%����m.�l5$��o��$�e����6�����J�@�k��m��a�$�9l����Ԓ\�KW�$�Xt�:E4ǉnCRI.r���%<�_Mn�o�����[xHC�%š (2� b$~CC���b�b�R�(q8 {��I%�?�Iy(%27$��9�K��|ϒ�K����6���4�m��`w��?��/�5dz컫�獘��^��ۦ�֭�n��c�7F��F�؞��ݸ��'�&���rZ��$�;v�Is����v��m�ޫ�'�:*����v��I%�݆��\��H�e&���rZ��͵���LrfRb�ԒK����$���MI%����$�۰ԒW8D�dma$�G'�$��ڦ���	j��\��jI%�vϾI+��]g���+����|�}罶��33'}���o���{m���wM���$�.����ݽ���c�GW]<��Ֆ���9G��T�F�5X�[�^�v�q�\݋v�����G�,�8��S_�;���"�Q��͡t�C��Iѯ#rX9�9�j8z�y���mDlC'GL���[&��C�(d��+�pz�p�mm���i���x���`�ƎZ1���ְu����ۥnu%��`�Dղ�,f��,a+�I5��t����郱&�{XZNnۻ���N��$�53$�f�˫.d���E�N�وq�%�,{L���V�u]&�=��뷨)�"<��	"����}�ԒK��|�Gj��K�%��I,:Q�(��Б0nCRI.s�}���G]�K�'���$�;v��]��<��c�	L��>�$���5$�8KW�/�}�ԛo���{m���DMN�#�Y]�i.p���I%�݆��\��_�v_)����~������Z�׽���}�i���bS��לm���M���}罶����ܝi��f+eq�=����z���b��f�]�,�gv�={y����Y;�c��m�����m�s���m��_y���������ߵM6��x����K,٭k\��3߮��!�
��E��[���^��~��P�m��w�{��,I~�k���?i�ܲ��%vWt�o�/��{m�>�f�����}���$u�)�$�0��/)YTPD�-�{m��'o��4�m��z}�I}�jKٍ����I,�<?i�$@n3RI|�k�����|��6���罶�'}�i����J/��8���n����s0����R-�TJ��i���=�n�k���w?f�>�G1`�C?��m��~wM�����{m�N�P�f�m�z���I/_c�x����?�5$��'j��ffcm.�l5$����$��ڦ������}�ַGQ-	c�{m��wz�����߳��9�IB%fq��P�D#3 ��R��P8>P�.���o�[����]��+o��OB��Ɔݪ�i��fI�����m����6��K�=��I);�M6��t��In@I����8�Tԓ��Ig~7��޶��ߵM6���}7��������WfT����$va+b�Q�\�qf�v�vS��h'غ���O��^>�_��4�8��q$�|O/�I%�݆�����|�,�#l������3��VXD�-�{m���T��~Y�Zu�����o� ��u�j�
d59�V�%�5RL�����Og �+�p�J"g������]Γ�����H�+�h>K}�����q����$�	JR��h�~���zD�aA�b�%*�
z�#��s���I;ߌ!�Br��Aez}'|��'����y�-�}�@���;�l��S:0�:�<�Oqs�րuٮ���ݧp�\oB����%�+�Ӵ����pv� w߿^��9��I$���)����8)-�mڠ�~����?,Id�u���V�p�7y��ɫ�K���q��岽��|��N������:���;>�V ㉡�L����*.��RJx��������u��$�
")�� 5��*�6�$*�������^�	��W s���>S��$�8� ҂S��Ϭ՚�i������.�Wi�;l7�q�1�{�����g��}nر嵋�ÝѮ��l
cG\\�v���� �-wk��.�6�m���ئ�t�8]�s�*p!<�8�ӳ� �"ZŲ�g�˸�nI@3Jrq����Lk�CA����Zwg��x��-ne]k�ݰ��3���;�����$vN�oTi�̲k�|�k[Z�C�j��=K.��Q|T�qu�F��3�����ӣ�&٭x�8������SU	�ۏk�����2<ՐzDdchH��}����X'�u�|����D}!�{��=)l�갑�b�������k�3�bRO߿L���`�u�lBJd5��P��Q�z1w�z˶�=��%޻�w��=�)��Zʉln�Yf��b�D%]��� n�Ӏs��8
'���Z-�-1��	)?5#�9�ڴf$�}}��O�}4�}�;��}��k�'\g�m���G�\�N�,th�<�ѵѷi�v��Ϋ�{����d���eհ4��u���>�]s�}=n�(_Hsi��.��LM��ۊ������BO<B�
�6�_p�*� 4#T�d`���t�v	]��"�d6��'�y�w}�7$����9���P�Jdr�u���M��
�w8%����a(�3����9G|��VQ�##BD����Q
y��puޘ�+�p5(���u�h�ʒ�mI50#�@����<�y(��3}<��Հ|�p��-��1h�}E���h�p\��Y�\�u���ר�TF�~IfW���AWYpvπ�)��O:� ��\�IG��0����.Z�n��pv����k�IG�%Twվ��o���u�l%';���)��������hs���L �  1Aq�D"e�H��D�`�"�1J�8Fa�:TЊ��f������{}���85�d�8� $�qh{?f~\��Og �y�X	%<�{8�����U[qJܦ��I�=�b\���`s��hs���T���H�gk���79�XJ��B��V�v�h {A&ݭb���Ŋ��ҴuLa"k�}��@}/����f���)���+JұXH��Y�6��M}��6s���w�@�s��~�ߒ;G�%�i����f��}~4�N�������ff):����������K∟�!��")�-������]s��;	&�,�B�F@�QJ!͑����|T�8��K��MjQ	'?}�0j�mU�ڠ����T����D/(P����x^��}�}�@�������Lj'1=���v�;��8��r��M:�J�nb9m����}�����C��!��nٰ9�_��v��>]��؈���'�k q�m��R���v�|��%�&�/O|�;ﴴ���_bI$����}���uX�Us5f����s�	(��7z`�ƀ:�S�v a&נ��dz!BU׾��;�~0��f�(�Juno� <�W��r+��S%�Wk ���`J!z"�߼p����s�WZZ����sV%F�	z��{��kO���No�V5��m���]ĦXZ���k��)�)�	04�  B(��"�����BI g�< ���w�8�+fg'� �כN*p�8E>J�{&Ϳ��}��R9�;p�SѲ>�c|h4)�D� ��L��l6A<�HD���#
ȁ\_�Z0�����4��1�H�!#R	1"H�X�FBHH�#B!D	�_~���J c���k���0�ɉ�I��6ςB0 䬦�H|��p�)��HBx��a� � ����*}�}5*K��ԻBP�����%�+fkp�HoF��>>�=	: �U`*�U�f�l8����!php��U������\�������۵��v����J��$�i���ͷQlg��l������q�z�'�S�9�O#6�=�IƬ������;=-�9�,<�����h;r� ,��kO!n��xmɷ�;r�b���v�g�8�������Y�z����q�nf3fۄ��tt����+P΃��ݛ��#�tm�bYc0pm�s��	�d4*�U;��n�(�j�O;�;;�\����"7.w&#�+���x�6,[=�>{y�v�cYܵ�L�=�\�wF1t�`�n���{l^��O<�@�����,��zxR��3e�=�.]"��:��:ȧ6�M�ٺ{�1�k�k�������w6��� :Ҋ��ѕkSKCMcm��E[�p��܋Z�[��6˹�.�ڙ'`nvBU�@�J��l�h���kqb\��h칙6�e��S]V��yb��U
s9,�WW8���U:(j��beݎɵ�!�3�%������
��H$ֵ�֓Omns�JW�55�YI�����WfIkt���i+s���[��v��y6�
���q����(���zX[Svq���4][A`�3Sμ'Z�m��6���=�vx�piJ�eݷ6{#��@`éy�SU&�I�ɑD�c����e���3��j�^�
CU�U!�у.���x&*���飍��������/4�Ͱ8����#[�M��yRsNwf���{9��eOWQ{sӝ��j�Pӭ0e�vx�(�j\�h��n|�.�m=���v����<��kr�R�9�mw9ODy$5��J�Xb�ہ.44�l�l QY�^�cb��(5�=i�\g����Z���+��i�Y��������]�����]E���g$YdKk�wGF��鬡:���:���P!:='���pb�{7c�] �n�p���$���NR������5m���î|�"�h�Ԛ�p��W�Ёp�p�B$�DL��}���w���~~v��M)]*� 	��P�(�,P4@>AM*}�0A�ڣ@ 3�EO�1�;>߅�̕2�+�{���郃��#����9���:��;_XGK��G�W�/u��:�7l���<�!�nm�CWek9�[F96{��:�#�m�G2�e�9(jͻi�鰅���ѱ��[hw9��+�]98m�P�9�eN�~���q��p�����ٲ�u.yz�K��ή��������"n,v�&�l��q:(\2u�8�a�0
Z\5r�Мؠ��7f���)�i�����[�n[W\ݪK4����/�|�N�t�,^� ֿ��x�����{\�_�o��`.�\�s���} q�� ��(��X�r�˃��]����K?fB�:�ذ����vٚ�%2oU8ګ��ʝr����- s����~IB����um{Ӏ}��TE�H���.�`jJ�[��9�z`.�s���K���4���G�<�R94��LT(�'{����X��� v:�Q��v�}83�y�(vqե��u�(�6�ד5�^����B���}�q�[o�7�� �V|���>�^, �z�У�r��o� huO����

�.�p�׋z�@�H�H�H4hЈ!I"��$V	��E�EDD�Q��M�[��:��|�M�z�P{I^'ũ.�)MԪ���w׀}��0؄�����9={X���bV�IRMf~��۾4e~��O:�b��{x�U��eL���pMـ|�M��(�u�|�����M ��*�$'�����ͱI,�ݶ�U㉆b�V���s;s��������ԗ-P��&�{���h�ﮀ���z"!z"(:����:���] ۷#�h�﮾������h/O�zo����b�!�}��,i؝Cn�n����|�M�S	8HP(\ȅ1j�	F|�����o ���D��W3RU�ݘ�	%�
+�sޜ��Հ�]�uj���4�j��@PUAezo�t,�����w��6�=�w(Y@LdL�Px�DM�2~g롷m�����cuZ��7KA�h�]MF��}��Z5�詗Okq�m��>�e4��^����]�z+��%�128@��$�>�m���L�ҷg ���`�]��(����?	qDO�9���@�s���&���u���;�����Tv�l�j��!/DBU��z�۾���]��@?-X2d��$"9�B�UJ��=ؘ"�~ ˯��Ǡ=߿-L,EQ�r;f�=޻�=�	$���x|W�8��� ����~U:���g;��7ڀ�qHO<ݘ�b�7P�c�Żg���{�./�'M�0I8���|���Z˶�g�߳����/|#ڏ���ȴ���<��%Tvwެ ��^��\��f~H<(zL`1���-��Հ�w��P�z���Ҟ� s��*LD���&���g�Ľ��v��|�����Sݬ��PNͩ���A�t;;�?ffg��]�k���:�ެ }�*�D(�Q�֚��M=�S�{;��\r�^d8x(݄�Mvgb�`^ŌAr+��=��/6�۵D�$�45�3��9�g��n���i��ù�AfXإ��1���5�O�AGR�ۮ�:�������Q��4�����ݷn��ɀu�Ki�+6���WrY
4��mmg��l<�Z9�8Y���A�3�"�ݥj��y�`��j��:�ƳŞZ�3�{��z�}ړ�S|��[-�9��s�f��)��M5�Ρ�w\+;��n�'��S�f$9�jT0r�ʇe}��l�O[� }뽈I}!�Og }��&5'��������:���2���27��	еH�������oo �k�p�J�4�ՠq_y���+qƈ�@�q�4=�O]���V��O[�Q	L�{x�{Q�A�DD0r-�>ՠf%��B�����=���u��al����(�ֽ1m�Cq�"��j3�����v��e"!$��f�T+����w?�{���w�s��;�4������
!��A����n��r \@Pz(\�k9۹'����rO���y%
�J*���A>��]U�������p�]s��J&y/v�z�� �|�cc��SvW��%�>iog ���λ��y$�T�7Ӏz硟��@x9c�h.���h��Z�}�@�8�\kBL2vB�fMˁ��ɧ��\Avv+қO=��p�������K1*��U�cv̀}�}t;]s�|�nuBP��C��k �tN�2����t;;�ٟ�3$�;�Ӏvwެ |�؈P����fK62B!��h�W�@�vע����c"�)Q�#&Ҋ�H$b�V@S&H��C�9�S�;����;�}נ�zѩ�8�v��bY<��X����u��B^I$���'�����_���b�q��l�5%	.�{?ͩݬ��u�z"!J���߆r��n1��eq�s�6[����J7�h�O[��ۛ�����Ikg�7�Og �ԷX����%������=��QLJ8��V��(�2r^�`���s��9�/D$��s���$P�����zW����^���Jg���ͩݬ�j�	h�V'_�#���ߒ���k�Zծס�A� 1�A��^�ϼ�x�~���<��#�I�s��h:���>��X ��x�(��gW�3�Τ�l��`�r��*�Z�6&�q�hLI�غč�H���bBև�Њ�U�d	l���}X��� :�aG�t�p�z�= ��ƞ(�z˶��g���X]=��S�Y�/(U@����D&����@�����9�ڴ��Ĺ毞��}�}���Ddj蝬IO]���R����� �׋ /nu�$�bQŠ}Z�z�B�=����X;]s�b�d/�s������:�y���<���Dӕ����t;H��^�7k�u�֍�SH���m�qm\��<F�x�{/k�ݸ仑��u�Nܚ06�\${\�N�
v%n�u�fV��Cقn7�K1k����"m���N5���oX)4�eݛ���,e���x����:�:���q�y9n��t� �^є���t6�y]t�S^��:؆+�:�����2�z����:WzAL]rw �[�j-HR��3&׮õ���x�bݪ2���4i�8�ʢ���#�pϿ~����\��C�R���]A:D8)_�#�/;w7ٙ�#��-��{X���?"L���Ut����*ʫX]=��S�Xz!L�^�`׸��Ւ�����9��3�碾x%����Iy(�]��N x�4~�j(����,�}呂�%���~_�Og �����Q�s2 J���?��^Է��&ۜ�Yk�2,W;{YLd]g$��'�7'�ѝ�qg?������q`v�� ���?�I}!�{��r[�����(L�U�9��=o5�IO����m6
��͛$$b��@���Xp�TLTnHq]�6�7�6�~ W\����]��ެ�l(��C^���L���ͩ����S��>��Xy$�#�B�X�����|���w�Tӟ�<r5eU�����:�`�u��DBS�%��-�G�Y�
D��H����R��og�9�=���s�}���
m&��눜=�-�9i�V�9;v��,�Xs��x�{t5��9�w��ݺq}��1���Uk�:���2����s�^J!r�۾ŀuo��L��e��AWs�|�npr�� |�ŀ}�ns�
<�����G�ԪT�ER����� |�Ź��`�}��ؾ�f}�G�`o�U��}��,a���qX3�Ѭ��@�I��K��u�4���GyN	�-�1�x���(C穯�C���Q�k���'��Y�4��M4��,�Ú~s\��am����a�&Tt�	!d�HD`rD��bBD)��b�H1 �Rs�}�xs/���$�� �6�Ei�2�}��d|���-$�ŧ�&�$�ʍ"����+&Ru���4ҹl����xX��4������h8�	!`E�a!�t^Zk�.0X��ǁJ���&a�����f�9���wd���H$�<����$�Fƃ�S�t���(|��b��GN��&�4��P�}@}U=� =Mi��0T�_D_8.�>Gh� �C�����@��������C��mš�DN��� �kvpq����� �}�0�c��J+�hr{�@|��o���{�M��s@��b��iBl�š�>i�j���dy*Sœ���:��wX.��=��2-�4-�4�1���_)� 9�� ����y%	r���� {�C�EI��F�R�[4������ ��m��%
d{���QVM�Ԣf���q`�78{Т"��+}:o���.u��j�mLM���%
'����9�=� ��	���A
@�AH�A�# �@	�{��h9T*�1�A(�E�}GڴID%=�����,��� �%ޣe}��nT�L�v���n�k.�l�/b9�r�2=���U��f,V+F�aLD�W< o޼��Ss�G�֯��w*���"6�(�ܚ�n��Ss�|�z� 9��5(�2rW]EW�uX�Ber��Ͼz~���>X��������nh{�`���QF7*���]�N���z�μX8�Z;�!TQd��F�N= �-�ވK�}���zp�O]`�G�D;����[9u��.��[؍�+�u��qV�d�.�=v�b-3�m̈e��ek�W��kٲ'g���p�vM���z(��.ӽ�@��g����:���I�	�@�7B'Y� �A�^��N)Į�X%;�:���:v�<{n�m���fK�Nr$u�KӞخ���-�8�v��^��ݠ6��5!�w<z�Nb�S%�1�f�/W3I��ݗ�����ؔ��If>o�;l�*�qWkσ���:�]dY�3�u���ً+vt��q�sg��R-����&�JI�?�����;V��j�s�hr���'F�ɪ��}�nsb��)���=���?~ďe��2	D0r-����u���EW���^���aq�O#�#�@�j�/;w4�M��S�-��S��jVSJm��Z�n���v{��9��-�}��o��?���������u��bv8&�fi.K�������|�.�V4v�E�'ˢ4Ber���Ͼz~���������v�s@/h0^�bn(��-�?~���'(XƁb��ĵDB�J�{՝��n,�Ss�s�QX�yĤJ4���9�ڴ���=��.u��@�|�j��rH&��A����mP9���@o��C٘��ڴ��_��F��173@��ՠ}Gڴq���s@9�:`�'1vlt阍Þ�e�9��Dl��lݎ�������یZ^���w�E�9�5���?�niOg �+�pμZ���kvp@׋��(�I��Z8�V�y۹�}�j�>��[��H;�g�@&@m<Q�-z���-�Oy�x�*�X�$,x�/�\+��)v"5+�ҷ�����s�_��Ђ�c���}�j�>��Z8�V��~���}��@��1�WEU���+�p�Q������X�v� ���&L9�1�L�<�tm��mҍ�l��%�j4���';���\F���1��1��q���s@����DyDB�|V�p{�u��waw5*I���jJ�9�ݜ�S��9�ڴܰn�d�F�&�hqڴ�]s��
&{�{8��,����U�d��AWs��򄫾3}8u��� ��J'�m� &��-Qy3$s�Z8�V�����}�οyhQ���B��LpMd���L5s��D����A���%�yو�5��q���G|ld��nE������@����-��g�z�w�$���GkUUk �����$�Tw�o� n�Ӏ^v�o��ى���qE�qh��>ՠ}{w4��Z/p��7ƤJ4�����;w��@����4�M��B�wL�N�zn��<��f�k�Z׷s@���g���w�@���rM!���
B6�V�0j�b,5C�L�i�0t���o?��ۃ!�vp��3X���CuiɮŰ�{9�qܻt!<����q�������͞h�pj2���9-��z��퇋�gB�������H���f�YLb;p���mۇu�)c�`��6��"ŕ�cw[����e��um���t�L��#=�!�)��N9�m[����:�]�{�N��M��6��,l�7 ]Թ��cȷ2�,�v�w�=ǽ߽��o�����䥹5u�����m�\E<q���rEt�[�]����\�p�ͻg�u�7/�BB ����-h��Z׷s@�ڡV1c��Q�@��u�~(�������)�͙���ɑ�2G1Šw��hr���;V��ڴ�t��L��x�������w~X;[��}º��B��;w��@�����6��X�s4��ZתS@�j�/-������f�[�N+����s�f�4�ԑ����E���8�]��#pF0R TNY����ٶ`�u� ��/DB��{�u�N��O��(�*�v�M�N��2*AR(�X$�_����ۚ8�ZתS@���
ě�H��)�yn���O��ߒ窞4��-�������9��v���)�s��h��h:X�PjU
��k��]�>��]����=����;V��zfq(�f�鎹�n!�|ڝNg\�F=[:1�Wm99[zcS	�B fE&D�4q������;V���S@9�JX���8܋@��s@��ՠ}j��9�ڷ�#˥���pR,h�s4u��@��u����0@�W�%@"$"�,$�H�� 8�����=����;�}B���rU�Uus������ �o� ��Ł���yh�zE7
C@��]`J;�~_����tv��rZ�q���]�l�r৻9�}7�����Ӕ�{M��o7{��Bݾl,'O�;����;V��K)�s��h�v�y���!eE�h�{�_�?ff)���9{��8��`:D��Eu8�k����@s��z?$�?bY�G��,�����=CUs7AB��VMف�!$��׵�w^��>�78Ҁ���b�B`��igs�1q�Z���OP*�#��sWu�q���<�/(�P�^{��;��Ɓ��נ�ECn�cq,��;+��������ת
��V�M�/onr�v�4�,���xё9��v��S@��l�1%����ihvy�o꣍�l��us�}��3R�Q2vz����XܫV�f~H�[�="�&8�P�W^���,=
�;[��u�z`�tG��:ݩƛv��I������g �Gl��(J{]{Xi�U�T�v��LJL�>�h�e4.v��� (�.cľ�Ĕ� o�bedpB`�`{�=f�\�/�i<<�k	A��1��GY���x�"N+1����!#�}[�Ӭ��04��j|��
�Os���:�� �@�dH�>97�|fc)(J2�2���>5L�f0�l"�y�ʚRI-�`"Vf��|Q��is����m�m��`B9[c]Z6�� ���p�JJ�LF�V������r�vޚ��wF�d%��t�l�wj�P��v�X.��u������,���'8�Ԏ���i�K��u���B(W6��[n��%i^�I�,���9�T`�{6%֧t��N#qr��m�{%�����:"��s���T�1�7:i)��M��	�N�mnn����yKn�ˍ���^���͵u��� x1�n���UUt	���@W*�X�$8���|�l�[G.^�"Ű�Sɥl�8<�kv��:�ϱ�}�֭�{r���b\]�����շV����ѓmk��P������9��pr䶝g��9�����У���ե�ӻ�9������'Y�ؙ��۶m=��z��q,lg��+�0]�\]���n��6v�mٴJ5�5Ӈ���+@�Bj��� m�Zk˸�ɵ9�&�rD��-���K���8j�YUM%����q�ղ���m���vj�m�&(�gM�զh	LI�M�[M�N���s�A/iA,�l�j�n��L��'2�dʬ���`��
t�:m����7/VM����c����˺��r�;6,�ĵj��]ہGE.�G\���u1�"8����^v�P��cd!B�8�^���7�kC��2԰mWR�WF��������kV1U�S�;6��iuEm�ps^�i]�-�n5�s�,�ZzsӇ����]<�z�n�qcv�0ں�lY�ѹն'�B�e3��v6nwr���݋�+V��ںӝx��Ĝ���e��*V�1M�K���:�=�u�P�H"���c\�=��Nbs�e�Ȅ�0��"α�,�.��v��B�T�xu��p���6n�;st]�����Ji�1q�u�in2%���v.��eq��̚P�'l��r�ɽ�H����/\6����3q,q��F�Q�C��ݓ\�T���]v�7��a�ٹ��3ڱG%?��w���}�UP�'�����?P��|ll#辘)���< h 
�]+@ ������o���ڑ财�έ�C��v0�4�BGp�����zb}���^�l��+�{Y"�{u�L�K�l��u2ՍE��*YZ7F9��n�v����ɹ��M�t�]e������ЭR���RP�ݴ\�!]����3+�ֱ�]"&�D�6��s����;�/-�+I��n�7���k��Eڝ��C��n%�v{YZ������{����;�;��� �x��/���NukY�-������/߾�v����\�dSC�tt��qs�����ߡ/B�Pu׽8 ��S�VM�H�nՓv`�u��׋ ����tv��DzUM��-XUM)������ذ��Z�,����נ���u	�8�#"s4=������9OO;^��g��_}��B^�M��q����K)�qs������v��ؤc���½���=ֱ{m�#�v���
e��l�sN���G_o���Y�Ёz�B:[M���}5�L��L�߽�ֱl��V%���n���&D�,O{?o��p��L��_�~oB?DXV�N4۶k"X�%��~��!�B�Һ=P6�bn%���ݧ"X�%��g���r%�bX��w6��bX�'�nd���l;S��bى��������IȖ%�by���6��`#bX��w6��bX�'���6��bX�'^���U6J�]N2Z��f&bf&b��iȖ%�b{����r%�bX�����r%�`	by�۴�KıM}�~O�(�*�Tv�ų13��{�siȖ%�b�~��"X�%���nӑ,K�����m9Ħ&b��m��?�$�����m�&R�ں��*9�]4�M6�C������q�ն��2�n�3Zͧ"X�%��~��"X�%���nӑ,K�����l?
�D�&D�,O���ͧ"X�%�}L��(퉱W*�-��������v�9�!��,O{?o��r%�bX�g���ND�,K���NAB�f&b��1��n��,��bى�X�'ޝ�fӑ,K��=����K�	����:c�P�uH��r'w�p�r%�bX�����8bf&bf.�}�6ZKlRT�,V�Xr%�`%��{�siȖ%�b{߻�iȖ%�by�۴�K���ȝ����iȖ%�b~����_��M[�.Rۭfӑ,K���w�ӑ,K�|�]��r%�bX�zw}�ND�,Jb�ﾚų131qv��c��D�qG����dzb�/%3֥қr�vW��v�X��ÝW�,d�vq\M�{���oq����w�iȖ%�b}���m9ı,Os߻�D�,K���ND�,K�{��4Ynhɫ�$���r%�bX�zw}�NC�"dK����iȖ%�b}���m9ı,O=�{v���G����ߟ��������i9ı,O���ͧ"X�%��~��"X6%���nӑ,K��ӻ��-�����������U	N��iȖ%��`dO�w��ӑ,K���~�v��bX�'ޝ�fӑ,K��sЖ?Q�0G��V4@�Ezr��@6��,CCK�h�­�%���N���Ȟk�?fӑ,Kľ������5.�����ND�,K�u�ݧ"X�%���wٴ�Kı=�~�m9ı,O{�xm9ı,Oʇu?w��v{IC�=��O�7jb3ێ���hg�����:��k����u���F0?dBa4�}�Ȗ%�bw���M�"X�%��{�siȖ%�b{߻�iȖ%�by�ۼ[1313~>�-%�)*v�+l�r%�bX��w6��� dL�b}���m9ı,O~���iȖ%�b�V�����$'�eA�E�թ�[u��r%�bX�����r%�bX�{���9ű,O�;�ͧ"X�%!v����)!I
HM��*�UswAE֋�Ѵ�Kı<�]��r%�bX�zw}�ND�,K����ӑ,K���w�ӑ,K����;MۭMM]%֮ӑ,K��ӻ��r%�bX��w6��bX�'���6��bX�'�뽻ND�,K�H�>�?vEvƧ�6\��j�v�z�l��gҶ=�Y��gv�G����r\d�9��:@�Җ�n���h�����vzq\��.����
��<��UWK��]���,�k���hݘ��r�qiI�2a�e����ɥ[2�f�6�Q�ά��"'P�˫n�v���Q�q��[ f˩:�ۻu�Νt�ڴ�x�n{��u�[�KB�����"^ıkr�4��Օ4�݇k��u���Wm\�ñ�rr�@��n�k� ���;���o���Kı>���iȖ%�b{߻�iȖ%�by�۰�<��,K���m[1313���~�YBG��.�r%�bX�����r��L�b{��~�ND�,K���m9ı,O}���r'�VdL�b_�_����sR�X[\Ѵ�Kı=�_�]�"X�%���wٴ�K,[�~�pI���KY� ž�?&� 5#���'b}���m9ı,O}���r%�bX�����r%�bX�{���9�L��]���l��dRT�,V�X�b�,K�~�6��bX�'���6��bX�'�뽻ND�,K�N�iȆ��ow����qV]m����\�m�7f�_�D[ӮE��yv5kA�v��h�K5�m9ı,O{�xm9ı,O=�{v��bX�'ޝ�f��șı>�����Kı;ӻ�g�0��jvU�[1313;~��ŵ�X��>��Dt�'"X����m9ı,N�~�m9ı,O{�xm9���2%����y��%3Z����.�v��bX�'~?o��r%�bX��w6��bX�'���6��bX�'�뽻ND�,K�����X[�Xj�Z�֦ӑ,K?������r%�bX�~��ND�,K�u�ݧ"X�%���wٴ�Kı=�>��#��\�k�L��L�߽�ֱlKİ|�]��r%�bX�zw}�ND�,K����ӑ,K������?|���.���-��=c��Y�œ�g���sv���1�ۈtO�u�b������Kı=�_�]�"X�%���wٴ�Kı/���lD�,K���ų131s��m|��YY�[��Kı>���6���șĿ}���r%�bX�~��ND�,K�u�ݧ"~��2%�����94k5��%N��m5�f&bf&b~�߮�l�ı,O{�xm9�>�,�����$�	!��A)"dA�]
q�<=��;�{v��b31w����-����������ȶ�5�r��k[ND�,D�=����Kı<�]��r%�bX�{��m9ı,Os߻�ND�,K0�a-��X�bf&bf.v���-��K�G�{�ͧ"X�%��{��ӑ,K���w�ӑ,Kľϡ3����OD0����h@�=���l��l[��磳ې�6ۇ±�c����>�Ȗ%�b}�wٴ�Kı=�{��r%�bX����؋Ȗ%�b{�׬[1313_|���5YP�]�wSiȖ%�b{�����?#��,O�w��"X�%������9ı,O���6����bX��w���-ԗ.Y����r%�bX�����r%�bX�����9ı,O���6��bX�'��{�ND�,K�{�ftՙ����W4m9ıB����iȖ%�b}�wٴ�Kı=�{��r%�`g�#�@`I$�,D�
U	����~NDf&bf.��m�ϐ�,���+�-�X�%����fӑ,K���}��m<�bX�'߻��ӑ,K���w�[1313�O����¦UhH�K��r��֥!֙^�-�U��m#uâ^w%ۘ���J��5-���X�bf&bf/s��6��bX�'���6��bX�'�뽻�,K����iȖ%�b�M��kGm�5�f&bf&'���6��bX�'�뽻ND�,K�{�ͧ"X�%��{��ӑ? Ɋ����?U\������X�bbX�'�~���Kı>����r%�bX���m9ı,O{�xm9�L��_g����6K
7T)�[11,����iȖ%�b{�����Kı=����K��*�"}��~�ų1315���G�5YP�]�vͧ"X�%��{��ӑ,K�������%�bX�}��ӑ,K����iȖ%�bt�,$
�AH1+�"�H�?_$�C�G";t�9SG�]���tN�;l���ͽ��1cm�n5*b�%�mͲ����v[vꛣ
Ѷ-�.�ݬ���ֺ�b�`�;n�d���FaT�n�� B�EeƮ��V[:�ZrMr=q�];z��.r�[6B2m�{�#�6�\ҝ+���_N�\�%�W����v�h�A�.�/�44Ys:�=��x��g�%�tM\��??�4&o�Q��}N�����B��d��T"���7Wg����b������G�����{��,O�}��ӑ,K����iȖ%�b}�wٴND�,K���ͧ"X�%�{=�3:j���ka��ND�,K�{�ͧ!��L�bw���m9ı,O���ͧ"X�%��{�Nf&bf.x�m�ϓq�
���i9ı,O���6��bX�'���ͧ"X�%��{�ND�,K�{���ى�������e��
ʝ���iȖ%�b{����r%�bX�����Kı<����r%�b�����Ʊl��L��^��M��J�Gm�Y��Kı=�{�iȖ%�by�wٴ�Kı>����r%�bX���k�L��L��ߟ��D�W*���˦��������A]<��+���6�Kv�X�Ҵԩ�,��Mڵ�f&bf'��}�ND�,K﻾ͧ"X�%��{�siȖ%�b{���ӑ,K����;MKsY�R�2Mf�ӑ,K����i�t�"BH5
����:��!��<�bw;繴�Kı>����r%�bX�{��m9�#�2%�O������D�SY���M�"X�%��}�ٴ�Kı=�{�iȖ�by�wٴ�Kı>��|k�L��L����R�q��5��r%�bX�����Kı<����r%�bX�}��m9İ?,p���!|B����>�
򹫩��-��4m9ı,O=��6��bX��A����m<�bX�'��fӑ,K���w�ӑ,K�� a�����?��@6�\�0�}'��!��sMkIq)xlx�tmv��Μ�a���=%m��,K��߷�m9ı,Os߻�ND�,K���șı:��2�)!I
HOƯ/�U5hUv]]�kZ�ND�,K����ӐlK���w�ӑ,K����iȖ%�b�w4�_��$)!7��4U-We��T2�k6��bX�'���6��bX�'�뽻ND��@�'��@���� ą�/�٩���q.�Qsl%p�n����`fd�<%5Y��I�, %]�
JK��C�C�:�7 �)���$�lI�����&��y�Ӳ:32ci D#�)��5�q�Y��1:� �$V�R�O d�����`� �Sxc�Dq7�25��Ã0���&��jNa�JJE����8�R�$�_Ai���$��ƭ�-��)��
B��J1.���B�R
E*�f� r�f�sDqԤE�)T�C{�M�9���a�ouG4�JC4M8���`*��7/�D<Pt
A4 �(t���}v��P�|("��� �= }A��)�#�U4(A�D�'����ND�,K���ͧ"X�)������r�����X�bf&~"�O~���iȖ%�bw���6��bX�'���ͧ"X�%��~��"X�%�׽�v���.��Y.�v��bX�'��}�ND�,K��}�ٴ�%�bX�~��ND�,K�u�ݧ"������x�'�E!TD��K�G\/� �Z�mN�����яZ���8�m�5�*��,���ų131vw�Mbم�bX�����r%�bX�{���C�,K���fӑ,Kľ�;��e-ԗ.Y���m9ı,N��xm9�r&D�=�_�]�"X�%�����6��bX�'���ͧ �bX��L'Ȳ�F6Aʵ�f&bf&b��nӑ,K���fӑ,K��=����Kı=����Kı<�W�s�I%��NY^�l��Lē0���iȖ%�b{����r%�bX�����r%�`q��	"D���+�U�HD E I��"`�"{��nӑ,K����&���Ii,��k�L��L���}5�f%�b{߻�iȖ%�by�۴�Kı>����r%�bX��~���?�f��dY���5=�ô�Fٴ��魬���TT�����?��t$^��]�;�Y��yı,O�w��"X�%����nӑ,K����iȖ%�b{���X�bf&bf.���>dr������6��bX�'�뽻NEı,O���6��bX�'���ͧ"X�%��~��"~ 2�D�??��?a�nk2�ۅ��WiȖ%�bw���6��bX�'���ͧ"X
6%��~��"X�%���nӑ,KħO{�wRiT@��i�[13?	C��~�ű,K������Kı<�]��r%�`~F(��?}���ӑ,K�?����CU8�vWm�ų13���ND�,K�}��~�O"X�%�߿o��r%�bX���w6��bX�'��`�h :Mh��D(0ƈ��	��KT �ST�g���Ω���Eೇ�c�h��P�i�����(����Ur�O[�sd��=�F�.�����n�Jp��	�x1[c�m�����K6ڥ���j�������[�շY�%�ʜ	ey:P6:�s����\96�b�6T0r!,�:n�q,��mՊ�蒲�ėnc��������-9�	�f޺z1�K���N.ښ�]a�LֵsD��: �^�a`r���u��뜦;V�&{j%�]3Ip���2"�R7]i�Y�b)50�E��1�e�O�X�%��u�nӑ,K����iȖ%�b{����~y"X�'߻��ӑ,K���GYs�ˑ�ZT���L��L�����bى�bX��w6��bX�'���6��bX�'�뽻ND��0D��,O~>_�ʉ*���-��l��L��>ϻ�6��bX�'���6��c��DȞ��߮ӑ,K��߷�m9�f&b��f�_+J�H(ݳX�bf
��~��"X�%���nӑ,K����iȖ%�b{����r)�������$����v�eZųı<�]��r%�bX{��m9ı,Os߻�ND�,K���V�L��L��#寐["�&ݵ�<]�|0m�^�(��=rY�N�OR�FC���3���cL�X�bf&bf/w�|k"X�%��{�siȖ%�b{߻�a��DȖ%������9ı,J~^���T#+v��k�L��L�����Ӑ���c�Gb�,$Ť2Ҙ�ad��T�ȫIP��mӃ�a�K)L�� ߀!�!�L�bw�<��Kı=�]��r%�bX�{��m9�����@�����N��X�abX�'���6��bX�'�뽻ND�[����iȖ%�b{����rbf&bf'�ߦPv��lQʵ�f%��߷���r%�bX����M�"X�%��{��ӑ,K�=����-�������*�|ۑ�ZT嚻ND�,K�{�ͧ"X�%��H���~ͧ�,K���p�r%�bX�����9ı,O3�fN�)
a��
����^�]�Ql]�@���tvQ^�n�\kv�^r:l��0'���{��Y�=�{��r%�bX�w���r%�bX�����D�,K���ͧ"X�%1{�3N/��D�nY�[131X�w���r%�bX�����9ı,O����9ı,Os��6��X�)����'ղZ�;S��bى������nӑ,K����nӑ,p8@�Db H�2Ā��� ��O���6��bX�'~�xm9ı,N����5-�f][p�]j�9ılO����9ı,Os��6��bX�'��xm9İ?2'�o��[1313_��F~�U�ݱ�nӑ,K��=�siȖ%�a��~���%�bX�}�߮ӑ,K����nӑ,K��ZXCrܲ�_�����A��lM�H�5n4����SM�r[s�'C.�P^�`�"vW%���18�'~��iȖ%�b{�۴�Kı>�۴�Kı=�{��r%�bX��ﱙ�]j]Z[��iȖ%�b{�۴�ı,O����9ı,Os��6��bX�'��xm9Ħ&b��^�O����9ezų18�'��{v��bX�'��{�ND�,K���6��bX�'�뽻ND�)������n�%Bv�Wl���L��X���m9ı,O����r%�bX�����9İ ��4��XD�ˌ�\�u*�0�O��&�6B �F�V��ު}�9�^r�8bf&bf/���pq|�*"��ܳX�ı,O���iȖ%�b{�wٴ�Kı>�۴�Kı=�{��r%�bX��E>�����2Y�-�5u���n��v4��rƜ�ܻ���<q�j񤖶K]Q�����131{ߵ��r%�bX�w]��r%�bX���l?0�&D�,N����ND�,K��_O�Vƥ���;^�l��L��^��۴�Kı=�{��r%�bX�w��ӑ,K���w�iȐ_�r����*
�*�j�
(N_�X�A$O~��&��'�����9ı,O����9ı,Op�����]L�0��\�fӑ,K����6��bX�'�뽻ND�,K�뽻ND�,���ͧ"X�%�{>��Iu�uil2涜�bX�'�뽻ND�,K�뽻ND�,K���ͧ"X�%��{�m9ı,L�d 0I�������?y��v�Li��3K�l�&�L���B�қ/U:6��we�b퓳d�b8X�{ZM�z�Ϝ���e���C�����5��so[��
�O9�Ig��4�E'=vJm�Ҫ���N0�r�Gb-��۷���=�u��mÂݥ{��vc�鞇\���]Vw�^h��na�E]���)1���6�M�W'X�:I�dM���Y�I�����w��;����֩6:)\��[�#3��V@8�X��&��Vѽlq���q�^G�*ֵ4\�j�>�bX�'~�{v��bX�'��{�ND�,K���6��bX�'�뽻ND�,K�ώ��s4B�R�SZ���r%�bX���m9ı,O����r%�bX�����9ı,O����9�2%�����K�D֦���5�ND�,K��~��Kı=�]��r%��Dȝ��߮ӑ,K��>��6��bX�'�Ϸ3�V�n�e֋�Ѵ�K���Aȟ}�߮ӑ,K���~�v��bX�'��{�ND�,K���6��bX�'W���*�r�����f&bf&b���nӑ,K��=�siȖ%�b}���ӑ,K���w�iȖ%�bw�!ۊ��IKiW"dU�{�Oj�.{�&�whzt��zK�8���I�[�eֵv��bX�'��{�ND�,K���6��bX�'�뽻ND�,K�뽻ND�,K�$����%�˓����m9ı,O����r��
ix�9"X�s]��9ı,O{���9ı,Os��6��bX�b�ϨKG[M��U�[1313}�{v��bX�'��{v��c�D�Dȟg߿fӑ,K���߸m9�f&b��^�O�%��J�v�ų1Y�dN����iȖ%�b}�~��ND�,K���6��bX�'�뽻NDf&bf.�y}��9P����J��f+ı=�{��r%�bX~ ������Ȗ%�b}����ND�,K�뽻ND�,K�����]h���E����<�ۆ�vӖ����,��i�S\�O/]�jQ�-D�E�
7,�.���������"X�%���nӑ,K����nӑ,K��=�siȖ%�f/t�����]��jvU�[1311=����rbX�'��{v��bX�'��{�ND�,K���6��bX�����EZ�� ��ų13��u�ݧ"X�%��{��ӑ,p{�k�W)J��P�JJB�����6�������� UuDQȞ���s�ӑ,K�����6��bX�%<��;�a�2۬��]kWiȖ%����>�߿fӑ,K���߸m9ı,O}�{v��bX�'��{v��bX�'�O�grh�S.L.�WZ�m9ı,O����r%�bX~R+�w���yı,N����iȖ%�b{�}��r%�bX����ft����.8i˥���WK�9�N�7��ٓ�|�&:;����kpc+w����X�%����nӑ,K����nӑ,K��>����,K�����L��L��ڽ��(�-��9-5�q,K����nӐ�$r&D�=���m9ı,N����ӑ,K����iȟ���,O�N��j�����j�Y��ND�,K��fӑ,K�����"X�ؖ'�}�ͧ"X�%��u�ݧ"X�%���w)���54L��e�k6��bX�'��xm9ı,O>��6��bX�'��{v��bX� �����|��Ѩ�-��u鈴l��L��]]�G�V��Yu��4m9ı,O=��6��bX�'��{v��bX�'���ͧ"X�%��{�ND�,K���)ٚ˭B������d����=c#��/g:m�I��ök��7��,K�뽻ND�,K����ӑ,K������%�bX�}�xm9�������辁۱����V%�by�}��r%�bX�w���Kı<����r%�bX�w]��r
X�L��\�>��*�p��]�k"X�%��{�ND�,KϾ��"X�R"w��~�ND�,K��Mbى�����ǽ3���i��Jm9ĳ�"{����r%�bX���߮ӑ,K��>����K��r'~���Kı=>��f_��L�kSE�֦ӑ,K����nӑ,K��>����Kı>�{�iȖ%�by����r%�bX�|��<X]�~t�8@%���Ǘ�<|�Ιp#��$(B����7���s{��Y�y����I�)n�ӱ,�JԳ�M�9���њ�T���.�R�an�1i��sbpR}ę�f����~�p��ɭp��5dԤK]"�#f�({>�kÜN$P�3ﵯ�_'6I����͏)GQ5�U%�L��u8&��i�oG���{�r��+Hl���m z油a����Fo�40\���`E�c2�` ��糄���r\�7q�Hh��7���WF�4O�)7�y������>�)�bĔ���)�%%�0��<�-Ř�M�*�`�s��u�m��m�gnZ�.X��s��[�[;rF��]��rn�]k��dƹ�OV���s�Gjq�M��:�*m[9*�M��Ƨn��8��-�:�qp�xo%:h�%�$���	��t<�+�V����C�\s�C���6���N�:z�r�%���7&`�Wc���[scc��$G��u����ŧ�N�1Y�Rښ���A�l�u*�Rڨ�d�O׊�AQi��su�e���FX�]�7n�[Y�s�\����Gm�lA��6zOdn��îz��\A�y��l]lM���������4c�Wt�*O&���h�wzԫ�m��f�u��+�m���\�\tFD�n��_9�ݴ��s���2싷����P!���s�;.�G�[.�P!m����9g�!�V{v]�Wg��<55�/jcO�o/C�{A#[R��%]�6���K��9+Ƀa���΍�qV�gdx
�]qUR�*���^��Ԯ�6d����x��d
P@e'4�\Tv,�֣�kh ���s��Nݶ9!4�.����Yˬ@�SK*jj�\��D�]����<i�����m�=m<O3q� 톜��Xt��@�9gkm��%�v��}]��s�,�tM��**U�c�z�n���y۴mJ�[���y-d���l�Ѳ����9��X,��sin�l�P�U�΂���#.���� ���`�0���cKӶ�\W��U1��͢�+y���qEx4�e{nx�k�m��P�l����h#c��g���3�@���	�c� gh�YZ@�Q�b�K%:l�Y�k��rö����n���#6R�vey��G;29�H4%�\7Lu��2�N��m�4���c��Uחh�� �F1��p{n��������,5�K"ftu�I#VԊ��v\��SP0=�ه9��5�<9N��asl*���5�Zi�X}��4W��T#ƞyH�+��I�kM��vi���n�N�[�Թ�3���lߎ�z{����~@6
l��C�G��?!�p4�z���A�)T@�D�HA�H�LT14"��Oǂ&x8|)�;��68���j�Yr>���O���M�m���2K�|%���G=���e������m�p26����#s�l��DZD�������a�Ll�PxN�d ��+On�)R����
�֮�m�$΄��3���ty��'F�g��p�sV�{Jv2�t�x�q�EM����w�1��j�tn4�a��2P�I+���G
�ĸ�ř��SX��]�ղ�r��nN�V�Q��E�"wTm�1p�I�q��,�n�.���R��O�X�%��{��ӑ,K�����"X�%���o�j<�bX�#�ݜ��
HRB��R��B��U�u�ͧ"X�%����6��bX�'�}�ͧ"X�%��뽻ND�,K��}u�b�f&bf/.�GҌ���Z�Y�iȖ%�by����r%�bX��۴�K�C"dK�����"X�%�����6��bX�%������ֵu��sSiȖ%�bw��nӑ,Kľ{�u��Kı;���ӑ,K,O=�}�ND�,K�|w�c�n�k��bى�����;ﮱl�ı,?*��߼6�D�,K߻��iȖ%�b}�w�iȖ%�b~@?����Cn�Z8�{gu��h\�K"F��z<�E�m��r�8��{����}�i�y묚ֵ���,K���߸m9ı,O~�{v��bX�'��{v�Ry"X�%���kiȖ%�b_ӽ���ֵnk0�Y��ND�,K�뽻NC� ��DPpCnD�K�k��ND�,K��{��"X�%��{ݭbر313��$_))$��5v��bX�'��{v��bX�%���bX�'��xm9ı,O���zų131w����q�
JY]�5v��bX�%���bX�'��xm9ı,O����9ı�߾zų131{�|�I���E]]�/�RB�N��� �P�������- �h����DI<L�$�9N��m]��[�drWNa��+��N�3��mn��{�w�H��FR"9�����h�V�u�~�����,S(ݫD����%�r-�j�m���h�V�bA����$�I(��H�������}�s^���0 ���bb	� X��@u��!� �}[�Z:�ZX��o(˻��򈈝�ߖ�[��7M��%������������d���X]Z�]�@;m���h[6�Lߍ��sv{EyW/�y�Z���T������v�1mT�N�iJ;-*�����}8������H=���:ƶ2榭
�˫���� �n�TBJ"d��ŀ_?yh�V�~�ďxum{s	"�����X]78z��n� =ݽ���T�9`�"#��v�V�~Ͼ��O~��n@�����3>��h(���	��@�ڴ�٠[n�k�hw���dP��ӝW7�,��R�!<-�(.Ɩ}Vѝ�,���Y�n����**>�o�����۹�Z�Z�ՠU�D
4�,JI$�-�s@�v��j��f�S��	"N&$(���v�V��78l(�����������I�pm�Ldqh�V�v�4m�����;K���4�5�E#qh[w�j[��/�{[��7M� �"���HM85iT�E���%0f��̻E��+V����T�'ls�"`��1��۹�K�1b����N�]y�i�U�\�r=/��+̼c�;��Ŷ̷^��,�%�  �nd%�c��v��(� {+��:6$��n�/g�km�ws��i��"�����a�B���q�vn��,۔����������w6��m[�m<��״@�����?����|�;5��<띱�j{����=�H��K1a�ssͪ����_�60�9���rp{�s@�v��j��f����*D��0B���;]�@�ڴ�٠6�,�(P�M�S�VL��W73B����~���f�m��k�hw�u�<�A
E$Z�l�-�s@�v��j��ʲ��i�X��I�6�,����np���6$��ߝߠr'�qB���e1i�\ƭ7\<3��Q]=K���������xs>���@�ڴ�٠[n��.�7��	�	��-��o~��D����#"H�؂@�#|"U�:d�o�krO-��k�h�ܿ�&�ƲL�(� u�x�^,5(���W�8����΀����`�@����;]�@����l�9�}�H��")$���u�s�low4�����x��W�+v�N�&<�)\�
5��sZ^����óh����\h�rr׺Jl�\'NE�^YM �h���k�hw9]�l�%�4�٠^��h�ՠ^YM ��,b�o%www�>���:��׵%���	)��(�(�d�6"
�B�*ҔD}"-|=�5�vnI9���9_�H���
&�h~W��Z���@;m��n��.�7��6�&28��)�����s@�v��?��ߏc��s�6���
��v�vy��(��B�
�vQ^�oc]�Y������:��9!���4����ڴ�)�v��6;�s1�8��/{w6米��΁�~� �{/�I�������m`�"#��_��-��hm�@����.u�^DH�Y�C߳1{��0����x�:�#�(p�	b������{o@����H�Vڮ�%4�٠r��h�ՠw�S@�{E,��It�n~~:�%�Ϋ�Վu�egî.���M6y�d��N�c_��l�}X��㉻������X]78xퟐ�} =�M ��?ށ$I��!��k�h���f��۹�ى�ڌ�6�M�Ldqh��4�٠r��h�ՠr���b��I�E&hf%wv�n�,���Ko~X�C���`�@�۹�v�V�����}�]Ԗ.ux,m�:�]r�9��N8��r�ڡ�ܚ�YG�^v�z�tP�۩;���i��۱;yg-�K8�\�A6�ܭ`���]�ԋv�kD�$6쳬61��=�y��l;l�6��q�N%Ѵ��\�߸�^��=%M�&�#u�Vt�p:@�E����j�a�x��4lF��x;GZ��g�:�I�����秊�3l7�`<wOm��<��Z1$��I�Y�\�G-�m�mݩ�q�׷������^��5��p���������t��ma�K*��}���}� :ۿȈ�\����`������ʫM	��E�^��hVנ^[��}�<k�X��ߡ>c��m��ՠ:�����a��*������`��W1b�7�rH��w4���/m��:������Q�8�$A9���0/$��� ���`���8����	I#��Ő�s5nq'N$ɷM��,����9���z��-=	�/J@��C��/m��:����w4���;����*mZ���ՠ:��ML�K� ���A"*�`�����Pؾ�Z�_J����L��Xz�`�M��cQǠ^۹�}l��{n���נs8���'�D)uk�D$�	W}�`�{��]`��h�Z��1ĤBh��@����]`���>nـz]�-��כ����9���:Š*#5�;J�wN:��V�#��J�����+mU$�g �����{n������3�es(�x�'$�@��s@��f ��,�޺ͅ!�����n�j��dլ��� ��,)IJ�N��=��\�D/��2�B:]�V^R�P�!m]� C��*@�hh����#<E��P��j@���4M��	m��<�hx�!e�aH,�!GB$R����9�H�m�B���|��]hY4&��l�X� hqQ����R�p�'	���Cdc�����<D1Y ���H�1"BE#Tt��XZ��XI	�S��D����BBI�hE@خ:�5G�
� 0~5�7_/YD}���Sl���&�&�Q��(S�Q�A�^*l]���l�E�D  �V z��=A(|� S�j��ھ
�U=Ŵ�:��4��ih�αG�u�.ˊ���[ŀ9m� ��,������m�b��s�2H��3@����n�k�h�h�_|�)1(N�vs���8��n�Y���q��if�6�:��V�Yx
��ŭ�t�V����m��� �78yMΨ������`S�a�D�I4�ds4_j������Z�����۹�_�j�iĜI5��;�j�*��O�����w�@3�WS�(���)���^~�z{�vnI����rC���J�-!�8L��ԇ��� �ｻ�N���TӤ�Dܶ٠9��K@}�b������-����r��\f4A�;Y��P��D���9�i���W��+�׾��[��$J$��R&��"	��y�-�V�U�z;۹�}��F4��pmݗws�}�ns���g^���k�[�ٙ���-�'1���nE�l���9޼XjJ�{Og ���;YL+	 9���&����h��huڴ��h�{�"RdS���f���V���_o��/������'�W�!I
1�iA�Aa!D��pb�V�f�	&fk.�ۣ��tױ�Ov�m�V�[����s�����خ��÷X'��rg������kv^-:�oQ����d;q�했�b��q����5.�Q��E��Mh'*ug���b=�����KNΈ�|�h:;��˥�8�lS\urX�1���ex��u�V���e�Tףv�$N١�t����Й�;U��kG���$�b�R��;��q,��.��CD��(� ��<gv�4\\���=1����Y�,qF�^�!�N��ͷ��~_���٠s���k�Z�w+�QA�G�Q�@�������-}�@��S@;�)��X�M�Ĕ�=����-}�@��S@��� ���U���)L�MZ��B�ݷ��q��9}o@�{w4�*1�pO!���"�>��*��@�{w4_j�*��<���\ݗ��u������A�f�h4l�l�v�1p���r�qZ$봜̧k�b]��_]`�^,�띄��C�oL��H|�-T�@s�����&bg1e�Y��,�}|h�ﮀ�+�)�"�4�ds4��Zݶ�6!%2>����,îӫ���&F&�7���b������s������ ϻ���qF28(��l�9�����V��l����q��Yg
թ����tt�rQ1�;(a����K��i�ܦ�sۘ�����K_m�����>u�8�v�P�!} >�� �ߦ|��Z�l��h�w�_%�,l��� ^����̈́�S'e�MjT�ZUk����@�}tw�B����P�0��}���>�Z{ہ�8��!%ݘ��2���oq`:���4�L;�cNd0iɠ^��h��h�S@/;f��Ǘ�5'?#ʗ���6�I:�V�3��t�����mc;�E� �0�AI�<R29��;�^YM �;f�{۹�_����ĥ�5*�p�l͈� ���oq`��o����r��y� ��G ޽��� �]s�>;f 4.���i�cNJ�A�,O�}�ր���=�=��}7 ����b�A*P$O�Pښtf�R�h� �JCNI(�i,�䴨��� p�fy�;\px������Z�[����}4[w4-鍦��cȉ��_���Q�mƄ�M�5���h|����h*�8��ݔ�nB~rE�w�S@/;f��n�x�V�y���$nd���Hh�l�/m��/j�/l��U��K�3V�EM]����+�p�
g^���M���,X���	)���� }v� |��Q:�~Xƻ��n)2&��Z��=������q`��8e�$�J�! ë��F�,Z+9�"]{s�C�wnwM�$t���2i7B�662W(��u��u�2<s��C��z��r�� -Zx^Ϧ#5��u=`�t1�S�-ښ�Ci���)r�Xz���8�U'�{\u��Z��1���r�Gn1��9�Z���k�����^;�]��x�͍&���=L��l[�\�ٵ�Mt;�֑	fӞ!+/�ww����;�}v�N6��n/,X=�wZ;<<L\]�)��8�)yv2�ut����w7Vt��x�x���$�I}!���@=�_,�b�q7&�{^,�
&M�=�^ޘ ��x �:��Px������Z{e4�h��h]�!�pl�����h���٠r۹�^>ՠ^v�5I�Y#�)$��^v�����������cI�bI�d���DOv���SSnJFu�2�r٦7��n޼N��I��f94[w4�ڴ��h�l�9��(�'�����>W\�_%Ԣ.�q%8;�ـ�w�r۹�����G�y�G�87�7���� :�ș����7��pq�7��,"r(���@�s@|����(R���Oelڕ62Kq7&��n�x�V���M ��m��w���M��G��[�I�fj�c�]��@�5Ń� ��n���W%���D�o|�v��<X����_�����M ��Ϙ{����ަG<�2��.Kk���`����� �]s�	)���7!�GRI �o��{۹�V5�A����%�>��=���/,��qZ`�871�
I�>���9����0<�QСUu��h�E�H'���f��>ՠz��i�;�x�^,��S3u7�4��ny�\d��V.�&��sz�xv������]�vr׺Zk]]����o���}�f�{۹�s��h}�W�"�Aȣ��}�f�~ď[���wӀ>;fy%�CP���U(�����S�@�}���}�@�즀}�f�S���hq5������|�[<nI9��kr~ *)����='3@���6���Q��-����[4�w4qڴ.u��c<B�)��.�M���f�*ۙ��7.(�.W��y�r;4�"[�U�I?�� |o�Ss�(_Hkw��u�x���f�h��h��Z�e4�[4��AՄ�O)Rf��>ՠ^�M ���������I�&D��@���8�Z�8�Z��+�أ&�� �)��[ŀs����ـq})	��繽㮞�.z����mѢ�8���ق���=
�0B���L�Mfn]�,!'$@�ڔ�CFt&i��aq4���y��!3[�"G;�u�k~��z󸠸ty�=aށ�C�C����D�|D��h<כB�e�qll�\L�h���.�������8�@��S�DAFX��s��Nl�}�5z�bZ��C9��F�!�5ť���M�Q�o�����l�C�>0f�iLn,�>�rb���pu�!hbP�k��oi�o�^0�s��r0�B/LQj� EX�^�C�5�������`|?���c���E>�O�xa	sc�%g�Ai)�T�D�As}��{�g����`{�3wu�RV\�oa	��V#n������UuT�m8���&��;{wm����q�vP�7T�c�v��m�ӹɺ9��;�mX�^ݱ�p�v;pd�f_n�a�ݺ��itp�͉�Nz��Mg v]�Ue�y��si�'������ä� U�J�t���;�������<w�O��O��6�6|78w!����문�3[;j�2NC���oZ[��jlh���t��c��s�.�iID^��ۑ�x���n�k� rMm��s %�K^n�0
����Vb�厹�0�m��ݏM��P�d���\��+��%puѭi���D����l�{cLN�jt�۩su�m�;����N;]v� �'k��=����t�M�!����.�u�PP;_|kn�s��8��Kvpe��f�d���Z�]����s���mvN�vN������[�v^� �r9�Dq�Xޢ��tbb��n��$9�怶�ZU��������x՘�:^Pv:�eZ�h(��R�Uqڞ��^�^���Lr�����f���Г�]����,���9q� I�WVn2�!��(��lr8ag6!5%q3�i@P��Jgv��!.ݮ����g�ط �灊3�pO�!�S����֚��<��OIytv�;�ݎ:7�����W۴	r�:�v����jx��6z,�fٛ��"�z�k����v��Z�j���	5�p6M�m��U]U@XFm���ĭ�x^v{viVx�� �v<6����b�\���+�� 4�Y%��t��%Ti����aKv�͒0(ݥUC��q|�s��=E�S�[���zi�C���p�]ekR6�1&�]�g6���vąsIl�aSb���M�S�أ"�u�V�v��&1ɄIn����l8���4vr�K��<.��nr���ky�yz"���zV �@1��۝�f�j�lz���J旚�8��#؍R�ö�-gdR6#l��Rq�̥��hv6)}B;��j=NͻvҠZ�s��=�%ix�Ҟ8���v����f3Z��5S�=>TѠ C`�U>U:�GI�Q](� �"��pD�� '��$,Ii$�6��'�������t��<c�C���phݭ�m)���0z�^�5ў�d��v��c2�Ѹ)9і+�n��0��n+jW���q�t��<��V��ٮ�[\OV�6�l�<s�ꌥ-W+�jy�dh�c;�͸��}���X�Km��/C]����=\����{��:�VL��H�G�������Z�M�x��{�9ѷ�;���$3�4���c���+v1�[C�n�UiX�j.J����*u���N�pd�]]����wS�۴�]cQ۔��a$6�8����4qڴ�)�s�ՠ�_��Ǐ(ۙ�s��h�S@��ՠ�����W�!�VH"�Ҩ[^���_��N���33=}�s��h��HA,��rC@�s���@���h�S@�+@x�"ps#_�#��f��v_/����|����WhFG1�����[F1���zz.%Z�ꫣE8�	n�v#�<v9�dOӍ���>��Z��>\�z{l�9�Z�rc��uW8�fkW))�S���4�踋����9��O<�u�'<�վ��ى[��ߤ��4rF�qv���@���h�S@:T�0aaZK�ޚ:{m��B�W^� h�F�rU�]PJ�RG�}�ڴ��}�@�^נU�������֒��t�\G[��n�ܝ[u������N�F��&�c<έ([^��;|h�w�@oݾ>���v{�@���L��Y#�(䆁�j�%
!)���L����w��f���������@�<hq��>D�JE�A[�?  �X��jߍ��4:G���$r��@���h�e4�;^�U����vL��1̉��Š[e4fq������}�ڴ����%X�)�BX��u�9�k�ۡ��I���2#�n�'[:7n�(�OŏR6�$���s��@�����Z�S@:T�0ay�@�ڷٟ�9��-���qs��*ΖD����b�H���Z�S@��k�-v��ۈn!Lx�$��"�����4��=�jܞ�6�#t��-q0B�X��f%�X������갣y#�)�@�s��^נ}��h�ՠU��Ġ��`�#��1�����K<swS��S���:m�u��n��k����V�dkR=���s����h.Z��:5L$Ȟ�mǠs���Q
ɻOg 9������9���$�L#pr��hܶi��߳�^^�z{g� ��\mX��Hcq8��[4
���s��\�zC��f !cn	ɠ^�ՠs�����@>�[4{V`��K�$<��t;�)]K��c9���AuMb`I��,iۛ��y��\N �dg;y�'3u�nܽL��巚C��nՖ
��Z�}v{hM`��Ukg<eB�:��lO��Q���ZT7g�$l&�;R]y�]�n$��M�^b��5?�?}kr�O��&���1�"�ڵܾK�DMe�i9ٵ�5�dts�&�ϕ���፲�qO\�j��]S4O��>���F��5ubrkY�&k�*��n�ルaݎ�(��u��A�ѳ��;[`��u��y�L~���O����@>�[4����ۈnbS���������ى3���*���9��o�3�G���R��GC�M �wޚU���e4�٠\\��8����@궽�� :ۼQ􊮧�^�k�xD�O)17#�9��hm�@>�[4�k�*�\m�ɶ��28,=��hlۣn�t�瞲�sd��g,�noajb�q��nC@;m��r٠u[^��vS@3�ŗ��$�8G&�|��䤠��BU#�n�s�� �h*e�0����brhU��9��0�Q#���.�� tr�dI8�x�"I#�9��hm�@>�[4�k�9]�� ��ґDХ����
x�� �wk �;l�o��??���6àW��獪8Y0o	6�6[�[�i��{[q�#h��`��[�q�&�}��h]���e=��������1�BG�F�X��z�Z9�M �h��f���Ve
� �N�^��;|h�����b�f'���|4�M��ک�S�s&�9女�>ՠs��]�#��6�Wf q�x��w�w���lD$��|hN�����Ib�Ȝ���l�/]�@�����f��r׸�JY��cv'�����6�-sGcU�u�Isz���Q�;E��;u�8^���o������ـ�ި��9#{x���mm��&��@o��5�Ica�����o��z�Z+����R(�
C@/m��w�h�ՠ}��h矴�U�+ee�[��31$�����5���w���BI!E�H��`҉⋠<No���$���1�rG�F�X���hw�����˽w�l(�����ʛ*�qp�8L�7t�rJ�o2K���sL]���ܽu���z�%�T%+���;m{����-�@��z�Z3��"(�&�RC@9m��w�h�hw���ٙ�N����J<i8G&��[�w�ՠ}��h-�@�p�Y�<����@�l���{)���g���[����$�q�Ĉ����{)����w�h��:qڰ�"@`��$����sK���n�-NUGg���We��q��=�'��]���CA�Z�%�1gpgC��;(�s���n��d�0̕ ��2�:�us��[q�h烙���Mպ!Ή�a(b���PݻI�pF��k�T���>zz:rw9�ݷM&+ZGT����ۇ���^�Î�XD)י��y{�wF�cn2 *��E�u�f�ʍĒ;c��rV�#3�m-c\����<AO@���5�!�s2K��\4h�[��T�ӻ=Dc-�Dm�&�6�&�ӑ�;K����Q��\C�����@]�{e4��M�ɂY#��94��l�;�)�}��h-�@�q�cn�!���@�l���{)��� �;�4�2�(8D���;-4���@��t����?,v�|h�:��#�`��$4�۠���@w��4���@U�t�=Qt���]f��0�z�i�c�Msvv�}WkF=\��v8�Z��3H/ �k����wҁ�v����@7����!��1�i3e�krO}�_M�S�D�@�0O �+� ��}zh|����;�]}��cg�����mȜx�#"s4v��{f��9�4�۹�r�qd�0j8�cR�z� �(�����Ԣ'��L��`ʬ*V��,�@u�w�@o����߻|h}ﮀ���Эu<�8�1��D�n suͥ�x.��.{\�Sz9�ױ6�H��1��=���h^�h��W3��.efPp���'�Z~���������}ﴴ�Ur4�c�6��4�������y�bs�_��d�8�;�����(yϾv�M��Ja�I���-�`�x_= W4�"�/h6���8�F6���-l�U�qH�eQ0.�H�)�bo���v)秙S_ >���N��8� f�DIp�L�I2&T1��
y����0-!)Ja
h�����@%.�S1GlD�О;4��d3��)�&�4O��<���_�ea��n{0��<��� �@�6T��b$A�<z��G���j����{�# @��!�e`���1�HSZ�dx�2!0�lM���\8{������*&�M��i��,��Д7�C =L#�m2�H��Off��Z�bH��#cbA�"U�rP���Mp~�6�(���� q �0�� HK�����ЉT�hD#�ڴ��}&�a��4�a�6���G	Ka�ݞ����|�P/�,�c��T�'�T R��(A�Q�WH�D����14��W*�����_9�yD�A�뻚�즀|R�j�$i�I8G/e�S��8���>}�`lDBJg���>M��BeQ�IZ�h�����o� o���|]���ă�q��L]\�6����,Xl�Zv��c��^�����v��F�*�-
�r��V�߻|`����:؄��C��,�{Rx5$DcR�{f���W�}��K@wݾ5�I6{ﾚ����m���]��}�������{f�s��w$q�f4���{w4���$���ɯ��c���_0X@�X�4Uк�M�1��*k0�*!@�S�_z^γ(I�<�������� ��w�v_S���ـlD-�75�h����<�=����:vD�M��Vn�,^�n�]��r�[�biy��π8���]Np��f��K����<�IchC�rh��[�
&N7z`]�w��T�sTɢ�~�cM��[<h�����4�­�*�XŎ<x/�Hhy%	Kך`��:�c���ـw���1�#DcR�{f����������o�qqa�b�`��FJ���ŝ�,�˓F9e�љz#n{Iյ�u�7<6�c8�<�sζvD�ؖ�[o���ݶ.η[C�s�l����c�Sg��]5��q}�ز����;n:̩ۘv�zZ����Ba6�c��SS�g��)Ɍ{g��DnUe�[:
myd�R�	j��<�n�X�[�۸��'���)�!���f�c��bvk[��G-�b��2h�&��{�������w�����.��'�ٞ���Y�y���@&����:�v�j�ۋ�Hm[+,�݁����h�����o� }�٠\�/���Cs�I�}޼X[�`������%
d��m�'�i��G3@��<h����Zy۹�s���i��,rC@>��@����;�����h�YA�dR14bp�M���@�;w4�)�^٠w�ԱL��ݙ�Ϫf���n�be[r5`ɋ��v��6]���ڎ/l��C2C�cX�r8?�����/l��}{f�z�E�ueYK8�Ǐ
j\ѹ'�}�����$bE�a�� ��J�HD�@_�Tڥ�Ķ�]��s��������%ɊcJF��R����-����-����22`b�DG���Zy۹�[e4�Z��{�72FLncr@����-���m���Z�g���W�ё�ibiA*m�gہ��+��%�39�&�����x�;�%��$�xF����|���@>��@���@�;w4w�\��<��$4��4_h��s@��hx��jȤbx��$�oi6I���sΐc�B�;C��a�(� �w�vnI9���䓞��� �%��$��;����)�^٠��@�ʲ�qc�,Q*��6��5�������ŀp�����e֙�,�<�[��K��aB����=t'7a�mm�hf77\\�&�jC@>��@;{I�w���m��9j�L�!�D�RM ��&�y۹�[e4�h�ܗ�Nd���9!4����)���@/-S@�s:��O�s��)��w����	BP�Q!$�"��R@Ta@!�E� #�$�����W"n$�I ��gu��{� }�� ���m�������]��-��ݔ.�GL���I���ƍ����l*[���!�f���[��μX�7;	} o^ހs���=�&%���h����78 ��x ��7����ei���<H�s4W�- ��{�$z�@�o�4�ISRDF����٠���/;w4�j�9j�B�UC��k���=��K@>�s��w�qO J�IL��B<������9{���W�j�nw\]5Ѳ�l���m��t#QD���˻]���^x��^{l�vSFN�LC��u��S�G�L��U�!�+[���e- ���[��nX���n��F�N�ﳃ�C�ëJ�nu6:Ó�3M&�\�<�%�\t�g���ӭ�p���t��cF���-c�q��)�5h`�V3Ɓ�u��vz�K��sزwOl�#�֤:��@^"�o9.�K5����5u:5�v;9-�Յ���jMб�ö]v<=�/l�V�L�܎Uj�K�^��}�-z�Zy�4���˙�P�	�nb#��^�V�^v� ��&�y۹�s���M�),nE���@/{I�^v�h�ՠ���n6��Ȥ�yڦ�y۹�^�V�^v� ���L� Y1,m��S@|�ŀ>�s��w��sx�!.����9#��;U��k��tWm�e�V�f't��^<��F�X�;;`�=�j�c��.f�pm{Ӏ�w�9�\׾�޽ŀ^���$i��"j8��k�2t b,����l�SF��+h�Ԅ��S�C`��o��/���/l���Uzd�2�"�H��]��y۹�^�M ��:w%�72<sc�@��s@���{�4
��= �w�	 '���!I����٠U�����h.\vI�4�79�$ı<�Ѹ�"6㎼u����t;�.d
Sd,Y�l�dM�RX䆀^�����@��s@���ޮ�q��#lk"rhw�z廚���٠��L���5����/-��/l���$	$L-�"C�B �F �l�*�h�
��,��<H�s4�)���@����/-��;���q��I0�) ��]��yn�{e4fg���HGRƬ�\�͔獪�qTnk�=��V�w^)���n�ǩ$����H���o��^[��^�M ��:w%�72<sc�@��s@���{�4
��= �w��bxF����^�M ��]��yn���;[�:�&�*U]ف�!(S:���ޕ�}��lܗ��Sx�21�)iR�&8�1��-	YW
e)�)��ĚK=�6�9�@�����Z�f�94
��=�����h�l�=������O�ƛrds1�n��Ź�&������!5u�\p�SƋ��F��5�D��ےA���nh�S@/{g�g�y[��Xx��Ŏ6,Q73@�v��A��M�u����h�e�F&5$Ĥmɠ��@�����n�^[4v����?9����Jy��k �ŀ�� w��@�N俚s$���q�^���$��������r�X�D(�P������把���***�QQW�*����TTU��QQW�" *?�X)P��B(T #P�$B �B	P�T$B@	P�@T!P�DYDYP�P�P���T"#P��,B,EB$B�T DT B#E��T"	P�@T!P�DX�T#P��T"�BE��(@T"��T ��($Q�P�P��Q �B$QP�P�1�@T$@T$T��DX,B Eb�P��DX �T"�E���Ab�Q
@T"DX�B$Q$ b��***�������EE^����TTU�**�aQQW�
����TTU�ꢢ���TTU�TTU���
�2��K�Z� Æ�����9�>�
�aRPd�� ����*����	DIJ����AHϢ� (�
 P�BTJ@J" P	PJ
���$�UP$QT�A$����J!%Q         �  O�gv{9�;��8����'��{�9��ܚp�����כO�HPa�����x�]��;�X��ܼڸ�r��l�ww\ ��r�]k�p̗[�wEp��.2� =�A@
 U �X@�oj�>x���N������΀Q�J��zh��ŋ�E��� =}�R8ώ���A�<mۛH�� Sr���7��a�ҩ�"� ��6탐�ӓS���+�x }
 @ N!�P��U�l�59��&�� �JŻj��������ԧ8 Q����{Cū� eriw��Z��}P}�W6|6!�W6�r9�� ����c{��{��e���g�}�;�  >@   p�P�)Y��c�`�1 iF&�  1  N��� 	� ���� f�AJL@� рE�� �  � 6PP0 =` "tA�w �   �)S  �
   P� 0 =�)�� Ϝ���sQ� ��V}��Om9h�m�e]ހ���L���l��U$q�ʺqu*� 3!��2;������ ��}��7c�cy�q���  i�
��J�@ 4 H@�J� 4hb'�UJU<SA�bd ��U*G�T5 ��)����R�  �!Lҥ����w���5�����ْ{=�^�>�������kW�¢���AAT�¢���U����AAT���2������I���?�?����O��Cf&�>,y;�_���rp�(���V��[[���ɏ׹��h��\�b%^�cf֋3���;���x��/�g��j�V�d��"Ӌ�g��o����&�MS�1�G������R�{��{�t7�r��ft37�~<�sY�i�؛|H܍��$"A�m%����
a������mJ��3�GN��{��s;�ag��o{fή�A�M�xġ�*���J�$�D��B���ZŬ�U�z�r��d$�ɚz3�7�xd�>�x='�1�ѩ\�H�Wßm^���<X�9&B��eP]�12y��]���Z��0jH^^_���YdN�{�w�l��Z���c�S;���� �P�q��<'����U4NU�����3�5:��n�L@�DX�H�^@�Y��!XP�2�0�,K�
�)����*J�i��R)�
ı1J0�¢����,B D�A!�E�@E	�ʱ��Hh`M��ba���@��j�]y���顲���qs���t����T�JD�T;��:�����	��靇����%UyF�P2jhl�6�%q��xOO	Y=.����5��$۫�h����5��-��@"���BYRFI:�Б�$}�n��g��8�<(g�T]_�j��ӭ-I��P�[yy���読O'E��7�GY�Q�6��j	��#62u	�k�y�����}��RiHoO����2*�xk=��^�p|nQl��{YK[+�9Vf�����hjYl�ǩ����o�ղlɛ.V���i:�73齻������sA͸�V��_�d�x(v�W�,`Q�o�B�+
�01&�T#v)+�hd+,��FB�#n�q�si�1��i�S����"l�8V����*n4�����w�\ٌ�{�o�S�r5"�E��5�������@�9�teI�\����^�?H��;�j!������ن��Ȫ�/��z�32Ȩ��5�H��,$���8q���]�=�{�7����E����L�Llj^i^��˰m����h��3+��KL5�?NoEc55�sv�Oyg������=�ؕ Zp�J
~;g��j]�w���15Ḭi�T��M��mW_sovߔC${�vW��ok�Ǟ*�QU����w���^��u�^{1��=b�m�uk������ń��WD�L���Ըj%IF%�\b�CDf;BĉT���@���#L��	 Ő�H�лb�qXHSL[ h� ;d-�F��nCG�C�y�7�ik
�e��);�+x��[����r��cw}g�YYmq���˺O+V�۩=�jr�4�{����Y�/C-z�3%��g�ݺ�)dsѶ2G%�eU9a%ٕ��8�skXBx�M)���Hg��0��H�0�	q%0x���d� P�Y"%�%� �SO��c-�+o�Rx]�m���C��%YC�9�9Ym�#;	�zC���R�@ʿ������V�]|O�>��L˒�2���a0��ڄ�j�Y~E����c���Վ�x��y�LK�%Z!��$�wUq3�h�����V[�����_ڧ�#j��7��rc���k��N�_���.im;+����T�B�hƐ�?$D�	���:J���~�'�H���L@,Yȟy��]��5ɯ�1=��Iޢ���ިrLM�`AAEIӭ�o��,�zaɐ�H�����j��{r���;�MW�Fia��2��O{����.�~���B��0u^��4�[�Ds���eN��_�U=t��溳;O{������1���
0�Hm�u|�L4�!�$"���PMW29F�����N��[xmoo�W ��<7 �(	��%�"D�Ѓ$�T$PčS0�H0�$0D��D��5rX��XH� % �ŀ�1"�%BH��a����3��o��#�hb!Bcc-A�4��ǎ��ܽoS9�w+/��izP��<|w���14@��45���Ŵ��=^aqK���V<��e�,�{��ÌIa�y�4�����z�A������=�/��_+�5X����z�ٕU��s<贚2��DQ#�#\)3zq����7����y�a�K�4�;V�wea�3r�C�;�yX!�j���Nm�|}��Iyٚj:����*>X�(����c<�#����k�۽������~�u������Og�N��(Ԝ�S��!Y �%�``F�4O�+����_�ϫk�r��ٞ����^V��WSa]��μ��/�L�xV�s�C%��>�/�u�#�&?^:����+�����^w}~��F>��%]m�<��D��+~\/�!������v9.�ɴ�2[�6(�Z8�xy�	���+�)�+$.P�g�@��c�f�f�qކ!`W$�5��B�B�(,*B�i)�0�2A+���k���acBHX0�)����B�ZE
 B��A�	�/I�H2�����k��@���o��)99[�0���M��g���C��;sm�kSpbR�0��a
ŗG�8i0�x
X#ɨQ}�K��Iʼ̇8a!^L��~=g8d�K1��$�"�$Ja�iBa�"D��cF!�fP0@���!��No��5�aW�b�P�"%0g�Ŋ���vf���L���+4ll�dL�d)*�e*8��.�	��i�]�k�J��Iz���Y�ʭ�P����#�)������G�)_�2
�Z��͏�׽kH�$�X�u��i���:�4��;���)�W���o�>��!M�|�V��A�29�6a�Yᄶ�q6>���z����u���y؜dlbr�AI�&2J%���6�"�1 Hf��p Yc%�5%4�B�D���CF�j��0�佛�C�����2����ܷSy�)IUW�{��ڀ�ʻ����%'��,	]ն\�V�ʧ��B���������J�,H�K�"B4�H`�#BR-�haY����d�o.�S�W�$lmŮua���t���lJ�#c��#<��Lы(��L�ݹW:�曘��Z\Òd�vIT�s���o/�,o�B����v8�-�2cQRc.�sWlb�;��eXR5#bX$t��L(@!�8�d1u�Ł�0�Ď�eIYF$�!Hԋ$24�,XXY1 ��"X�"5X�j�h %�cB�0Rԉ�A�Z{S7j��U��zF���=|�m��`z��}��37�]I�J�K5i�Ǳ����<�Zp�
�L"Ź\N�r�R�egS�ޙŮ&)ws�z��~�~6����e��uzI����*<٩�ow;2Ql�S���SDo��Wcoպ�r$�p�-p�9������pv��d��S��fi�����S	��a�<`،m�q+�~H巴��E��eU���I ���6�NA+�g�Di�!A��N�0� �i�81���$�w ��Hqy���e��Sm��J�ǎQ#
p�<�B{Cm(�Y^�����K}C�"�ח�L��a[�l���헐�Fzm���F�b�ρ(`{!$`D����rkX�%���W��86�����{�x��N1�Ѽ�=�!����e14A1�1�������6q$ @�1Ѿ��c�-�fc곸��V¸�L��)j��UE��n��c���g�4��R$�4�a�P�"�L�8g���z����ep�����N��#cN'J׍�����f�c��Rݰqțm��4B��#eZdTcD�����m��d1��I�C�l����F+����hvR*۽��MV[u=1p��0(�`B�$b@�p�4$K B0�R�� �6㒬��A�l��CW\���+,i�pLtD����n`��NQkV'T�ѕ�Yvn�2iܡ�'�����FI�g�$�:�X[e�"��B�9e���ׇS`4Ƹ����WDaI?,��&=��`�xƼɅJ$9%�:8aZDf���{�����5��&��~�M92�s��yٗ�����Q.����x���a�'�Vo|��}���ۨ��l㞸8q�Sy����龍�E�I�Ѱxl�,Lp$Y\6���h��cm)!Kc[>��m�Os��2B�q���J�`�Zf1u�C��Ą	#��f��e{��/������������a2!HԁY����'�ֵs��}����p��^j*V��!���#�������+�]An:,�B��ˌ����Hē3V\Ԏ��=��l��,�|�2ے�L���N���11��m���'{��l��gG��6�Q��;de�!x���oO٦>��av�fB���e���4�
B��#\tJ��%�*Ơ0t�d�)]��e��U/&�7�p���4�I
[L��+��KB3@�D
�W"T� X�Ԅ�B������¸���j�0+.1�)��5�B����ԑ!2�D��!LqmXUp���D0f~#�����u����B�1h8'��B��'�#H�@`�i6T�i�m�ndn�Ɯ�����_��    �l   m�@UR��l[m�V�Tސ�m;m��	 �d6Ӕ�@�[n�	c�h��n�v�8m�eR���6Q���x�n�`�M��v8��v���D{U�mPcȴ��mM��8�YY�c�mv�*�v����Wgnٳc8���q���`:�V�Wg)�ӡ����Z ����G�t��-�]J��Y��檵M{g(c��dׁ�@�S�Tں�S6�iU]#Af	�3��1�������Pݸ��q�-�W���Z���Z��\6�1��
�&�XS�=jiV���PΞڹ_1��T�TvQ���yj�=�3S��ivB��m�#���-��*�=:;m�[aR�]����[R��U+&����j�<8��q�n����� �dJ6�a�8�wLH�;����Hl���%�$ 6�		k����@-� ���q��d�k�MӒB�m,�m�m��(�B=9#>�*���q�kA|����3�睙�ll6WF��Krl���7eq���gU�L�*�om�%v��}����Ų�[&��nN�<�qu�v�N��X6���w*Þ2�݋K��w[ �Q��e#,f^��z��"5�vBZ�;��o����D	�F7j��kʫ�i�Pn�Gc��$µ�	aSD68��qK��zMlu���&\U�;�Q�*��®�G�[����[r���c�Kj��m��=۔��I�̮������E�m۶ڶ�c��uT�ܦ1l9X�@�UPqF;k�P��UU �l4 mG\��1�8�+��=vZ4[h�` m������g��{vmJ&Z��4�v�"Z�9���楓/I�4�� ��6Zm��%P6ڀ�	<�RLmU�c�����ݶm� ڶ-�-J�xඁԒ�f�݋n�������$d��i7I��
��W������r���ʼB:� eY]#��.�Ā�` �u���S�m���{�n�mdI�H��6�[m|�h��6�6�մ$'��-�u��u�TT9S +���T)`*��U�iI�y��  -��c��P���t�Pq�@R�z�VWJ���P[D�  �`�[p ��q � �kim�^�[@j� �m�[@ 4��i�_kh��0  ��'e6H[��kn�Ͷ��m�mZN��  m� �`m�mm�[@  ���ofU��eH��p+��[G k]e�sv��~^~�%ڪ���ڪUڒ�H���[@ 89��l�§m=�ƶC�HOK��@Wm ��G6��7e�6ٲд�P��m��lm -����M�mKG �,6�M�;u���&��c�������� N� �H  m b�i�DPֶ�ζ���	��q@/-Z�m�g����q�û�ZT�
�IeZ�-��-��B:��۶����H�m��� �$�u+Z�6ٶł�V������ڻj�y��8i�<��EQҔ�M�5��w`���<�5F��ً�q����6+iu*�+��V6�9`�T�ڇvA6{+���+Ԣ�=-��p>�mɘ�y�,���Llb�vHufj0;f�q��g{)���mx��Cb�r.���"n(�sE�R�sw;��9km����<� =N���U�ޖ�LR��X�rd�ܲ�٤ܻ@�[E�Un��*�<���]�R�f�2����ѸBe������4l�-X�s(����>Uw����u�Dt
���M�5<�,T�<ꛎ ����sJ۵��e�k���p�t���lEE�ͽ�a�k	��Sd5*۴���om7�j��qn��tF�ɔ�e`���0r3�l�X�V�,6x���[u�UT�۲��쫳̔@lYj���+��X�h
{M�+<to��4��U`���WQ�X��V�@WWmP
s&���Rܳ�=g��hw�n��T�dD�b9%�%d��,r��,��,q��h���`���Ѝ�[Sl�v�����`kC�I
:��n#v�3M�q�7#���/�;e��ܴL�R�$���ѭy�An؀�2<���v*L��n<k[W>�v!q��: �S�MƳ��� �5�aU:n��s�Un�Y�q��<��{#Wu�4��I34ƑhEԷV�G�Z�1ؕ�=�2�1R��HMF
h��m8ȏiU*�Ul�cfZ�]����i��vذD�  )jT���UU���j�ݜ����`��)����[OK���Y�
��F٪�֠8��sne'��
t;sb�*hг��zWm�f壇S���dA͵��Y��T���˄���rD��4\�ױ�Rsk�� ֙�'a�+�#�ny����b�����Y�)�<��v�W��&�ki��A�*��u�];�p�)�5�s�����u�{�t��;5)-�=�7]�"����c�[��&!9�N	����,����Su�]�3�C�f��tݍ���#���/v��l�֏<s�뫊J�@���6^�n�v���tE�eLA�l+i��=Y�
i�����囪���%�]��rc2P��e9r�m�ո�nN��^����T6ڐ�0��DӠ	z��m��U��8kղ���T�7�
����nHş]p	�~�}�}�M������  :U�KY���q�0ѩ((�U*�[J�ѱ��%�ն� յ�D��n��L��m�` $[@ [@�d�m�D��l	 �J�`�mY�6�A���6 �gZm�  �kX[@-�	  kՄ� J��x�eZ��R����[m6�$�WM[�*54A�<���6�e�&װm��$ 6�n�Bv� �( ��j�m۶�!��� m��)�l )@$�  Ul��l�@UU�*��ANm�H  -��p��uU)�/�r�WT�M[<��V�lmkn  ���  �`ڴ� ��   �`6CL��f�& ���M��� � �Z� ���nk��)˱jj�����/ �nҬ*��sr��,0��		[]��}6ӱ:a �g��q��e�  �`T�.��T��HU� $6Ͳ��� $&� 8 �� $Zڷ������n .�yWm"ʰ*�UT�d��$`�`�pJ�ڧ�o�����[eZq��w�I�Ɔ� ��׈^�m��h ��3��[�W��ڪ�I���lgK���	9�kX4[i�Ā�L��xݦ�֛"������ۂ��\�Bk���f�A�.�*�p��R�UcS�F��i���TJ�8��3p1ĵ@U�	xx��u��A��4�I=V��uI�2���%��ml[N��8��:�Hd��"�P\�Nʵ*�;�9��@{f��Jtf�N�1hW����ie����K��x`�l]\/���J޻b��M�H/Zw+�ڮ�e{b�n{�c�|�B�۵F���6�J4�S��XA�f�U���V,F �ڪ'֟I�I�`(ܽ��|_N�3�'[l=J��C�ic��uP��hS���Z�����⪩�UT9��h)��A�������f��穪�����<n���i6���� M���$�t��@Tq���卛کZ��ѡ:ی��jNؐp`�ۀ�K���z[x�Y�m��� �A��+���+&I���v��[iڇ&gjڐ��R�lڶ�� \��0�m�mZ$Mh�����9�Y��$�n����g������fM��^����N��Ļq�����9W��*�P�s+W:ێ�:�坥��8m),N{`A{�20H@>U�y"wj5��`*�K.�b��nSn�I�ѝ�f��  YmC��U�gv� UmU�V�J�K�r2�{����H��Sl
Sr�w5����݂73v#ܷYF�U��m[eq�!RktcI9�WjZi5l �[���u���b���U2@X�q��@W�d��-H6���UV��T���� ܜӲ�4�E�yP8&(iW��n��j�6X'���qm�a��mH�X���jT�&�
�lÙiQ�iV���K�;4�U\��"�&�c���m89��Z�M;�H6�`���K��mH   ��[m��%��t�8��b�j����-U�v;!J�}�GԫJ�U]�U, ��P
�Q[���U�U*U[J�r���*�K���=J�J�Uu) 6�D�Ym��I>��"F� �u�ړ��@��DI�ض��ۀ   �d��Ѻ3i8�rнv�p�X�J�a�!wT����`�)]�]�9ݲ��R�-�m��  ^�GK4� �[m����  x��$6x����UUUU*fiyUj��W�UꪶZԆ��`  ��'EJ��m*� ���u  t�6�\�&�IVڥ����ʀ�xh )yk(E�s���Pvp�Jt�{*���_o�MRUI%��m�E �� 8m�6�ͅ�����^��4�)Ѯ�R�ۮ�`%v檪�� ,�@��ռ&��<~��w��������' [@�6�km���d��6� p[��H� pi���\p��9�� �IrJ�gH5	�F��lհ6��>�v�!n�ִ�DLP4�К��B����U?�������A�$�0 ��dGp��)���R(E�;
�hB�����]�M�� ʰT".�P�(��1C��EM*!�A��>(?�v'������l6�I�	����`�d!�GC�8 ��
�
G4�?"`'���U� �
�TL=U<� �)��SC��! � ?�}U}U���E�C��>$�$��"1H��.�Ч��(�#�}P�@���lU�Q���C����@$����]�>
��@�M��D�?��z�@$D�Q��H�DB q4��/�=R�'���E�z`�؈�C`�4�PaA��Oʸ��h�m5�?��D��`yU�� �PD�D �CH�@�A�T�j<����
�B#���/��b��4~D=��USԮSLVA?z�R���K�!H@�@J*A����.�C^A
��1<6'@<�� �p���$	%E�
PNTKX�~<@xp���*�����$!E#b�j:T���*x:�l����%)PU�))aJ+mi�l"e�������%���)l��V6��ma5,�R0 ���+($�1!J�z�����b�$d dU ED��� ࡊ	��x�bD��/� +�L@0 n�4��b��������	!�VD$R��*!�#aE
@ PR6
�����TdZ��v][n�k�����:���6�$9oW3k��ayo[���u�^-��	�n�v�Ǉ-+�os2"��ν���dۯ#F��ohS��|�<����e۳��Vg%�����=�v�k�����[s�	�CZT+c��
E/+ek�ĉ���/<g���2��v�;�lGD������@ۢ.�g�uiļBq݋l�
�]�ѭ����.'��']�p
���99Μh꠺uڱ�-H���q��@����n�UX�<Gd˱!��[�����W��щ�9I��Mr�R	)�ݷc�P��z�x0n�v���Z��tn����3v8�z�a0a��������ׇ�f�*�	��IY7N�d:K�I�Eqn)���k�s���Ӝ����˕�T��dl��& ��v�G�E/n����d���[Μ�nn)�c=q�s�;U�vٱ9�q�����wvl8�/<g�w伷��������m�&��qJC�I�ݼ4�pP���9��-5gd�i;k='�Y�g�&�z�u�ٻ`ރj5ίh^݌�έ��:�V�t�ȴ�z�&*����˙y��v�x��41��c��������e�g��iM��k����ܠ�V����V��U��A$��I �����1v�-��vaU�j��w%��Ii����`r��^S���!��n!l�/[��1�0��=v׬���/V��&��n�il`�n�av��'<
bh��8���ł�kQ�5�v݌��;;<V%�Ce�{=��Y�� �SK�݂^��G�f�}���xޔ�e���[m��PG=Fo=;��t�n[���q�r2`G�s��%��l���]�9u�K���q�ʚ����g�:���W�̃�@��ux�F���C�մ�X�%6��з�1�$�v]�U� ��ӌ�NY���5��v��\p+íc<u�ZɶC�]-��{"�qz98��X� 5S���f��e�LշF��k54�x.mW�O�W�|�؏�v)���E�T��J"�T_U�
>��|@_��+�1��@�<��YzL��am�[h��p�H�8�;A���{W8H�@35�N��JN�r�Xs�U�]�����k�#�-��l
�*Ǘ;�����x��+hw;�� �ѥy��s��'�ɇ������bG1��hV���U�� �.�[;E�ۧ����-�p����d6�v�v��l��<��*'j34N��^�m��3�
58��k2ꖨ�B�Q�l�29^��]�s�L���n�eC��@y�<#�*c8Pi0Mb�}�ڴ��P��>�3? ��Ɓ�?Q��acY0mŠ^;E�^�S@�즁x�Z��@'�'�DڐZ�e4��h�ՠ^;E�w�U�V��DE"p�/;)�^YM��-����αԦ�@�m���h��hvـ?�ـt(�ֲ:�M�e*��pd�K�\�m�6�.�bR�
ŭ�aE�6�Q���P)#rA���lJC�����^�S@�즁ye4��\ei)�I��-�K�'�y�f�T=P8P�|<U*8��S	D8��ٙ�� ߝ� S��9�U�F<NcI�@�{)�^;V��J����=l��λ8�0M�q��ڴ�Z=���^��|�z6L�"CɃNW�=���9e4�)�{�%����$y��
ܺ9�f�A�R��U.�(���6�Oev����#�U�]���4r�h�S@��jzz�X���dDR'�����9;�k {���	(�>��6�T+*��� ��� �w\��Ȉ�B $��E�X��\TE�}�)vJh��8�p����F6%!�qw�=���9e4�)�w�ܸ��S��&7�/{)�~��/,���{S�;�D��H���2{e�������m*&�n^^�����ju�=��n��z��$�hNcI��留��hW�=����,���
������
!)�g�M`��~��9],l�&D�5��4K�5�=�f3���v��}�6�O�O�#RD���h��/�u�ܟ�����T���Et��_'�wΌj�0Ȉ�N9e4�)�qw�=��p�(��-�.z7�m�g��]�d� ؖ0�M��i���yꌺ�v��v��[���l�>��5�=�gD$�Hn��l�?H|�C#��8�ڞ�{�M�����;�r��io�'�X��� �m��;f�{k�p��k 9�ӨNbX�sNϾ����|h����������h�,�VL�☒����ڴ}�˶�O�z�� ��`(D%(P
NG�0��¬֫/�g[C[�-�K��p�!v��Y!^\lְ"ɞ�w*�� �uR�X*�6�;x��v�G�Vۥ�n�Pu��L��6�렷S�:��ׇ��E#��Z��A���5[��:˻m֥�Ѹ̙9���ֵ8㰶���s���n�������͓;�n�.�9��t\�\J*%�ʹvv��̮�ֻm؋�	�������w�������d���Tp�̼�:^�^h��7m9�ܑz��Y0��u.���벱����4��h��/�@���Ņ��w77w�=�fyD������ƁWWl�;֨�4�����w�S@�즁Wz��/;)�r���lɄM��4=�/v����^vS@�,����뙍�21�)��٠^vS@�,��x�V��������������v�ϐ"m�^޻g��	����q�z}$�ζ��s	\���ʩy�	�������YM���ffg���= �s�̘�%�'2D�h����K!��H!JFZ*��	�R�1���p*$�t+��"6J�ݜ��/� ׯ�w��H�L���4�ڴֻ^��n���M��U��$�,dʴUU�B����Հ>�ŀ7���ڴ�kHs��ɒ7$z��`����}]Ӏk�wX�Q+�޺,��HWK�6��:�pp��̠t�,�ةnLIm�#=sp��gn��Nf�y�M�ڴ����n�����9�&�rm��g���=����/;)�~V�:�0$�s*��� �Z�m���!DB�"�b%~��
�Ie�� ��f���[mn1"Bi���w4��h�ՠv����v�ܘ,��<�#s4��h�ՠv����w4t� �2|	1��1�NEl��,wv�3�vx��!RJ>"�n���kSӰ[)��ڴ����n�y�M��U��>k�Lqh��=����k�o�#�~�I��"2d���}�nh���;]�@�}����Rm���LPR9��e4=�}��y�y�rb<D����X�C�_@���3��nI�s��EZ�fn��]78(���_����4ܲ�9�F�Y1ĂLrnjb}qn�����u��I���k�H�s�� ��r�c	1��F(��/_lzm���YM�ڴ�r�[c�cD��]���Y�L�o_���k����
�0pkɒ73@��)�v�V�z�c�;m���Xu)F	@x�����Z:�c�;m��/{)�~]��|�1/���W�������k�0t��GȈ��*V#��}��\4kZ�]SkB��tcls�q:9�ţӎ{<�˭�8�V]d{����pl<��\�n��� k��6TJ�qȁ){&m�-��ݻ1D�兯M��n8�9b��������v��>�g���7�Üt��V����Tu/3;ûJ�����]q��t����j&�.�[�W�=p��^5�t��m�ف[V�Չ��[��t�&vE� �x"��`*p��2]C35sY��P[�Y�8:�W�k-/mvw�.�(�@m�ˮ��=s�q'��ɒ7$z��M��h��=�t`�)���"p�/;)�^;V�W;^�{�M�k���2`%��/�@���@�즁y۹�qr�:�8��b���@���@�즁���h�ՠ8i�QJ�*��̔M�`vـz;o�g�=��-�v���q���DF��rݣ��.��!\vz7���;�^�{�G�Ką�8L��ڙs4���������(�_�wb��P5]7wn��ۧUVco�W�L� 1"T�b�������7ɻ��=����;�w4.�U$���>�4�q^נv��h�n���V���X�N1�n=��s@�;w4��h��zz鍉�0���&�`�ŀk�f ��^�X/��˾b�X�cԓP�f/����d�����@{OL;�x�lٹ���s���lʙ�_�}]Ӏ~���m��7�x�+ps$D�b�����^נv���7�x�{l�IL�5>�"�i\�D�� ��,~׋��
(a��s�=r�o 5D=�r��u(��	4%�N�Õe]H�Q��sBn����7������0�^K����6�]ۻ������'�f����U�k&,Lc`��i�nU������0��&65HWB�-����͒~���lG�����P,V���|�E�ʕ�n��^зu>+6��67*g��~���P�Ul��Y/+Ia�<�ֿo{n��$��Q�L�d�?+���9b���K�fVdz"B���� r�6>5�b`2��i_?U����jxj�5�L���3O!57�I���ShA]��t^r\�6A7uӁ_0S���nh�ɚ�!F# �"��oK�-����}u�a`���ї�R5`�$����g�2�虎��A��'*�����>
�D����h�b��0�E�!v��q�EH�����B��R
�"?�!E��0��X��6T���WUV�9%
%��� |���u��I/$���w�X�Q�W��T�6Tլ^�0P��ϫ��b�7����ﳏ�_F�j8���#	�'=2��w�g�f�s�=� ��%f첌GNf��\T�H�wg�>�}X�x��^.��ߐ__nh���8��FDd��@ׯtz���ŀw�ذ���y$�d�~1<l�aAH�h�ۚon���u�k׋ ��gaڨ�U��Lݬ^�0ε��^,	B�"%*D��1g����:+�� ��A��+�qU�;��x1�̑LS#��?Wڴg�">���_b�>���>��Tm
ԅ�u�{3)�N�����*���ܯ�`ˌ:�܃����s�o(�
?�o�����`��X��8�Z� >D�L�ڙs4�s@�}�@�_j�;{w4�c�71��4�h��h��Zon��v�h�:��E&5�FL�h��Zon��v�h��h���$L�Y �qh���DB�������pε��F"<}hAb��-\#�e��3eӹ����v��	9�M�;]G�}L�T�ܙwG]���ذÌ���.��?������C\��r9p���j�8e��6sz���;݇�#��.�nn�^�9�,v�R瓵gY��ۊtf�� �.��ۨ�)���pquˑ�.�]�V�7n,q�\��[���+��W���$㶻K&U㗷q$�^&�Q�5��j亓4SX� �U^S|��#��v�77.d��wk��h��2���\(��9�N^�p��v�,Sw��x�u�pε��^,󭪜��<	��%&h��h��Zon��v�h�����F4�L�RE�~u�pm��7u��5� �|�=���"R-��s@�{w4��h��h���0Pkjdiŀn�ŀyDC�~���5�ŀo��~=�=��g�
�EΉ{ٻwo#;,��q�˺Q���#�^5Ga�R\�[*��^,�s�k׋�$����h]�/F��1�&I���V�J"#a%vK�`��X��g(Q�bG<�q(��bY �qh����v�h��h��Zz�H�����4�s@�}�@�_j�;{w4����c���0Ĥ�����s�k׋ �׋ 舄����E]�Svm\��*#���h��"�Λ"Ћ��.+�撶?�����7O<�8���{Ӏk׋ �׋�H>�Ӏy�=����O"m$�_������-���/���?Wj�}��~F16Z����6��m�T)�̢�H!K)	 JB�e�2K,jJ���_=Uz���.�{���~��[�LcD����'�8�>��^�X
[}�`:���1`6d�����V��ϯ��/�6�����	��l�Խ�Ƣ�x�y�l<��k�f�O:
�S��y�����|�����������?�X�X��=
?H}��8t���T.�.I�nn���y%䢫����;�I��_�$��{�7����uP�e*��b�H�I%}/���%������������$���jI%���S�A�b�ӗW7d���~���I$��ߴݒOW�ʛ���E	�h E �R�g�qP�/@~�?{��[o�ON�N�
t�U$�nd�O}�ݒO�������J�_/ߒK��=I%�����Bn:n�������K"q��n��۵d��\�B�t=��6����#?���ok#*�*��R������RIv����IqYG�Ͽ6������$�ց{�8��4@@�f����n��#�H.�}?���I$����M�$�{�}�|�K��E2H��&��~I.�_�33�_����!/(J����FL��z���� ��+�]puc-����y��}���$�����I'��}7d��!�"����=I%�����ǄB��L��$�Z򌙙�(�^J;߻ӻ32���ffu����$�t�x�F;�7"M���c�:vƝt*�����>C�Wk\wSn�v���+Q�a8�Z�"x��He��`;n��Z]����v��:��Yy
����[WG]g������[�a�����љ��v�m�E�4�`ւ�����tJ撖ݩ˴Nu<M':@���#�	�9�Zۣvw�O0tWE���d��;I@U��N�v��\�.8�ի&��]
��G`��[Na�L�����]g���ѡ��ᶥ�z@�]�����-;H8�<��ٺ�k��ل�5���$�{=��~I.+(�$�oo��}��4�w��I$�{?y�k��8�q1�� G����}�T>���7d����S�$�������UO��?���&��ԒW�߳������O�%U_~��M�$���	�I&���_S%3!s&�e����|��~��v�{�����Iޯ��$�U_~���H�������ƈ�Ԓ]��~��^�3��n�d�}���n�'W��y$�{�����3�έk�6������)p��[�l5���Jn�^N�����9X<�e�� �c����I��G�I=���vI:��S� [U$���_�$�}"�dND����Ԓ]�{Ü'���"BI�E��B���$(l��`���I0	M\M����HK	�M���o���pT�'�(y�׹���n�g޿�M�$�_�~I$U'�;�QG���rܹvn�#�}�^I$������Fd��j5$�����?~I.���cx�18�����}����/ߒK�{Q�%=���vI� S���y$����W�.�v9	eӗW7d��dy$���#�����I��MI%�;W��$^�6�$A�=si8:sÌw^x]����Зgq�嗏1�uN7~�����0�y�B�Q����i�$��;�$������.�{����I%�*���,lBy1��~��G;)3� �BWw'����7d������O}�����*o�����K��؉����~v���<�y7n���"�KZ�b�Z@(t%S��_�#�$���?i�$����w�I;����e�� �e˻{�O� W���O$�{�ߴݒG޿������߷�ݒO~���K�w#.2��uu2I'{�ݒO����~I%�����Iq�V�$���ְz�t�*�v���n���V��8�p%K�#y06u�܌�߽�����|�"��I�����'{����'J�ҿ!%�Q.�{�~��W�1��a11��$�����*�zWߥd�O�}�M�$����~*�����W�.�v9	eӗW7d��_~��$���i�?� /�	]����9�$��=��~I.��F&��<���"��~U��q�$��_�x��_���_@*h�����ߔ5���{���:p� ��N�����g�sۛ��||���$�-��2�r�g�5����+������{�I����Y$��{�7c�s��WaW�=�q�k=��.<���S\�|�Y�J��\����������}nD�ɭ��_��}���7d����VI$���O��uIl�5$�_n�d���6d����%�^��?$	*�O�}�M�$~��;�$�������I"���]���ʻ��v�uY$���~�vIz�w�~ U_~��Mؒ�w��I.�fT�0,!AE&~���O�GY�y�����w��[o��=�ݷ�C�Qֻ�~��-��f��3�e)4I������������+�{��쿬�~�����>���$�Y���������J�#Jg��*Q@]�ە6Fa�΃@F���+\����}�H�Q0��2��U�$ͪh։sF���"~Hg��X�c���(��L2ª��H|*�Uf�U�(�+X��6�+ xB�wt<��9�'?e�5*b_�kZ�\#�Ж�ۚ���m�P�����0����u�Ԯ�����}@�ٯ����q�+Z��H�=�Fx{���8�~6\#<6Hg�D d$F`A���F	Į�ib��@� ��x��FI"��BH�0 ���B0bD�XH��0���'~t���v��"�3��˸�[�Gv��*�;�:�/�-v����t��'��`-�#���qD��'<����/��d�<�H����Y���9�v�I����I��ݶ.�˰:��rt�67���6��v��8St�-�$9�6v����X@�9�@�c�h�6��]���HU�9lXv9�B)�\��Z^M6z)�H����5r4]�\�Um[�Y���  t/(d^(:��]Eͳ�����@7fm�l��֩�u=��O;A�y���~�~(�X�u�d�(uS��/-��2l�{��Un��k�&^:i���l�2O(����7��5�\�����[�^rO����~�^�Ͼ�:{�8�K�1kL�������(f�Hs�CWXU������X�h�T�8����z���<�m�wj��]ܷn�v�Fك�K��։n�f��S8�����ñn �ޱ�;��Zg�r���^h�q^�c�������:�{���)�2�Ϟ.|���q!:��w<��ҥ;lln��GM�ɡ�NP�x��7n��Z�ݘx���,��k��KB�a��r�<�O-WzV�����1 ��N��w>��@��3:ڬ;�d����l<h�m3�#Z��X6,�*��S��ȵ]�Y���Kyy�p+mP��PF�%����Pg&�l���L�[[/nKֽs�i�[v��<�q��()��gppu2��RMl������9���c|��l|��KƲYY�6��z�Jzzo9:m����V��r�t��uԬ	'n�_.X�>F�F��g�dݻmp 
�2qp�y`��T�ۄ��S��W+\�=�f˷l�%�@{[b�c<FaN��je*���[I�B�vX-����Mf�%21�0q�ѷ�me��Sd`��':�"M	������f��`Ht�{A��ܗ*�\%����]*٪J��S�D��֜�Eu�(5 Y�pm8��a᛫u�f�L֬Ԋ�Sj��ӊ�P�*�D�8�X��@�0�D����T?*���g�r��FS5�WZ����Xh�9��f~�����<�\D:Qv��i��k8�[Y9�fM�M���U�̩�O�O�'-g5q�0�������us<	/]��nH��=�ܶ��lW�tYE�q��n3n�ټK��!��W mG��W�V��fZ3����|�2��V�����b2qq����n.�k5�Z�W.f�.!c��a��\�1��5pK�^ � ���s�.�Mj٭�hF�x'�]�6�퉛ƻ�;=�\*��km�����t�s���l]8��� �/�>�I����H����$���}���7d��Oå*aL��T�uu2I'���n����&��=ݶ����y�m��kܻ��4�2�y�bI'�Ng��$v�T�{���v~B*�>�βI'߾���O4�r51�Qȵ%�3�n�o��z}�d�O}�ݒ~I�����I"����L�16d����%��G�)? ����wI$����I$����vI$����3UV�M[�O`؝a�y��V�f6��Q�mt�RK�UW]���{���䆃tevL����wb�?}��[�y%P�%���� �Խ54 �\�d�խ�?~�^���#1IV",����%YQH�R�F0�!T��"D
EN���7��8��V��Y�興�;޺((�̩RZ�*��;޿啕â""e����;�<h�ˎ̓�#�Ĥ09DDO�o� }݋ ���0:""%�o����?��EN8��w4���^q��|`��s��������W1t�[qB�b�u�Lu�dw�ۮ����'�sq~����6��n�`�]�kv��ծ|��D/�;��,�ic�L�6Q�@��3�m>��v,��l�G���6_#�6��1T+EMY�k����ņ�p�a�
��=Qn����nI�;���9�{]Qsur+�]�uw8Q��]�{�k��koˡ(���`4�ɚ�(�!AH�h��@/�}�����s��h��h�>�q8�_'��5&$]����۵���gy����V�#��1�$\ZO�{��g0a��11�~��s@��ڴz�tD(�!��� �yr��v��L�ں&�����9�Jd|���� ׯt(IL���U�y)E�T��� ��,��lÔD%2��,�Ӏ}�L�B�e�34nO�~L������� ��k�.Bi���P�`@h���TA��|(��?�������$��aE4�u`P�<�!k���{�ŀ~�m��}���>��]���� ���c�9�/9#c�H�ogh�&5t����1O������O��N��+E]Z����^,��l�K��������qDd����;{qg�G�%F��{�� ���Y�B�E��	7�@"�f����@��Ň$�L���pϱ`��T���HZ���Uf$�K�ߖ����5�Ł����8�>�\���SV�bm]Uk ��k���!.����}~0m�h�ٙ�d9��$ۮ%��R��Q��뇳+����krbf��:����cm����^�ݤ�q$r[,��
�ۋ;vu�;Ms����s�.Ȉt�ז�7lv�6w<a�:��Gf㉹v����ܝ���������Hpi\ꤗe㝶�m��X�QT�mӬr�a����B�Bl��N���V�9m�I�"�9�A3N���I�6�a]����u�x���YѸx�d��i�Cu�v�I^�����9�b��KG �����s�|Z*%VQ��������1`��f��9$����N�C�8$*Bf����~�e7�Y�ޞ4u�-�������H�i\�L�6JE�_?y`��s�B��}݋ �i��N�;�Wv������p:"�����X�>ա����Z+��dM��wv`���<�$��B��;����-�{)�~�>ߜn%xb�&$�C�gi��'CNuӖ�M��=��G^�rq�N^����ﹼ�o�	�A�&~��-����ֹ�
�ϱ`���ʥ�)Vh�.j�I��s�����[���V���k\璄��BJ�s��U��M�3E�7W8�w� ׯ�BK��-��-�����c��a#j9u��BJ+���`�ޜ]k�DB�BP�o�Հo�A�$*B����լ�ֹ�5ֹ�?N�^�X�*�}�n+st!�u��]����ϳZ3�uٗu+u،�4�k���ww���@:��lAS���pӺ� ׯ(Q	~�����:�E2H�4@�h�{^�}�/(I$����� ޮ���\�%
!$�����q���@����?w<��i`�`A$A��� ��$@H
��,#�Z�%�X+�P@���|�+|��n@M�.L&%��(�������>�����(^��U��|��%J���)-J���]k��D$��}_�|��V��?�>�}���q1�
B̆LU�2m�������J�Pt���5�٫�[WWjfWD�\�����5�ŀnֹ�F}�~A|�^W���i`HڍǠk׋:DL����S��?Kn�В��F�.��J�
��SsV���N����D���Հ>}� ���N6�>l ")���1_K�q{�z�|�f����Rg� m�=�~�@��d��� ۋ@��u�k׋ ݭs�k�s�z(���n,^�����RٲanA�M��\nY��)�s��0��y��������]��X�����w�`�k�]7<���O>���UT@Z���n��V��Q
d}]Ӏ}<��m��(�Q�QC�Z��R�B���T��ޯzp���
"e�v,�0����v��L�j蛻������V ���m� �V�����,	Q���w4Q����������P�BXj�Ӡ/�4�71��AA$�8�v��]C^l���hj�͹�[l�`F�lTt5�̔%����v�r6�Hff-$�0$��p��4m>n�۲r\���Z�v�I鲯���5��m�Ն�N����I��b� ΃[�i淁�[`����!�����=
�DͬgL��gԮ�E���@N:z��/T��w\�c �g6+LR��������{��>���o��Z/cJf����=m�q�������
�Yv�.��S ��챳�BkѼ����Tڛ���y׽8�np����~����4tj��cO�"�Šv�g:!D�����/��{���΅!���2A�Ɖ�r-���@�sO����]��/����v�ȣ��HL��`rJ������N �78IB��}��<���UPyR-L�W7k ��k���]��?��u�`�� o���渻:�vk�N���pn嶁뉜c��vN��ۮZv�����	�9����M��k�h��V�m��Ͼ���9�|��g��c���}RE�~��[���	R�L��4���q�
�%`H4��	P��7Fā��v�n��O�W�Mo��7������9B�
dj\�TJ�6��T����݋ ��k�<���%	U{��N��Ӏ}5jG$�HUTڛ���~��� �k��ծp:��=�ߖ����dC��DB�8��j�=�B��^q�ϱ`��s���urM�G����zW��M:�XI�;.�j��&�u��5*�u��?������}��g��p�6�7|`���?mk�B�BI}Aޮ������RE�
I��s@��ڰu�p۶��B��J*�O�ª�<�-E]լz�Ӏk�s�����IC l�����2��ו����pֲPˉ1s���$~��5pۤ�F�܁E��;�Vr
���h���3%q���H� �)1�@10`���|yZg�u��T%�;	þ���R*��)�/��3j�hk�o/��d �,���R�
�v:Hh����X�q&i&�4��_t;���kRB�+� ����%��~Z��#�q'0��wV�њ4@�!\j�@0������-K����㨞�|No���	S�1 �!k��_�U�!u�� ����$�BRF0�+0�p+C������6��#�.�Wǂ�H�*mC�`  �4�8&�ҨqD�U�D��C�U���x�*�����]�t(���,�^�yh��Ʊ�B0x���W8���N�w�����ֹ�?+���7���F%!�~�e4g�}���_��w�@��ep��v��Y�����m�5OQk[��8n}��n]��n:���}���=����jQk6�{���Z� ��IB�D}A��� ���1�@�6���@��ڴ�)�~ݶ`-�Έ��>eur�Ԗ�Q3rM��� �����DD/(Q]>�� ޮ����s5j�)Q*���՘�)��� s�Հ~��8�B�"�# � ���yɹ'�3�XE$HȌ�RHhVנ{>��Yz ����� �Ky�s�QE�\�������M������$�m��T�≃s��9rd���ɛ�M �Ę�p��Ӏkv���%�A�wN �܁I��<D��qh�S@���h�ՠ~��[��8����x���1)�O� �m�
&~t�p�|`��l�S��USWw8�I/DEu�ެz�Ӏkv��ֹ�?GڭH䐤�1�$�?u�����}���W|�[w�yBA���BS&�Y����۫[�^�a���p���uj��u:��S��˰{q=���>�*N\�!&^^w�s��^ܚG��7iQ��ԫ�q\]ە.����8�1�N\����q���d�Kn���.횤�cR-��)��s����R���?7c;>��#����]x�T�� �Z.���)݌���+�F�瘫v�:۱�����=������?��;^bK%]�d��l�L�t�X����i����*V{�2ݟ���o�O������ݏ��� ���p[w�~��8�tuI� F,m�qHh��V�3�zh��h�S}���{���$������?mk�?�=	Uw�~0���w;r11f��&����hݳ ���p9%2����bUB���n-��h������4�}�@�;(�DdI��q�&ݟB��z.��`�;͔�{lm�F����n��|O���?u�� �h�۹��=�O�w*?$����h��of���a ��eX�⡛�f���,�����h��:T x���7$�y۹�v�M<�<__M�Z�ߦ"d�%�rf��?]� ����]�o���y�LP#6�8�4��� ��y۹�v�ՠuv�lU,nH�Q��ĤbF&8{/�S�;mΜ:q]��mZ��v�(��	�@;{f��v�h��{�y�-�L�y	�0qɠw���k�Z��V�v���E6ƽ�R\�M��S��?:�8J��DD%����"@��Aj�P��g8=��;�nhW�50����@�_j��٠w����_K�{�+��	�����@;{f�������|���� ��P�B4��[;Z8ɚΛ��qŷ�=�3��or��bY<F�(�X��Cō����;�������ֹ�^K��޼z��z-Y2c�N93@�}�}�$s��h���;��� �z*�10�Xۘ�qh�k� ׮��
e��X�}8�S�p�8�&L#�h{1+��^�nh�\�b��D4�E}5�p�������0qɠw���k�Z��V�v����ی�D/�i��b�E�l/lGQob�u�/b��KS��k�H��ܮj|�b"MI�k�h��Z�l��I$�H=}� ��\�Ԗ]"�&�� ��\�D(�wb��� �M�tDDL���:�隠AuU5ws�>�ŀ�l�;]�@�_j�9�q�K�&�������h�ՠ~��h{��1_{߳@�h���!23�X�@�M��ֹ�5�� 7�w�|��!D@
�h@"D���-ks�~o������/���.<<�d0]'k�<�n{u֩�A���·��ژSl3�o9ㅮ����r��Am�۶��M�E�kG^*���6�#����l�3�W17A����ڴ]r0k�c��{����&��(��vݝ:"�����s���&�+e��泹�7P=N��G\�v�Ϝ��9��فZy��-=C{,��jٝQ@BP�=߽��O��O�h��ӥ6��٥�3�#�%�����;Dv�t�̖`*�[b�K����Q���;�v۹��l�;]�@�j�g�&L#�h��o�bA{}4��-�}�@�r�k�I��1�&hy�4�j�?.v�����.L�����D&��;l���s������Q?k��6w��ڒˢ��UBr��נv۹���4l���~~��C�q�<�
)�Z���!�\j�������"�q�n���su�u��ΰ�v�USuW_���ŀ��xn��D$� ����;���=�'�`�@Q9���{�� `�c `�0X+��Ԕ/ߌ��`:�`�ŀ}�I-�y�D,qɠ[e4˝�Og�f%�{ۚ��M �s��LL&5�9�9��k�-�s@?s�h�M�u��S"Hj`ۋ@����f|����{�Ɓ���h��~q���1ӧ�	���1q���S���qشd2�Ue]zNnu9r51'�cI0���s4�;f�oe4�}�@��s@�ː1��<���ܚ���?q�������k�?.WqLR<i������j�/�{�s�H�(H�a"����0"0a�P��_=�h�}��\G0]Zi���qh�=Ͽ,��Հ7����8��-$�%�<��s4˝�@�}}}�?λ�v��h�oO��ڄ�G�O��mƋ��Gw�%=�c=�t/V��v�"�{�}�7~YF$@n8��_nh��V�on�x�V�w�E^L�&5�9�73@V��/BQT{��X�w� o^,�u��&24�����on�x�g(�BQ^�{�^��|ժ�)��"�&�`tBP������,�^�w"�EB�&�����$��4ݹ��bɈj7"�-�ŀyz"!G�{���{ ����7�xcuF���-��2c��l���u�<s[�ҙw[�p��%+n)+��<��n;UU��M� ޼X��=	$�H>}��\G�YZ�M�6Ғ-��s��$��uw� �w�`�ns�!L�VSؒx�&�73@�w�@�������{k�pϱ`������ȦK��p=
�}�`;�X�x�=���/��^����cXӘ�s4?7X�x���pz�` �Wf��M��'0c�Q�6->	�E5�Ț�B�G�	n�]s�Ӑ�^)JҞ���jFIX�@w��H����,�-��*a(b3��ɗ!%�
K.$.�?�h�Î����Bs�q4�?O��P*~��FdS�c��!t�x�z�a^�9��$��Qg����L�y6��n�U[h��l&���qv��ِF�qT��u�z�t�qqQ6hh:��u��[��l+�a5�4��㳺\�q=I�A硜�K]�,��Rݭ�r��$˛(m7W����{D����c1=�Ts���n4n��mط��&�>��\z�Z�Ƕ� 7q����x�x1v-����Xe����b�-�X��y[���\J�'e�Tv�C��o:큦�vj3�i�ͻ��N�[U,��8m��F�U��Bved&�RMč�
��
�N�� �,j�mf̋mj��� ��6j�L�į���ص#˰�N��w��^��g�t�����c�sZ6�<\�z9�[�ٻh�C�&�\��N6y���<����,�WZ�pFI.��z��/�MD��٫��8��F@KZ޺&�C�zI��vL���5���,���t:oB�!:� ��e�h;sv���nm����jP���whMD�N�����&S�C83���n�d�u����ೃ�)�Z�x���{u-q��o=���3��q7��Ų�۱�RSl^��ɸY��s��`�t����]��}Fq�8���mt�NP3D�)b�cB�s�n�
�v��S��;Em�t�2t2M�pW-�#�يU@@c��x�4h�	�n���lS�!U�en����:��0\�Z�m2������oX�AɆ��c�+RL�vU�#u��r��ݙ�幰e����:�%�vۓX�݇��g�)���9ݞ��
�W
�� `3ll�7m�`��8\4�cvl�V�8gۺ�⁡�Y�v�k$^�܂�Ͷ�9�䛺Վ�׮v��	Ѽ��l)��rn�릮��m3�7�v�c�̬��7S��祤p�'r��j;��Ӂb�gEQ��
�v�7d�n�fv�t݇\`v#��8bj���;�U�wT,�+p����5;u�d��t��dn,�:d�I�����ҹbṀ'<htg�dV�l�:���a�x�Y�������wn��j
���Qҡ_ "~D
D]��W�	���F ���b�	U�#�'��Q����Ѷ�^u�!�b6���[�3����4e����n�v���B��eH�3Ɇ\��������6'6g
�g&�]7.�L/M�a�q��ݗ�����mvxA���½B��z;�v]�`����x�mdD��9'.ng�q����+�gc�����2��^Ŭ��W<N���%::�k�6[���"ɬI���Rе���?�����s7������68���<�)̗`�1^I\�y������������B��"j�}ذ��p���B��Q���Հy?+
��L��4M�Z�ֹ�׋ s�u�7�yB�B�w�D��S0Ɉq)�������Z�{w4�ڴˊ�&)<l�Ńn,�սՀw>ŀ=�s��%/�~Z�{��4�#mG#�;{w4�j�;{w4
�k���7�ja��0�%8���v#Xj�u1	��י��v��Z��_�5S2��®���{�ޜ^�X�n��G�ϱ`mH��*��q2XUs�k׋��U��I/(�Y�����;{�`i����uuj"cXӘ�s4
�k�;{w4��ff%�}}��~��p$Ɣ50N]`���ֹ�5�f$�OV�Vr���גl"�f�z�V���}���:w��m��F܊]Z��Y�r1\��Tj�۷��s���}��w%pql��l��O�8������LC��h�S@s����^Q
<������ �s�"仕J�����0:�g�D(�wb�9��6�脔�Ԝ�eOT��T�]��݋ z�JIj� �o\)�����nnI���נ~���A&ı'�nf���z�|`�|`u���D�w~X�R!�J�t\L�MY�6��.��_���nh�S@�N��&G��>M���qjn�hО�h�K'h���%//'ZɆΌ��FLks$R]��۹�^�Of~A}��@��&!&�	����Y�&Nu�8�0:�g�$\��4��M�I4�s4W�-��0�%U���X{�ŀn�Ys4J&�Ȫ�j��""_vq�t�u`�Œsd��ņd���*�IHP�D:����Қ��AM8G̞��鍽�����[��q��.��n�m���� ��%�s��	��d0�7$Q��s�	�c�U��t]t�͹`ǘ ��#!���C����ڒG��{s@����)�Umzﻏ��4bl��s4
��}�fd������� ��,�Ԉ�r�]�1" ��@�Vנv۹�Umz�ʜD��4�H�4]�@����k�;l����W��I���m��Vנv�M�l�2#�B�D&�Q�S��.���σш�/��5"�:���m������`.����.� ;��#�Ԍ[�la��n�.GCF�l:{t��c�ѶZᵮ���nz8�x���������E8�C�MvWguNZ��v�uFI$��Y%5`v--t<ݥ89ix�5v�����v��59��mŷ9N+�5��f�W+JӫV�V�뗒�\:��������{׹M����mnט��n-zW�m�ɓB�۰Թ���\밽Qdǒcl�6$ґ��\���ـ6�� �� �칚%i
�Ud����3Д%2wu�>�ŀUm{��>�#���� �#h�ō)���[x�q#n�nـj�E��
���,=��� ����5�f�m��?}�}($�d��9m�С�g���� ��,��u��z؏r�۱�FD���0�f��������O���V��y�pkl,����v��l�o�G�>���ެ �]���Q�sR�S{�}���fjH(9R7]��a����~�����H^����S�\�]Ғj��uv`�{U�zm��-즁��țaR�$����Z��%P���z���� ۶h��h�nhF�
|F8'���(���? �� 6��}�ʛ�\l�=���0���X�6��0��[�mlm�e�A��6�'h�r�nـko 6����0��b�%��/�6�rm����{�� }�� �x��/B���\ǂf�H���������x�l���Aa$`�@� H��e`I42��5E!(��GO���1����4�hزd��&���Ͼ�������Y� n����䛢�UV����oС'Ϗ����M��h���u0Ɯ�$I.�jyp,p��]GK�������zKw5IL�A�Q)�"S������*��[�rJ!~���ŀ4�ʪ��%P\���͖�-��B��u�wwb�5�1g�"&F�,&n�*�Ȫɫ������`�1`[u�~���s2+�r"�\ݘ	Oww�w>0ܓ����M# �B!ƨ� ,P�����BB�(Ud`���E'�w�=�ɹ'���S�R�f�j�� ޫf�J=���� ����[n��Į7SYFd\[>��G����m�A���#۬�GW<9�7
��"� N,xщ��$4
��@��f �x�/���0�̇WE��R$@q����-�s@��Jh6�=	(�%T��U737E�4UZ��� ���X�V��np{l�>t�`�H/�j`����}s|h��Z��`y(����`>���t�������Uf ����B^K�߼|��Ł<��^��<jF|��)) �!@hq���.��~��l���(^9:[�C�@Y,<x���`�,Kٵ�
�����6���Ls�'���3��Yx�VN�k�9�y��<�nڽ�-�ͬx�[f=�������KmN����KcC;[\wBt�"ۦv�vL2��ԁ)��=���2�vnы���`���l�q�>z9�i�{\��T�fU�f���Q+�u�u4]j�L�j��3�z<:4Ma�^e��Д�� ����9�q��v5�Dx)�V�Gq�sk�IK�4q�ݺ707:����x�z��_�9�t����#"Ȃ#D�4�w7��H�j��9�t��\�djE˩L�uT�D��3@��<h�ՠv�ՠ^۹�~΃�X$��$Y!�^�L]k��x�9D�k8�>�����&!" ӆ���V�{n��ܔ�/l���T�M�"R)�C22�Usۮ�m��r��q�6��q#�4L��NO۷�}n�I)���̒8���nh��M��h��h�����bM)�ѹ'��kٿ�	)�0K�ĕDV�~2�[0�78�x��(�2\���g�'Q"}��@�}s�ko�2ـn�A��J�HW"���5ֹ�5�f�2ف�/W{߼`\���d���.E1sv`ݳ 򈄡F�3��>�� ��ـr��{���7����{e��-˯,9���^J�(�����y��6'9�P��:������x�4Wf�������0��ė��O>�?y`�ƒ������c3�d���>�� ��-��ِt�d����~��;m�ӿ}��%�5�XCm�[e�Pd���V��I�	Il�iŀ��U�TcH�!e%�s��i�o�Ĕ�%r!qVښwĻ9���. ��J�$I1"B$eeŸL�7�����r�P��h�,SY��F�Af��!��ٌ��;�c�[���y����rZ�5�����l���@ٶP!e0��w��F�%����h��L˙���#.�.�F0�?$�0!%e.��b��?Bf�Xse�Ma!1�̵(T�J#��� ���0t�R���ٌa�:��T,�b�)Lk�(9)@6U�%Ӕ%QXT��r%�P�gHm7���!��h��bm�4��U8$��T0@Oʋ���/��(�
<V�UO ھ�?�#�	�J*@�|�S/�~nـk���(�ō���}�~����v�M�l��κ;�HmH$����[0(�%������ko3@��v��j$0DQ�cDQ�a�+F�[/��E"X���7:�^��x_WGe)��m��?v�h��{������[}��,��Ȍdn����DDL���`��0nٞIL�;��"$F��C@���4sj�;l���YM�2�x$���q0UV�:!N��� }����ف��$!		Y�"B$P"�p`*T�'�q��^+��d�Ga"����ye4[w4^�舏�qU_���VZ���&��/8�s�ǵ[��Tx_kL���K��Nmx����6���Te2XQ5g�w��`6�`�[0�)��U��#6�8�4[w3�B�5|`��k�fy(�����5�q&��73@��O{e4��	)��|`�ذZ�MTS.B��uu*���]�Xs�0m���^ID*��~�ww��lR��Ȩ.���ـy$����sW��������ڬZ4jE�eH�ULR'�A��$��Na/�jD�l����uk���	
�D�s%����콒xC�Ʉn6�s�
J���gQ��E��C&�ɱӯC\d��}EsY�kd�r��$���..�^�ۡ=������u����vqo"��]�5���B�i��ZȎp!��t�/X�g��e���&�����sm�N�k&&�ܐ��.�jѱ�M3Ʋѹ�����[����{���fv��e�\M��N��g�v�nO'=;]�r\t�79-؆�#�n3	[q�����.�-˕�B�~m��߰��l�6u����|`�Msđ�M|�`���[ܔ�:��@�m��x��%С(�5pWzQ3T)�RXUʻ0=�V ��0�BJg_vf��\�4ˉw�LBDӓCВ�=�8�5�b��l����ꪳ""#6�8�4v�����B��~��w�x{l�����-V���]a�Ξݗ^�3`Z�j��̮[HPޢ���A����S��� n�xn��J���X��)�����躺��pu��Ј�T�!��"Hd��L�$�	�Y����i"a6�� ��$Y �ROP�b���L� ?����y7$���f�k����ḡ�$0�x��@m�0�x��P�{��8 �u����jE6M�Ir)W3v`zD�w~Xu>' 7[�BS��� ԉ��3":���
���7Z��<�!N���w_;n�w����Bl�8�
D�I{1����r���c3�t����\�;W��]�s��vf%���o�4l���۹�gߐ{��ZR���<�b &���S@�m��-}��vپ�H����Y��2E!�v�ۚk�sX�D`�?*QB(&�<v���h��ư� Ě�8�htK�|N k��l��BS����|�&g�@�̎6���hϾ���?��� �k' ��y"�]i��0]�ݍ��c���y�0�qv��^KF��N��&8���϶=�Q,�#��p{�� ��f �k' 7[���Ի��	"R-���ďy�@��l�(S#R&��̇MLM�UZ�;��8��xyD�wv,_v-�t�M�!���h;l�o����k��ARB�PLĈ��OãZ&�c �)$JZQ!ia�K&7��c1HW
Q�=�+ �ze��Wv��,&����ŀy-}ߗ�;��8��x�(P��:�K�- ���,���v� ��x:�.t�\;�9�Y�s�ֲa�;�������L���o�����@9�g�������4_���D�I��� ޲��n�m��>�l͈����^m4chc���M����vt�={M����qADF�h��h��;{M� �m��޶�b"�DB�'3@�l����b����5�� ��!A�A�J�~c�����U�U�Q��GY7:������v�m��終�t��l�z�v�S�,�[<�6Zݵln\"�'�y�;�7m�j��k��x;�������;bP�ŏ05��.Y譍˛����L�G{a�v��(�b�k\lY��y�g"v��m�Zq�'�wBVӅ}6���Z���M��[5�Ȧ�4ѓ�ij�M-,M!��ww�;���ǈ�B�H���t}�S��U%�ݤ|]�c�<љ1ֶ��F�wm�/�,��8oi���@�s@岚��X�ك 8�3@;�o ��,���f,�2};2���H�H����/�����i��74��h婬��I�̐���Т���� }�b��� �����;Ȝa�50rC@��74��5�� ;f�[FT�J��a�33��G^<s��۶�nsŵ��湹��\�uR���s;�K]��o���M�����h�nh�n����q�����߾��3��	���B������, {��ӻUMP�6D,�9���-�74���#�����X�Dӥ3!.�.h*��Dz+��, �{׀6�,��`���H�ك 8�3@-�h�g�{����=�{ �nq`���o���=@�nڠ��;k�#���̽� j�C�ێ���[��s����N4�bKv?$������w4�V�[l��SY1B&��2'3@�����H�}幠��4m��9]�Ț�bML$q`�� 6��G� -�(JDIA |�D`A"Ȕ�XH�y|D�v�KhЀb�/}�߱`_�`�j�9�WFI��k�-�s@����չ�w��##��-�s@�G����|��8�:�`|�t�����m�l<=c&��KA=ю9��&2��R�ccm�.��V�Jh� ����x��s� s��DG���X�.�3!=D4Uk 78�Т&C�u��ذ���P�S'ɇ_)�J�,(��XϺ��Ň���ݙ�{����?.����Fb�LI94�ŀ=o �nq`JJ�*i"�
D5�w��䓾w�.�u5�Mcs&D�h��h��� ��h۹�uw��4��œ<����3k�ev��Ci���FUQ���e�tIL�͉���	��G3@��nh{l�-�s�gߐw���[��fy�A�3 �o �x���X��ŝ�N���D����������4v�Xz�ot��5�b�?N��4
UE+�ULլ�}ߖ��8���X
<�W��|��^^�3!>��&��`����,��`6�`�R���uwhuY�a�gǡwX&n�%8��X�M�3f(�h���e)B/�xvf�l*2��E0��u�~�ʼ=@H㗚��~ё�	�S�j�B��̼ڳ[I�%�tBqY�~��^p9OP���2me�]i����4�5�0x��IsE0�&��%��	,(�
�`Ga�����/G D�)b�b��lB��6@rݗw�9V�
󯼏���C���j�4m�]� ���.�T���rۻ�S�yE��'�(��S�C� ~�� �z�w�~���Z��`�D�Bz@�{����i�I�ܞ���!���p@�D/�X���d�RL�&���@'q���!s�m8�H\(v[��va�븲��E�u�Z6�X�۰��;I�=tø6��v�H���k��}�c�=�jI��Zy.�i\�v{:7;�slj�dWX9��;��&�W�p�BKn��V��{"��獛��t�������=����mb9�کQS�^�-�oR�\�[f���;��Q���hwY���hl�͔�G*�7��F0��m�D��n��;C���] ��pl�Pe�iU;B�j��E�rgGJ���%;���	��ZՎ��n�Pc�
yj݃S)q�v;�ը��j;y#�ɵ�&����w`����5�.ڷ
��q�Y�[s�\Y���v��5gR%v�[�jvq'��n6�6����%q����ͤE�弛����U�-Ȓ�%׊���^������`p��'N��r��됳��\̛X97v�m�bz��j[����nɓW�y5m狰�����.����m�[�z�y:�ʗ�݂���ɝ������ú���q�m��/6d\�OBO<��	�;m1�<9{[��:�@��Y��qڰt�c��k�e��um�(F%��V×T�K��Й:i�Z�VI�u�g���s�WdɹK"fm���V��ʴ�ۊ�DuU�m*�A��0khq�&[�ӍeW��R���ǭ\�ҏ&`��lB��]P����-8��ppԤm��:I�' \�mǬ��yݧsZ������v�����^�[)�	�{x��f�ǐ�V�ם�P���Tl�bԅ��1�]�+���2�jH�t!qj�a�<248�+�rLʯ$U��^��A�11�9��;ܒU��on�������d���n�@`68+��Լᖆ�Yr�bR�GjPu��8�B�<�A]�-�tLn� �-T�^�,�L��gw�� u�j{�n�U/�[Kp���T�T�v��g��ђ�i��K�TƗi�0-CI���!:5�3Z�u����Q6��W�^�"zA�.�=Aȁ�Z�ت1���$=q@1T�z��^ 4螀M�j_��3�7��Zs�$b\��P�n˜�rƸy��R֠u��mt��l�x��Nc �֭��H�ܷA�;�����,j�M�$��h��#�Lt��G^M��ԉ4�s<Ս��sW\�u�	y�r��[�9ۣ��!!O*��s�%:��R3NN������8��z�zܕ��cN�"<�����qT���sٙ�uA)�"�r���{����wwz>._��Ʒj�=��n��㱱AΡ�`�.箜��Դs�K���]�ɭ�%����`�� ��.Q�C��q`�_C$2Fb�O��4m��;m��/-[�m��yjj`�#Mcs"��X��`�����ذ��X�ʝ�E�	��73@��nh��h۹�w��h{SLEC�+�*���o�	%���~_v,�չ�{>��ܗ�8�I|�H�Ll�"N�ڷn�b��6�l��a^��q�sF'��}H1\�ItȊ&���{��,�o �nqz��Hk�ŀ}.e� T��(Ք�sF䟼�ݛ �pT�
*"�u�q`�x����B��5Չ$�0M��=�幠s��h��h���?g:��|�1�h����^�XͼX��,�z�, ��w��������r�F��by���ӑ,K��#��}��~�bX�'}�׆ӑ,K�����ӑ,K���]��/h��onu]"r6�ջ'��nu�E�4k�q)�1�����w���杢��y��tm?D�,K߾��ӑ,K���{xm9ı,O}�xl>TI�&D�,O~��ND�,K����Ʀk.�Knf��f��"X�%�����r%�bX�����r%�bX�w���Kı<�{�iȋbX�%�rY�2I��kZ���iȖ%�b{�{�iȖ%�by���ӑ,b� | ����J�["�1�D*B+�qg"n'���ND�,H����4�kDh���}�oK�Q�75a2]kFӑ,K>Q`dO~���ӑ,K�����Kı=���ND�,��9����ӑ,K��;e���5����sFӑ,K����"X�%���p�r%�bX�����r%�bX�����Kı;���q��M���pRՕ�z��nH\6"�ػ�8�a^pцV�V�>���������ѩ33Fӑ,K���p�r%�bX�����r%�bX�w���Kı<����Kı?�f��\�e2�KsWSFӑ,K�����Ӑ�@�DȖ'�}��"X�%��~��ӑ,K���{8m9ı,K��N�5Ma�d)f��Ѵ�Kı<�{�iȖ%�by�{�iȖ?2&D�{���Kı=��p�r%�bX��~�.黗n��U��՘�h��4{���ӑ,K���{8m9ı,O=�xm9İ:/�D !������h��4~���~�]Ժq�3D�f��"X�%���p�r%�bX�{���r%�bX�w���Kı<����Kı?xk�sY5���snσF곷<q��&�n���"Ø)�1�r����	L��;fwT���w�{��ı<����Kı<�{�iȖ%�by���ӑ,K���{8m9�F����=��ۗM��v�ݘ�h�,K���6��Ȥr&D�=��m9ı,N��NND�,K�{�ND�r�D�<��~>�\f�SVS.h�r%�bX����6��bX�'����iȖ?+��;߾��Kı=��m9ı,OL��p���3WRff��"X�%���p�r%�bX�����r%�bX�����Kı<�{�iȖ%�b~;�fY�nk3R�9ı,O}�xm9ı,>H���~6��X�%���}�iȖ%�bw����9ı,O� ������Y��ڒ��SD��{u��[�Y��+�nw]�;D��aX�-��8��S���SK��{d��r�8�GM�L�h�n�ء5�D��.��<u/.�>�m�r���\��p�c]�M�:299z1�P�J��Ӊ���~�����#�Ш-Ûv:�w`�V)���/;�e�J��3��vc+R�*�M�6U�'TPO��������oh�ѫ�xH��E�8����N�j�����F`�%�v�6�a��[���q�%w�����{��'�}�ND�,K���6��bX�'{�{.ӑ,K�����ӑ,KĿ���MfMd0��F\Ѵ�Kı<�{�iȖ%�bw����9ı,O}�xm9ı,N����O���2%��tO��CZ���S.���ND�,K�ߥ�r%�bX�{���r%�bX��{�iȖ%�by���ӑ,K������$�d.�n�.ӑ,K�����ӑ,K��{�ND�,K���6��bX�'{�{&#Z#Dh�����r;r�q�ܻѴ�Kı;���ӑ,K����"X�%����˴�Kı=����Kı>U<��$̿X]h��Y��U�3r�����9.:Sڇ,�v��f��0��>ӎ� ���[�oq������Kı;�{�v��bX�'���6��bX�'{���r%�bX��N�)odf����ND�,K�׽�i�pH�?	�Y��A�$�B�H�<QL�)��O�,N�~p�r%�bX�w���r%�bX�w���Kı<;:o��\e�f����K��Kı=����Kı;�{�iȖ?��=��m9ı,O���K��Kı/�%���.��[%�r�Fӑ,K��}��"X�%��{�ND�,K��{.ӑ,K�����ӑ,KĿ���MfM0��Y34m9ı,O;���r%�bX��]�ND�,K�{�ND�,K���6��bX�'����Yu���2]P�S�{]��ȹP�ջ=Z�7j.V�g�M�.�z18��kں�{�'��u����{.ӑ,K�����ӑ,K�����ӑ,K����"X�%��;wr�ِ�5��%�ԻND�,K�{�ND�,K���ND�,K���6��bX�'��{.ӑ,J�=�߇��v��n��wf#Z#E�b{�{�iȖ%�by���ӑ,`GK� �� �x�S"(�Q|Eb��ȞD�����9ı,O���6��bX�'���ӳ%�d�V\��6��bX�'��y��Kı;�w��9ı,O}�xm9ı,N����r%�bX��N�);��WRff���bX�'s��ͧ"X�%����"X�%����ND�,K����r%�bX��;�sk2
3���6Y�]�f�.�*m�r� :���;�����mݳ�Pa�2kM�����%�bw�}�iȖ%�bw���ӑ,K���6��bX�'s��ͧ"X�%�y��R��e�Y�.�m9ı,N����r�$��{�&��	���fБI�=�I���bX��{{��Lɣ&Z�33Fӑ,K���6��bX�'s��ͧ"X�%����"X�%����ND�,K������d2�D��m9ĳ�Aȟkﾙ��Kı;߾��Kı;�{�iȖ%��b	 	���.��ͧ"X�%�ｳyے�V�C4I��ͧ"X�%����"X�%����ND�,K��}�ND�,K��{siȖ%�b|?|N�����%�2d[�����p��z�6;sn�a\�FM`�X���c�ЉAF> ���g"X�%�����ӑ,K���fӑ,K��{���|"��L�bX���p�r%�bX�gl�C.e��j˫��iȖ%�by��iȖ%�bw=�nm9ı,O}�xm9ı,N����r	bX�'�C��-'fV��L�jm9ı,N��ͧ"X�%����"X�%����ND�,K��}�ND�,Kó���mƗ$Է-֮m9ı,O}�xm9ı,N����r%�bX�w���r%�`6's���ӑ,KĿ��s�պ3Y),ӗZ6��bX�'{�xm9ı,O;��m9ı,K�{��ӑ,K�����ӑ,K��z@��nf'�̧\��`.�#l�����ݖ������e��.�{`{��"V�JDL�y3(Y1Չ��\���v��X�ݎˋ�xwH֜��p��zc�����F���.��ny�B�fm������}��:8N;lʽ��Sg<t��:y^9���x���։vm��4�F��@�JXv}�vn.f�5��
��:v׫�f�hsZW����{����s�/���홎kaxӫ�Kۣiޗ���"�WY^n72����n��u�.��j�+w�������{�N����ND�,K���5��Kı=����(D?DȖ%�����ӑ,K���>�������S.��kSiȖ%�b_;�涜�bX�'���6��bX�'{�xm9ı,O;��m9�ʙ��y3�.VjC4��[ND�,K���ND�,K���6��c�\��=���6��bX�$��������$-o��\͓6��5.��iȖ%�bw���ӑ,K���fӑ,Kľw��m9ı,O}�xm9ı,O��/N�.e�����fh�r%�bX�w���r%�bX!|�{��r%�bX�����r%�bX����Kı?w��\֝d�&��5Kqk��v�s��Ϩ�m$�^z����0�GSV��3	Hk#uu&f�6��bX�%��kiȖ%�b{�{�iȖ%�bw���ӑ,K���fӑ,K4x��2�G*�#�������5�4H�'���6���`��P$E#`����@`A�C��A�?D�9����Kı<���r%�bX��{��ӑ>G*dK��>ύ[4f��٧.�m9ı,N���6��bX�'���6��bX�%��{��r%�bX�����r%�bX��;���.M0��ї4m9ĳ�E�)�=��}6��bX�%�}��r%�bX�����r%�bX�����Kı;��驚���S.��kSiȖ%�b_�����"X�%����"X�%��{�ND�,K��}�ND�,K�_~�̿S35bϚxIu�8�kJ��&wffM�p�Ϧ�ۅ�]����f�Ay��u�ʃwV�����ı,N��m9ı,O}�xm9ı,O;��m9ı,K���5��Dh���}��n�%��Nܻ��,K����"X�%��{�ͧ"X�%�{�s[ND�,K�{�NAı,O��oN���f�j�5sFӑ,K����"X�%�w��m9�!�����2h��w�t:�H#V����pe!���ؐ#I D�$K��b�%�# ��c�fP^*�oTwP9D,h���AD���LX�#��?_ĥkf��"���ә��f�@1E�a	xJ��l�J�-�Ą�	f���d��C��%%3A.kN����RᏌ 3�����!�0��T8R�eB���ue��).3Z4h�fK����Jť���!����;�hF���ZB��u-�6ͥ
CBF��u��sDH��N(��(z)�SJ'�?�F#Px"EX��=�����?�� ����& <N(��M���ND�,K���ND�,K�!�ܒ������34m9ı,K��{��r%�bX�����r%�bX�w���K����6��bX�#�?���J�Q)�n;���kDh�'���6��bX�'��xm9ı,O;���r%�bX����5��K�7�������:О�lA<�ɹ�x�Cq�L���w'��������ɬ��ٹf�����ı,O{��6��bX�'��xm9ı,K��{��|$�L�bX���p�r%�bX�����D�&��MjjL�ND�,K���6����"dK��~�m9ı,N��m9ı,O=�xm9ı,N���W�ܺ�ʅB�wVb5�4F��;��5��Kı=����Kı<����Kı<�{�iȖ%�byޗy3�܄���7Y���"X�|$�����iȖ%�b{߾��Kı<�{�iȖ%��x),i�#>�$ĂA�Q1`o�7���ӑ,K��߻'5l���i��ZѴ�Kı<����Kİ���}��i�%�bX��{��ӑ,K�����ӑ,K���wٚ��t=Gn�����Yu���]Ot�sm��])���l��: ��7=�n��"X�%��{�ND�,K�罺�r%�bX�����r%�bX�w���Kı=2��)K�B��L�Ѵ�Kı/�{ۭ�!���,N��m9ı,O~��ND�,K�{�ND�US*dK��t�I�.I�u���ӑ,K�����Kı<�{�iȖ?$2&D�~��ӑ,KĽ��]m9ı,K���:M\̺3f��Ѵ�Kı;�{�iȖ%�by�{�iȖ%�b^��n���bX�'���6��bX�%������)��˧*�F�F��=���m9ı,>c�{��[O�,K���}�iȖ%�b{���ӑ,K��>�@6�$0��D�XE�;;���],�6�{uY���4 7bP��mȁƵ1�7��?N���{H��r����*.ҏ�[Y�-�.����U
q���뤊�NL��c�n������5aq3��Â��Y=�;���,YsI���[!^6�cn6^�Ցbn�Y��sMu��竷�\/6ʯ^ GZez�6`��5ɳ�&.6Kk0�������L���,3����>����{��9�}/l����\�ܙ���{dR�5��l䶡�h�]�GJ�9����׵�M���v%�bX��{�kiȖ%�by�{�iȖ%�b{���ӑ,K�����ӑ,K��ޗw-���і�Zͧ"X�%����"X�%��{�ND�,K�{�ND�,K�묅��$)!I	�ȩ���mH\.��iȖ%�b{���ӑ,K�����ӑ,K����fӑ,K�����ӑ,K������.d�5�j˖捧"X� dO{�ߍ�"X�%��u��ͧ"X�%��{�ND�,K���6��bX�'�yON�J[4X]k%�Ѵ�Kı=�]�fӑ,K����"X�%����6��bX�'���6��bX�%���̝ɩm�:��Οkm��J`㱥���,nMn������u��:�r���5�������x�,O;���r%�bX��{�iȖ%�b{�{�a��"X�'���6��bX�%���>Թnf��٦f�m9ı,N����"� d|ڨzy�,L�{�iȖ%�bw�{�ͧ"X�%��{�ND�,K���rh��hɄ��sFӑ,K�����"X�%��5��m9��dL�߾��ӑ,K�����Kı;���j]dӔ�h�ֵ6��bY�@ȟ{����r%�bX���m9ı,N����Kı=�wٴ�Kı;�K���1�E�&]k3iȖ%�b{���ӑ,K��{�ND�,K��}�ND�,K�k���kDh����򫪹#�Dwe�sDgfu�V{D\��;��S"���F7
��sF%/L�&�.�&���֍�"X�%��{�ND�,K��}�ND�,K�5��l>I�&D�,N���6��bX�'�����\�&k$՗-�ND�,K��}�NC�D#�2%��u�ٛND�,K�}��"X�%��{�ND�Tʙ���i��Id��[�d��ND�,K���6��bX�'��xm9���$HHD�A��� @���I�lX��T
DGf�r'�}�ND�,K����"X�%���7��KL�,���k3iȖ%�*��߾���Kı>��m9ı,O{���r%�bX��]�fӑ,K��y��2�����L�h�r%�bX��{�iȖ%�b����ӑ,K���s6��bX�'��xm9ı,O���t�'�֪㦓��ȃ�����p0�y�F�.��.�g7Mnp�:�\�i�w�?D�,K�}��"X�%��5��m9ı,O{���r%�bX��{�iȖ%�bw�;��R�&��SDֵ���Kı;��ͧ!�"dK�}��"X�%���}�iȖ%�b{��iȟ
�TȖ'�����,���,�2�Y�ND�,K�}��"X�%����6��c���;���m9ı,O���fm9ı,O=��s&j��d�55�Ѵ�Kϕ��>��ND�,K�}��"X�%��5��m9İ<ê� �5p�A�X,h��%Bd�� q�&)4��`���~�'s�p�r%�bX���o�as$���VY�4m9ı,O{���r%�bX��]�fӑ,K�����"X�%����6��bX�'}��ܲ���-�˫;c�Nt�m\�&���V���[�Ĺ|��ia�b.��v�+�r�.��U��h��4��}�fӑ,K�����"X�%��{�ND�,K���6��bX���3�(�HU:��ʻ��kDh�'��xm9ı,O;���r%�bX�����Kı=�^�3iȖ%�b~��e뙚3f�K�Ѵ�Kı<�{�iȖ%�b{���ӑ,�$2&D��ٛND�,K�}��"F��'ޟ�S��n�:��J��,K�����"X�%�����ND�,K�{�ND�,�dO~���ӑ,K���>ϵ5.�VL���f��"X�%�����ND�,K���}��~�bX�'�}��"X�%��{�ND�,K�=��C�����{�|���䈅��8Z�(k��9��c�W.˷d��2<��X$](�&��385p4�a.�ᵜ�۝n*����8,��oFs=β���a���r�r�f�����5��m�P�2F������Z�X�,X�H���vL�[��N��+GN��Z��v��nu�jw8�C<يuə8W<�]�ppD�n���k�	�=A���{���o��wL,:�cF�Y�۰6׬Xk���uK�GU�	Q�m�N����k�vu���{ı,O��8m9ı,O;���r%�bX�w���"�O�2%�bw�w�ͧ"X�%��{��5���f�&����r%�bX�w���>9"X�}��6��bX�'}�׆ӑ,K���wٴ�Kı?gm�;�$�a5%&f��"X�%�����"X�%���p�r%�bX����6��bX�'{��6��bX�'{���f�Me�)u�33Fӑ,K��{��iȖ%�b{���r%�bX����r%�bX�����r%�bX�æ��i�2�Mk2h�r%�bX����6��bX�'{��6��bX�'��}�ND�,K��g�"X�%��������7��[v���0Sx}s�y��ۊ"7x�	f��弪K����^V���Z+|��bX�'{��6��bX�'���6��bX�'{��ND�,K�}�f#Z#Dh��O��cr��(ueӫ���Kı?w���r?D^ wq,N����r%�bX����r%�bX����r'�TȖ'���>�Ժ�Xe2�&��M�"X�%���}9��Kı=���m9ı,N���m9ı,O���6��bX�'w��]�*h,�������$&��fӑ,K��}�fӑ,K����iȖ%���L���}?m9ı,O{ߎY��nj�j\�M�"X�%����ͧ"X�%����fӑ,K��{�ͧ"X�%���iȖ%��{��w�����/]u�ٱU�g[��9�ד���|��� �9˖v]I:��I�;�֨
�E��WfB��$)!I}��	bX�'{��m9ı,O}�}�!�$N���7�N�'gL��5�ܥ�d�֦ĐI�}�i7�,K�}�fӑ,K��}�fӑ,K����i��bX��ɼ'r�fL�SZ̚�r%�bX����6��bX�'{��6��c�y��H��S�qt����M���m9ı,N��g�"X�%���ݳ:�ѫ�,ѩ��M�"X�%����ͧ"X�%����fӑ,K��{��iȖ%��ȝ�y��r%�bX��ߧƤ.��LѬ��M�"X�%����fӑ,K��X���O���Kı;����Kı;�wٴ�Kı/�'{%�t�nL��r�����*n�]��9��n�W��=C�ѣ�������j�6��bX�'{��ND�,K�}�fӑ,K��}�fӑ,K����iȖ%�bwΗ}ְ�	�MZ�Ѵ�Kı=���m9lK��}�fӑ,K����iȖ%�bw����O�L��,O�ߎ��ї5a5.f�ӑ,K������Kı?w���r%�bX��{8m9ı,O}�}�ND�,K�N���\�&k$ՖfkSiȖ%�X����m9ı,N���6��bX�'���ͧ"X�ƕ�B	
D!�_¾ ��s�O��>�ND�,K��Ӧ]fE���fL�jm9ı,N���6��bX�'���ͧ"X�%����ͧ"X�%����fӑ,KĽ�_S��=���ku�6^�l���1�{q��5�=��k;��i���z�yv�.�iȖ%�b{���r%�bX����r%�bX����l>b��dK��ﾜ6��bX�'�v�d0��2�����r%�bX����r%�bX����m9ı,N���6��bX�'���ͧ"X�%�}��55��f�d�jm9ı,O���6��bX�'{��ND�K���wٴ�Kı;�wٴ�Kı;��Mj�f�&L���kSiȖ%�bw����Kı=�}�m9ı,N���m9ı,O���6��bX�'|�w٭a��$�5�MND�,K����ӑ,K��}�fӑ,K����iȖ%�bw����Kı?q��t��ș��c�I���n��w�+�$���l��] ��>:ˆ��!*��d���-����{�ӄ�^i��4���+���?���I6І������n���������`��d���a%�,R�6����?y�5��=�!w�7��n�bs�eS������Uݴ=Y\Ի�6�(l%�R���U+�	@��@��&6���Ywegw^	�3�~�"	@c��_|�Qm�n猬���4X;�4L#��V8[��1�\U�r晚#R���q%Ĕ)E��ŭ�y:W�l��p��!"R�^-���1m����ם�n�B���#�O��=��0����P�Nx�0��Xa=�{�,���4ȷ`&�jő���k�j���������b�� �ȧ~?_UP宭�y�@�bϖx����li����۩�x��M���v��=��V��3�����\��[wn����s)�9Mb�qÏj�m�ڠ�ZL/;[k�nܭRP�nL��n����k��g���d�w�i�m$MeBӨ��|���ׄ���g�\��.���ɸ׎����k��S�[�;n�Ǝ�����	�v��/]�:�ml��d��m�e�liUw��|㞐L����i�+��v���`�eR�ؙ3V� �(��`]�J�;�#��r�Ѷ��l�'+�3�"E$��qM��Yyj����i8r�,�-̼���3��\���&9}tq�A��E�y�R���u�7n�m��KF��l#�����nM�u���[.^6.ֺ��k��g�.8�)GF��3���0q1���ί,�@�ۻ�2�\�nϴK���/�<�[C�;��sc=`K���J��.N3zMs
���GWP�����>��2�!�lR��ΛN$&����V���O�;v��gˮd�n�8�$jݗ�v�=��ZE�%V�s�e8�4�@��!;���8YvN+["�M�m�eZ��v1s�^i���UVv�#_4�kL,2��V�1���^U����^j����5Ukh`�%���ev��V2(	�5�EB�9tl���0һK��N�\�N�ԫM�ȁɩ쐧�#���Гk���M��l��s<���h�t�;ڼ��綟F4�{gq��e�&��.�m՚k�K��qa[�ێ!�6�w>.sv�rlF�#�H��,:6� ڶ��b�l�Ș�z��ܚ0	n9!���ۗ��S7i���8�۲����ۧW�sh'/�u�1�P�@1����5�z�s+KY�q�J�r�=�%Q� �X��	Ƨf]���v0�����t�Z�n2i��,�R�ݖ�U�F��'`��j�ֆ��I�6IW������-r�rQ*T\�ү6�����Z��ۧEnh���֍]j����T4�	^� z��GN����.D\�=H*��T��l���]�������󰺡���n����	��[�7g�k[�Z�:�Λ1cK؍����2~���}�P՞��T6z��'k��¯i�1z.҃�X����	���-�e�
y|��\�捃\]c�N��n�[�k�9�n���}�OX*V���ch)�r��������#4v�QR�� �z�V�9�>,���l�� Z����743[��=:�,ΪcBVW?�����ni�,��we���Ӫ���a�s[Ůԡ�v�lT!r2km���Eu���Y�	�.k?��Kı;��m9ı,O���6��bX�'{��ND�,K����ӑ,K�����{K�$�d����jm9ı,O���6��bX�'}�o�"X�%��{�siȖ%�bw��iȖ%�b_}����,�5�3,�jm9ı,O=��iȖ%�b{�����K�	��<���m9ı,O~�M�"X�%��ӷt��l�2MKs.�m9ı,Os��6��bX�'���ͧ"X�%��{�ͧ"X�%�����r%�bX����/\.�\�f�Lֵ�ND�,K�}�fӑ,K���fӑ,K���oxm9ı,Os��6��bX�{�w�߬my׶��uŃ*�j�ѕ-Ƃ�I��Ǯ�n70����vv�:�y��{\٭jm9ı,O;��m9ı,O=���ӑ,K��=�siȖ%�b��d/�)!I
H\�wYw3ur"��c��x�h��4{�O�b5���m@�@� �?�n%��sfӑ,K�����Kı<�wٴ�O���,O����kE�d&�4fj�Fӑ,K��w�iȖ%�b~���m9ı,O;��m9ı,O<�����4F�}��J��e�#�˃��m9ı,O���ͧ"X�%��{�ͧ"X�%�����r%�`|��ެ���$)!I	�����T�I�,�֦ӑ,K���fӑ,K���oxm9ı,Os��6��bI
H_7�d/�)!I
H_s�*����.��u��vM��R��864��k���:�v�n������L������ı<���ND�,K���ͧ"X�%���wٰ�V~��,K߾��iȖ%�bz�j���-�3$Բ�֍�"X�%��{��Ӑ��L�by����Kı=���6��bX�'�=���O���,O>��o�F�L�t�Y��Kı<�w��r%�bX�w���r%�x�_�_D�4�'"{�ϸm9ı,O��~ͧRB����,踛.�H�R]ً��_��ŀl�u�~ݶ`i7c��#5�	$4��w4������Ɓ�e4��F�X�H�i�]�6��m{Y\�Yiv�����6Q�ܕλ������&��&h]����M����t��yre�"hȌ�wX��ftB�5��|��Xӭ���X�C`(����4v�h�Sŀ}:�`�m����N�jf�#6���?w�w4�ڴ�즁��]���h`fI��8�x�o�ޚﻃ�μ�o$�����즁��M�{�s@��C�7�2�V8�ƹ�z8nu����:tm�uێ)�s:}2�M�狴����������7��ـ~�O��u�}:N�.&ˡR-T�v`�g$�S'ͮŀl�uh��M��nF�G�Ƀ����`O���$�^�� ��� ߪ �`�a0&)2L�8�k�;��h��?^���;˗r<�a�G�w���9�)�~�˹�qrנ|��!�����*�|K���v\c�xa�v��fCk`	��x�W�U��6
�`,�v���n$?��|�ɾѱ��˄�C=��U�9�n;S�ٺ��=s�Svێ�^�9p��}l8�=��gmi��j�ήX,�,2v�\�4;͍pdc���6��%�y���q�7(��y�7(4������[�*rm�Gg���u�6^�Q
�]����]�+���pJ���kP�%� 9nA�5����2�ެ.��;<ɰ�p�cm�5�E�I�$E���;�O�ܻ�-zy�M ��]�^Y!J�jn����g�P�M���0�otB��a��+�H�$�Wk ����7�`|�,���`��j���dl��mǠw���9�w4�SŁ��k{� �d�L����T�T���9�w4׹w4.Z����v������[7lݞ^�ɞIxGl�Ԙ�N=�9-�iM&�tt�gNsW2Κk����]�����즁�YM���u�L���&h\����[
".�۶`|����7��4J0Ȍ�#�;��h���}�%�\����y��K�U6�0�Q��w��=sۚ;^��vS@9�3��(�A�i���]��DB�������?|����T��g�]�]�{[m�bN�n�Cδ�k��Gc�� ���s	t݋�콇kz��O�� ߶ـ~��9G���ŀ}��ذ�bQD�7#�;��h�e4�Sŀ};��Mne\M��T�T�����f��x�Ա	!APB>���Htx�����k�~��;����r528��L�`��� �u��7�`rJ�}�h���`�L	�L�4.���;e4׹w4wo�9�>3g����1qv��Gd���d��P�{��^;nh#Q)#@D��ȰR=�즁��f��x�(K��� ݙ�D�F6�
7!�s�S}�}�$s�=��u_y��e4��]��i(dc��R�ܻ�mzy�M������2ۙ5,�ѹ:���3��0���>�l�j�B�@u@�T�(OD����Gxh�a~���$��,qǠw���9�ـ~z�,��� 腵��u�RXU��q!F�^���wvݸ+<�,^�ݡ�%k�p��(�1��Ġb�Fc�c�$?���@�-����������r519�k&Hh幹�qvנr�S@�]�:"�򛞺��H���V�}ذ��0��0��� ߵѸ"�ɋ�4^�h��7��,��u�~X�C��骕4"���9�)�w����۹�r�Sd�4������ 
����o�뿼����Km\����$c#kYdl�����#-���Wh��3��pS���\��.W6�9<fy�V��7\=�!����s�4��׎�ۨ�]�Ѽ�=6z�^ȑ������̓���qۗ���N��t� i8�[XI�cavKʻ�������Q�` 磸�4��9���;�2&^r�e���JSZ�ӛ��M-lPN"5jɫ=������w�%��,�p��B\�r:��V۲Ykk'Hq��E���~�}"fr����Ü�]s�H�#$19
����;n���M���>�5~w&6�l�jL��s��`=�`k�`�k�\ɰ�"ВNE�9�/e4v�h幹�s��hv�21��;c0��� �[Ł�y�� �K��&' �L��/-��������{e4��;Y���Hj��v�';�m� 3*6�/=������Q�m�\�bq���a0&
L��[2�rt�}޲�~�x�}��+w��e���ܓ�<׳~���ā� �C�Wh���U@����nI�����n����y�Y�X�E��C@��Ɓynnh��h���*�\VFǂ�H<br幹�q�� {��R�g�*���j�fi�MI�4[w4��h��/-����M��KN5l��H���{n���x��*�F�ln�����juv�nr�n��v1$�.�`vـn�f �mb�>m���U���x@h�{e4�ss@�s@�즁k�ؙ1<�T�E]ـ?�X��x��Z�E��w�'�o�A!qqCAX�C��{��~��l��]�2�yW��T �@`B��
���Ȅs7���$�c4k|�Q��'����)�)�\�����x��$*I��!x)o0�
)ٰ�%eq�%������5
L��V3�_f�e�*��9�A�Irk�40�����334�A��vm |2TV<߾K���[L������MY�!P�U�3�AS��_��2b}t�3�j�:M��� B@��?%,z	�A��s1Qp �C�~ǈ�P�hE�+��B�u��j*FS�L	��5)��e��mڞ7N�� 6 bŰ�Jv�4�_z�w���V(`l���	����X4 U��i��n0���!I_���dX���XQ5���M%��D��04���'���+��s�Z��
@��z"i`��m@����t ���
��'��h�*�T�Wb���}��3�\��/�@���px6`H�&nլS���`��n�s��!BS�ܿ,��DخA\��]]���0��8��� ��ŀ~�Բ��Sd\̌c�鍹ݗ�Ǯ�,�*�(��M�뚹�[5�<�.�]���k}�v�� �mb�?6�r�����t��/H��P��QŠ^[����h���-v��$w�c^��#I�WV�`��`� �M� ޵� �m���(�nD����ht���X�%$�\�&�D:�
����|�A���B��S�(P�?gj��z�ҥV+��aSsv`���X�m���ـr��??7���H�;l>m��z�۱��L�,M��Hג/@��ֲa�G4:��ru�����ŀko �vΈJ���-ݸ����ɚm���!L��|`��p��,w^"�2 Ɉ�H�h�S@�v��74�w4ե�u6,l"�"�����gk� ��,����qYk�xĤ4����;mŀ?�ـkv�҈�(�St�t��l��m��NJٮ-��E�������..Jqp\bT�`�X�<�����l�I�r�/%�@B	m�%t��G 5�A�} 1I����b�[�8�J��N:�r�q���Q���BE�q��YP9�,���;Hy��<�J�\���y:��ڛ�֜����7h�\�օ۬=;g�DŅ�b���cG�����<
M���P\�*���{��w����ﰽk��p'�l:{c��u���B�ζ1k�����z��u���{��}Zrk	]w��?�����/;)�v�M�74q��TLX�m�s4��h�S@�ֱ`�ş�Q!�.��R��H����0�|`�k2�����^v�ɉ��cY0i�@��������m��/;��	���>�JL��v۹�^vS@�v��74^�2�LpX� 0mL�&�ꇷ���u�nM�*��S�H-��g�f����&"%#��^vS@�v��74�w4ե�u6,l"�	)!�v�V�D��b5�c �R	T�FW� ��t���޶l�;m��/;)�~W.+#C�F<b�-�74�w4��h�ՠw뎳,ƒA5&L�/{)�^�S@�v�����9�[i\L`�mȓ��{�M�ڴ�ss@�즁�3;K�q���8�8��Ȧjp�GegƸ5���� �J�"�n��,�n��(C�����y�nh���/{)�r�U��@�5��Z�i��^�S@�즁ye4�p�TR..�j��L��0�lã� BE�<��(z���@0�����r�ڍ��܉a�2#"�8h���/�@���h���?V�q�ر�ȰȈ�4�j�/;u�e4^�h�n����md�5cpO���f8��X0v����ܔ��� ̉cI�)#C�F6%!�w������/e4�j�9�q�e��BA4�F�{�M�����;��F�����q�M��p�9{)�^YM���h���qu�G�1�P)!�^YM���h��ܛ="� �
H*��*�,@���J��USϾ����w��F�<qƲ`ӆ��k�0�l�>{l��ـrP�}ߛ|���i�Q��xm'���y�Y�=�����)��nFMvU=s�{v���r~��0��0�rJ���M��� �D1H�4^�h�S@�;u�e7ٙ�G<Ҹ��Ǒa��4w�Ɓ�v�4��|���4��Ɓ���� � ؔ���v�4��h��/,��߻��,b�	�"4��h��/}<m�{�1�4� �AF��6@ĭ 0�tMM@W��%�u.��L��5�9�K�r㡝�.�8w���ˤ�:&v��k�Ō�&wV���ٝqۨ=���Cy9��r1�$965�pc$�ۇ�뫚�ܲ�1k�[��m��wZ�<��WKh8!�"m�8$!9���K��^'k*�M�n�l�kV�q^���ٗ� �K�禊�[uF
-vLֳ5�f�h�a�?QO@��������!��pp�\�O78Ӳ6;]�tm���cΗ�\=�����%Ա:r�;m̉8p����9��F�{�M �[Tx���r��9��F�{�M���+�Q��DĲ`ӆ��������9�)�^YM�u�"���|�Lr@�즁�YM��h\������"�E"p�9�)�^YM����/{)�g�{�|5	�0m�m
(8輗���ӝ�ڎOd�j�:2C�J��f�͔����E�#�����@�����h��8�C�x0�H6%$ܓ���o�mZW���	�<9( ��CT���zb(� �ɮ�[���=<h�S@���Y�
3O ��Ǡ^�S@�,��ye4.[�@�*��ۘLQ�������ye4.[�@�즀p�����Y15�rye4.[�@�즁�YM��[�rI�&2`L�!�D���;��S���>ݝ�֞��FˢJtᢵq�f�d������9{)�s�S@�,���:�`�a>j&71����9�)�w�S@������0�E�jK���0�;f�;fBd!PI'�%�`�Ӝ��?�'��׍�b�:�ĞF���;�)�qs����M�즁�Ά; �a�lJC@��n=����e4��0BIK�j���VM�U@Z.�J���g�[pYuq�\ձٱ����]SG ��h�k�1)�I����Y�@�즁�YM�ۋ@�*S.6�%��4�^�S@�,��x�Šr�S@8p��Q(	�C@�,��x�Šr�S@�즁κU�&D�5�5f$�����`��=�f����#/�P��)k-��\%"�HU���0�s�Q!L��H;E�;���ܓ��֮�4�'�D� ���h���/,��W;G�r���"L1<��28�m5��Х��h�oJ�&up#���:�^�0����`LDR'�z��@���\��3? ��Ɓ�2��)�@�m��ڴ
�h���h���8�C�`<�H6(��*��/{)�^vS@�v��+�X��$�	�°:(�o8�;]�?�����89Te���D��sN�e4��o�����캒y�����EE_������ � ��TTU�QQW�
����TTU�ਨ���T_��(� `��R��"�",���B��,H",X�,��"�b��R��B(�`��X�,B� ����"�",�"Ƞ���"���*� �A`��b�
���QQW�QQW�����h����TTU����������EEE_�***�QQQW𨨫���e5�k(8 ?����?���u������PJ  �e�	(��%(P$�� �� s�   9IR�	T�"(
�
H�J(�U
$P)Q�I�    `j�@ X��v��ӻ��p�_}�^��l�;o�ч���<����+����Ys9w6��q׼�:���>�9��7&�Ƌ�x� P (^�9Cm�J�����_jݲ����{�+���}��m}���|�������+O9��8 :3����hݽv:9�����zx�����c��.wB��((P  X����ݻ�G]ϸ��s��e
�6އ��=�w���{�=^����w� {��u�w>���/��v{�w�{��p*�糧T�>F]}�zx �(�   ��C��3�2=��`���W�|�{=�;�um�;��k���c�ݏ[�{�� ��C]�;������v��A�p    ؠp[t:5z�����޽H���"��Х���̊;��Js���<��uUf�  I��ͫ�G��a�{tu����V�����Udx��ݎZ8@H��H�@*�MLT�!#���=G���i�@��@      �~=UD�JQ�      ��U*��R       ���aR�@      D�R�S�S	���h�44 ��b3�?���o����ҹ�9��	 ��C�DKT��O�'���PLV�����a��:"� `�)��b �)�+dU@E$]A��P���R�����6�϶�������_���_�t��ߙ�>�~u�0�2�&6�XB٩�e0oQ�&�SF�ވ��ۖTwgR��	�;��c��d0��	iP�.���ɖ���K�U]�!z�Q���%U�
���2t �HQc*����$��$�F���`�Z�kl.o,��a9t�@��!bJ,�H�����+�]��d�gR�1h2Qd$h�cQ�H3�2Eʲ5e!S���eo��k��i$��$���
b]��\�t�$H1# ���6ӡdm���\
"��5OP�(�"U�պ��Qnj�n�M�* D�� F%�\����Lq�B�0�Т�H�E�t��#	S�+�+z��"@�l� �n�6��bfà���uӗ�m��wW��D�xdi!Dh�-aQ ��+縷�0"��r0�Ș�<�T�P�"��"�]I��l�	�A�f��w2U��J���k	
���j�F�5DFdi��!D��J�]�ʫ�;��!�\e\��R;��4Io}aZu�np�7���H"�"F� �c���ogfa	p"G��=!o�7���}m���b�A�$� J#�ThbP��VZ�(#D(Ɣ- 5a(�����%� B-�ʅ����$!W�.��!�!�(���h�^�a�1�����`h��IR�8��c��H$!x�@�PUF���
�̂Q���������	�J�*R��RV��5zQF��a	
��h!u�Q��8��2��S�yB*�I"FB(�d�Nu���'vi�	\ܬ渐�F;.�Am�"R8�QN�ݰ�њ�Äh��D@dF�YWMT����t�)�P*-a&�oUh�0��F0�d����+X�3A$��U���Y
H�
H�� s��a��=۟r�#�ø{��"T�&�h0eQ�]S�ʻ��՛)nY2�6��I� �FU���t
��J��G]��B���$��B�Y��ZB�X�lܣ۱b@�Y
.j�:�Z�������dU"*Y�[wl��� �E�&
4�2�&3	6|��E-듐Pr���c.��4��d��Vl����n��T�쭲4-L�rA �2� ���]XGhmM���/
���e
vt T��L���QL*��Ԫ4]�Ql�V�U���K%F]\)�$aFD�s�ݚѭX��ab��.��D�͕�J��e�)��]�Q�z��$$ܗ'I6S�Hk�,���(%ȥ�*�:�T{7f�,&]�W����C*Mc����Q�v�\ ���*�Qi$��paD �J%@�ZE)#"4Aj4�!�(!KbB���� �"D(b���Y��00
v�� Q�6$,,�:3G H+�
egfu-ݖ���ˀ� �I�bq�\2cH�9��;���D���&2�9�]A��� �%:IMIb^P�L�!+ro2�������7�/=s�n�3���B�!GB�j,�$1�Hc@�4�
K�#Q�!(�k�(!2�/ejYR�\�R��ҰTA��6p;d�-��F�M�BD���PC �2�d�j��frh-��9�RJ��
%�D`B�2��xJ�/s;�oyP��Au���Ό&j��^�H�bF�e���o9�jM�*g/u.��!Q�$H�#L�c$
�xL�Xho��B���85�% `(C,LeHʉdn[a¥U�6裥6��D�#wF&%5��Y҂�me�!7 �)�5i(�s*Hl�\ec�rew��k�5�A	�(YT5��f �Tjns	�P���e����U���{�B��8�@��e�����) I$�X���!x�ڰ#F�Dle0*A,��*�E6@� ���WChqq�D���aAi�`���
PH��l�01[����k^XR�jEDR媨�C�,E�/`d��z����w\���F�X%�Ci����T��KѶ#��*���	T��P����J���YЂ@"�[�F4]ie6d�fk��EMԬx����B�aI	"B�0�j/��9�+Y���e�,bF?	Y_sP��Q	��$�BT�E淐�́�2@c76sv�Y �8%3t4fٱztHLf��2M�9.h��͛k��s;�``1[!!�`m	p%��4q���zn�\	I�ʐ�nR�N]X�0Ɠ��iV��u*�lFc�&U�6�0l�� n�S��f��A�#�݃,[�8�/��f����"��H1$Va�ݲ��e�KÒ��%�^��Ad#L
e�$$�0��e��aBI��^*�E(�CV�%^:)(*Cf:#L(!M��$ Q�+w�-�o�����'Ƙ�H��4��և��;*BBJ���u��w �Uc���L�e�M���^a�����1I!	"�I�THں8Z^��˒oBVQ*�U����hsV�Vl�I�R�j�"�2'q�Y��]wg�w���z�@�u�6�l�5�UL�t�a����*��0�a�h��y�ޓP��HU��N����#5���Xe��I7D�Q����W3��e���(��)�E�.a����	RF��l1!D���bCn�[�0��Uʺː�Y{�"PơVf
$�H���(��M	r @�D�!#P���J!.1!L�0��P�Jmd %����,�RX��� ��V�%2�B��ȭX�Ȑ)-@!0�F#Q�p�)-�i-3AD(*�B)$(�lV6qI�{Õ�h@���LEfa��H@�e���}ΙU�і�f��<3�g�x���}x�I.�         �   � ���  	        ��                                                                            �C�                                                                             ��   �M�A[yl4����]v���sU��A���V�l��6�-���$&�$��X6�m�Gh��LPuTpc������uŷ�mJN�t��r�cb��h��d��dY/Wd.�N�Η�q��djl��m�7S*r�ꪙ����Lݶ���W 6��u��F�U���OS�"�9��UL�2�@�u���k�a��$���.��e�e�Bz�mٖ� �d-�V�2�bA:A�%��E���+˻7h r�j���ڮ� u�m$p-��al�mze����  I'p-�k�� ��h-�m��L V�JͲt� H�m����VUUU�
����;i+6m��`�H'Ju�TF/Z4P s�V�Q �`�n�f�Z�j���`��q���I]��ȸ��
��Z�u����!�� ��"���U«����snwLh�֚E�m��K��lW[R��A���w6�i���<l�nҫ�$�Cp�m[ w$�W�=mm�	�[v�kcK:n��H6��쫨
���󶚪U�
��Z��mX`j;c�a����I�m����7��m.�X2��;:�0�V��'g���NXب���*��*~����UԂ&�USi%�u�Qܱ�V������  6ا��i�#�&�&�U�U*�C�MOF��u�d����U��l��f�x���Gm-�m�f�6�-�۶�XJm� Xa^M&ͷ7^�� %+�UT��' ��*��[�z�s���W�1x�$�����h~��
�q���v㧕Q����E�m:*n��;nN��0j8��HN�s����m��O>�4�8�����qs��f���6�tj�VG�=��l�e���,����l�
Hlm��-	nNr��5Cؔ�뵶�5s�H�e�z��n���k�v�IWh
U�`�N��H�f�
km��ѫ=��N���]ejVVBz9�}����n����غ;j�y�_+UUUWb�'Z�QI `h-�� �c�s,�5�
��UU\jk����l��@�9��@���������+-�K ���ĩ�&�gT�U@@S���E�c�q���V��D�K]�!6�]k��.H��P�r4��8}�8�Q�Uc���8��Q����@�0�s����!�H�0}s���d�)���/!԰f� �L�W���:7H�n�Q]�X%[�UV˲�Ъ�ź�RjF��%�6%L��<�댐�<�rh��&vdt���ld��`�ڨ�tM�t�ie2[W�Kh���-�j�ڕ٩�p ΕV�bޭ"F�[D�{N1�t� ,3��9c[n�&�n8�i���N��M��iV��
��/�L��nݙ���u�kh�< 'O6�[\ צ��l  qi&v�&{S �u-�[*�Ҷ�v�` 3����ٗf��v����R�*����]-�6Z-��$�m�� 6�˭���-TjBJ6��ﾪ�X%A�B���l�G:���z�2��8[�V� m����6B�bYV�
���T������ *�cTgp�^�
��UWv�lq�4Ȩ�l���Iz� ' sPY-��^���G;�vjR"�
3V
�c�k�H�l�X���
�SJl����gӃ��6U;�/b����x�z�Icn��tݣ̸�Ĵ �gUuʙlU+ht�l������t�<fxc�g;:ܴ�T��<�R 	n���g�eh]�]<�����T�*'�N�Bv	�U��s4�7��N��7[#����=�ү%�q���,�����bUSv�u̫S��.��%�se��-�hS�u���W��-T�TIU��컧�VU�t��P�P��ݠ�;N�%.�� 8ǩWT��j����۴�Z�I�� �����ň�Yt�j�6ͤ�K�=H􁖀��f�$  �f� A:�[UK���iЫOQ���s-�Xn�t�8-�    	  ���m���$ :tUUT��RW�iX�T��4V�lh $[\�`  6� 	$���@!�ŵm�R�   H�h$ =��k�;i6��mp�[\l�_��o�^� �À   ��eZ��iV�ق\���lʰT�UUUUR��x��^�d�:U����uf6�^��m����:�i䰙��v�N�U���x(�0*Z �����l����`��]JP+��ԣ�W�c�a�K�vX��;b���Tm�Y���RK�j�����H�h��`�����m�� @  &� 8h
�褕�]I��&F��$��]/l�[����`m��kh Zm  -���N�`�a 	e	����f ��݉Z��Onb�k��K�;�51Gf���n��6ѳn�m��n�^����5�I �u3�+��R�-UV��"���h$�� ݶ$�k��\ؒ��$u�_wקz^��nө�刜�f�J.m.3�y+V�	����^K��{g3R����Ъ���Z%� Um[pm�m��� �$m�e�����5�[u�mum��*YlaX�Z���y.�\� �o �jΜ�o]  �mN�I�N 6� szޛ}6�)��<�C����#m�-;kz� x  m�6�   h�Q͍�n�&I!��H�ոp�	��̋i"I��m��KUFG��J����!<��J��]=T� uPQۃ�	���.�P]�����8������+MtS�]���6HN��
]z�g �i6  m�+;;5��r�Q�q���ꪙO=Wmr��J�m�� �` p[@m��I�i�l �  ��  �[N�-�-v��-�m��o ۫`MUVp�)-ml�u����APO��SqQ����������Q��<QF��H����D��@��b�`0!M	1z.�� BX��\�B�$ \U�S؊pUX�� b�����腸-�q��uQ �@n�1v�)�8�GIN�T�Z�Z�C��`��C �&�C�	�ĕ�P-W����G��!Gt�����b+�8�q_��#"H, Ǫ�^*|����@	�h0�S�`��O�z:&��i#�6T4%���C���Q�	N |g z(^�H�pis�4��@�"���@��"�Hlbh���u2-����
'@]�;D��Z�:��)�x�����PL�h��V#O��Ѐl@�څ�W�0V���(�_�h<�U*�`^�! @�Q>""��F��Ρ�-S�qx8��C�G��¦ FI�g -H����@�(i8� E�!9 �I��b�C����mT���T�U
���bB�J�(�C�*B��/��FA�`A$"�#$!H��H�&}F����G`06���G�0V��>`Fd���'ːF�R��S@l�J�*����]�"���)2��l_��H ��)JP� �"H�+�k_U�����w��[@l              ��              l8�ֹhn�F���!;����6�<�����4�tY8�X&6jl�mvҲ�=`x�#itP@�J�����\W�j���.˞�����Jۉk)���:� �N(�fD���{ki�L6�A�[mn5ʥ˚�[qN���̹�� v��cn�آŗ�u�$��h�艒Hv�:�vz\�yn�1mQ��ið��J���/ƪ��۱��]r�셡�G�����e�[8:��Փ(�]���8��v��]��qմq�mn������������G*�(����� Z=�n�[�h��.�p����M�U2�`*��maX�cS��J�j�V�;'���Gn�t�Ʋ3%S������U�G�8&���uKdN�[�rb�B��z���N�h���n��u^��9ar�[m��9������t���L���J�̮�*�yt��h9Bj��M��2[��gn�O \s�Ny�gk�D�K:�i|����UJ����/���y��n�u����tgT�J�촵�t��TAn�-�p��ڝ�AnΦQR0n��4��{C��`'�jmY�����[N4.����1H,��R�4��v�D��@�욜m�g���;y�z����i�����S@i0�>���y>����<!!�)�T0"����j�  6� U''a5 mk�2�'�q]��d&ź��}��>^8�V�z�:�.��_�i��ZG�{kiwr�-�N����y����;.��+�F�WZł��T�ն.�,M��{#��VQ&]T�y	�.�+0^�(X�>�U2�Ϗ&�&����s(PP�C����̩(��*t�{�|�zB6r��q��Nd�SD��7��8a�sݮ+wx �D�B�u��wk��B�9RXe6�b�y�����8a�Z
8K��j��s��A�0빏@���?~���u�L�v�'PAz��b:��ڼ�6��dKr��A�0��b���^wL�R����n}!zn>�p^���7���A��HA�ZM���b�u�o �ީ�ʗ%�%�B���o ��5}����s%2�%��A�0빊�����;�ߗ�����r��y-�kP9�ĝ˘K�:=�Vx�L �D�c�:�b��q��Vb�*K��RK1y��f��A�>W؋=%c��Vh��y߭v�E#�T0D	æ3zث�:�NdKr���8a�sݮ2�Z���YIP��f1]�~|�����M�v瘒�.�fɍ���t<�����k�a�6KI���Vn�����7�R�䶨_w?D�oy
:a׼�<Nd�SD��7�g��y�c/��w��JA��n��0�1���*�2DA"m��79k�.Hi�$���Vf���(Ꭳٍ��rؔ��
2���	;;���gj�`�z ��)��A�.Iˡ}��7���� ����ӐR��JT�_^uC,�=�o\fgt�) �����:�~�o���A��HA�ZM��@9����3|�8cz��#*\��.��s��1GL:��<wy:w����m�     ���:˵�]�j4�ԑ4�\�Nj���M�vl����s��97&z�W����*�i�x�8:Od��6rnÙ����W��[�Н,>�1l,�u9�u4k6P0s��:��ȋg�
�NN_V�"��_�w��w|��U��c#�y�tr�v͸۹箝Yy�In�f��[�#<���ra�]�Wv����P% �D�B�U�~�8����ʗ$4ڒY���+7\f��]h!�ˆmP� �{��A�0��b�t�%9�-˖�f��]�Wv��pl�Ͷ�2�l��S%F�.Ϋ'Y�ر=�ٱ�X(�NZ���YIX����{_���l��l��$n]��u���	��S�&5A	kx!�Se��A�1ʗ%�%�B���o �u��o86��l)`�Ǣ""��3��P��}���*
���	8�O��1]��7��Fsm�Zi��d�$����ƃ�>�;�&)ՙ���SI�*\��jIf/;���q��Q���C��4ڡ}��F����{�U�cw*���K�[��
��7#F������y�%�H9,��Y����q��1w��6KI���Vn�����/m��H���f=о����_n6�J�� ]pq�Z��2��a�mX�{�3ypî�y���KaK���4t�_��{���w���Ph�[�g�:�b���o!Y��.mI,��s��3y	�bX 
�5�.�PC�4ڡ{����o(f'ܣ�{�$�A)L*H�&��:�� ���)OC�@kRg�0��e�S�ܹi�o �u��wk���Ԥ�RT,�W�Wv������%�ً��+7\f�������Xr\���3ypî�y���ÖN3ypî�+�\tG @=קy�����o@     �^��D�6ɓ��[�9t��-�l!f����m<�9��Xrb�8�÷7d�[�	�K�ې뱇Zط���w`���l�h�u�B;9��[�U�
b��+$���^���i�]4QȐ�jq-�l�&D��h0�A*0<ܒI-�S��+m�[��]�]i��v�07g�zu�~���u��o��o!Y�d�䆛RK1y��f���(�}h!�ˆr�_w8��b��w|�\��Js"[�-8��b��w|�wk���Ԥ�QJ��0�������Ϯ�=���iλ��h�Y��J9���G kG7Ja�6KI���Vn����@������K�yuXeL�ѿ{��< ��F�$PjHP�17bA Pj��:a����fCaK���Q��q[���d��d�t,�w�Wv���b�R�I���,�����37���=W�m�ٔ�6��D̄�,�r+�n���X
aJ��0e�9v3����(�w�UΞd�2%�rӌ��(�w�Wv�@�F���Z���e�a�w�ߖ �W)7f�^�w��J���9Zֆ�N5L�.�*k_��F#aH�$�A�	$$�+�-N
F���9�Cw�o4w7�ۖ���.jHp���^�i�$,��A�rW!�i3g7W�-�	.TBL�BA%PJ�8E��a(׬o&����|J @�K��5,�e�dP�� ��k��ME�dc	4�R��T�*�w����s��B�z�� jH]RQxh���SB�B $1�X0�/���QF)��"�Px�O��	�M�J)�X(��D��	>��ZT�h~J�<ڟ ���@��Pw��E�����n:���r5y�b�u�f����1���je�?L���}��^����������-&ܾ:Ѡ�5^<�)q�Y�t��-FZq��ں3�^�}w��^}(_��7�����L�B�����/��{���>�����d��H�c~��Vn���w�Y��h!�ˆR�o=�i�>���E�/䔠xA�(��ij!j�-*�z���h�	�޿C���F�U%J�3�C^@��ֵ�y��}Gs[m�Z	�Ԇ�R)�2���س����Z���y��E&�4�L̲�V0񇗌W���"�ō�fd �-&�_�������y�{~B�(��[�n�]T%;��~���w��<b���<�fCaK�: 7��,�^�4@�{�3�����L�B��@��A�s�5�v,k~���c����     m�6�GU��ڱ�L���,�=�䶌<�.ܹA���F�i��琺���F��]��:Ett��'X�Yw�(Q'kn�%m��=s�\ �ʼip�is斺
�����]�Y=��on:�]:�U��C��+�$�������z��������\%��ۥ��h�(}�x���ls�%�@��*�L��jIf=�s��+7�D,��bh-�E:�s� ���xïc� ���Js"[�-8��1��|�K��{�׽ر�{�K��ꣲ�@�>1w��{����1cw��,��w#Z�y$�!k��V��CoϽ�߾���43ny������6v���c�K����7]w��{�	N]e52ÐS����V�1GO� �BB�Z�"���K�NB�\X��B
|(tM���
�磯��5�w<�GRAF���uj���u&�5�kSb�����/u-�L�jIdt@�w}�/{�V��@<b�؂D0�N������9�|k�� {O�ĒI��؉�&klv�yA�����uq�ڼ�����}��`√3���:b���(_��/��Ԥ��(�B�D E���s����67y�y%U�{�{s��7d�HB��:��*wy�����z��W�U�Q-�� g{���(�" �k���m9 �.,o}������k܆=��Ԗ������[��`��X�ڞ�6�:��Y����绸�����ɖ�7銬�+��  "���w%ʫ��Iv9KZ�'�@����-w��= �ϱ4�a�����y� D}1w�b�x����[�-1�7��7>���a�m��@��jP(�Z��:���r������e]��e�Y��.�h_��+w�}�e�n�e��^���뫕��Yo*C�O-�����ww������əH�w�1Y��~�"��1���˪��������^�Q�����Xǵ6 ��K�T��T���v{g�GP%Z׹{݋:��UXݒ�n��������5�wȾEk���;�]�U��e�q�k܇��\�r���{j����~w��    US�\�L6[�'�p��d:��1���6�4��� �M ��p�h��tF���k\c���]�$Yx�rc�2�mպ،:�p<c���i�9y4�V+�w�ޭ��s��+m�[�$;ڛ�{r%��)���GDx
�d�cm�ܷ%��I��gQ�9��CfK���D�%�g�N�D��a��÷�8��b��@�]�X��<�E�-˖�V 6x�ߵ����D E���J�L̲�T0��Vc��������fD�&e[>	.�W9�C\�b���u$���Z�nSS,9:�s�@���P���vNy�f�tT��K������kӣu�t/���{���%�e�i��y�:a��� ����{{�U�Y-��L|q��hF#�Ԥ%%JaP��l( �,A�(���ý���}�xAIϾ��U�!6�%��w���c����y�<a߭���a�.��=�T^w���p ���a�<�E�-�ۊ��� \�׊v/���$�D���P�� ���S��`�ױٽ��ɳ΁^�Ӧ�L�fYE+|a���k�^w����Ȑ�d̤b���DD�{�3}�t�Ae�hFSR�rT��y�^��)�	��(�0��)-�,(,Uaeʱ[
._
1y-uƻ�r~����B�É!�w�Y�׌h�~�TooxL�B'&[�g�x@�͡~�8��1B���h��T̛uM�mc�k����1�� �Y�����|7lԻ[߯��b�u�^��E�k=�k�C)t5��x�[�OgS`��>��ݹC�9"ι�ct���g��5�v,g_sR�S3,�� ��5����y)���b�"��@t.	�(��4	�Gٽs��QE�����|���5��+[�{/YԒK������?����=��g�mᗆ�u��#�ϻ�޾����ҝ�ѿ{�c;�1�:��w[�_w�$q�
�9qc;��BO<��u�c���I��z�^H]�xL���s|Ί�3����/u#��%6�d~ � "���7��,g~���$�����9��{܋�y �}��ҞΡ�(2�:zȐa$`HH_���	*V�e�~�:��T[��Em)I �bHA��WIU#+f�Gbm!�Y�td$�@1���V:�J,�P�%2��BAi��BB��%!E�S��C���$�	1R�aam+ N�E�7*��HB��A:C��$��(t�ReNɽ}��6�p�                           ���    U[O@^�U�ms��ËRf�M��(5�P�"��*�uns��*�6��2�.��δ9:0%��.�b5��U*�'f'+.v�8h�҃K��ӻѰƉ��î���)�іlZ�v���Ӹ�X�ۮ���_D��[>�t�Y��5�a�
ZyX֭]e��-͑˺Y3�ٽ%�$`�:2uq�˸ܪ�&3Uuy�!c�$��콟h���v��9\���Y+/l�{�]M���
:��.��������=�3�$F�;���_c��ۀ����gK)7<�'h1�*6Վ�k��M%p*:#HrWk��;@(�X�m�v�So�~�}�^�૜8�f�4��[�Ļtx�3���H���x����p[]���������L��s\9�O�):ٲ7(3��p�5�3�B;�&o�<�]u8C�ֈ%GHQUX��ڰ��M�,�I���a�j�M[��N��\���'=��L�nC�g�/�U<��d`�ʴ�Po\�˷UՔUn-��U1�\�g6��$�]&ɵ�N��,���p7�tdKl"n��%�8�'J�g\:�l5M�R�'C�ut�rz�[٧,�E�R��Cm��r���-�䗋�Hm�I.��T���_��""$-I/08 �b� �M(R�!�b=�?�>CBuC�oh|
��|�盻�����9����o@     ۞K�ڷ�Fnq���! ���JXs�ŮJ5�i�\�(\s��Y�r8�P�[�ׅ�t�q�6��Z1&8��י�m�z���Ĺ�����]�G��� O5:�ݛ��8P1s�'%����?d��-�h���Ys*�ffB(�v�C��f�װR^:�]]u���n����&gRg�r}�wN��Qrl����m�?�<"(g��/7�jn�㪎��5_��<�!�{�c;��D�̉&�S����p��8����e52Ò���"�ި��8ۓ�I��:��I#��UAˋ�a�	�LW�X�{\P�}��m�e9r��䲄�b�mҡ���`�V+`��DM:��$$J`�b��Q&��Y&��;�����|���6�kRNW~���"�VDҒ�B$F)PF���2�
�>A����ԓ���Ԓ}ʿ��!#��`��a�.h��}�Q&�z���'d���@?��P���a�y���4�\�������ISH�����6���^K���=y�Ԓ{�~���3��;Z/�l�\ʇ;��a#�������w�I�d*)�T���@z�ל�|#�"O�(�w'x#)���.h��}���L��̀vM ��+�F��T~���$�rPr�{�}�6�5V�hAĒ� ���K�d��uQ$�o���H���a�$ x߹V��o�y���7�����;�0�S��I3D��(���3����-ݴ�IB�R�G������q�=ِ͖�&^�	SB�4Cd�.l���lfk`s��.o%�5G �L	!$��g7���!�4��=ݍ�D��^�RT�e$�:$�l�M�䳰"f���/w�љ��
�A5U,?G߅}��F������~���i��@�����q�s{�\�k����u)�S���޹�c� <#}ﵦ��*۞�ʒ{�?���6p�ɬ�m�'en7�Q����i:I)DʁR��̀m����DC���lszD��JL	���H��K$��z��{�Uz&N��+�_�UB�`l�JטٿD���`\�@z���TBAU*Xd}7��`^�6�J����٫�%
`I	&�9�?G�}�"1~9���c`4m&�U+PPX���}���      .�rTk��N+��6�MC�M�"p۶`6�RL���u1�^Ե���֖9�����aѸ��Ǝ^j=�.����_sы��m�3	���H	�͔U�,v6l�\������Q7.���	��]�T~����;�{��^�F��Nל��#v8��E�r2�]��f��@��5*e32�R��9>(�sy(����">����ߙ2�J����(y����lN��}2��EJ�P��R���lfkg}L��@\�J��)$ �*I����{�����(2>�wo��� **)D�0��q�o�HK���V[z���6����~�����K��7^i��ܻ�x;=�FJ�L��qS�u+餪��6w� �1�=�Ϣ=!s�yWQ��D$R����n�}"��� �_�;���I=_DI����8@H��E�-�ۢN�~lN�tG�77���v���eL��3(�)�?�Z�(���,�_}�D��������o2d*�IT02se �1�=����Ҁ~��$��BE*��ץ<)��܈n����MA�9RCx)ˠ�����sd����������B����Of�HALL�ZtI��U}>" H��Q'gzco��$�
���x�8Yp�&|�K�n��ɉ� �AI �ĊE	��"A�!�N:"""7y�*�;��Q';�\�Ħ�Mǆ�!�_;Q����o;�q��/@-I�և8�����M��U}3��d��I���I�"#�?u��l�e��I�$�vx�ܠ�z�0���y3��$�z=�?>�����@z}s�>�r������	��&�*�ӥw�L���@{�[ל�� �";�}��Rd�H�'��K$�f6l}7���.x�9��J�E �u�:%s���$�~��$�}.O�P���;�e��ٴ�R������lN��\�޶���ݝ�P�:�WD�8��Å�;�v�����#<~}�U��k�\U`l�(>�@~��}���l�Q]R��J����]2e���`\�_�#���J��J\�'���@z�[:&rt�=7����Q]R J$�b&�{��(>�@w���[�)3EI�s��z�%�ל�O�?}z�}��w���^���     ��sV�3i`��:�Ze�J��F�ϧ��ۢ�������
3��t�uG�on�ί$��%<yiV�p�ͼ�Wۧ<xx������Y_�\�l���aRC�:�m1�@�U�ƵlÐ�\���Jh�i%�Q �"���$T�z�ˑ�W-Q�)�Fl<�ߟql�����n��(��`z�G�2t���EJ�E �R���o��d��l�(>�_� '��y6�a0e�i�'7�TI��Gﾙ��J�����T�@�P�RL:"&�J�y(�ca��:>�������a|�Ħ�D�D���d� �u�&�y�=8P�Ř�I%)H���*$��k�_mr�UV4�s��H�T�)5�AU*|gs`z�[Ӈ菡Hzo%vj��)R�$�&��k_��P�%��H)A����E�BA��W�TSC�Q���?M�Y'o�U� @�9��I3,9�FJN�9<Q&��Y�"pB_oު$������k&B��C�6P���o7������'.sB2��%K�_k`w��D^o{�\�@9��b��������d�� �x{m���t��\t/�����)�	(/{���(O�z#�r}��noB�

)B���(O�Y'����{�U�D${�0�)�M��f�>�},���TdpȰNUt`!���"�ByG�T��MA�Y>S��C|"�$a
H� ��E
�:6��)$��-s2�ؑ�cZ�D�ҧ�A�q�5�rV�#Ԣ�D�+kî|U�2^!2���A��h�H!��C8'1v]��j�,�4���H�%V�R�hM�
z��FJe]W�l)�[E8B1 p�V�T���u�8ā1�j0chK�t����U- O��BmPN�� mT��W���%��H<CHl�B�R��غ@�@�]�}TI��7�Е�'	�����s�������@z}r���U�E"
P$�ٚ���]h����{��=qSڒI"e%T�R@�D�"����[=x;7l֤��t߿��9�eB��&����Ҁ������#�}�]w~l���!T�J����(�c`{3[ӅtDDL��7�D����R�>�z��{�T~� Kg�vw��~��RnC��KN�� ����ԓ���&�|���,`� D�m�$���`��a��s��}���:�[ٜ������U:�(��<�9�7��gvy1k�h�l�{���}�ٽ���`t��@_�ٟ�}��(�UXE/�R����������@z}r�"d�5WA�R�I&��`zp���f��P}����f��T�M&�����b�ݭ��3?6�3Y2H$����#/w�s�TI�҉?� �U�I%���m�    ��k^86T	7���,O)�]��5T�g:9�86#>Z����`�N��&+�m�:7'gW@�1�3�Jz�����] �w�sX,�r���)[Ԡ�k��6�Í�]O�3�lH6JD$T�i)BCO�| 8ɫ�Uur������s��d�탷�^+Z�u�5���������p�*)
U����_�/5�=8P����IL(P�@�02�[舙.t�2�{����C7z(P(QJ��$�,�T D%���O��Usy�t�)$U��=��y��}7ZP�QQ8��������s{��J�V =��I�J@�u�mX���(OC��ꩬ�fu��Ν��`z�|���שN��_k`nV��3JI����I7]�f=�WaIg��ƅ~�}�q��v�`e�6�3XLH��������D���`\�@s�&�J�B�C��������l���+;�T�
D
�/9�=8P���l��wRI*&iR�] �؋��K��wnS���N7�w��똒9��{�\�@_��{������l�QSP�*�����l�����]�����QHIP���l��ȇ i
�)ý]z\��_fI7��lH��	$���lN��A�����oL�4���
����@w�k_k`e�6�7RI(J�e%/�I��EP�1s�б���G1�X6[c.�m���ƶ9{�D����@�b'g�N��e5.)
U��[��"d��l�(]X���ʤ�(R �����s���3yX :� �΄�L�R�)0舜�(�� ���qC���Cɮ�f(���)QT`fֈ�ۛ����:P��I$��R�J��j��.��ɍ�p �cV��)�K�*Rp�.Sh�'=ު$��Urx�!�9�K$�k���Ô��9���DU?�6�@?������3+L�4���*i02x�=ub��`^n��f�d*�IT0��?}]���9��No�TO� @�.I�[��)E �C߳�`~��7��'��[�$�!eФ! �D�%a�����'�;�_/y���<�m�      9�빤��j�����՗9�p�<<j��w]!���<��L֕8s��g�o]m��c�-�O3m0����mu�ȝI�v��H�a�L+�,��jn���=4.
��i�BCFS���%BY�p��":�UUUu:us�M�/L;���n,�"�]]����>�����E��w���:P���{z�fj)��R��0.t��/*��9�/;[���WR��U5@��h�yx����s��`���R�����l�(?����Y�a]_��LT�UI0/?k`\�@z����RO�'߾��uhnYʋ�[��㶇\!��G�����2LҒjd���2x�=u� ������"?]��́���!T�J���X+��	E p�kO���޹�a�s� �z⊡T��	P����uQ�	��I��'��ԓ��
KR`{�[�J;P��'ݝ����B��T��I�s��G�����lvk`n洒IH�P��*%QE�QPۃ����g�T��K�iT��P�yx�����ҀWj*ʕ�*RP������y�2x����%�[]J"�B���w��z�;~Ge�	�M� ,"��!�TH#oJ������{u�=u�2LҒjd��â>��V��齔��߳[�3Y2H$���@t}��x������~������L�y�ҞBU;	>6=.���u�~��z�O����O���lnk`\��"��d�:{6��"�R`{�[��B�|�;m�ʍ�{^�:"��o���.[XI�$���K��g`G�@��}�Uw�}TI��'[*PL�>� 8���7��D���Q(@b�c ���x�Of���p�-JsD����o�߻�i���ܭf�o�~�$���l�`Y�3mv���W���y;y��3v�ݛ��L����ҀR�{興r������̧&\əN�9<W��H��J�o������}&ho2d*�IT0.s� �����D���l�(���5R���*X�����Δ�G���=�UJaD��PJLvk`\�.��I�Ϊ$؏�#A �LR�)P�-���L�>eh�¡y�jwG8�o�&��ԼuhJ.�Y�����B��	%�L�1	C�p�H�^��!!GS�-� Ȭ$�D"�c�Č!� �FD�$	"�2E��b c ��E"<�y'N�$��-�� h                                 H9���x�I���B�۩yb�!y��3lbv�y�8%#n�7s@�l��bƶm%�����N�v:���G;UK
�3*��ưD�<7N��9�rۙZc1�*���(iN�t;�xcy�h�Ź3r�6�ݘ����8��ŵm�*j�Z�=Z�%٨���i8`u�����Msl�,\�MvM�^+��D�eݗm=��g۰�h������ќ�ϷE�5Lp�/s��@��x�s9=��F����0mջ\I�Hº�I%�e�mX��2n�p[+re��Hlc���h�bK�}%K ����<X�����Q�2�4v-���I��e��3�6r�F띶�;�P�v�^6�lYᕤ_i�ۂ����A9�F�K�6�p��fݦ�v(f8��R��á�n��[K�t u�x�j���-r;���A�f�U@	U�w�NW�9�j�В������rW2�ݣx��+ml;g�'�6��� �� �g]k�Γ�&��Z.�}��j��)�v�7i�8i:�2tl���zg�l!m�*������ؕVJ�g��m�vٮ�=AuJ����KGF'�������)`�	VE*�s�̽�ƨ�-jѤx�XNVo�>y�y�y��"��z!��2��P�A����>K���X��R� :".�KC痻���~o�d��     ��v"/X���6�.�명g�l����e�{v���s���{qB:�pf�:�Nn�:�hŸ6�Գ�l��I/OE�`쑜�v�9aI���Z�d�yɻ9t�����˯6�;1���՜�z���\�uR�B��F��dH���d��Q.e#`�!��=�6��;l�|�(���NWl}'J;P�{|�G��"�3�~l��E~��)5��T ^6�5�.x��|F��\T�M�b�;���$�n�Δ�(@{�el(��
�&�D�oy��� ��g�D����̭陙�$��f��J�C�p��g6����ԓ��|��r�s�yV�mtq�U�k�۫v�͌��>���2H$�<��@;�l���D@$���M�͉J[�?M*IϹ�b���ّ���_;�c�W]�ӵ����(%DʂR`{s[�D}5z�$߷�D���X.SXI��r���B��a�>������(��)
j)^�@tD}������l�(ʻI$�JRRTTD�)3�y��6^�Y�o"UR�EJ�"�JP����5�.u��ŷ�r�����eF]B]ɆM��U� L��I��&����L���L��re̙�蓳�.��q  ��Q�Ego=�I9���I9�;��PU ��a��M��@{3[�5��DNW��"j�)QHRJ��9�/s[�J;P�Ⱥ�I%	D�JE1Kzp���rm��X+&�9�[4]�et��Ҟ������ԅΔv� �����R�(SQT��J��d~�^�`{�[�H"i
j)^�@?^6�5�2t�ڊ��|��B�a�y����d���ɉ�B�� �b��62͙TI��T�m�xux��" m�I�+�A�RÖ�o�́�� ��@=�l�ﾋ�SܒI[W���d۝��u�ٻb�&ϛ����x�(�B�c`{s[���
�U^�]2{w[�y�=:P�뉪��E!I*�����l�3s� �� 6z򪔨%EJ�4�o舊����?�_� ���fj%|$����&�J��`{�[�5�O]��y����޽�m�     �[F��!a$�qV��NwM�l't�ϓk�a�,��z�jM99�uԓ�'�E<��W!�ۮ�ѩC��p8�^W�a�����OO<D&:ͣ�whˍ�ڶ�ݜ��s:��cd*��X%�v'lh譹���y��w{�]={�3�G&u��n1�Fwg�s�H�<&lђuȻ�|�{����6�k`zt�ڊ��BJU
����o�#����.x��#�"d�+���DR�$����=:Qq�ϽQ@=�lM����PL��z� �q�=�����L�R�f�`]��c`{w['J G�Ui(J�n.π�/��'H[=������N[	�6.Ԯȶ�ܓ���6�u�2t���C���ͪ�*	E����o�}�a� �pCJ�4+�:P�� ���}��2�Х|*QSQI&��(@?w6��`^�iMBEE!�}}9����l����Ҁwj*�TBJU)�`z�[;�����k-�I�`Y�m���JI��懮���=.^�AI�u��k(��vh������Ҁw�������	�0J�&�02t���Oe�@z���u����p7���T�J����ٍ��e�GF6��!�C�9���ԇ��z�q5R���)%C׺������ ��;yUJaD��Q*��u�2t��B�u�.&�I$��O7@������=���gT"�:��5�W����=Hd�@;���`^��*6�IP�������"&O^k`gw6N��QV�J�R���u�/w['Jߔ �u
h���T�������\�\�%#�@�� @�i�s�әQ�I�'gJ���n�����l�I$��V�˶�|a�pJ� ��i��ky�� �0/qB�1�/w['Jz�q5R���RJ��5�/w[�Jߔ 6v�Q2������s� ��2MvuQ$������tO�N�(e�@>�l7��s�����]4������(@<�l����҂oi�d! D�B ��O��m��6�   US�ۇ��ɱ�Q�F�b`�	�n(̘y��M;Z�]d�tg��r\\y��Ev���b����Z@n2�Ba۲6NٺY��㵞�`\vQ�7F'+vƭ�1���nL-��pT=tH���E�[��D��D :  DNݶ�l�I�*Z2�����ɍ�pl�9��i"���e��NRӔ0���TI��l�?�!�]o!M0�J�I�}��艓'��j����L����Jf	�f�02x��B��`^��f���!D�P���w��{��t}9\P��&�R�	B�T0=�́{��:P�� ��I$�J��笛F痋��<
����]Ėe�����l�+�t������Ҁw����ff�Q@��/35$�}/}"N��-HI!�a�l8�����P���|� ��ln�٤T$(�0/qB��g}��ws`d�@;�`�	T�SP��g6��`\�A�D�-��[]
Q��i7D���Q'� �Œkq����߾��N�$�P�D���H�@�q�g��8ct��_L~���)��*f������B����}�����7�ʪ%
&j��/�'�5�3���J��q5R����U6���m��0�/8�!�:�CT��Bw�	sF�"���ꛫj۟P�&�Vk{4Ť�0��J @!	$#�� 1��%$
���E04$"l�I����BF62��x���z�A�@����D�Z52�MX�f5h�Xi%X"����E��V�B��J1�Ү����QM2�� �2`T�dX���TTҍjR�Q�H$`CFAe�Ԣ���n��[�.[��Bb�[=AkX���4�ˊ�����1#a��C��#���mqN�@��� ���6�/§x��_�xR�` @	��;z�$��jI5&XR���~����'�;P�}|�^j$����&Δ}��8`{��ݽTI�ަ�mː�-�BCD�O<q�&ܝ��[%{<��dT��QP�����������Δ�QV
�J�T0=������}��<P
�� �[]
h���URL����ҀW����]�l���D��`\�@+�����>�>�	r��Q;Q0Kϯ�jI�N���U2�5Cۊ��5�.t�o��;�U]9�z�ϮP��Hl�-���DOhϮ�����5)J��I*<��`^�Δv����UJ��*	I���o��'�� _7�>�����T@������<P	ڄ~��g߳�`_o6�Ul�
)
TR�P�yx�����DG� .I���-�h�(�o�D�����䝯K�f��I4�l�W���bF�]24X�^�uU����    m���H���g2�`	�J��)M�b�����.ث���"��,9t;b�d��'pN�9�sqVzj�g��3��93�9r[��ܵ�4�ɰ<�
a�,�;U��"�n�	�:�8�Ag��3�{r�;���wx=���|�UTU�Y�Ag�,(`��z���v�w?�{��3�
h���URX��`\�@'V~����r������)�&��JL�(����������;���eT�L��� �6tD}3��'�Wx))nXi�r��� ��}�I߽�0.t�����UUJ��*	I���l��}��}|�d�$���4��t�K�'k�G2�瞈ӎ�k��-D��r<��:P
]�����zB�y�/�WM).^L�/&���}YA����QKj�����!A!a�I) 5 ��~i{����I;���s� ��U��$R��,nk`{s[�JK�@?VV������tD�oy��� �X�}|��͑R��iMT���Ҁ菡�`��g6��TI�/�m�fJLJq.e���ޜP��즼�;Lg�|�5$�H�B�U40=u���`{s[�J���R�
�H�`{s[ۚ�:P	Ո�����3**T�	����$�}.Y�ĉD��"1b"��2N^uQ$�w9p�lL��tΔv� ���=����ժi)
TR�P���=����́s��z�S~~���&�ыz��S��5Q���ڱ-ԁB)P�0=�����l�(�B����|��T�ۚ�:P	ڄ�����l���JR�R`\�@'jo[ۚ��h�MJ*�F�7��$�f�o������(��%��%����!%�U�B@� ��$��
J[�bL�D���Q&�z����]c�� p׾m���:���!��8�5�ƶ:�"��-�.�q��mv�OrO�߼�:P	ڄ���2�T�!M"f��&Δv� ���=���}���FuuMEM5�P��Z@>�l�(v��!"�	Cۚ�����Ҁn� =9{
B�IJ�I���l�(�B��`(�"*"'��	�i4�<(�wrI$�H    ��rӢ���<m5��j�1,��)+��]�^�Y�	�,�	u�;I����7n�d������b���u��dC������n3��s��ali�u6�7!d/^p��/:�ۦ;UU����l��ʡ���t�qGw�ߧ���%��vN�T��d�&���vn٭I���1���*���Ҁn� ^��u�3�ʚ�(USC�T �6�u�.x�  ��𤥹a�$�I߽�Q&���� L���Mް�>�f���XR��I�� x߽�a����1�F�=� ��R��4���I0.t�������l���RI*�P��	Pu���h;=�wg�u��>H���M���)QH��� ��=ۭ�s� ��U�D$R�(d���  � �b� ���$������R�JURLn�`\�G�f�Xd�����x��4�I��ʤç+����́��l�4r�j�J�h`]������Έ��&���a�SNe����T()���1峪:�[A��*�T�P*Q$�X��6�u�.t�������
*T�)0=���s� ݨ@=�l/uJ�Ғj�$�}.I�s�[>�BJWĩW�ZF� "�DJ�R � Y{������lf-SHP���ã�3� .�[ݺ�:P�EX$BE*���`w�_w{�t�@7j?�j��:hQ��{Y�=�&�V9�7I�1_$�T�ۺ�:Pڄ���ŧ�Nd�NZi�'���@�7z�$��6�u��>�3��ʚ�D��������g�3����{��RQ*�I5�����Δ�&&b7�%�T ����$����wu�at�	I���l�(�B��lD�����k�˪�-�gnǵݹϋV�h�nff��P$�:Pڄ������V���HQH`]�����n�Ε�%�(�H�BP���lf�Q�L���N^��5k���T6��~����'���2>��W�[v��
��JR�R`\�@z]���`{�}�I0��i���˛4B6��@uh.`q���|P�Q���� �!D�U�,� r�E@���T:0�؉��4Z��B¬�6o{�2̂Q���X���vU>
J�,��Z�*�0��54BW �e�eh�6�e,*1�Zd&bc[̺,�HXAl����p�DH��"Nr ¹��@n��m ��}��
Ε�M�P��h�3�k5��n��� 4��I�O;��{�w߿-�h 6�                                 H9e��ܷ+N�y��u��Ū+st��l6�r!�j�=q.n*�(���0F�u�OlAl 嚨mr��^�;q#l��"��.�0�nѪ���0]��wB%׏(<��l����m��.7�5�,�d�zT�Ӎ�f�'E�lѮ\�#ۇ@���m�uԁ8�AN3�s��Vc�!���5�!���l�s���gq҉����Fz�ضd�3���%����cŹXu�[n��Ő �v�wI���h�;&�n؃`n��	�fۂ����S���l��5u\�Y�"q
f@��gF[*ʴf�'�#�xԺ���1�؊���� Nim�ލ"uv�]��On��c�\݆�9�Ѷqsv�^z��#g
���g�u��\���r�\�@N̒�k�-H�q�LlZu[Q��leM���J��Hgp�٦ڀ)bl�ʖ	����4;$KRd.�]�E�c�჎:81����=.�e�4�[r:JҮ�J��n-�u��JZvɑ4l�������2�1��8}l��Mg�V��[D��d�۪�Z�����$F�s��M�:��
�m^YS��E�պ�n����-ϛdܕ+�<Y�"�Ѣ�9u^��Fsֻ)>��u���y�"��O�q��x���C���R�DH�dA�M`Ё�*�E�|N��ʽ^���޽��o�     śKZ[l����2Mx�	�J�û16����j����8gp!Q�$q=E�R,��vn�e���r���]�-�u����3�F3��*��ܑ��{C�z�b�XR�X�`��Ů�\��X�;3@.�uդ6I���N�m��e����ܓO���1.r�EjY��ı�Dȫ�J���I��|�'��lf��Hd�@?^C�T�J�SR��g6�u�.t�=.�t��ٵSR�B�$�L����ҏ���7>�@{�� ��T��4���)0.t�=.� ����7��`_r�4�	
)��@~��ۛ�}��:PFfg�IV9gL�¸5����,���DGc�sp���������4�K�$�����}�TI����noe�o/$�m�I�$߻���4D @�b 6vx�NM��MfmW�2sW�Jd*��R`d�@9w(�́��l�4r���*�h`\����`{w[���(w��%�D�P��g6�����'��P�sv$��..�zɠ^�!29��������]�����.��)&R��́s� ݨ�C��g6�ܩ"Ғj��J�P�{z����G�%�.SHP������&���R!���@Ġ�Q  " U��$��D��aa-��ND��菦�{�����Ҁn� �+aHW�)UI0=���s� ݨ@?��}z�}��~����αI�.[��ۍ&5m �Z��v���I�)��R�R�<Pڄ�����a�9SUH�U40.�B���}����l����Ҁ^�êT�J�MCۚ�����Ҁw�����@�J�e&��`\�@;� �!��!x�c��m���*��Q)&Δv� ���=�����~>�����\�t�W����.�ݒ��Vv2T6ȨHQH`]�������O�VD$R�(`{��ۺ�:Pڅ�2z�k�HWԐ��`_w6Δv� ���=u�¥2JU*L�(�B��a��՟�~�q߇*j����ި@~�fo��s`\��Gw��w������Ͷ߀     �d�5�s�ƹ�t���0�#eU�uպ���c���&���[��v�l�C�|�7�ٗ�n���@��i�C�ë;�]Fy�f��
��E��\�F2�<��q{��{��\����[��0�V��޺�zǝ�z:W�9��u���M��)ں����z���a�R�I��i�2�w=�Q'�u�.t�!H{ء�ٴU)RL���n�Δv� ����>��������Q)&Ov��}�?6�s`{uj�@����ި@<�lf�a�NW�(��P�M*��9�/7[�J��P���;J���d�6��ʈh�G+v�N�����>d*���s`\�@z]�}����̈́�����ʢVe^]検���(���� ���B(�"��-J".^J���=����f�T�R%UM��@;�l���7�́�� ��U$�*Q*jX����n�Δ�ܠ6v�(J�fR`{7[�J�~����2�5$�%���j��Y{7nN]xyg�s�Rb��^u����vv[�cԓ���I��{����y���Z��B*R;��yx����s��`�
r��$�oUs{��G�`L�0 Z@.,b! `@y_"u`�ng�z{%�jז�$�M��tI��l�(M�Po[��HPJ)���Ҁ�ߥ ���/7[�2����Zyb��t#K�%������63��LPJ�*�h`d����`{7[�J?\8�I(T�T԰=���L���:P��L�=yEP�BU32����.t�=.� �����D%�f�M&OI���I�Ϊ' F�� \�����-SHP����ɽ�����oUrx�KVcm���2�ET4��h2���r&
�M�]�����qL!B�5*|��`{7[�����{,�x�x9%Bl���M�s`\�@z}r�{z��/+N�Jf	�T�L�(O�P��ٚ���2�I�.T�D�""yw��ow��7�͇�����U$�JP)�`{��ٚ�:P�\��>���fe$�I     Iwf�������,b�7L�jT��kr*8�C�▿�����4��H��ӌ�]�U� �۟k��O\nx�]�\��pvK�n�2�h���#��be��.X|�D^˯6��g�pө_/W�/=���\��=��~��;��������2룛x�J�:�pv��pk���A�a�(�BU32�����:P�\���ϻ�I��|���LL��:$��D���@=�lf���#�����"�!E#D����MnmQ��-��Uz~(�y�,%�iʗ4I���/w�_ro&ޮIPۖ��{������4�L?��,�[m"[nPl�D��A�.ٳ��|�m�jL���%�ĩ!4�q}�Y��}��fs��ޙwwy%e]^���K��T��@"�8 %xk>Ý�߾�Ux�I�Ķ�1]��fk��B���_f�ݸ�$�����B�Iｕ�z̼j��>q���h0ؙa�q}�Y��}��g|y�y矝�����B�F���I�����rd]p�GoV<SN���,'�Ǿ�{��g�������0ӕ.b�y���܅��� Y�����-'C;�q}�u�� `���rgJ/�лfPT
�+����!N�m�hܔ5ƍ �p(D��ɠ�Y��K���D�3EBI"��HP�a�M��a,�(�RB���h���O�f�14A��@�����;�&�������᭱��!�yĕ)P,P�*�00_����ނ|�q�#�Pv �: �4E�z	C�6��CJ�?k�a��'L��Bi�����Y0�9�D^��3w�3-)d˕*��釙�Vv�����m�Y����X�}նx1�U�:�:%�홹�S�������/���ُg��H�XmL̺��� ����{0��q�͔܆,9N/�5�����q[���%�,'Co\�7����*T� H��,洂�S�r��V�1� E�uF{�Y���~�@IK�k��k�.\��t8Ⱎ�Fɮ��\f��7]!CN\�B����!f�a�ss��Nd	����^���{|�g��D@�#7{�2ҖL�R�q�L<�} �s���uxI��LK�1^�1Y�����Y1�١��3.��s�g��ه��"
eƭID#��Q뻰     �!��{X财����5���p8���[z96�n;=���fKd�cmnn���ۮ�ɋi:�s	�wW#��;t޶�Knc�ۍg,l���n�Wh/\ь��wn�Ւ�r�O��xa%0Om��D�q]��w{���|�UN&��aV^e �q�s����cs30�e���S��!f�a�y�����̲YA��t4�L=�b����!y�,%8a�*\�v���/�5��W6T�C聝�Tg���ɇ��s��Nd	����B�d���+;\v�m��h$�9w���w5� �9-yn[�5��4�)lB?w�_��3X��~��#=�(^ha$�I�r�+��(� �i���f�c�'4"r�%���/�5���gn�a,9Lx w�C�ÿy��k���fY,�\��9��X��q��e�6�m��*,;�볆��n,���j��v9�7
͙�uB9���+7\gw�@c��fyx8����t/}��@o��ه~�� �N�2S�(�̼Ǿ����_�� ��b"k��ny�^o�e�,�r�P�����+;���8�r*�0���-)���/3\grs&=׀Ϲ��\�-�a;9���r�����b�]]D��9L"r�-���܅�ɇ}�3�e�C��N3�z 8wf+=�/3Ϡ3���l�a:{��X��8��/-����R�z"�����o=�� � H	 �V4@hF  �kf.�6Sn����BϿ���߮��|����αI�-�n;v��ƭ�N�^wi��[%9�!6�q��Y��w��fs��ޙ���eʕCN�ý�+3�gr*�4QH�r�+;���c���sf=�ЈI˒���^�gro$z �{�7���,���'�C�2sf+=�+3�68@�T	"�	;+����33     qg.�	�d�FuA�I���:���{V��b�;�nF���=�����!uƩ맬(��Qfy��k$���4�7O=�O[.<9Yx�ڕ.؉`v���$E�HѮ��ٲ=tY0�������ֈ�x�=��p}}UQ4#�s��v�c=]�J6�m�򳱕�:��B�νz�ηk^����l��Eil��nT���y�@�y���Y��w~^d�
)�B�y�w!f�a�ss��)̉	�ی�B��þ�+3�e��̴���T�w��Y��;�t.V6�v��^[pvxZ��;[��W��d{F}u�%��^��+;���q��Y��������*Kj���f�4�v���Ͼ�s\�7�瑆��[E�ؙa��}�,�L;����q{���a�a:���W�ǄA�y�´�Qm�T���y�3�
�������ߠ%b��[�Y�vӴ��yr�e��<�a������v3��3����Vr���)̉	�ۋ�B�pþ�+;\e��̴����W������sH$*�HT
w��gS��B���)��Vw1Y��;��DD��=���I�aImP��8��y�������m����JbQ)��F�*[��g�1v�\	M�M�a�2��q��]Nw��gk���C�\�����X��q��� kg
��	��R�^��Vn��rS��.bLʆ�mн�q��]N�0tF��|�˝>d�2$&�n3܅��}�Vwǟ�����^�yd:mt#K�n5�dћ�lv|�9+�K3,�T7'�;�b���o���R8-�����q��]�����������܅��}�/�e7,���ӌ�B�pþ�*�^��re���f�y��^s��B
P�B':.��x+�$#�=��Fg Ry�5Ϸ����G՜�Z���J"pN-t`� EiCDf+f��0bB(s7a%U�efH� �����wI0%ѹ����s5�i��& (�S0�˫����N���#6h��tNG#�@��
�\��8�Z��y�X@����M�ƺBN�n�� }U.;�J+}�ۀ��$��pʟx�:#�`�*�����W��+�=�����N���߶�� �      �@�                          A���t�!n�iWT���7����K*��G�z�:�mF�2l�$(}�S�h�d$�j��m@7t�;j��Ҭ��JD�Egz�N�6�*Ƶ:-s�g���gj���v�Z��ݹ]�sH����-/���][C�J��p��p�Z�׈7Fp��	�è�AjT�k�5�m`��W���C���-ەא{cx�C#u�!�\kaN܅�d���`|�2�U;k\:����q�e�xq�m�$r�����rclpk��]���wm��ĵ �y��:p��<�ҩ�����gg�6��KbS'������9S�U���kH�gW�s�k/ǴN4pt�]mۖ8��)[��)�0��sM��n
N�u#��\��֍�;[V�"�ў��ok���U(^'+j��
kAb�d
q *��[ms.�̪�UR[�і�/ݺ����X�t/-��
�+Vʭ�i��f���v����)�Sz�L#X���c[@ !5UR�mXҙ 0�c@�W;ڝ�d��ۭ�6��N[:��"G�;�ݶ6�z�$ۥ!ж�W*t���U�@>���m���*�5�KYv^9� �o�,��V�v謎�A=�[[]�ItS����ʳ5Y"^-��޻���.��j@�ȃ D?����T>�m+�LCp��CӢ1jo��n��      +����v�Y���:�}����M�4�ÂG�u��g�M�'r�h�]�:{M�.Ƽ�#7N��٪���X�;^ۭO��=�<m��-���7H ���/2���6�۩ ���9ӧ(��&'��Ǽ������l5g�n�y�8�nMӝȘ*�1���3E2�	��R�w��U港rs�����h����܅\�ݯ�ogO�)̉	�ۋ����#`�������*Y�eJ��<a��y�+�
xR�)�h�wsy�+�
���w[m�ؔ�q�n:^Q�;rm��ҏ*Z�-��j��;e��j���>s��B�p���ٲ�!���'ܮ)G�LaE�~R�����r3׌U�@�ooxXe���oO�<�b�<⻐��8�e�EK#� ~����q^�=�i��^peCE$�^o�Wrs�v���km�ɖ�l�����k�5<��j�5�2�L$T��)̉�ӊ�B�p���D
����	�*Y�eJ�{<| �Ews���^��)H�b��b�7�?;	B���mu�z��}�'4"rXR[_��  f��B")�z� �	�_f	 �&��bj	 ���rQ	
�K���m�m��M��0I�5�{PI�;�hI;Γ���:~�����[�m6ܴf�۷O-�=�=j�6��՚���*T�T.ab�_\؆�\�ؚ�H&��kBH$��z� �	��$����˗Y4$�H�ｉ�$�o�}�	 �'}�L�H&�}�$�H�9�_��n\���n	 �ｭ	 �'}�L�H&�}�$�H�罉�!����7r��I*LlCh�{i�I�/��I\��5�:�t�H$�0�� �N	�����hI�9Ͻ�*�%VK��n	 ���0I�5Ͼ��A7�}�lCh�{h�Cb��$��ێKst���K9ft�%��8��
ݠ��WJ/f�Z�v��7�{PI���ZA$N�֙$@�ZX�H�L{gx"�h�����$�����V5�>��� �	�_؆э{�b��򤌄�V/4$�H���2	 ���`�?�&�4g~�F��k��0!��\�<9
�#��FX��ow�6!�c]�PI߾�ZA$N�֙�M��;XJ�32�&��I}��5�M���В	"w޴�$�owقH#h��fF���rx���$�I>I�   ������vgex�5�R8��Sڝ���<�[����u����V�=b̈́rQ����h��6s�ln�U��3YymSn�n�s�=��n�f�Ol�x�e��6ݫҽu�v�s���F��(��x���N�����]����{�=�'�{�	i����v��)�]�x"vMZ�s�7$�*ܹy��z	 ���{ZA$N�֙�M��0I�5�{PI�/��%�QE�U�hI�;�Zd?�
�3���3�z#Cb3��Ԫ�6�o��U*�:���؍����	"k�}��$�o�~ք�I���A$g9�WwvVL��$D�}�MA$w�hI�;�Zd@��u8���6�{�Ζ�ܷ�%�bH'?}�hI�;�ZdA5����1��#Cb2P��I$���%�z��A*^��q�r�i:��E';:�Jz�:N�;�ZdA5���$D�=�MA�����6�s���*T�T�a�H';~�� �r	"w_kPI���$�H�}�L�H&�}�eˬs/.L�A$N����A7���	#���߭2	 ���� �&ϯ�2�B��#,Cb5�{؆��z� �	��$D��ؚ�H&�Od��E�L��В	"w޴�$��
[�v!��;��0�6#>߱�Γ��<������7j.�Mv�;G'ZSY뱬i/*�
����Y.�I�$�v�,I�3}�&��	�w�В	"w޴�$�l�:j����%a�$D�}�MA$w�hI�;�ZdA7�,I�=�W:\�����zM�$���В	"w޴�;5�2#X���#�X;5�YbH$���������T�7p���0!��}� �	��bH$����5�? �����7��Ò�r9P��e� ���$�H��wPI߽��#bF��Db��x�I%S��r��c/cIì6CC��գ��s�n&'%�gG}��ݢo��&��	����$�H���? MA$o�$D��~��­²�I�!��=�%��!�s޴F!�\�؆�3�Da�lFu}~�ܪ*�e�f��I���A$o�bH$����5�M��ք�I��J�u��%��7��*�B��V$�H��9�!����m`1l�x�@�iz����2	 �=�Ʈ��˙�u�$D�{PI��}�	 �'}�L�H$�jĐI��Η����m'6�vn�oQD�n'<Y�uumͮ�79��BS��1�߽�`CbF��FA$k�bH$����5�I�=��8܅T���m�m�lC��ĐI7�bj	 ���ք�U	"o��%8�r�s�؍ם�lCh���0�6#>�1��m�m�pM���˗X�^\�4$�H�ｉ�$�o��ZA$N�֙�?)����m5�ߢeE
�0���׹�hI������MA$���$D�����$�@0��> �D~O/N��;������6��      z�mv���[��r[g8�9���rc�0Qz�&�v؜vK�F����k�l�p�v��뇃���L��ܧ�H�izYnְg�rÞ��bn�g��y��0/7p�\�hc�3W�Ղ���;�ς8ٞ��PR�0ܤI� |�6 &�n��
w\h��5����p����;���m[0p�o3�H$���֙�M��I�3�bj	 ��}�	 �'y�x�ʺ�U�����H'}v$�H���PI߻�hI�;�ZdA6s�5wwf\�Y�$D�}�MA$w�hI�;�ZdA7۱$D��\�r�2�e�7�N{�kBH$��z� �����6�����kވ�؇���H�rPu&6!�oݴF!��؉�3~�&��	�w�В	"@>����^ck�cu�����W�����T�6�m���V�F�d���h=� ޷�A׹��I���A$]��.���ʙZA$M����: xP�#'�����}��ZA$Nw֙�M�e���T!�`׷�*\�2�6'{��$�H���2	 ���AD�{�!����7r���.���đ;�ZdA7]�$�H��{PCa���g�9�{�T��꣺�&��	���$C�uϾ��A�=�lCh߻h�Cb3�U7$�M�+n��g��������i�����v�:5�}�$D�}�MA$w�hI�;�Xxxb���m��|-��B�e�7�N~���$�H���2	 ���؆�3��a�lC��rTnB�	Y�A$N�֙�M�e�#��)TT�x��E�@�M���rῸȡ�:�nt:��PACL�67�.��"�	��f��$�M��"^`Qh��v�%�p9��#�ݙ�,�'qc�[���eղ�4��'�J9�D4��4:{��]�Y����E��Va*�Q����(����P�(`�X�"�J>b��B4f���

��p�0�j&
i�%0o��Ns	��U��&�D>��)�x��
��4��yP t0Kh�h���'U�>�$���c`' �'6��Z �G˸�s�bj	 ��ﵡ$Dk��J��r9P��e�o�/��6!�c[�F��g��0!�:h�i�I����wWX�^T�4$�H���ؚ�H&�ߵ�$D�i�I��B"0:��[m��RjX*L�v�gp@(�����ь\N�rI*\�2�6#]�q��"w޴�$�n�,?$�H�׽�!����7r���.����6���L�H&�ĐI7�bj	 ��}�z�Ch���R����������y؆�6���#Cb3��ؒ'}�L�H&�s���2�L��$D�}�MA$w�hI�;�Zd@�F�@ ��D!�A�Q("TʦE���Z�tQ43=,I�?k���˺˘Jr^�!��=�lCh�{h�Cb3[v!��g���؏]�s�J���;<ݹ9i�͹۹v�����`H2�h���flI�>��� �	��$D���xI<��׹�`CbF�����ə2���n	 ��K_�Ơ�&��Da�lF��c�7��#،j�iJh�ӒY� � ���D@$&�ߵ�$D�i�I�vX�	!��**(T��ߒ h7��8؆��z���f��CbDϽPI�/����ˬ�	 �'}�L�H&�ĐI7�bj	 ��}�	 �%�����	
F�ߝ��     ���v���"s�x�ܥ�J��Ev���v.�t�����\�3�c��b1n�]&;f]yݲ[���%!�����+3s۝u���g�^�i�m��ݣ�����յ+<���1��.'NqYK�ɮ3p�'R�h���BY���$�ԷR:�1��V ��`={'�[6A
*S.T�2ʕ�8��:PCbDη�!������LCh�h�Cb4o|1WE�)�-�CbFw�Da�lFy�c�7��#،�݈�BG}��wu-�S�0��$���ZA$N�֙�M�e�lCh��b0�6!�]�8܅TfhI�;�ZdA7]�$�H���#Cb3��؆ўo�*8���/4��H'k�ĐI7��j	 ��}�	 �'}�L�H&���s33.L�!�n�T��}9ܙ⅌�:[!3�4��"z�	�7�{PI�{��$�H��֑�lFkn�6!�c<�a*I�n	 ���֖�$H3��@��H|� 	j���$L�-2	 ��KA$Mo�bj	 ���=�^UyYu��$D�޴�$�n�,I�5�{PI߻�hI�;���VU�J��w��A;^�$�H��;��$�o���$�H��֙�M��MU�teL�sBH$���ؚ�H&���В	"w�ZdA7]�$�G����$�nIVU�e\*;xmH�8ۈ�B�u��J��B�]Jp�伣LCb7��؇�z� �	��$D���MA$����8܅TI��m�m��M�e� �&��bj	 ���ք�Ch�7Ε%2H�Y&�!��� �&���j��R��]���(&�l@�����5�$DϹ@d@$@�[�)M�rK4  ��߱5�M�ﵡ$D�޴�$�j�,I�5���1��³3I�$�s���$�H~#��Zj	 ���� �ь��b���I$����r4:�7D=�`�'�� -ԙ�ܙ-[0p���{��v����ZdA5]�$�H�߽��$�o��ZA$N���VU�J+%��7�NW�� �&���j	 ���ք�I�z� �	��髺(̓+.hI�9�{PI��}�	 �'~��A$U�bH$���\�r���S+4��H'=�kBH$�߽i�I�vX�!J;"M2�4�U�ȕ�،1�|��InB�\���H��֙�)��ĐI|��L1�Ͻ�`CbGP�p~���Kr5�9�r�vn۱�R��sU�rMzxe�г�]ǿ;�r���mη�!����� �D�߭2	 ����.]�B��ɡ$D�}�PI�~�ZA$N��L�H&����T$��{�[���w*ab�{����6����$�b3\v!��:��0�6#:��F�Ur�˘غ)����1��q؆�6�gވ�،���8$���ުʺ�Ed��&��	���$D���MA$~��В	"w�ZdA6u�e��$6��D�u��     ���{4��\/Hp� f�quّ�&B��.^]M��Y��u�)^]b}j�2�赫vW��̼<g\اvrJc	p-�F]e�ح��W/%�w.Ԧ⪗��mn��ss�vӮ���0\XvSN	����!�T4 l�J��33ː��:{n��sӺ\�湦zx+v�:9�n��h���v����9�Da�lFy�c�7�Z#ؚ��A$O���K�u�0ʙY��A9�{ZA$N��L�H&��ĐCh�{،1�|��\�����0"A$N��L�H&��ĐI[��0�6#=�1��m�9��S�9VI��A9^�$�H��{��$�o��0!��|�1���7*��˒T�4$�H�ｉ�$�o�}�	 �#|�1��m؆�6�����ޒIXi�ey_Y��8�n����V��nL�Ϯ/\�2�1�߽�`Ch{�l��S�1���n�QRT�qk|���K�
o�EGh�����K#`�n5���ǽ���r���J��0������xR$6K��^w1[��7�goT�eK�Ò�о�q��3�w1D�m�:Z���h��E���W\n�<b��tvfF槵q8��7�g:�b���n��Kl�A�xì�+�\f���Ғ�)�$���k���d��(W?��z�M�u�AF�p�M��s��A�0빊��̔�D�.Zq��3�w1]���=���7j.�i����l�����@��=v�=��X!-"YIX����{\f�]�iH��.Z1y��n��A�1�Sx�.KKj��s��A�0���pM4%3-��	߽f�c����x+��Đ���D ���W��}߉l��urfh�����q��z n��m��fQi�2���km�* �Z�pg��6�	0���ܩ,2�rK1��1Y��7ވQ�~�xK��j����F����{�`�O2S�ܹi���g:����q���.T�"YIP�Dd��^��k�� ��������w�Dg��v�yk���ͱ���cm�� �T��� ��~(�>h??����I!_��~��L)�Ι��e�� �؊�=�H($���� �,  0�
 *	��I�Ϗ�1/-�?�	�������8�?��#�L��s�݌�S_7o�hs�|�"�ɰ�L�$4h鿘�/�/��� ��Fl�BG���B���g�����#�c;��C�{�s�~�� ���G�3��`�AB�1?���l�?a�J��>�D��}_���3%*li?��:���e!$�)BQJ"���" %D �E�EE��Q��p�
�,����`�_�~i	_m��>��p_�Bb�����K���?q�H?��_�?`0B	1��\�/���>xDϵY�P�"���>���?g��Ө���~ߘ� ����>��_��D�����kS_�b�̡��$�>g��$3����3�2�s_�:죧��ih64�-��BB)���:XR�Q�C�AR��d��.m����#A��W��0A��}���S���>��<A��������}��>(��4Pϧ��?��3� ?Z��~��d�	�!~(����>'��>'�>f��?��y4�(�I?��1�)���}�>Ol�ޑ�|���x@�BG�<��������}B��I9��:S�W���AS���|D��|� @!#�>j}�B�6����0��cLg�R�1���?�]��BA�8O�