BZh91AY&SYҳ����_�pp��b� ����a}�T@� ��DJ� (�( �*��T%(	U"������ �)T)* �$*���R�)@QJB�*���T��U( R *��UB��%)UJ�R �     �    ������{�_>�>���}_]�5W���y�1��+��Wg=�� �=q=q�p�  �\` ��P7�Pi��U8�]'TP���n�h�=K�5J���(\��Q�ӭ
q�@ }�  @   S��zU5s:O��w7�ۼ����nTs>櫋W.m}�/R�@r�[�}�0�] �^���ԫ� =<y��>��C�Q28z�x�[֕ͥ�9:��͡8� 
 (   �d��Ic=�9e�NZG-��/� Sn����˖/i�u)� �z������x(����^�w�J�p ��W.�8����>�}Ο���z��Ωqe�gk���\ >�    P P@ =�_s����,�n^}���=�T��=8�X���qA�Ɂ�>�G����e\�t����t���K� ���[�T�L��q9�S� z8�d�j������׭��\z �      
3� }Hf��.X�\�.,%� CS&�Yi�,��iW8 _g�Jo�����7 y ��Y.m�ʰ He�0�y��ܼ�w��0��� Q�'nA�k������W@        LC�
m�R��0��bdb0�ODCR�SI�=� hɉ����z�QO%@      D�*�	�R �� �� S�S"�j�R�  F@ �	R&MF�O(�dz�z��!��'���_����^���a�ﾎ���{��U_CW�AU]
*��ʀ���Uq ?�Uo�e� ������t(
���_i U��_���S��?�~�{����f�:�q���j"z7���	�4AްL�2�bwe�V���=�s��݊�y�=��Ƴe��Q���Z�pcd&4A�c�&��1���ba����Z�d/���ޣz	<і���M����{,)�ҧ]�k�E|O;�$�u=��v�B�n��[����A��fG�zN��w[�V��w�f��K�S���G�Fh�nA������;�]��bADC�MAޣ �Jd�[�ɥ�(J��5	Bu	JW��<�W����5��닫��wv�L��8�nK���AYU�8��.z�/�|v�=�~;�'�s�]��5s|ߖNi�؝]�������F��x�Y���+�t�o�BP�%	Ho#G��0�H�&y�aPXaG���S����D6`e�=BP`G`����9rd�*��'$3(�F�Ga�K��%	I��}u[�r��C2�3�c�i;�4�rCYb	BR�d�۫I��w�!���!���c���)�[��CV!�쵙�o;��M�4鵉�KΒ`(������vy���}u�va^U�[^I1R�L�YO�=��{��&�5�XS�e�����7���t����畺ﹼ��\�uQ�I��4ej22GD�NZm΂mtZ��"������ɺ:c4mu�u�q��k���o|���P�Fo�:�)	�}Aw�]��ʜV��r���L-qw�3�}�Z5�(��*q�d�N�.�[UK��
�N�0���_�w����Ds#F]��r��,��6��x��{%,�Z��R�R"����*@���w+u��c�=�:��ʢK�{�g;�\DǙ|C�1���峱�L��t�uA��z�x矗15����
�%���,�b�S�z�����8٣4yg.v�(J���E� ��-�h�h��(<#S�ż����C��0��dC���i5��5jE	�'(�wpT	�D�`?�fnZ����s�s��A�s0�Vi,4�5��[c<� -�rsNZ, ���	!5`I�0PZ�ַ��e�9asx�2ִ�!a��|�η�q��"#��yG1�4�\*��T���:�'*��bkm��R,W�!ם��)�xN�g����<��4U��t�%���9Bw�٫	��^Rڜ�V{z`�L����u��+�<�ּ���8v3�6l�Y��*3"e��)p��&	�HjUiX��]w/�ğ4|̧T�MEȮ�	��h�{��)K[��/b=�|N��14S�sl�!�W)<�_g���W*�;1�kG,X��V�W�ڰf��e�K�&�+е�}�p2'շfqN$"�Ő|�]�}]V���� ��hj�)5�����ؚW�(�P@�+S�`�F�yxƝ����s[�@�R�um�	bCLdK�^@����֝�I���&P�YHpt��ւ ��9ۘsv����١��	���m�[������T�f��#��F����$&N1�N`G��S�^Z6m�2����]��Y��:�7�ƶsRNEX�d�q�Z��?t�&'|]ū��X��Ўa�j	�$龿Y�FU�%������{�=�mjMҢ�����mP�!�����&�4�(Sm�.���W^�c����{�ԥ�y�Sw��i`��8���}�J�ke��G�yrܥ=��0�5k<����7	��a��Z��4�e���ݧ~qE�ԭ��2�ȗge{��BlM�f�[׶���FcD��\
��2�ߙ�����_cfP<J�j.�ua�U�+
�*�%|��2u�)�l�3�|���5��h�K��:�NN���w�h5;&2tZ�cV���k|W
I�D�/+k�GE��<Xk��O�D�t�3���_ZH�����&�=��Yns���skk/P�|*c���ˁ��l23	,8l���۩��[�!�2\��"�	T0�Nipw�MI�q���sm�R�$T�â�A8�4`F��5΍�J
���ɺ�A�@���}���/��Ń[9�K�����(��;�u�CAj�5Ez4���W��̥�Б4ؠ����s�"�D�|E��a@���[ QJ�8���9�؊��1��^W��q)t���R.e��WcH�R'&.�4��i�4��*�H#%��]Y��_O.o5Д�Ef�V��D�R:�B�B1ܵ]�q&jb�������$*4hFu=�n�~oy����q��K�[+�EF�����o)����r��SB~R�ҲVePĄ�)w�+���l�����vر��/y.���㦲u$9v<����T�t.n_};�ū���ю�Q.�LO73|�|iuSĦBs3s���|�җT�'��ZE/[�2�0�;rqrB(�U%0�UcWU�Zɕ�y�+��r�]���{���O�.�;.���)��M$*ِ�m&A8i	��+�]#�(J�Jp���qcrcÛô�!�tN�0ܛ����!,��5�%%2�%ӒP��1M>�8�0��4�vٓ�{���}������B�R
su��)8�sV,]f%�Bior���e����͏���V	��z.xO�Թ�lH�G�hQZ��d������buf�s�L��I���Rt���<�J���Q5
q��������9���8�ñP�E��i��l\�,S{N��r�3%r�Qvs�伾	�N��+ˏ�e���2M^�s��X��nį)xI�!H���1�C~��*��r��]Y�r�K{WlĹJuyPC;��v�Кe7�BLi[�F`�E��	���"��.��ć��׳3�\����,q��{���!k������]ֹ�Z����rnq�}�Z�}�p�#�r̦֓�0�CA>���%�G73�\����=��;3��1��!���5��{�8��M:��8�.�_Sb\����5+�M�Yĭ>�!�}&.*�8�_���qQ �wB٪>uAΖ{o��s7���i�t7Rbd��3���a��\�{�ε,yli8��@�Ǽ)��H;�aZ{�u�[�f�c�a�v,��+g3�(yy��\Ĝ��Ԥ!,KFwm�	BX�D�Db�� ��r�#�]�A)B���|��ӭ��!�f5	BP�C���l�,p�C�e�D�w�����#|v�/v3����P��	BV4�b�dY!np
�^Z�:,7�5��G'��I�d�FXÕ9F� ՞���=%���[�!(����J���m-��sV=I�<�:����fJ�U��0�خK�x��Y��ʨ&#��5L��4W+�:�'�T��\�J�S�������-Z�i(bD���iZj��O�Z�yX����#����hN!$Skk��8N�p$�Jqw�m��b	�`ꌌI�p2�)�w9A�KA���ѨM�a�1F19�(p2�^�����&�lNF�
Wx�..���$aВ�j�m�w	C�d�S�#����;�%y�<����TC�9���\��<�Y"hr�B$E�e;�;����;��"�H�S�q/aNjV.��gWĬ 20�*
�� HN��eU���f�޲ߖ�ӫZ$�ZB@V5)�iX��^�����u]�5���cnĶsq�EV�4�rV����r�f<�jX��Ȉ��%�hp�cy��Z���Cy`t��V�M�K����GY�0�hrsNh�X����޺�'�FD��@Hbj�k�WJ��wpQ[��J�|\9H��x��$wJ	�"br&�Oa�^����k��AS���*-��Ђ;"����w�8�V�/(Y-$��D��(��8v�co�Т�<@�����x�:���>���58\�'Q�'Lj41�~��ӷ��r���w�Z�Ģ�	<�4|�I�q���q�B,��	����q��w�{��&�#.�F�f����jĈ����T�^��5�ׂP���L��|(}�ݓ#!,;�5�uLdo-G*��:\'�#�a]�2Ԣ5�"E	�.�R��v�0�L���"Η�r�8�_ �,|&�S�q�rr���fv�$7|�v��r��I	Mq%8����K}6.�����w�a��T�����p��J:t�v��a�+�~�u��N��'�,�ki���I�Q҃3j�Iq3ܛC�М�&QQ&�b�]�\�����PT�Pj#�V5+�:�k��Ԣ�]�&��� $�ά��/) �<�LB�1�ݜ��^�v�Mk5R0��&+3�����ʧ���k�33%�{�<�����U��k,	�շpF�#r6��OQ����V4��i
E:b�
�Hl�w�)��]"�bW:�8�6��LGD���_;���
"f'-��̊�T���/���hH)\)N\����[@3�����-X�#*�����s�-(�]��)2�	>)�E�	��+5f��c��!������s)!I�m��� WXN��'Gw#[krc����;�.��;X1u	H��Y�^+3p@"ல
���E.����13Unړ��;3C�V�����a��w�:�"5�e��d����}{�dki���jLF*M�Q�G Bjz�M�]�s=`��Pi#^�����,Tň�j�Eh�176��e	�bːN�4Jg�]1e=��kz�y��Z�k�Y�Ap���%	���{�t����*fa��p���h���E:��8�ΗQ�`�mXh�Q��q٭�̍L	A�u�2	�Z4e����� ,����ј�4ڰ����*x4uL�*� ��6��؎˺X���� �2-%�BweS4-�%�u|�k��4Bb�.�v5}���HHf&αk(�]���ǆ���CI;���Me��Q��T:�*qy��nw���p�&��bmբtI�Tj{#C`�o|�5�@C�WxʼE1 ����$tI�g��R�,;B�Q����;HV��hӨ��]����|�X�GRճ��ba=N/f�[H�N$w9MRC5�ca�%Ea���OC���ӑ�4w��jŋ1"�P�Ļ��̭C�m�c�lQw{��\YQh$�S�Eu��-X�((��e�ϛ��Ν�/���ɫWE3��0`08f�V�z�'T�Q���ӲmX�l�0j	0=�X���g)`.y�Å���PL!�OrdMa����ε�1α^R Ɓ�x��i�3�+Y�|X%��$Rc���]�\���4������4l�G4��9��5���DTB�&$	����W��)d�n41��(⮔�D��ӯ��{�v�_��m�          `      9��  ���Ā    �A� ��    :@   m��JB�)C� � [AͶ�8       � di!m����c�-�p     �2m�� I��T��7ok4�b���U�u۷95�v��m`:��U��Ҏ�s��s��ɒ����cz�[yJi�`ٺ�[C@-�Q9�vxə�v��Q]�7BAS���Һ�.��y��{�:X(+�;���ͳ��J+�=]U��UPԵ��=�0�*�R���.��͞�۫gvݶۀ	%:�ܾ9l��V���U!;��qm;;L�X$*��
�Qr���3uW*mn�� �Ye�l�^���%�2�\:�b����齉.�ր�m5� ���k��\�\�.Z���68��i"U�'W�UF�k��BiV�E�@��}�溪�T���m\�\��â�WS����H4E#Zt$��*����]���Wl�1Z{��/a��9��˧9[i�΀by����X��`*��V ݊�	ڪ�P�ڠ5s�)l �]:�o/Ui; 6�e^�c��iV�j�L�������ں�VT����ou����  7%��B@۩��ZmO�!c�Մ�Un��PZI���7 I6�/=�7YXbv.���[�p-S�xv���r��Ђ��n��:�;� :T-:��óW��bLhwmvr����(*�؍��;^h-�px�V�#��������2�l��V��Պ�.�Z�ʣ	��9U����ݻFs���^{mφ{\N֣�[)�c[����t���8���݆�iKm��m�c=/��Ŵ@ .�5��Um j�ua�d%d{5A�dw@s��(�nQ�����k���M4eo-{��R�=W��,�Qy6��r�:B�\��Ҋ)6ʫ�T�R��Q�T�2�R�=��eC����ݹ]�����؇��e�U�jw-J�]]Om��^a/G[)�sm�]�Z��L���UTpU���&�eV�+iI�,���ݪ����RC�80���)Snr�e�Bez]�4�NP����[� �k8']ס���y������&�N�m��A��� �&��͵	x\�R�T�WO.l�we8,t��v�:@R���������K�5�j�o0�m�D趀U�i`�\�J�UR�� h��>7���EZ�����]����buŵ,��[pmpm��9�-궅�0,�'���uU];\c�Ш���6��ckwH��[$t�܃(�6ڶ;m0P�X�m��8rMae��Z�&VB�
���  m�h6ت�b�)܆�]�AJ��� {uC��l�]N��[#r��͛:^���$���� 8��Q¶5Щ�HUP<ݨTt���V���5Mcg+��@I��c�&�6��t�ݴ�j�"Z�v�1R�n���;��u[�j���M�j�1βg�]�s�L��v]�w�ͷ��\��z
�4P2�u��[Κ8�f�*K���t�iKh�WN8�/V�@��v�֘����,��L���Uə��}�ꋳ�k�7�5�n޹�V��
�.Ύ��%�g�3���M�چŪN� �kMME�Kj�q�JP�֩�u9v�;:�V[��'�<�Z�㗚�^vjn�Pj���NMS&�.˳R\��9�[p&�K�cu.h6��mg+�mÅ�r�k��̓D���iamV��#�s>�0�̓�.G��p�UU@mUt�:8y�\��n&۶[���okՀp����KT��+^�J���9��ruuӉ��ꩇ2�k�� H]#�k2�����V�v&ݭ!)��������J���UܫJ櫈�6�:�   �m�4V�]&�b@�l��%fu��A�m�Z��/i[m�L�I�\ԧW2��+�
�յP �[!!z6�E�@ֶ���۝��ļ�R�����qQ&(�QB� �r�Ӟt��!c`4Rg.�#!�L����Y�z�u�R�۰��T趋��y]�:^N״�e�]���f���K� ���(�n�6�Qn&嚺��^2Z0ګ`��X\��n���%��4�����m��+Ars�Uyy��YY��C  �]�]Mu�������B��j��@t�#m��n�hs�휶�m �]�Nն�lu��Uu5%6���8�m�ej��F�K&؀��h��;-u��ڒ����jRZ��Z8�Q��d[M�p$6ؓ���k��sm�l  ���m��+��lÌ5UF��:*8��u�Rr�2�B�i�[[l l  � URJ��ʵT�+�h�m�h [4l�uݶ4IG+̇l�I$��[v�� aF��yz�[;#UUUU��f�6ضCµ:L�
�m� �6�j��[( At��2X����I"�$�m�G���{4\����WKq����d#��A૪�K�-媭��
��YKd�$�� -o  ���H��g��m��l$9�����i��!�I� �m�!&�F�*�Uj����cb`
��[VVg(�U/.րim\�ni0�h@UJ��V��R۶��b���s�Bn� ˻f8�=��@.��; Nj���N�p�l�ڄ��`A}9��p��bö��ہJ�k�W����rNY�t^81��u��`���=�艣n
�m�T]��zbb�g�J�a�n��j�����F�Kf��t���i%��]H үJ�:CmѮ8 ,\�M�G�6�m�V�*�Z��
�g���kdG��Z���PK�.s��7^~���z���v�+�@@yy���D��� �Z�qM�ĳ��t����i���{[)���a92n���I�c<4lv�Xy䵐@�7;�96��Kz�`	C�v��"�m	�ے*�e ��}������k��D
���m�+�#N4M�6��6¤�:[��b��U�뤡W�kcv.�]#�p�]U�hV55R�C���eZ��#� ��lj�g-K��*�UJ�(R�7< ���V��(�z;]Z��Ԇ�l,��%��7Z��� `Q�-n���ԺX;Q�J�^̬�umT�n����6zL�wDʵ��tF�s;U^��r�~������  p];I�l�2A'h�ɀ5��,KB7��Z8m��  [@�Z��ڗv�vZ��ڥXa�   ֶٶ6�2[sm�l  +���{bZ	�W�}��N�N:v�5&���P6�V�\���s�+UHN��˲�v�R����T���%`�wD������ZE�V���Vj�`)V
[�Yyj����!��S� �6Ƞ l p�ݸ�#�m�ض�ZXm[[m20m��pr���R��	b�VfL����UTjn���ef�Vy[H��n�	�M��p�Ut��V�,�Ut$O.7�*��_*���B�x�+����J�Ϊ��3�Pn�i�m���5�p7NZq����YÞJ�G@'n�mwM���^��ٵO.ҹ.*�Q2�Afv
�h֩��G����U!�ݻx�.��td���U��I�p# 7^�"Vۛl��bt��-c!"��״Q��$]\���j�j�3�K�o�Om�@We�"�@U�[T�� �V�����Z�UeZ����v��i�tӧ��[���m���`�6�um��m�[%m��6�^��� *�iUVvWeS��vi��m��P nZ֎�X�HJ�� V;q�N�۱mh���	i��eV'R��UmE �D���{kR��͞cԜ���q�bU���<�����d��UQ�FN yW%Um i6�  ��lYݕUpsC�mb���pH�(�  �ݴĂUJ�9�va�+��v��h2@�.� l�JO;J�.�B�m  [c-JZ�*�] � ��6�7��ʿh�UC�wi]RmUuf�հ-[D��/ s���	n�k���[\���Qڋ �U@U\�6U�v;'�)-z� kY�j�F��[ErՉ�r+�UP](+h�3�.ۈjyZ����e[Th-6ְݶ P���F����j^L�����UV�
~W�[��� [M� �n���R��l�n�+��ے[A�6�� 9΀���f��m��V��[WYvm��0��㝲ѐ -���XY������mΎ��4M�Eҩ<��H;��CU��q�m�J�U��<LQ�=�S�g�%1��S��EP8�Rdڠ!�P@��Z��y邭�|f��-�
n]���ƃ`����  h�ղV�a�5['�RtZwjŻ.ӷ/mk�  ,��  �O+�U*��J�*��j�T	Z� g.�����ץ�$`�v�bl�����$ה�;v�@n�lH �M�����+W�_[­US��q���X�U����Mu�FWLy���mm�    U/-T�P�!n�ĭ@&�"@��kUA��`
��R�������I	rfͱz� �kvS�d[Cut��0]!�v}�$�UU�yRP�y+bN�v�����ԨpԼ�@5K��SjNM��lF�zQ�6��p6�6��ku6�v�-���4�Vה�Z�m-��5���[@A��2�ptv���V�r�+A�W��{�0Mn�H��Jm]��l��AӶ7��=�s�ԪjUUiv@�.Pj�e��(5�ἷ�����ݽ��@U���(*�����������|����xӯ�?���� ��4����!��hO���� �BR T�bC ���K5 �	$)�|1=$T�z�A �'J��'ZD0�] �J�(����Et
�(�t�#��&
����Q��hסA6'6��#fIHD�B:���@]xv��)2��ad��T�������`{ �tb	�=G�Н��<qA;���@�D��U�D^>��
��h_�"B@�M
���9Ʉ�P�=Gi��PO`�8 ���=/H�z�u��lE��C�a
�S�,%LL'@�+� ����C��;I		$H�a�#�@��U�C�¨z�`�!�	쪧x���*���� x�=QS�Л8 b�!��"0��#,�T0��+�	���E�;CFP�Mz1���=Tҁ.�`qP��E=�"�R	N�C�W����M,BS+&@I�,2�R"H�m@0�����S���
/h���&�>C!U��LTL1Q_C�"�	؁�x��'h��h�d$��QT�!�4��3����!��U�Q��2eL�`bZ'0��E�S(�0�2F�I����H�`�2"�0<;EЇ�iB�2�I(RP*���(�6���~�&��i�Nr.�L	v��K໗�� U�I��������?���j?��Pr��SL�̄(		"�S'(h+2X�r.�Dk�(H�� ���AM$�	D���y���ѳ_@� A�^l=����h-�'���|���-jR�v�'�"�fN)e�Qh��q�-\oeR�zͫE���2��Ա4gat�i:F
�M�%��u��&٬0����Oo[L-ֳ��.��������GƦ�<q�;g[d�;`���V�ܮ�����"Х�<�vz��nel��)�8�4X���X��q��6�.�=��G\h1��X%$eG��b�C;���@�����M�5�Y�q�=�0�M�[l�]��$�j9F!�:�J�k�e���B�Z�H�=�5��:$�U�yς���)�y�b{&��׳�Wqu����{<E㌓RX�H�煰��.�]cU��q���.ku2��:� 1�V{l	�ncN�u�.�e�v�ڮ�R��t�cC^3ũ��q�m��p���V#֕��aB���.��yhq.�m��؊S���������&׭�l��� ��-�vsR�z�n
a���6煲��@c��@KQ�c!���v��{=�⊺����V���Y�{���d��7 �:�X���= ��-��c��1f��ȩQ�IWZ�Q�MC��j����cBm�vW��t�m�-�J=�W�N)�#���v�nY���t�n��y˗�g��v��B��Y�Ir����]�7c["���▧D���&�m:ItͶ��d,�J���bX4Ͳ	�$��]
J�RΊ�4�d�O@�]�vy�U�Eh	x�N� �6$��bu(�+m�puڸ��>��<��h��Ҟ-bZsq[%9q�i�y��B��k8��]ƗuÈ��Y�M�+���Š`!ޭ��*����LM#U9�ͬ��tη��M��7$d�2�@�88��s��qr�V{C֨�b-��M��n�s�cO/I@�!��.�)�g����U<!<����t]R�ڕ�m�V�['-m�n8�k UUշ;(3��#��́���[�V�1����룰،�v�-WM�����
��CiV�����T �\��<�"C�����D{�/J�HT	4 ��=@� ��!�(�T����L����;�r�1��*�f�i���.۶7Z��7��Uk�6^�&��I���lc�̧6���x�ܶS�#���k<�푥����6���em��7�J�1�Or���j�n*ڗ<�3l۠L� g^�%pe��M�;JE�J�$�D�Eй��45��5ړT�8]W��@y�#\�Y��q]l���ř�ٙ��̄]��.�*���!Dd")$pL�ݶ��>�<g�p=���AGJ5l�wqXn���zՁy?z9��� [��2�iPC4���ܗw�owqgʩ������~� �}��n�-��Վ�V��ܵ�s���}� �}��owq`�-���v��6���}� �}��owq`��� ���jU�V�V�ܗx�����ŀw���}��J���ѧ>��٫���o�&��d_N�X�\ˌ����xv�1���[ӎ:gN���}�_b�;��x��� s���y�G��r�v从�wk �g�椴�)Z�N`�b��|T�+�{��Uߞ{�A�ݕ�pY�(����j�m��� Ϸj��������{ڪ�>�M�q+����m����ݼ{�� >�����x���]`꘭4����{�� ;�m���x����I�w��߱�m�:��A-�n�ю!��c)��J���2Y\�u��'m���L�+�4$��Z�tx��< ߻��we`��$��-�7WhI� �{� s���owq`{��*��|}>jU����;�.�����7���)yWH�F$IZLFS�vXz^� s���:���lD�թhM.���, �}���m�;�x�tsP\�ݷ%��wk ;�m���x�����ŀ}J��S��q@hpy�{M�����<�\ۗ�um[����mq��\����9,�U��ma[�I�����@�wo ������x��n%w�3UU�g۵i�ݝ�䭬��X��< ���.�uLV���I7�w۶���ڱ;�uU�}���ck@O�-�b���� >�����x�{��\W���{W�bm�{�_s�*����Ue����BM�{��{����, �}��k�M����Pqs�����{i��(ENӶ6����i\ʘnm4��wK�N�S�m&�{����+ =����U�� �Y���6Т����X��o 7���o����������c��X�� 7���8��0��, ��օ-���V�x�U�� ��"�;�� �}���-ĮErI#lww�q��6ge䱰��V��Ձ,�� 	�X�D�8
��k�)v�N=������}�}���� �7�
 �Zݮ�����X��=r�e���8!fT�me���Qn�Ҁ���l��/�нNu���l�Rvi��5�C�g��s�Jgm!�h�8:�X��{gn.�������5u�.�si�@����3�w�5ͱn;�t媩��6PqJ������������,�K��ؗ4R=����n�q��~�]�{ս�V�-ۗz�����qu&W�4ո�ځ�'Y��p<ŷ��g
���~��`{� �{o ����7Q��R��jY�ܵ����$�}���~�`�vV�]\�%eX���o 7���8��0{w w���
�ݚԫP,�ӗ%���ـs۸���� w���:���m
Z�jZ�0{w w�����xwf�UK��������;����lm��qגfcZ����d,�!�=���va��,n��mր{� }�s�6��R��V�}�e`�Y������j�o ;��w�_��i �eZ����C	u�YĪ�Rt������9�}� 9������ڪiU�ZIYm�o�r�9�n, �}�����_�m¬�; ��Ԫ�>�~���~� �}��m��Xu���4*hHu����}�_ ���0wۋ �u��Y��rx��6wGR=�f����o77����kg]��]B�|bځF��s���8��;�ŀ�����Z�j�Zr��8��;�ŀ����������ڻ	`@�s
�=�ʮ����Ā�$FS��*�T�uyR�Ja��x_�f��f��$��n��Ӭ ߽� 7�s�5��0wۋ ;��=�]��v���;���ـs��X��o �i��8��8�Ǜ*P�p���
b���X�9y��Li����<(�����ـs��X��o 9�m���ߗ4~b�lE�I�~�ed�������~�<�d�s�t��ݺL.��� w���;� �}��s��X���Ĩ_��ݥi�	w��< ����W]��V������⧦�Vm�^ WV�kR�@�+N\�x��o ��}�qp�߯ 9�m�:���vl��1�(=�d%N�@۠1u��\�N3[rvѵ����Nzv"ä��9�n, �}���������u��bL�۴14� 7�s���������q`t<m�m�[���ww��������q`=�^�j�V�܎1�� s���9�n, 罷������!W�rK�����{�x��o 9�m��O�4b�b�N��3�zk�̭�+�vٮ�n�+��I�ۭ�u"͹�D]��x���6���h�p뎀��E���
����J���+��o$�mP�=^�Zyͳ�1����p��d�A�KKT�K�-ͺ獗]Dv���P�����JR�����ٸ�#�*�'��c�%�� uv�H�, ��v*�2W��~����������`fϞ���6�E.����A��wo^��ɠ���,>�J�n���iCRe����sx�ͺ�m�'*S��fGAonx��%���O�}��;� �}��s��Xt�&2"S��rIw��������q`;� �.�إZ���.K� �}��s��X~&��~� ���<Ξ�+�-8���wۋ 9�m�;�x�{����uv��ěv�&�`;� �}����wۋ �|�d���&N�۸ͫ�N���u���r���u������tI����8��f&� 9�m�;������U.1w�����q+q�rB1��s���*KEUI�G	D�q�O��������t5z��U�; �r��s�۬�}�\������k�WV;R���s�۬�}�\���9�n/.�ij"S���w&��>��'c��O���o��ӧwff�y�R��i�1����Jp�0��^v�Kl�p�W�x+� �Y���>������]����+���g;�����cwe�*bX��|Ͻ���o�U>}��۴�݆���֛��,r]�ے���s����(I�T�y;�f%�Hi�_\�۷�+����'D��+�$��>�Օ�J?<>��pw��^�zG�u�޺�����!<�#FgwEp�1
c�Ξ�:``���{8F�s1���	K|��_l!��w�ϱ1A_W;C+��/���R��QY�z����:0�oE������(0�^ƫ'�8���8�:2ND�Ą��5�%��u��--%!9;��#�p����y�����BaؑSD���e��s�|#B{h��sY�&��9 E2iHp /�Sr�bg[,<
��5L���x�L(��O�{{����6w���G����'��f�
��}N s�jfB�qԠ$(Wpd���Ɇ�(vv{�68�+2s(��M�����ǒP��JhbC����t�#��O|�Q8)�b	�; $��Qq�	��@P�>DH@J�
�p=!��1t��a��R���o�R��w����)K����m�m��ܷww�H*�*�}�ث�R.����JR�����R��!.z�U��;�3���*Y�&*bfI����z��.����JR�����R����w`w`gϽ���w`wnnm�j��s�t��֞����y	Qwn7�;�y<q\O ʛ:�%�q�ޜ� -_�{���N�����)K�=�|R���=���[�JR��߷�)JO��F~�kF��խ���R������rR��=���JR��߷�)JN��߸=I��%>>��p�i�7o7�������)Cߞ���ԥ)w��o�R��w�pz��/<���JR����u��;4o4ke�s|��JR�Ͼ��):��~��)J^y���$ ����44�����sZD2`��?|*��s���ԥ)����YF��ykuj���)JRuߞ���R����.>�����~�/]���|���Y����fU<<Zm��65��N�N�*U������Үz�έ6��š��N�?�)K�=�|R���=��ԥ)ߟ}�)JRuߞ���R�����_m��ܗ.]�R
�
���U©R�Ͼ��)=��~��)J^y��┨{~��r�J���3.^b�H*�|��qJR�߼��R�����)J����*�T��k����D����s|R����=��ԥ)y�o�R�>��pz��;���)JO<����Z6�z��ڲ�o�ԥ)y�o�R�~TH>��߸=�R�{��8�)I�{��JS�����BLތ��EBRA& -jҨ�Ț�ݻ�����}�3��"�D�N�!��.s-�j��/Eܾ�!��[�i�W.^�i�t�<�ݐp[��pp)ٴ+ؓm�q�9�=s�4�<v�z���Ks�t�Z��,Oh�n�Mj��N��4^�s�kc��-����b�cf�FH���X�ݞ�Gqr�M�'g��Y��h�cqBqH�}���� M���w}�ۏ�j��cY�`[æ�Z��^��\����Zݸ��\+:�Mź:��ݹ{�ۘ��M�F��\kҮ6��)饉x*Z��&�&�]�������R��<��qJR�����R����yT��..���E*�V▌3/1W%)N�Ͼ��):��~��)J^y��┥�����)O2��vQ��ٛ6eo{��):��~��)Jw�{���)C�~{��J��ߵ�)J��k7�V�X�.�۹x��R
����\R����=��ԥ)�y��┥+�{~�\*�U.�����ӗ.�仗�)JP�ߞ���R��'�{��qJR������ԥ)�y���)I�~���̽�qr񋋆Ocv���tF㗷1�^:�A�u8��B��u���|�=��`v���|��)@=���)JRu������;�=�\Ȣ���{��#ԥ)�/��~�A�Z�ڳZ���)JR������=C�6 ����Mg�}�)JR�ߞ���R��<��qO��d�)n�C��+�;[��\*�U/=����)C�~{��JS��ߵ�)Hv��J��w`wmt��T�4�L�UCL�k�R�=���pz��;�=�\R���>��ԥ)�y��┥'G����F��7�5���o��)N��~��)<�Ͼ��)Jw�{���)C�{��JS�����ֳ�[��՚5�2���'�c��pS/n^:ܜ[\�
5.�x�j����flٕ��])JR{翿pz��;�=�\R�����ԥ)�y���T����߭[�c��[WiܼU©'y�k�R�=���pz��;�=�\R*�R�~߱W
�K��ރ>N�N]ɭk{���)J;�߸=JR����)N�X�+�3 ����I2|=�*���u�}pz��>�~�eR
�
�}�K��W#�$�̹y��)Jw�{���)I�{��JS��ߵ�)J;�߸=JR�e��a�ޭf�Y�k{��)<��~��)@~Q�5�ߵ�)J}���JS��ߵ�)�m��{��~����Q�7Vi9 8�j�%�ڷ\v�xv2�q�Ul�ñ�][�g6��nω��͆oV���7���JS����┥�{���)N��~��)=����*
��_oū�d��ڒ�eR
�	��~��ԥ)�y��┥'�}���)N��~��):>�>��4�ѽ��35�pz��;�=�\R���Ͼ��ԍ)�y��┥�{���)O2��vQ��ٛ6eo{��i=�߾��)Jw�{���)C�����JAy"��H"�"�|H�ԗW߻ٕH*�R��}����v]��{,��=JR����)JR���}��R��<��qJR�߽��R���O��������;�[�)����v��)��mu��ۇj7&벺.ː�o����qS33U56����ιw[>���{Tۥ)I���� �R��<��qJR����r[�\��1��U©R���0�,9)I��~��)Jy���\R����~���-)}�zg�h7�Y�VkZ���)JO~��=JR����)O��~�����)O3߿k�R����|�娓�;n�p�@����L�T��{���)N��~��?(��;.]�σ��(��4L44�P����)JP���}��R��*K�����)I��~��)Jw�{���)I��)�B���>�7�FoX�o2����qÍ=�T�[ok���!���/S�������N|y��z�=Z9�!p4�l=�Z9Ș�g��1�]*�)<:^͹�m\�i���u��Kl.x3��= v��1v�+X�����$�$�7i�hTc`��nyl��+�[�n���q<qە(�3�*L�)ۇhr"�n9�G��L$gh�]Vҩ=��L[.BU*��U�J�/�8�컌m�i�65γ��n^�}�Ǌ!S�׋nټ#rr;��n����h��"�j+��xܼ�_H*�����┥'�{���)N��~�
R�jVσ��z0�UE4SS@Uo\R����~���!Jw�{���)C�����JS��ߵ�ZR��o>��]�%�,�����\*�U.�ߞU �T?}��pz�JS��ߵ�)JO���W
�K���!�'m�]���v�?�2)�������)O3�k�R��}��pz����{�qJR������V�Wv7	��f*�T��u��2�QB�{���)N�׿g�(~�߾�\*�U.���x��J�n�r]�-_6�v��n^�<�.�ʻ6���&�x�ny&w��w��P5�RLQ$L�Tۻ��Z����R���~�)JP���}� �R��=ߦU �AKw���]�Q'pvڎ�pR�����5��E�@����8����7�0ֵ��7� �*��;E%(z�����)J^{��┥'�{���iOr���l��Xe�l���R����~��ԥ){�o�R*��}��pz��;���qJR��Q��Z���n^b�H)R��~����)I�����JS�����?�.C��߿pz��=3�?~�c���[6j���R�����pz��? ���o���)J�}���JS��ߦU �AK��Sah#\-w��m��H�m^��Af{[ 7nr\���n��{��;X[t�Ƙ�������T��qJR�߽��R�����k�J-�~�p�AT��ob�v�%۹z�qJR�߽��Q� S%?g�k�R��~���R���k߳�(
���\�q+�ݸ�3��\*�U/����)JR{��}��C��"E蜕RX2`�S*�L"�O� w)�k���)Jw+g�݁ݏx��&(�����wjA)>�߾��)J}���8�)C�ڕ������j�w`w`v��@�4�ެ�a���=JR�}�~�)JR�Z���������vvd�+g�ݶ�������vβ�B��[[�Tڙm�.x��v�������.־�y����5��[ݽ��y�)J���=JR�g���)JR}��}�N�)O�׿g
���y���U��'e�r�p�@����k���'�{���)O�׿g�(~�߾����}��n�5��"���j�����ԭ�vvJuE�O�!���~��)J~��~�R
[���7,�Yn+��wx��R@��~��)J���=JR�g���)BHK�A��4g�7��q�ZHu����G��'�tnNu����)Jw�cz��N�d�w 9k*�U U�o�b�JP�U���~��)>�����)O���R����O�ϵYfZ0�6g'�v��f����#d�g8���������[<F:yF��wws7�C�Z'.~�~����{ݥ>Ͻ�\R����~��ԥ)���Ê(R�>���pz��.�/��5N���ff�7�qJR�߽��R
)���ÊR�>���pz��>Ͻ�\T
��|���Iv�;���wx��R>�߸qJR����R -)�}��┥'�{���)Or���l�kQ���{�y��R��0*�C����pz��?g�k�R��}�pz������~�┥'���~ѧf��v���s�ԥ)�}��┥�VA�K���݁ݻ�[[��:^J��w)L;Gv!'R�vG�S^�'��b2�����)U}���K��,t@A��I�c�X�a�P8'�儘oa���U��m��Z�z�aO6���z9Y�y�=t��7������ ��79��x�Ƶc�DmM��GaK_|�w~�s�'����ݺEU%44��������� �`f���:Y0�hB��Z�e)&i(*��)�%(I�&4oCD��#YPёHX�ߤ�5�":@��$�AML��D`c�R`���C� �{prJ0�����	d�bҜ�ul{4)��`t&��1e\�LKj3��f-�e��
���h����b`��)����� ��@�Ab
�ZXj!��M�d���<�@�,����O�� -�כ*�,TV���NSH�ձ�tz�$�[�.V+���,�p�)�n;��-��)��F�X�4N��!����v`�A�k;	ڞH8���;l���&�ʶ��ͻ�zj}q��a��˧u��8�:�(��eȋI�ٺQ�9��,�?�D�?t0aE/m��A���v��p��k.��x��*c�������Vɣ�|��m����)���k+El6��'&Sf��������q�zc�e26�.��K�%��M��7U	�l�M�p�e&�� ]EP��zu]�9ٵ��+��F{]_k��� .ǐ�9���γ�z�2gluA�&
.Y����$�A�y&��]�&�8��=�1�[�.;3��rFq���a�ה���p���ΛxwXݞ1�@�*ۧ�B�.���o>��]�1�GO]5A�Iw�"sŀ���V�^����$�6�l޽��}�*Mx[*���m��.,*�sqV�|�O�,r�H��UP��;%�ZH��J��l�Uj2t���p�ܯ&�vj�K�)��o���{)�OA�N���8V6�H1��ո�7OZy��i׏W�g�R��p�A֝�q�� ��p�N�h�n`P{M=��|��𝒧WK�u�q��&����.L���^��5ع���n��.�V�[v)]�ε�'qpJ;�8-PJ��HMM=Z�j��ĥ4��s��&Q�B����ض!�(lServPt<-��Z#6�
��Δ�9x���y����0n]I��d+n9�۰g�]sY䱱038��[��ojdUj-���;Xwl�F�m��	Rq��<�J�zK��4�T���"����A�ԫ#�y���̫&�S�r�V�͕�%Q��T��;�t��K���n�H�g��v�\�J��q�)r�t9$�5AN�tU�:�4�����0���W!/�����ܪ;liX���e��L��Hs�pΣGh�����;�ݳk`q��v�\�f�Z7�ݽk[���^���!��@�C��b��_P����}W�P����@�@�5*��w��`D����Gݶ�5ˌt�p�F�͞��j�`�dJxh۶%��D���U����1�"��p��۬+�-�vr�Ƚ`�zܞ�u62�3V(�gl������g�^:^4���r�����;5ts�pqZܯ:�a�iX ��vLF��u�]�H��
�,i��$]o!�U��c���v�d�8z��h:�-�E����C�b���������޲s5�y�zN%Vݺ�I��R󋶮ޘܛ\u��ɐ�-�T�+�fX�K�iڵa.�U �D�~���R���{�)JP���}�\��B�6�����z"h����۽�k|�)O���P)J���=JR�g���)JR{�����D)O�T� �����������vv}^K�ԥ)�}���� ���}��pz�۹u���;�3����LK5PM�3��s��)P�>��qJR�߽��R���{�)B��y���)N�!���\����T��-�w��)@~�߸qJR�߼��R�����L�AT��}�c߆�r�V+wFZ���S��N�/NG������q�r�vj�%�|�g6�s��{(����j�o�ԥ)���ÊR�>���pz��>Ͻ�_��VWwf �YG\ļ4�%ESX�����X�%I�8�dD��`c�л�F���C�g��j�u%�Z������"R�����TVEM]�
��>[�0gwp��V w�&hVJ���`�Ӥ��;39��Y�%���7�J�9����yt��Q�D�EQQ-OUQY�%�����~ԯ P�M���Y�{u��.��0`�����s�B��u���p�l<�ռ�bke��Y��{����>��c+(�M5��jX���l���wg���;�[X�K��If�	���jbj� P�M��0-՘Z���U�:���k�=$SLET��0�Y��݆�g{�wvkT�р(�S`{��J�������f������ٻitX˯�G�M����I]����VȉLrӻ����� ��_}� ������l��$Z���;�`z�e��'L$�.�ڕ�Zأ+���Νɵ���q*Wx4�ȝZ������p���/-Y�}�J-���[䱰􍬪�y�
j��������ݝ��JQ`-�X��ڦ�����H��)���j�-=�>��	ޓkJ��T�tX����(��ۻ�&դ�w��_�����c`�l�0�s�4<;�0���2�a�xhS�EO�|IW�$�����w�~;�D��\n�5m�z=�lgf�ggn�]���'zM�����lN����iؕ*7��Ëtgp���n�kvg����0��;�����������Yl?[EӻWm�N��� ���vg�=�6�ca�DM8EL�TT�`G���q���;�� ���`I�7O�UA��cv��:T�k K�c`�j�wq-՘����4����WNӰI�h��W��&����S`��%䱰}k*�i���$*�l�V`��3��{�����l��S`E�7��-�ecAMMA�n����4A� ����[���gu۰\��q����.v^�WA�.�.�u�ܜ��wow��}�3;���Ӭ�<�����C�Z*��lv6��s�Ʒm�Ơ*^%U[<T��n���s�8�0�nMv4\�El:�Nt�%!vwa���펤8������.�tn�Jcm�nv.̼LG�X(˗/$���Y9#f��l���"e����������}��*v0�%�L8�خ:�ҹ�	�RΜJ����Q�/h˾���[��޹RN�RO�K��K�c`�j�wfyj���3)U۶]�M�I��;�!�z��`Ӧ�_�Y�����-�*��:V�*f��=�6�՘;�����[�p�$WWr�����ݫ��~�ON��}Jl�V����6�ca�DUS1U�Mf�y)�?��ᛖ�q��l�0�CP3C�1QC��,z�]��a�v���n��H�<Ὃ�ہ��Q�`���N��I&�	ޙ�� ��6����,��EW�ҫff��Y��uW��k�@�؀v*��%�>w}��([�`/��g;���;@-��uQ4�EPHUT����>�%6UF�2��'U�&��`�U5���JlIZ0G�M�1��\�n���R��l��i�M��IZ0��Ӏ$�f�y)�5z�������e��7k�p�=���LF�ٍ�/Y���F��־�{�__U��[7"DEMـz=�l�՘��ݝ�Rd4��%Y����ݫ����79���ٝ��ot�wu�z=�m�ݪ����Ի���m+n�4�@��"�:���դ#A#J0�J� @4�@�
!�D�HRX ~S���D��O��7@���cv���4�Z��vgvc�F����7۫09١����ӽ�`&������������ �{T�;�;��u^�y)�1j�h�U�?�)/�n��R��!Z� �c��rt��%2cg�Z8�#(��eCs�c��5PHUT�R��>�%6-K�ٟ@����$�R�ݶ;L)�Z{�}Jmݝ�Z�6����7۫3�������.�斈��&f�jfj�����v6����gvc��Y�}Jl>�QTҪ��B��yZ�����>��y��k��.
|�`x*v��@�>����?66����S�5m�����������Ա�G�M������.:f&�6��R��ܵpn݋�����vq���Ą�6Q;V�[�w.]������ĥ������3u,l��Sn�}��0h��Ye�M5V�X�I��W�����>�՘���ٝ��g������VS�6����:�,����,{�����R2�'M�ajƚ��>�՘����Ա�G�M���򔭴��0���{�}~�`���-�G�M����1���ۙ�ɹ��~��a�b`n�ь�k�����c6�ݱ	�X�^z�{ u�;bG���Bss[�m��A�.ע�ݹ�
���V�U�ic���V�:�H4��U��MT�wm8p���:b�T��pa��^Nv/X�MѮ Kڝ�nq�2nx;l�Dmz���u؜�O+�p)����L"�pv�5��?t�s	c^��Uv�]�:���Z	^O���{��߽���?�2�~S��#�m�v�v�m��]p]6����v(ܽ��\&����G����_��,*m4�m���M� ��<�������E�����*��N�����{U^<;<;0n����S`f�g�@����:(*Hj�&*���K� �<��W�{�C@=� ���Ի���m+n
���ݾ��l�V� �j�wff��ـ'I��$�j������F ���UX�՘еM�̽�o��sEg�z�Nv�ݮ���#�s�뮪Q{��7����p
�ɫ���o��n��PMT�O�`��`o�V`B�6��d�����we'M�`�m7�w���?b	$�XJ���5��xi�4�B�T�U2��
w1���L1:�[s�Mcg]l7� ���m  �>G��Y1������ o�U�����l�V�lv��-=�>��`:d4���3�4��`-K� �eLBb"����i��m`U��C@;��UUR��~x���]�)]�[l�w3 o�U�;��o�U�
5)�1j�`�~?H����2˺��C�q@�<ܷc'e2ฝ�L�;a����L��w{�;:���x�!� ���j]��JlZ�7㳎���.�<�\DS�S1U�Mf -J�Z�6 -J��ufs43�� �(:�^	�j��&�l�wceW����a�u�`�Zt,�A�Ra���L�WFK��QM���|�-f�Ű2:7s��,��a�o�q�u���u����{��s�{!<9�B�H��l,�)2�L����<N�8Y�F-8�Y��&&x��
�qޓ�Y��P���O<4jf�3a�ӑ��1>Q���]pځ�j����U:O���Û�ۡ��ќ�`o2HH
�	���ƃ�8��ь�����vf4���g ��0�EzWԎ�M !蘊����} t>�	�
J�b>��1P: p]>���{ڂ��:Pht('hv /Ⱦ}߾w�U{�{����D��*�؛Wkp�*��:G�}��t	}"�7�d4��;����Ӥ�i��UUK���!��x�z��U,��IYun��E҅s��Ͷ��fj'��j���\�����V�w���^c��N���i�/�X�%��R�gc�$�0)������M;N�o ��6�t� �����UW��H�%���hWm<� Z�Xn��9��vh]�`|�v6�J%�g�l�V����G��7J���ʺ�߾��RX dI�eU�'H��~�Wo��Vݍ�{�R� gv�ԭ�jU`}��0w�������a���m��z�[���'h5�.����A�D����n��{����W��4�1UV�u�R���X��:G�J�"AN�[��ڻ[��-J��uf �R�7U�g�	�;��'�:-����n�/�X���!��x�Wъ�M��WMӹ���wn��6�u�R���Y�}�+�V;e��M"�����ٝ�gh���.�BJl��ݪ�*��~��@��e�[ro	���g�.��,#�쑣�|t�3�:�:#n��1���{�pm��Ľ��\,��3�p;��ٷn{^��Gc�hM�E�Y�����h9��q�J�ڲ��s�Z�^g�
n�=��Nw[f�l��wh�[�C2\�m��c"���gJ�t�ն���M(����h
��W����|n����Kq�����P	���� ~��DC���f�u�f�l��5��#�ֱ�ǡ-�r3Х����B�֗�|��pk,��U~�O3����MI,�����#�>�t�\�`��
R�Zv~I�m��wMҪ�$� �t�`IU������4E=13QT�`IU��{m~���V��ـuw[�iՠ��ڻm�~��h�<}U~$��]��T�:Un��hKp�	$xU[�t� �G�o�� �����;�X�wi2�nK�^�9^#v9T���^���Og��^n]�3��]Q�:O�`�m7�o��tI�wd+�� �G�Ou_F+m66�]7cOv���|�^��R�u$�IA�b��+���uY�^�몯~����M�>�ܫ��I��Zo ߻�� $�X;1�{V`IU�b�J�!��պJ��������䉁�{��w&���ݵ�}��t���E��[o ߽�tI�{�րI#�7�>���Ut/��2h������3� m8yx���sk�۰��צ	t�WǞ��޵�%mK&i�I#�7�t��	$y_���7@��rӫAV'I�i�}��h�<~H���=޻�D��*�U3�`IU��n��障gfl��wfvN����f�����1*���WG�O�`�m7�}���"�7�vC@��I#�'���R��lL)�v���"��U�{�4wG�o������&;h����uLƊ�d)�6�����#u:��,�i����fR,)6��6��7�t��	��{��W�a���:7�l��b��*�Z`������ݙ��{V`ҔX����>�*�g�l�V��=���J,���jX� �UXy�����T�UA5Y��������ڻ��n���{vmd��ת�� ����M/�M��� �t�Z��US�e`{�n�/�,d��Y`�;n���t�ƙ�KP�<cC��R�n��N"��)ӊ�;��s�~;����w�*_�*�v&����'t��>�t�G��gvf��wc`���5T5PL�ESX{ufs3�û�ѽ�`}�ݍ�-�m|���3@rM�3155331UDMfѽ�`g�Z0������ ��Wr�v�I6��6������C@[����۫09����ۧ{��>𻩢��&*"fb���y+k�ڗ}�_��k�u�s몸���4�W�bSJ4 BЦ�P�$�P����_o�%q��C��w8|���o�m��qЛ��U��S���I�Qu��v�q�)-�l��t�3��"u<^}L��9�:�7M���:çnѶQ��,Mω��{9o96ݱ�m��<jc!��Y��ݸ�VKl�<f��3���p�bvZ�r	���ň1��p��5ʷ% �N���{=Ul8�m��,v�Aq`�{g�[\ڪ����C-����y����gǲv�:=077F�s��)���Ε�c���3���ŷ�IAQI����.&�y�"�&�i��K0��,�V�n�k�2}DE50�Q0�D�Uf�$����u�%?����7O���n�WK���m1'x��C@�镀}���$X���"��ҫ�bi���e`{�n��$�Ý�݆��u��&�y���J���>�t��,}�!�wt��>��)_�V]&�-R�Jؚ��F�.�u��l��ri|X�����xկ�w���9�Y4��[4�h\�`�2wL��wvf�hԻ0)�悢�����i5�o9W^}�>��ʣ "�~CY���Y������IM�|-T��!�X�%n�a�wt��=��U]�;�l����>@ҡCM@�2EIUM`�{۫0�%6-V��wU���@�Yn���n���@>�<��?ܻ8��[Xn�� ��� �$[e�pݸ�6`�ֻu�99<q��ۦ�����Y8����i^��N�����.�X�-�V����G��W�#E-.�Uӱ4�[��;�V~�=��tzG�l�!�~�D�K�n��+C�� ��Y�$�Ηa���a݇n��J�a�2�$�I�P�#�=P����uuW�}��$���i4�6$�@�����L��;�V��7@���%X햒M;��M�:d4�]�2��t� ����n��/ʕ�Uj�L���qy]�tK�2b��7{n��9z�$�;j:����x���&��%v�a�N镀w���E%�:d4�R�.���H�X�T��ufs;C����>��� ��u�zK�D�t�[��7m��R^���gwv���[X���5	X�j�_�N��v��~�����2wN��}�|Q:�1e�C��J��|��׀zz��
t��ؚI-� ��m`s�;3;>����=�`f�6�]w+��wWh�t2�I��
��rOcp��n�j!���=h�;`G&�.�ť�T554�TU5���Y�|�(�3RX��߿~�;�e`��v�I��j�:�ot����;���@}�ݍ�y.��7�ՙ��{f�UKD��ECL�ME��ov6�궰fffs}�Y�o�TXxZ��������"���ݚ=˱��?�@�.��UUUF�I��}�JEt���E����>��7@�.��oޓkB��~�ʺ^z�ؼ��l�"/v:���&�	�2'C!�����l�L�B�N��	����V����۪�9�`f{�o0�b"ۻI�-�KM]ٛ��*���=C÷^!�2����M�d;}&��M�������7����a)�F�a?���Ww��׻�� �`6����!m�$�jP֛�& d+�fj��l��K���Wnt�R���un�9���h�'�\^g��ی	��ڝ�
�l�rk)g6�B�g9�Kω��ʹ�f�"�L�seE�u�ѹziJ6
.\�l�R�vg�Y"��l�P]vd��u�B��=��{F��W�v�c�����u�4aɢƵe��:�4���d���-�ɉ���m�4�P����'�y��nctl��؄�.Ma��%�-�ͤ�f�s��(�$���gv]Tv$��Oiy�\�d����
�t��]������V�u���p ��L��a�;����x�
4��\`|�܇݊��%�;uq�㣑ظ(���95��������;k�8uaFV���1u��gm��[��^۱c�v7%*E���3p99Ж���"�k̦+{N�k4�nv��Z�"�8iDݴ6N8{kl��;-]Е���ɻ9��6���)b���F.[7"��#T���ܣ{.�3P�2��ۄ�tʁP����[3؈��C�R��=V&ES=�/I��=m�̬���X�t�6�Y'�';�m�v:��ٕ�z�'9M�q�q�:���ĒոθZ��I����]�����M���u^�qX�6�������g�4=���i�<�&�ԧ8�'�9��d̤����kṈĄ���4�SҡQs܍����:2)*���
����ɠH�]���P�k�U�^rĄ.ic]�ش��L���I�ю<�F�؊���8s�]�q��5;v@�)�M=�0i��m�H�k�qO[.�	��i6[j�[W\iY-�ӵ&Ú��6 4��Q*�O[�M*��2QY]�.������zl���z�Q��d��ggb}��W=�]s��m�[I��dG�� �	@��T=�6�l�誗vZ�s%s�^P�b�(2�H�Xm���m�bBڵt�b�r@(��jz�W���q�َ7��;��:�cq'Fwj�=5�>|�&"�ٴQv��!�b��'�:�@��N�\�=QT�������`��{�����o���W�נ�=�]��l��á�ͭ��-�wU�x�k�l��xz�5��膂��sx���4n�����I�5ćr�!�H�+`�scv�&���B-������e�=�c�S��]k�WZ�^��TȎ6��sl�u�e��97/nn�C���m'��tV��[��R��Ů#�p�n�'U�d^6�bu"u���������uo�v�����*�X�m�;�Kx�n9�nڞ�㛱e�v�or����{��2�Ӣ��M���@=�����!�|�[s��3<��� �w5�EL4��5I�-��7�L���镀}��n��]"��vx�`GT��5A5339f�u����՘��}䱰��B�I�Sb�V�:�����t�yIx��6�
�S�e`�Wt�I���m)���(�3�K [�����՘{�~܇���c������V;v����l�6m���ݲ�������:����F���L�i	�xӿ���	�2��O)/ 7�H���&+V4�	�2��! ��!Ґ|!�Ùy�~�0�R�>�X����4�t��R�@6��t���R^Q�zM� ��x�r�U�!������=�%�����zG����t�q%bv��Et��ۼ~��Z�ޑ�}{�K�>��F$�E�C���T ��tu��Ng��Q{c�n엶P 8�;=l�vɭH��j�I$��ޑ���7@��Q�����{���w2�SO4��Q5V����fgwf�7g�,��|`�#��@OH�i6���i'�����U�{Ϯ�h`��d�&*%
��MH����z����*��:n��Vt��V�m۴&��W��~����|`�uX}�Y�{ҔXh�:WT�jƒI	��H���W��L�=�%��솁%H_���uj��#[�a9��mi�_3��9C� ���EՖܼ���i��Tշw��V�m��۠{ҔX��C�36 {�U��6�	��)�5m��)/+�~�}��zG�}�t�q��4ա]t�QU{�р�U`���}�����7g�,�`�x��A����g,����#w��y.�ޔ��3�3�8�5�3X�E � ���r3Q8ٌ�;Q���@�|*vf���ٝ��� N&ޘy��	�)�x�wM�=�%��L��{�<6�w���￈������ssj�;��)�����V�{%mi�vWq�1�� kG����pW!�ն���i'�ܿ�� ߽2�H���M�>�Δ���nݷm'x}�h�w�ggh��=�]�ޔ��7��ҿԘ�j� o0�{��>��f����Ｍ��L�*��[,��>����]/ ����>� ��TJ���4Rc{�{Ӫ,�Jрy*�=�%�;����U_=���B����,Q8�M��\��E�dĠl�ݐݜ�W��H ��nZ��s۬��� �����cN\ۅ��b�RԷ����xa{uŬ�@7+��G9�0vaw�ֈ`V�[W�8�����!ܹ'��up�U] pQ��y�;��j�`�&�]ɓiR�rg�U�S Y���M�p&tkn�l;Uaʌ\g��&W^���'3�9e�+��r]4Ҋ�}fu�Um�����t`�77� �5�:ڵ�	�	������3�Z0�%V�䳝���g��]6�:%��*%�����0�%W����f�+���������9��j���*J���7w�0yt�=��߽&V }���E�]�v]$�,�?}��^��� ��<����}�(um�ݻn�n���!�UN� ��&����	:TE�A{:���#n�vB����B��D�*֏+\��#��ݤص1�5uHv��V'�hޒ�{�f��Tv@{������uD�r����{�ΪJ�P�V+�zj��%h������h���C)1�=�=�^��d4�tx��7@�t�T�eX�7m'x߫��w_�]V�� ��TX	��UĆ*(j����4�H�����ws���d4�W����۠wh�i�sIng$lm�")y��uv�Xsκ��<gC���W�7N�hv��=�I���0��!UZ�H�	���#j�i���MV`ݤ_<A�w_��V��7J��>�Δ���m;n�l�>����W~}��v<@���(&jHeb�?c�X:믷�_����� ���uHv��I+�4����J�{�f�m"ã���0NOqD�S$Q UUX��������F��d4�H����5Ht��f&�j:��Sۗ\�ɱh^Cvl�۱�68�[�t;n�;���AcE*n�{�{��}�V� ��U�����y,�������	x&���&�g3��������m"��wwfw����L�KJ���{Z�� ��&�w8`}>���A����]�n�.����I{�f���`}�����w��pgw�*Ih�V�r���>�������.��N'#���;��%MU*������t�x�I7@��슬MSj�U���[v�O]�z-�Dhp�Q�S��,ti-�P��f���um�ݻm�ـ{Ӧր}ܪ���,vw|��E�{E�e�J��j��yZ�tx�I7@�s��-X����������b�G�i�$	��V�f��E����`�UXI��6X�J�m=�+�{�0�vC >Z�Ù٣V�}�w��*��p�i���,�j��9ٝ؏r�5ovuW�{��U迤� ��P����F @JQP�@�����j-��Ǳ�n���sݺ�ڜksl��Ld��7k�J�.'Wgۭ{�f�#�)�.ó���&wM��F��k=i̳��]�p{%jץ鉍��ɭ��p�������������u�X҄��9��;g�k��a��î��d��6�;�t�/!���+x{T��u'`��a��糎L�n��.CkWn�y�J+�Y31gF����~^�|~7Y�uj'Y4���,�p�qJݽF(^[>N��b�;B8�[D�$i8���6 or��� �m"��j���%H��n��`��o �zM������UŁ�˱���V�-P�dUT�Uj�"�����6�����I��Y*~mջm�V�M� �N�Z�txw����p��u�����]���4����I����vC@�w+m��b��v��ll��d1m��AC���ksc�݇B�a{'[�O6�)���t����;�&�w8`I� ��<�QRU�`U��*i�o����~��'̅O� �A9��L��a4���IU���9ٝݚ ���CUD��55MSX�W� }���7@��e`�\W)�(j��fg,����7|�`�V���Y� y�����(�	��j��%�33;�������-U`s;:�{�����1!�#���NN��Fֹ���fp�7,�,N��vwCƺ��f�س���_|����m� >Z����-������T�U5US54������G�{�M�=�X���$���7qG���}�׀{�}�8jK�[MTA����B,Ѣ ���7"��ΰ��l� �p
�H������Y� �E�e��fX��+Vcj4�FXa$�F$Q6`3�j�����ĞFĊdN���s��qk}�p�{��r(�0#�*�0��0h�,�f
������c ����& ���3:����F��kRF���[3i�Gz�0�&�$�>u���:��$gd�|���M!n5��T���LŭDERĔ%��7�̜0�8rJ5���q��[٬�ԓ}@.������u��8��� �!IX�ۚ�M;�I���N�m��-�ޤ�7��؈E��I�Տ1�t9�p&��oJm$��M�$�j�B5�8��4����l0̰,̬�0#4	��kznY��a�����N� ���d` "x1�ԡ�:�d��N�,�O�0#�9�>(Et�|'j�Ѥ|C�1�ā;E��> ��*������Eң��{� ���qp�Q짪���&*`	��b7{�0����$���#�>U�e������=�V�;��w|� {{����Y��%��1!��6ʻj����ۺ싄�ۦ�V+F᭻MsxXg�lj��nӻu�{��k@>� �I7@�t��;ĸ�$SUal۴����� ��ݘ�����X�80ktw�6lM���twL���M� ��x{��+wm2ت�Z�i� ���m`}�V� �R�d�Ì��D�	(��3�*v�u�����$�����e�;�'��h��*�>�%��U����������'�B���Ą�0�����[����28ɋ˙�d^՜5�9�3�j:������{�ED���ݟ �{���|�`Z���솁:���W�:.�wzM����U���[h�6<��;;4A˚��&� �Z�jk0����vу7�����t��t:xʷj�Ӹ��k�rY� �{��ߵ,����S+ ��q\n�b�һm$����jY�{�[X-�F��=y��٢��DVX؆G�o72�e��Y�k����w��:�'n#N5�K��Ei��3Y)����WU��lA�\5G�:�D$RU{n��8�]�c���T\��ہ�d{=���9��H���q��m�v}��λ+���*>x�Q/7�ñv`6��!=��䶻*{\mڻ<Xd-Ѱ�x�ݼMY����<5N�s�-�0�q��Q�6��8���n"�\-�߿{�{����s�������NGrl�gqq]\�QHC�^x��Ƙ��gk3���w;�U���l��X��tzLk�h�g�67�lI��DEQDU��BOtzL��N�h�H�w���wwf�wwh��UMSQ3UTT�X\�����vh����w���;����(\����;�8UU%���=ޓtzL��;!�IJ�JM)R�v�ws ���s�$������ ���h~�`+�D��ue�t�<��N\��G	n��9��E��]��%
�oa�E�ut�]�AV[�����wL��ݐ�y)�g|�^]ـ.sQ�M�w��;��|q���B`%G�K0&'D�#>��:�]@aF%�I�3�Ц��p�E�Wꪤz�r�;�M�'t��=�\W�Z��Wm���K� �M����A��+ �Ӳ�WG�`�M���vx�r���k�yZ0f�yE�}�����.�U�-��>��X;ﷳ�����`}�՘��6!�RI��p��8��nخݓ]�\�(��N��n]���1�{;K⬫���]���?/���߳ �{T�|�c�����h{T̳!�1RJ�Y����E�}��ޓ+ ��M�?Pt�|�&���+v�wm�+�������%x>���HQDBئ��y��U�{�������h.
+wr��t�.��q`�,lcڦÝ��٣��� \.,MX�ei�4�`�M���T]?���wf �����w}�8�&Z��I��ݭѶ��GYz��y ��ر<vν�g��n�d������rY�mhc���~/���{!;��{�V=:mh��w�6��6"�k ��7@�镀ON�Z�j���>�GAD�2CD�I15�j�lzI��K�E�zt���?6�ci�M�4� �N�Z�tX�����+�4���c5�f�5��V�a�L��6��\�%�L��栙����e��,�w>B.��c���o���2�%I4L�$�U� �ڦ���Y�}�X� �v���߿�?�~z�r~ ��v���;��uɜ��:��97k�4���Α�rI�"�~~/���>��,�K�ݾ��j�N��*?�O�XЩ����s��Ic`G�M��f&f�9�TIH4L�12�������@}����m����/�+��M�h_�,wI���zI�����&���[M`�M�>�8`�M���ߵʃHĐ0��=��G��o3bL�����svRz��`X����'͔�{�q�Hݳ��v��C�Ў3��Cq�I�2��=�!��6��^�`4U��y�φ���+�7N�۳�i��˴:�E΁2,Q�2�'g�bA"K���oX�a κ�|�����1��.��RvN��c�Ɗ���(���s���NJTE��ƌ�u�nxZ��Z��V$^|�����{�{�?t�|k`]#�pjΈ�EȽr�l4ÜT jw�ޝ�qv@ք�[�v��.�U�Z~�;�K�'��Z����n�w�@�݌m;I�M7xzI��z��`�&�yIy�A˦e�J��������l �]V���tG�{��[������RTļ�LT��UV����˻��=�`o�M� ��<��)Q,O�Yn�6�{�}�%��k@=� �t��}:�}���'']��R^Ӣs�;,j���ȃ��w`�ם��dK5I��&�$̽v���k@=� �t��}�%��\W�wK�J��{Z�ty���Uk3�Ӵ3:w�k6W٘ޔ���jX����#_��0lWm7�}�M�>�,�wfv�Ի��uuX���T4��uj�6���)/ ��鵠�G�o�&��Z��v1��[n�n���X��j�>If��(�9���&��;��p�xmmlf�n
l%������n��v��z�J�嶯��t�&T��o�7WU��$� �ҔX��c`)_F&���+i+.�x�$��)/ ���k@=� �u�A?�e�UEMV`zR��-X�'vx���K;G�c ��`����H����l�'ׅ,���� 0�C��S���a��}�Vj��iL�RQM MUCU�Ѿ�� 7WU��-Y�}�%����q�wt�Ƅ�v�ր{� W�:f�����{�&ր{�r�B�Uv�W��^�b��HJ��^qv���v㊷Q�p:оڵ>F�Ր��yj��JQ`{�3> {ڪ��3y
jJ�!�Z&�f� �Ҕ_3�������`{�Vg333D�����jj$��*j���wv6 {ڪ��������>��|"J�;IP��o+@=�U`{�V`zR�ކw`vf�`��@��B�{��U߆�߷kz���+i+.�xޝ7@��K�=�I���G�N��wM�%uE���(�c]On�sd��*/u&��<�=��҉e�u���v���*cM�����{�k@=�+��>��AH�41Հ�wE���jX��j��-Y�}�J-�����,�V4&�I�h���zt��)/ ��&ր}TN��䓶��SU`}�0�)E��V6<F���=��_��!�]Z�M��@��K�=����{UX�0����:t��0��J�q�Z(
����#����v��Ǽ�.p���I<�����$�PE.(\�6:�g��+� r�M����ݣ�X�X�tX����Tu�E�o�-�������䩨��l�g8z	�Ѝo|zc�8��ʳ̜Öh��b��9������-F�GDt�r,�v�dD�E�����jmN�g'"�t���Pp!�ц!$�=�Zw�7L�Qks�R.��M�>_��uX�.!%=�\MK�Nh=�h��a���A6�Ak��,�BQ�b�=wҹ�^s�S6o{�f��,��É��Q<�9����e��oO��k,C��{�=3�{]�U���fj�F6N]�fu�Gt�/��4������y&M4�;�Yk���VD�AQ(��鋩��6Y�N��;�$��G��w�]��z0�jL�:�=�  �` &�0HH���Sv�0 ������-�s�]��]+�\lt��{]ڻw9��f�L<Y���2�ű�.���H]��.n�"N�u=���dM��[m��NݳM��\j�rm�ŉ�m�x�vڬ�q��8���i9�=���n�,q��%m��Y_m���fx���S�3���la�6ނX^6�gs�%��l�!0�a��2p�;rK˳E�r�&4�{�Bҡ�=H�d�f��r���R��Y��7*�x���rG����<�����
�ǀ4�jZȮ��-vN:y��G��l�=^�m��b�8GE�}��[��Nҭ��V�:c&�A��-���WZۭ�z1���%�����pt[�mn��v��my���gr�����H=Z$�Q�Rů\�:oer�<-/9�%pDm�He�	�l��m����u��Ө����Q�=t���p��G=��<S�m����UU!��rA��W��2����,�e��vj[�e1ɵ�l�'ivz�*rU�vQ<�0�hE���g9��n���y���t�	d�$�s�m�v��Pi��0��[�z���<V���@�^F�!6�Ƶ�qŐ�rshw#e��f\�{H�ulH��ъ�XR6�g�=�{F�v�p%UlcS���T�N0��c�i�9Z,�$�؜ʤH�Ŵmr,&׋唲\h(#-X�%�/*Zmm���2��˄�H��8ol����,��A/��Xخ�
.��ƥ\�Y.��ݤ��O%�k&��pvx�b��3tl�'YxV��l�s*�F�mG'*h���!5J��Uh�cu�=7]V*���K���A:.j�K�]��	D���wH�G$Yɸ���ӻ�[�)��͍$����:9�t�f�EV���*�E8h���X'd{�n.u���WW^��6N��VZ.3t'X��N6��EՖ��-vs��v�z�&�oy����@>��^�N�_E��E:=Saӱ|OV�GBhUS%T`$R\�S�>��"tv�����T:��(��ޝ�'��w$��+�ң��p�3�ݛ���z���\n�:g%=���p�ش��:�^�V��.�:u��1�����y��_^Rm�ݛb�����a�M�[D(n:m�)��
v�y:唝n�n��ö��)�zr8a��'m�N�3�ͮ3h��V�7z#vq�;aa�˻v�D�g�:�x�r���iH�J���P��m��2k���{�������Ƨ��<��tp�^],�FI��V�n*���A�Zs��]i��C����������Vyj�Ѿ���tX���%T����%i<� ��<}:n�����{�k@�����;iR��}��t����t�Z�tx��]�O�Yn�1��@��K�=�I���G���Ӧ�.~m�M�1Q`{�K �vh�]X��f���<��ھ����eأ#r
Ԍ9�V��gv=�9enޣ�ە�bc��s�~~�||�ӫ)U�V�m'��t�xޝ7@�Ҕs;3�d�.��9ɺe檢()��7��u����^
 {(�Ҟ��$�i%T�I.�ݟ������. {���盛Tn����Zm'��R^ﻦր{���7@;��6m�V�n�}�6������}�%�׫�IU'j�4	+I�h�������=�`{�Ս�kn��(�1�s��=�V8�g��r�/l�
�c��[����a�	'u_}X�u;��#�~��-Y�|�(�=������@(K���#���.Ӡ�1��@�)/ ��&ց����M�=)��M�ݼ�߾���~�v���_4��T*_� ��S%�..�Q����w@��K�;����N�AM"�sX��Х.�w�f�Øh��0�rn�i*�"B�����u%��Ix�L������\��wVWWY�>l��%��:��j-��;�\�{X����3�u�>;�;��D����q�߉���t���,�$� ��T�!��[n�n�t�������얗M���� �JQl���Ԧe�j&f�bbf*n�cuM��If���������@�J�1�~�N�I�M`jK0���U��;|���^]���*��K����>�ƴ|7ve�+ot���wL�����I7@�3��}��^���\!�&/�^�9;�I��/M�掜Ɍ�͸k�x�ǅ
ܫE�^2.�ۼ�&C@�� �I7@�)/ �_
;ub
��mn_tY�vywv`��۪р�YL��A-R�UM���� �JQg3�F���.O�{�RTc�.�U��{��_��]�`j]|`�l9�˻�����M�nմƛ���!�u�E�}�M�>�K�5��S�8;�*���/7d�q��SmU���W����\��`z�V:Wq�9=dYC��ˍh����q��W�Mm�ű�q�m���u�7L3^��&�;���D��{Y��PG�G��Aùn�v�s��HY������e⻙��7Mc�[*�c���e��.����[p�����(:����v�Yx�	Zϋ]R�fe��M�))��#nYwv��I&�,#��pP"a���ܷ]�rv��y��ټ�ܻV�˳��u�@�����X���$����J�J��$�x�$�褼��!�t�}�?[�m*V4��>�&�E%�� ��W����ZDU �T��T�f��=������%��J�)���X�v�x�L��wtx�I��Ix|z�Q۫⭃n�����jK0���+F���w������M���1��ܛ1�=��T���`��c"-թ{{WKέ�Z�"��]ݘ�R�ڕ� 7z<�⤨�!�]Z�M��@�)/>6!D� Q0�Fj()U�����z��u\ٟ:G�{����ʀ�6ݫi�7x�L��wtx�I��Ix���UI�Iڵi;Y��wtx�I��Ix{�C@�蝴~N�n�!����7@�)/ �t�hwG�O���ZQj�*ai*m��5��6���>�9մ�e���,Y]��Ƚ�c���?Yn�6�{�}��t��� ��n��$�[I1��4��ۼV�Fs�DK��\�� �JQ`/�\v����`۶� ����&����%*v=�j|3  )*��� H&�Q���$ZQ�D�z"�+��7�߳�}��� ���J��Ҧ��xI&�E%�:d4���>���Ch��V���@�)/ ��!��Ӥ����ի�PX�m�*)�۶�ɮ�^óEշLm��=m���aq�C{5�m+vƛ��L��wtxN�t���x$�/�ݤҵm��a��u]�I��Ixw>0r/��h����cI�I&�E%�$�hwG�}ǿJ��t4*m&�C��=����� 7uU�3;�oC3�ӳ����;��`�Ri���)�����m`$�hwG�t�n���������n�f�d"f�!��j���N��#�a�:br����������=�n-`��b.4�AUQ�� $��I,�>���3���� 7��:e��`������I��$XNr^�wtx�⤨�!�]Z�J�{�}rE�t�%�wG�t�7@=���m؆�Jݻ���:s�����:t��I o�Z��iX�&ۼyz_tXN�t�#�:s������Gv&���.�����.���m[mϳ��q�����W��0�j���h�8����m��o̄�N�KӪ�F��E��t�\�/���즀�A�������i�âwK*�v�[���*��Yێ^�B������)p*�n�m�UW�E�VvS���l���^W,��y�N���V	�fT�tc@=/4�ҋQF�ܱ��FY�pm�Uiv�%�QR�Z�_�o�t�}@aNl�6^0�B��nyʀ\��q�;>�I�y&vS��,rB��~o�f�$��մ�~���@(K��ڝ������-Ҧ�ot�H��� ��<�I�AIHM[VU��aU6��� =�Ug3;D.]ـz7��`��J4��Eݴ6�q��{��:t��}~�`H����#T��.�4[M�:M�+�� �E��G�zur�hUm!�Nյdq�r-��^��s�Pͻp[^���"wO61���ZV���� �E��G�t�7@;�'�bnջe��*��{���H��"A24 t� 'Z1d ��Q�_f��3H%�Հ��Y�}Jo�� P����_�4&���x�- �� �}~�`�-�/�wn�7v�Jˊ���vf�v��ѽ�`j�j� ��<�K�Wi�4*mZ{�}~�X�uN {ڪ��� �vf�(���M�ΰ�6͞7ku�nbVA��Ѓ�k//�3��kuד�f��������Uv,�0�[U6�K� =�U`-�Y�}Jl��F�X�;w�1h����&�G��zV������U25S4�TT�X|�`G�y��_�m���2�����'C��W��h�C��a�M:�,0>O˧�wӐc�@�����D�A��{H'g�jZ0��b:3F�<Ѧ+4�X�vtf�[֌�k5S� x��`o4�&�ʌ'f�f+�:֫M��:bF9;|���^t��I0��}Ax*u�`���O T0�.,�=�C�z| �!SbJ���i����0D8��9����<�Ut#��uj����� �.����*����޹?��v��[m`�9/@=�U`/��0��M����jnn�%�	�t�V9L<&6��<5e-ɱ��K���QmONq��Ro��}�|�ԫ�5{���O���`/��0��O;�c3�w�_ ��%�"�j�&���_y,�wfh�F�M�۪��-U`{��
"Z���T��@�� ��6�ӣ�:zL�<��SPMT�TET�s�.]�6 o.�V����sC43�8�3�sPkSK�P*T�v��]43���EwM��S=3P4���U53X�媬fe˻�Q��`j�Xٶ߯������-� "p��x���&h���x�"�0���[��t�mPg���|�ՙwN*�U�M������,�I����U{����t��[ot�H����˻ 7�U��R��gvwh��w8�4�15DUEUS`w.�l ��Vs3<Gr��F�M�j7TQ%4UEZc-fe��G�I�n���'I��.�K�~m��Mۻi�N�t�%6[� <�U���٬��4!�xh�<6�,� �1 �e\�rT��=ϷF��ݘ;[�4������$]hQ;Z��uݕ���c�<t��q��=�Gj�L��\��N��Am�%a�_�b>:��<᫅❛uMu/#�+P�m���� <����O.ӳ���6a2t�d��S��[���S�r�Yݹ{�����Fw�Wl&���/8Ԥ�.g��VǠ���Y�,��3�Ah2�]Xrf�v	�roy�w�����������jE��V��Q���� n�D�̠pǍǰ��T�2u���ݱ��vZs�	���	=�k@=:<Ot��\)LvU��wwm�OI�����7@;�<|�D�X��`�m7����t� �H��}� +�=�>r�j'n]��I'���`��=�V� ��V��ʆ!�V��N�{����d4ӣ�:t��}�e�hwN����E1n�.!yLH�h��l���-̶v�/=��<���iիM��Zm`:d4ӣ�5jY������ \.:������n�f��]Uy��o� ?A�~n�M�>�H��d4�2� _�wmSUSU`o�,�6<��������ƀw��x�:U�2����-��C����t���� <�U���f�s�)�l*�ӻ�����!����n�w�x��.Y`��m;�B�l�c1��֓��q�
&���3�W>G�ӝdr66	��ub�wN����4ӣ�7ږ`�*�vv�r�� ��z%�A����j���Գ9��ݢouX����-U|���}��EU4�0LMf �{���$���f�v v�`fX*��b��VE�?�hgvv|?'��???7�0l)N5M4LMQIU6������ 7�U��Գ �� '���J�:�mӻI�h�G�wt��u�E�}$�ZWW�g�3gn\��\�l���6����9�������,.���ɧg͢�M|wI�_�X�I����:�
	j��*�����6<��;��D������`o�,�wff�7�GQAU@�MMDS`{�v6 yj�}�f w�x�%ub��6�okC��;Do.�j��c�M���̙�ٝ���  �4��14#���iJZFQ�P������P4	f{�;:�<��օ� ���Q5U`o�,�9ٔ�t���� yj��S	�����y�X1��K���َ�0%�]����q6��:���!�h��v�$�@�� �t�h�G�w�M�	��SN�;M"�k �t�h�G�w�M�:�"�	�:�$����vۻK0�N� �jY�3�<B��ܺ��>��
&	y�v�ݫ���;�&�~�`N�gwh���`{��A/AUD��`Jlg�.�> �]V�R��D~dq%`c�_�.��էZ��ݜ��q�H������^�(�Ku�-mv�ڛ��l�<�UzΛ<�&x7[g<�t[AQ1�&;�zF�^\K�1������Z`�fD-����#���o9�b!�dc)Ju�F!Û�8"�E�ɘg��b6������N6W��Nl��nJV���fȔrn@�̩%PZ�&8ٸƣ��:� �uA�Gj\a����0!���T*���&�f8� � z�t^�֊��]�by�쪼]v��Zٺ�t�k��kvͮ`�n3Q�S��~?�����`���7ږ~;3�;� �{���:8����`j������0��W���-]ـz7�l�����ZТ^�U�i���7@��"�>��k@=� ��u���.Ղ��_�XӺmh���~;�tK�N��V���i��};�ր{���7@��"�>���T�ݗv���ݰN�p�����<;V��l=NrWKمÐ���v����vۻM�h���ޓt��,���鵠}���v/ɻ�����;�7}���IUZ��t���y��L���0��W���{��c�������"�k0F�M����0g`=�U`o�K0���:m�X�v��>�솀{ڪ�߼�`s;;G�{��Ztq=1MՍP�N���G�wޓt��,��`��ޖ�Q�C�D�AO5�Mr�mЛ��:�q����0{DxV{ .2�F���ޚ����zixih������0��M���d:��;�`{�x��)�Z�����l｜h�#�;�I�S��	F��������	"j���n�0+�=�|�=�qT,� �b��^��}h_�X=GT�]Rt7n�wv� ��U��� �<��s33���ݍ�yqPt��DT�T�DMU��$� �h��V������U��o!Lą5�8�;u��(Żp۬'Yr���uh"B՝'/]g��g�;q�����k�����o���=��^�}� ��M�$%7e݂d��6�� �����UH�~��$� >���gh���tOMI�,M1=yz�� ��M�����鵠� ��D�K4�UL�X;�3�^K:���~�*�Ͼ���؟� %�ifgN���ה�2�dq���F��$��+Ot��ޒmh���zI�����������
�k�89�۶+l�t���S�n��[ ��a3�$���u�n*�n��M�ޒmh���zI�ߪ��fgo��j��M�S�LQTUT��V�}� ��M������k@���h��&�؛�e��zI������zI��{��>�\�X�:,��Wi����<ޒmh���zI��u�v�Rn˻m�N�[ >���7ږ`G�M��O���l&�m��8��9kLS�k\њ�6o�Fz5�n�q�6~�#)*C�\Fm�8u)�q\�"R�dQ���`!��{�����
�, �#1�o3��05"L���w	�o��tI�ݰ/1��eR��2Foc���1h��!��
֍.�C��{�s�8��4�&�s
�j �['n�]t��M�d0f0��X���5�xw������s�n� ���kV�f���ctgD���I���m�k}o�4u�L)�r�]���q��T�tJ�� ��$���Hh� �C pƳ�Dk�d�ضȴo��w�DУ�R���=�[Ȋ������(:@�<�&C�H���3�tN�:�;��
z#7��A)1Ё�� v=��a�p\\�
��ʋ�c��9�-�N`���8�,�Ϗ~��� h 	���A���`�a�n�& 8Gce-��m�*�z��9���sm�F6q��A�#nۅN�S���&��b�P#�5����e�:�W�`� N��7#��N��;�Kcn6��]��L�v����ae��kfݖ"���6���w9]юl�S��YL��kFz��i��8���61DbEΰ�����]�6�[�e���B�X���q��z�;i�69�Y��P�p���Rܔ�a.�g9�$�ݶ����W���v���z���x���inI��<�d�
ԑ'<��h����6�]���粐ͺ�K�FwV�$ܒ��q��F�nŉ���K�.�/!v����%�:,c�u��O82v��]������ի2i���P��yeE�����"��cjcl�xYN,朴��ۄ�Jt�OiFU��.d�i9<iݍ�h�\9���}.q��N�J0l1>�u�����SA�ز�W-�v�M��*�gXt��"�
뛀�s͝�Q��K�"���\f�;j�ilݭ�aq@���#��j��4�ĚUq���F�=��˄:�Y�WoXm�r�6R���;��S��[��7WY˅������۾v"6�M��g�����#�j�Bn5;B�1������0$]AS�z�%�4;*��%θ��g1Us�@@i	�RvP@�M�Nu
�U��mg0A��h)1�Zc��ųÈ��J ���D�ڶ�v�v���m�;����lt�:�lH����hS�OZ��e˸\ɠ�	s���Uդ��h��ew;�c���t�&�N�gn�˞�gXNY%���HlJn�Sa��v4j�%�5*Q�q�݉7;S|���˸��i�q�r�lM�f]��$�L�[;u0u�Cz'`jr[q�/i�8�w����m�r��T.Y��W���bX�V��瀣
	�m��.>�vN�m�B�jBM� ۶it�35��N�\Lph^{�Ʈ�[[<0�FN7Sp!��禚�;S�S�����]��w���w��CH	�_;U4!�������(����$�v�,T��,�S�YA�m�c]�63���Wv�-��$l,Mg�ꋔTݻ=\!�Ft�s��!7��qs�l���-آ�0�q�t�o��>���'�����h��������`.��m��AZ�9�L�6vv�|�v�h�T6$�UX� K�g�:�s�	�:���m����ofpqշ��K�93�8�7&��Jpv����676{XY���h.�v.qKJsYG��[�������YI�l3����:�>'�䃧S����p�y����f��]ю�'H��	��yZ���� �� �=�l�K �kB�zixi�m&��t����mh����a��>m4Q�Q%T��$HL�`�]�R�Ýݝ� ���j�� ���ӫn�n�ě���mh����t߫�]/ ��R%uI�M��wi�h����t��^���=+�x��[tQI"���-�T�V��n(�]��υ7<sZ��=^@����l9ǚMTL5X�ݘޝQ`|�Z0�lxҎ�����Luv�{�}���~� ?���v'����2��~�р	r�}�fs;��SuT5EP4�UPUE��]����U���f��U�uZ��$�Li���?�_��O�]ـ}����������rh藦�������wR��JQ`|�[Z�tx��:lAb��ؚ�졷CWю�%�j�uκ�t��ۭ�QѲD�;lbE�E�Z{�}�%�I&ր{ګ���%ݘ����������(����cg3�4@n��j���JQ|�����:b����jj"&��uuX�K0�}�q��f�Ӽ;3S5?��3�c;;��g�,�wc`j)$��USUa��B�ݘ�{� �wd4���J=~tX��WSY�}�J,�j�> �]V��	>~����ib��env�tNrg1+���<-�ð{n�4K�i�Y��=��^��$�&݁m����h����I��R^�\i�ZE&	�N���J�x�n�f��>Km �0Z�Η�V���I��R^I� ��<���1�mV��$�C���]�`wN�N {ڪ�)���ٛ��g�g�m� ��y���h���������')"�?Q�tx�&�yIx}��p�<��<]��;��7�EvN�1����It�������R�~#_�yѩ����h����M�>��	��Q(�MD�US3U`/$�9�٢�\X�wF /j�p7[aJ�)�&j)�*�� Q�S`-�J0�vwwh��uX�ݘ�U�U4ļTMMEL�X�d4{��$�7@�� �ėaV��'M�� ����T�%�
=�l�Z0o�ٝ����ʢ30��[G�I��/Y'�I҉����`��ݍ�̇o�I���c��\V���ls�"k��cp�y�a����:���:�uqy����n��b�z5��j6n-��n��ùs�S�g	�Լ�]m^�h8#v��J2li�9� .���%N�����#�r���)BtR��c�yݥ�@��lAܹ^8d���I؛�V$ό7A��������o{��¿����ŞKC&u�k��L�	�\��E�c��q����b�;&7:��m��}s�"k����G�M��Ս�ڪ������J�"	bI���{T��3���_ں����vh���LT�S5UUL�M��Ժ0{UXV��{��>�T���m;m����	��Z�f �j�ffa�9O.���!���l�iwm�t�'G�NS��	:<pĶ��iYeX4�-��s��s�"�c��KyǱյÚS'Z �i������m=�	:<r��I��N��t#J��[���-�U`%+T�3�ghgyv���Y�tx�T�aWk�i�t��Z&���Y�33D˪����V 6�*�Η�V��+��t� ���}�U�	j���6�suIU!,I5�ܺ��wv�����;�U��vn���vZ�S��e4*���J�)�=��64q�	l稩�\�9e�9z�Ψkn�cM&ƭ۴�.zG�tx��ߩ��f�;�U��9�GK%AU5T]�Ǡtx��tN� �ӣ�>�h����[�����:t� ��|���IĻ��h�S��4%M_�N�؞{s�~�ֺ�����Q�K�~av��Wm��W��s����8�UXs;��r��`���H��ݶ&X�m`���G�I:n�t����.YWJ�m6�4S����E�c[�«϶�nޛ�4Mϑ�&BQ68�V�w����e��Ӧ�Ǘ�:<I�0��y����t`p0�%�ᥢ����Ij��ggg�r�;���@:tx�Y�6��P�'��UX	*J0wV��If �)������*������wgvh��� \���Y���fgqوwv�vlgl��� �%wD�~C���^�IҬ�Y�	j�)IN���8�j�qʝ�{G����F:�d���n^��	,n;	GH�޵���}�|]c�b U��ݘ��S�N j�V�l%.����N�]���K�'.�h�U`/jY���.\�KL�TU�5UQ`v�� ժ��`�TXqP��?�Z�t���Zӣ�'rY�j�Qa����]�8 �.��ze��U�i�wI�����H�}���]���" BRI%H$d%O�d% 5��(�˥�x �rm��07\j�U��'�i�����K�)��̷{$��.�t��&�:۱��M�j�륬��]� �-�\�M�:2ϴ:�ۻvx���m��u���3�yG��z{W"`�ըcsr�]�lnr�=k*�	9tޜ��5Ӟ��c�>��0Y�x(g��u����rYQ+�Ǝ�Ӡ��� �[\���kz�+{�f�y�ˠS�x!����Ɵ����$��C	i��C��Λ��f�@d=Bܜ6�<%��Q��Nu;ēW�}ӽ�ԧ �V�K0	p�(v7m�n�w�NRE��3Dr�9wv`	N��w�P-S-?��m+H1<Z'G�N�n�"�x�$Z�Q\�L�Ͳݤ]ݶ��Y�%:��JRS��˪�Z�:O���H�V��.������h�'I���zݱ�:�nݽq�Y^��V�۬�=��W$�B44�W8�bi���t����,��}�ﯻ쁻�{�����������{7���k������k�B�,���T�@zL:��}�U}���9W��k��A�2�8��)婢������ـ%:���ճ`�ڰ1��
����S�]��@�t��>0����I��r����67m�;�;����}�M�$]/ 'ޫ�X�� #s������Wg��]�s�Z������Hlj�2ٰ!����|��[Sa��� ���=�M�:��`9�}��|�;�ͲƐ��{���u���:s� 7�� �]r���	+aI7�ǵM��kK?U�Q����3����T�C�INbѠ�Vf8b5�B�!@Pm���_�]pC�o���՚D&5�'�N㳡��uMk�A�	�\�A���]���)���7<��Dcc��AG �"���̰�2"��(�FH��
���<[�����-�Z���a�YXƴ� �(��8zm����P��fs��𸐼fi���W�RMK��i.�\�Z��Ĥax��s�*��h(����� �������Q��	��3[ �n2��8xyu��A̴�AHgQ��8`�NEa�� e魣�;��`OtI��GC3�P>x�5aB�t�vob�c6'jq�"��GA��і���$i��!�L�`�MǑM\HjQc�������Ɗ.�::��*�a�7�c�N`9�Ԟ=��Km���� ��A����{B��(�0G��H=��x="&��"�l�(� 4*��Ф@��x�� ��(�t�Xw�vf�1�Bߪ��|�`��D�M�LlLJ�&���� }��zt���3�;�B�����*�h&F��jmk4wG�;��_�X�ό6���~����Ҙ�b��ڞx���Z.�.$=��6�'��ð�e����N���:��o ��n�/�,����W�&���DUTKS�3Y�(�S`}�ZX��V�K3��)�
��m6�uv��=#� w�� ��t	~�`~������i�BY��M�V�K0Jl3�ɏ3�ó;|���H���	;�LB]cb�@�i<�F�u�.U�z�Y��o1ۧm$]���?�����E�w/u���V3;|���&a�f�*jh��k�N��p��W�(��)uk���-r���$�㰴��35,AU_|F�M��>ذ���ݲ�Wfܨ��!�&������7����3�D�U`wj��y)�;޺�1�*ċ������	�'�n�/�,�^��
���K��&�����f��]�ѽ�`f϶,7��}P�w`4ݪt]]���H���ŀo��`-���/�f�C�o�u�(n�{r��n��^��������v�m�ݴ�bюu�2v�n�8��Q�[�I5���7[4�Onz�:��� T!&��wp�ٚ�غ�%������pO��Â.���Ř3%6wc���m�ۛv"K<h"�v��ⷤuz�W���6���P�jz��ʹR7d��;M�Cv�E��7ض�7n.�cu���Q�a��:[4�H9➌www~{���<�?qe���d��u� �`
����31�����jy�q�V��m�
j&)�*��f�������Y�(�S`u��:*���n�V�2�wG��՘�%6�>ؿ�gx��ؔUD=STT̑UU�ݫ� Q��ߧ���<J'R�
��MQbOt	~�`��^ w���=�t	9�J6?�lT�V�k ���x���H��]_Jv���Ӷ���i�ڸ���A1v͝]����m���/�h3��:ը*ċ������	�'�n�/�,{=� Ѻ��V��+N\�x�{~��/�1!�1����W`|�����]w�U�k�x��<�u�e��v��uv���"�;�� �{�'�n��:�:wm�ݵn��X|�׀�s�$�M�=K�:���K��wv�tڵ�q����/j��i�>ذ?*�]�߆�C�KD����d�q��:M�+�6v2����h(㗴�Hy&{eb��%LL�0EU|�����<��`o�� ��� ���)`�I&��'��8`��^ {��IIΒQ��E��r�{=� =�����J��gb�|��QT�z�o��u�I���;޺�Sn�e�-�Wz��|�X	{V`[H�7��ŀ7���a�骞Z�&�j���0f�����e�{���R+*����:�ճ���lC�䗞��]t9�:#�k�l��w]�� kAηv�`4��t]]���H��{� ;��Iu�)�ӻm$ڷWm��^�����{���"����t���e��ڵ����<Ot� �����^�}�m2�&��$("����0y*�7��Ň�]��܈R�`!�rT{UM�J�j\O�x��z��.Д��%� Q����� �UX��0wv�������f��:�ۚK�$D��"<1�����sx^^��.�P�;V��fcu�6�����zuE�o��`r���fo�;g�,y29����&�i���� [����0�J,�}�|��� �Ĕ�K�M<�4ML�Xڻ0�J,�v�^����<��+�Q�E$��t]]����X��b�=�ڰ����`
7���CL��&նZf�/u������0[H�1��Ì�0��1��0+��6���kz�Fۣ5��3n7Lpu�g�g��ݫ$۶�3�� ��q	�D.��=bn�����b��*)'�[%�/F�p�c����m��m�n5S�Fd���v҆ml�(
�����)�<f�yr�OGCcDlh�<6CZ��t:�%/Jg�C�{n�.9�mf��񣉍ӻ��VCD����,u�%��VI@����V����G��[�Y���Y��_UT�EG�=�;�ߗ�N�ۧ< 0�6�9��s��yݤ�m��vq�ҵ�F���F*ݶ�fe����{���K�a<�^���[L_�CV����?��n�/�,�^�����PT���[e$��Ğ��"�;��?��]��<�����*.Ji�cBb��&��/u�{��	=�t	~�`}����"�V[t��V^�N��	=�t	�%���^�~�q)j�P�~��"�6�zsu�u&X�2�֋��Нn�ga��b}�����)婢�f� ��ـ|�(�7��^ {��}
�F]��
�$��]����<�t���8IE'7�0�@*P.��_u�����*�����_�r�2۴�V�ۼ�^��{��	=�t	�%�}eN�n��m�����	�'�n��R^�/u����~M;BHV[o ��7@�� ���<}G��nӷh��n���؃����4��Ң��n���[�݋����;wt��N��*�MQbOt�H��{� =�s�$�M�$ArRO��Zm`��^ {��I}rE�}�u\��H��Һ�Yz��|���q;<UXDv}Ϸ�'�K�
�㻕����*um��'�n |��~�lXs�F=�ouD0���:*В{�I�/u���x^՘7!5�t�T<��LL�CA1Sj�{������%J�7/XJ:�(���PۢKt�i�ݤڷwm�yt� ��� ������}eN�n��m������U|�v�� �wU��O�,������	%v[o ��7@>�<�^��{��	*_R%�I&��&k09���#��V�� ���aq��a�96���]C�ŭ��
G�むlG��s���U��+?����Ƅ�i]���/u���x��7@>�<~�.��t���e-�Cil�8����v�
=�f"���U�����)��l�2ݍ�E��n������ �{V`�U�͐zuE�:IT4�IL��U3U`w�ՙ���`}����<��Ď�hv�h�otzG�o��x��<}u�)��.�&j�*��w��Z�������	� o:Rwwm�i]#3/@��ݛ����7�������_�b�����`A UW?��
����'����S�]�9���DD��k�f(�������� ������?�������O���}�?����?��E��׿~��O�_������?�_��������I*U_�}��������?ހ
������A UV�?���,�����������7�PU_�����<�������x������������g��?�����ހL�P!�I��Ie F�JPH�����R �Q&IeD�Q �	!�RQ�YQ!	Q!I�$YQ!FIE�Q$DeD��H@TITQ!T�RIQ%HHYQ!XQ$!D��HYQ!Q%HQ!	Q!TI@�� 	 %D�@eD�E%D�TaD�T!D�@%D� �@HHHFTIHID�HQ%R@I��U��Y��X	��YT��		��d `I	��IT��@`  ��BU	�� ��d BP�� $	B@���������B		d$` ������� XH��BBDF@P��Qd!AHBX��H �%��BR$" �BIa$ 	$!$!$! IIFB 	!%T��RBP FB��$	XBBF@�!!		B �$!	FB� IeP�$!RB���� !&	d$$d!�$ $B��`	T��XB	a����$��P���B��		�"P�	� ��@��  %IB�H$	BE��U$	UHBUYd%IF�B@�BXa��� !		� �A	@��%� R@��&B�1!	��)�%�$e �$�$	U�$QXBa@��
���&��$!	F �HB	EIBB@��e $P�%�a� � $PD�BA��B�� � 
Q�P�$HFFQ��EhFYFXFFV���a�d!�dVQ�Y@�R�$�eX@��a$H��P)�
Q�P"$!e	@���@�dB!�
	�deBP&A�	 B�Z(@�X���@�@?���������� UV?��σ����c�����ި����������w�w�����8s���5�?� 
������}�����~�U_�
�����s�p *����a��[� *���������9�v�?��������gb ��������DU_�˳#��c_�G#���� �����b ������&�?��!��~�W��w�t�����'��]�_�s��@U��g����h�8����_Ǽ��w�����������������ސU\��������k���������)��=�P��	l�8( ���0����f� l�PH� �>�   :    �t E �� b�| ���@@   (Ѡ(�� 
��J h    Ѫ �  2 4x    �q�@*�hА 
��Zo��o`{�s��0:��A�x�+«6��=���9�:w��]JJ�p:ͻ�J��8  �,��s۪���Mꪬ�Pu�nf�ZU�]5K���R�f�����{�<�w�k�緡� �}@ ]�  ��J��o�J\��:n`
[� �
�PP3�����(�@���f�JR� �;:  
Ss  �������JR�YE ͔����R����J큛������h n� :Yef � ���z [	  h � � bhR��}���=�zo0�ZwT-�@͇�N{y�6�9շ��z�Zp  /G':��P�g��s����ћz;#s�u��  >��e �A@���O�Z�A�a��`t��M8��v9�;���vPrzx����a��px���<����;�Ԇv6�����xs ��n`�d  >�x �P�  �m���|OA�ށ����`�z�Af�c���빀�tPy<fzC   C��&G�x �3�;��eͥ͹�����{g�w����`t�     O�iM�)J@  =��*�S�  U?Ǫ�'�4   ������UM4�&CS��R���@ h"$)��)�@G�|���������������I���u���**�����"��DTU?�PU���"�����DEES���?�����4s�~��7��ƞ��捱Z�XB�$�i�����9�C_~���M�������Q���!����I����ZS��~��*�gNP��>��[��T#�}ki`�w>�y��v���w�;G{]�[�	n���T�o�_b�ov�(W�}�xƾ�ՙ�3������ס��nֽ�����g���o.l��}� i����a�����������߹���s��}������Q��sf�&Ցe�oO�0�o���g�oZ���7�ٽ�����>�6�w'�}9>M7���\��[
[Ȓ�Nf��
��Y���#�>���{�	/�s��
�W+��.��r���KK�d��T���)�!klIyY���wϙ�L�?}ݒ�#��K+��+�����k�]�_֪)c��F����sm���\��?g!�p6h�wd�wM�e'8~!BL4M��.��fk�,��$�27K�G�)�j�&d��e�K����\	BY%3.�ٲ�q�޹��WF����X0��:=����twɟ��̔9 �a;$h��$
���k��d�G�	y�y��S4��h$cBcvpq�:W�4% HԔ����55��L?a3�>L0:럍l��I����>�{��	��6�3Y���:�H��܅֡�]������՟�ЁH��� ���sFȑ#"ot�he�31���З36��]n|������>���2vą�rb��T�~g�~��s��t[�BR�`RR]k{�}}��)����E��-g��]�i���yAJ��S��J��_gʮ���k韭��5\i	*S�Nh.kD7�ne*��X��6S�O��cz[�Ϫ�+yֈo_�t����஝b�t����kk�� ��A�RbGH�Ѹ�P�`�`��j0+$H�� ��!p��L����Oߍi�i��(��m�ٻ���_:8
�q0���S5!t]İ��,�C�"��0��7��K۹�5�cC���>d�H0!��ܿdsZ���3�|�0�#\7������B�	�L�?p�a�����Ы��P�UA���G��T��mn��*ӈWQy���Y���R���/�u\q��������ݑdl
S�wv�5���'���zg�2D������"��)�aK*ZCs��ֹ5�g*QJ��2mjo{X�QJ�/��7W�}�����޼�}���[B��ʵu|Y�&�_�%u�|���tQ�++Y����/G�E��T��ǔ���w[ə�ۋ>�����R�}ߋ�f��΅M���☻Ws���}���߾�-��<_V͟1�%e1�\`@��b�a���\
4�:$��qb ��5�d�����@�ke����,����+����w;�����Ue�_~��@�}��%�����?\>��<�3��O���p�<��j�ߴ�|�t�������t,�q6��U@p*����M~.#:`�k{se����j4�Ip�S����I��F��T�12:Я㱦�E>�f�����R �J���c������3$�@:�FĦ�0%9����\_�Bsq D�X���Ҙ0+)
�)����0ֆK�Є��HQ%k	SZݼx�KP*�k/B%r��9.Z,��B0i����v܁f*JD�c�71|��sM1�Ĭ4t��N�	B�,�`StF�kv�Ԧ3��f�H��T��f�|5���0�X�?~����dd���O� h�|���� B����d�3l!5��z.0!!�$!HIc@�6`IL���aX�RF6i��2��p��l��R4��%q�B�������C#�D��@�1��#�06I �yg,�o	��RY��i�!�T�e6hȖh��3��+!+��!��3g2�����)���r�p�?a<4lؕJ0����/��aH\%�BXR}��d5�͑3�p$$�R!$�6A#�9��MD�j&G��}4H�`@��m>uI���B�B��c.R6HVX�Y:�P걊Κ��4���'ܸ�B.�HBv��9�̹ٺ�ԛٟ�1��?o�}���ѹLө��7
lԄh7���F۳|���l`Mri	�~���3L���"�H���(@�1n��X�%�h�nib0 @�`0�5&[4��\4�HP�f�8��㨗5��T��CT+u��~�d!��a�}���݉qc"B�,!��	>�s�� B:.���et��뙽�#[��Ll�@�,l��Ϗ�l7۹�H���p�%c
��	8�pLM��%I$t�����s�9�P�����>��C�u�2! ��D$u͑`I�17�Cl)��8���8~�5� ~a����:���T0���~����@qeo�ߍ��Ƣa CYM7Z�|@�.�xi��e���4G0�$��`N��3�%�+�����$����Piq%�$#�� ��ru��c*dHL	bI[L%�|od��j��F��!���c �k��ʒB3D4�f��c����IH#`�u�!3F$6F�n�¤*B��Ť�� �,���	/��C�3I	�RYM��N^�a�p��}�yJB	���$��`�%2���3�Ǥ�C!T����?H��a"O����s�s�w[���
@��	l֓?@��Ga)B�0.�&B��~��LntHeĀS5�}�;�6Q8����S	L#B^@��n����nAִr��O���#]�BX�0�橉3y�1�)	/��ˌaD�B�#.浜7�l���`�1#\���#m!G�odo�00�1%!	L��B�HV9)K�&���`�SFϥ܄)l��۝����,&���	w�������"@���2F�@�)$		Mn��ݦ�d��o5�L��R)N8ᎉCF����5�f����Xտ��@�bl���4$#m�@`I1#��rRh����9g E0�$$�$c D����D+���k{��V�Ns_ZRY[�u�]�(B�b	$X�b����)0�ԅ�7�e�� �L���rj��k�`Ѹd���~�f��w/8t`ӿ�H��m	;��%�<)��5�亙�[u�Ԅ��gkiÁ��{NK��Bjܤ&2�Hi!m!��U�4C)5������E�!��;̓�aso�iJa��.�ٓ�~䱄�	-�k�+4l���aL6��T�]��\$5 B�i,���
�0(�J�L�)�\.kd�)�7������A�)�)8h�Ń�g3�������$��i�$$h]r�o3|'���Qe�͹�.�<�L�LǗ��r)Y/�.%圳-��!���% Y%���(tD�
�k
1 !�\���\�
��>i�Ka�+�4I>��O�@�3Z�I��%��6�FCn���~9�Iqwꜣ5�QJ�����ͯ���¥%��\���I���na��!�T�$e�䙲}���o�蒲�)����MҎ54��[���fΐy��R�e����ĒG_F� G9���������r4%�w�38e�w�Wl�/HB�F��cQ�F���o�i��4��K$�~-�9�K7�K`]�aB�;	 ���\�	e٨F�E��e�����E�0��b!"A� Dk�)��k����#&�B @�F���,�D$��u����d9ƫ���?�(@�*F�a�a��krI)��éх1��Wp�@�F�Hb��!�P7�C�2�~�Ϻ|��۸���&��jf.��%>	%�Ê��+e2���>��彷Y��]���Nk�:&�og?g6sZ�����>��,ˮ���$B�]oF�p�&~}��M��m��4`F��I
����N��p��C�g*�,�n�԰����r�����	��n~�&���0c�`k�~m��pbq<!$0b0H�H5�h��ÿ�����+��w�����6��0H,lX�0�f+�a4�e�DXd..$ƌ.��n.k���\��~�������B	!�!\��޹߾���}�:	sB���R��\�'w�9�N�2��}A����h7�����\	�����7���$	�C�k�A4�Z20�H`��� ��8����$���GccHϷp��s�Co�HK7�<�y�y��!|�ٜ7�nr�Ü7�]ȜI�yg8�\x���WG�Ys���۩?<d���ӣp�)�.$�ˁ1/ڥ�!94p����ӧ	g�g�)�C��IB�*�H��%S��ĵ��KbC.�w����ĺ̀P�C�i�jI)�I#xr��4���k��?Nk\��HG�n��4�'����(dj������F#�r%L�!��l���������E�1H�!8~t�$�B��6%�H��F,b�ґ4h�.2<$nfE��)RP�ֲH\B��$&]1�`C
F5�D0+��ק0�w�����[�����K�M�9�ߏ��Jp:��\	�h�H9L�R��|Yh�����ЙY�L��vo�x^Vp�-�
����n��np�mm�S6v��o9�t��,�o�a�(�k3�ᙽ^e��`I����jMg�~�O�.��o�K�}μuK��
(��p2����/3�|�}ߨ�ʪ*��`Ua�(�WKtt��r����y\�eP�����+���s��&��HI�%P�R3�y;<'�o:It,��Oy����� 	 6�            6�                 �[Cm�       �` p  h�[@ �      6� ��    �       m�                  �:$  m�	
��Y�Òڣ� ֮�X2�t�5�V�ԍ�n�v�Vıj�a�UX�V�*���A,���la�m�UUZ�2��v4)-^;u5�UU�ce�D5MT�z��\��UO0)//ۏ-�Eh"�0�P���v����O [g3>� �������$�M�8z)0�HS��UUU@UU J�e��jڨ{-,pa��\�V�^�@�R��5U��Z�e���
�Up�*�ݪ�Z*��[`*ۂ��V�T�[�k��%��`DjtmүPN4�A5��=M*�VRPvuE�nUBuUm*�X����3��r����m������r�k��j�����+�u�b�F���'v�izӑev	��6Q����
��M��t�J�	�ʵUU���v�j���ꀪ�N�U����v�V�U�3�f������8���P i��
Z�
P��yk�J���n����*��[ XlmuU�f�vWNðQ�q�'�`������*E�� 	)@Æ��)awfj
�#���Y|T �]4B�\��UUJ�WmUOk�0��UU*�j��ڪ��u�l�&���'F��@R��CV�WQ��j�Gm\��ͪ���v2
��f�/��ڴ�c���0`97-V�񔞣��,���Z8"ܻ�q���H5�D�ֆ���ƫS�1n^^wdϠ �������tiI-۷4����r��T�mN�.+oX���͔��n��h�EҺ9.��n"�v'��9�m-��f�'�b�
꺩�6T.n��Ү���e��u�T��T �UU"宬!�j��K-P�ݞyjT��u�dU�p(-��OYn��8�2�V�<�l�kl�s.�uUG <�El9jکWj���A���-�����癖��
�q�a�u��AȺ�GplrX-3hv�g�L�*�
���Q���UUU�PWf{*�uJ�[[U@�UU�������
ej��j����V���^Z�
��en{	M:㮹T��(J�R��� ٝ��Sj>���PA���|r�P�� ].�j�����乴V�J��*�U�R�T�#
��)-�c�誩W������]V�@6��U�Z����vU٥Z�����-*�U�UUWR�W+� ��PUmU��J�����dj���UU2Eҹ���S啪���`VyUUiV��Z^Z������Ԫ�UUT��R�X�[��UuV�[UK�j�U�N��
ܖ��m�TNs�x���U��UV�4pT��Uk�������>hj�
�iV�ꀛUF�����wV��մ����v�୥Z�����U<���Jl7 2�"��Ώ���j�\fU�l���b�N�.l�M*�]3�j�MO�1�&��E��ETU[UUU@UWUJ���*�s�ٵ8��[[U\���l�X�̛�h��� v�VE���`�j�(nU��U�����z�)�	#):�j���\��U++\�U��UT�a��vMO)�s�F�ne��7] X	���j�Pp�
�<�G����C��ݬ��.l�%%�m�&'pp�e�P�<R>���lr�gE�H�K�V-$����0�p®Xk��UmPIټ[�n6�i�Yy����t�t�Q;`
�eP��:0�1����N+�UPԲ�W R�ە�j�M���V�:g�u��:휗�WU�<�q��c3P7YT�c9�GA���}�,���x�km��9���M�Ġq���F�;4q��w2����Sc�`�d�(p�P�Y��1fk�A���c��AѹӴ������p�\�y&W�-ٟ)J�<�̈́�jcl��"�p�5��X�n�MW.��O�9�l݄�H;m�v%�R��Sܭ��{F�N�ب�(�L��&%7m*���R���D��9��`�Y�UE.Km������p��P�ɹ��@�$l�;8�"��6�l��Ic�<�Tuq��]&�EUX��J��� �ĶڮW��&����9k�5���m���yZڪ^t�Ed���j�8Wv�Z�����M���.���N�}U�ڄ�����Q��jZ�mPq�UR��C��5� �-*nk�+PuT֩Wf�yEU��kg��iV�[wj��v��j�vAM�Ob���n�U�`*�0M\��U[T�J��,{q@T�j���U�.�=+�sW7(ʵH��UUUGR�+Y��SU=����M�TVՖe}�1�qtl���q;�앸����|���F"�����Se���uz���n8�<���z�%��۫6�;*��zs�
m=J!�/\���(y�5�K��;;Uj�Q=��v���g�QP��Yl��QV,A�˩�b많�UR�UUpR�͍�[Mc+UJ�� �Ս�����R�R��UUR��J�uu;�z
p�dCi���XrX8�tTm�FՑ�q�����Bn���%�����P6ؐ  �ª���S��YxT�R�V���u�����8ڕ@�"fUmav���J��	�Z��@���	3��]V�����Z�bT���6��Լ��T��UU@R��I"`)3l���ƅj���<��U[:*���P(��mSj��i#[I���@C�Z���Tk���mڗ�j�ګj������nERaU��UU���!U�Z������T�_�]_T���0]M�����B:z��&����]�e�(�+<�p�U[[]Um��7\J�WumUP��-�q�UZC��ú-���"ݻ$��U]�Z�U�:Zr��áB�@�+nW�V�`[�)�Ô�Il���Z�pZl㊱l��h��փ� E\�m�UT���p�*�
��+�T��.�v�{VE/$YV �����b�8
�L�X!�m��MK�z��/꣙v�ƃ#@�a�BUupt�R�.y����U�U���_}�l�C\]�svO[���x▝��5mR�poU��ط*�p.h�5��*%��\�$��`�U���mѡs�ƭ�i���MU*�K�� U@T�⫶ʂ�l��	�b-Wb���kn�ة^j����Y^���V�	�UJ�UUe+UJ��P �]�\9ـ��	����m�2 �J�@*�*�j��UUl����Z���<��nv�V�V�������j�h
�%%��^V� *���U���YUP*�������V55]�9ye=2v	�G U���� }UUr�mVҹx]��������	�Ey媛K-T�UT��T��ܬ�`(6����Vk�UU�5�W�	YW�eYx�Ҷ�T�U�u;cc"��;$���[i}'<�T�U]�𕑭��)^\�ӡ<���fk+%����:ێ:�5J=��]�08�{ó�s2�\�Ptd*�v�: v+�ڀ��q��`�r��A�[���|9��"��v�UԦL���U�e#����UX+h-���;RUl�\9ݥj��ݪ��e9�UJ��}o��Ǝ��gEEV��\�L�n�Yj�����&
��
 ��s2���m�H����f��v�	#�m������-�oJ��: �X��[<��Rک[GUmUR�+U*��6�����ƕU3�U��x������ګҼ�.�@-UUR��q�PUt�Q5�KUWUR��UX�Uﾾ�����*T����20  8�-*��*����Y���	iV=mu[T�M�<ڰ�� �V�6��z�B�r����X�$�9��Aڃkѝ��͙�I�lKJ�\��!
C*�1c���� �����u*�T����^TVVU�&��V�� 獭uT��UUU�qK�
�Y]��eM
�]u�]Z������^[�s5Pq�]�+2�OZ��,��jC��r�UU�m9�,UU�pUmM���d�U���3hÍvtUP������.�	GPMMUm ��Uc���:�.�#+UUUR���C��V����wd-����[M[E��0S7FAV��%����]���UV_��g+hX���uv�uS�+R����հU-C��G�'�ڬ��=Y�����3�"e؁m�\5)A`2���R��F����@7b�RZ��.�`��Lԫv�R���;�r���R�5T�/;*��LqB�[WQ�+,��y��s��T8���F+�� j��U���CT�`{k�jU���󉕪��T{Z�T��4ۀ�鶰��A5U ��!�eF�U�*�UVÌٝm6U���%�u UR�������Z�*�2S���%�uVy��U�T�r�UUR�TUT�*���▕m�[ʮ��Z�:��+46��z�j��mʁ��M@r���UUUJ��T���UϘ*� ��N���l.� HH^ ��6� J�J���V�UUU�,�4�ذ��hٝp�Us���Z��Y0t�-#l�U�[T�u�������U]�\���H4kQP�>�Z�y	��W;:B^�U��6:�jYC�Z��Z�[`t��&Ԫ$tAs�T��@6���ဨ
U�V:�@Z*�U��,�8(.Ȫ�m���*k�SMC03�����^����&IٳIZ���U�|�|�?s;Sr��) *���Zֵ��PDTU4�`���x8�h� ����C��t|�jB� �A6]#��$E� �"����"�ި$
1Sj����6�O�P ��P~� � ��p� �4&�'�X �����!PU��H�Xh*"�	,6�����:Dz�ʒ b"� �a`ȑ؁�)OT>j� :8���N�T?*|��Ù���/����π��`&υb1`E+�T�WH#�]D�����H�� �Q�|�A���ٯ��v���� 	w)�EB��~D@�z�?�X�"�УN ��Ez)�{�0�r�`�C�TC�C��t��p �P���"�	�>PG�
8��bH�2"�$�^�~�D?"x�`��)�L�Q���:����1AM�m_���Q�RE?E��N�	Uc %��ZP�J�Hb�Qj+I�Ps�H8�� H*��M��|(@�u��Q�$��`#� �`�'^��Sj@�� �f�l���ioôO���P6��lD�P��ҕ,���)B@JBElT�F�YJB,@���`6  ������)�'1"�X �/��ld$S�v���l��H��6%6(�����T��_�u���^(��?��`�-��D(FB �!�>��\P�B�*.�(�EU*��`C���	����2��
����    � 

�x����V���
��ڮ�������n]����[�3�t�{84�ct���6���p1GVPJ�u�t��\�*VD72�)e	6VPW5SPɣm�ܫ�Q�C�� P-\��ӳk;v�:[	n��t��l�X&C�xI6�6Γq<'nʡ�6��9�I%U��4-���$�v&e����3f��+b�x0p��N5��U/�Wr�=�6(�y��f��8^zvy�T��l�#8���5�6���t�E6��Vk�	�v������.�ڨۭB��e��%ƥ�a�2ڤ AB�T3�<�m�28��6Ս\n�	d���N���:��. �n�ș�k���*��U�[����m��9ؼ��*p<d�I����}7���6ml���q� ,��;5�{��X@շ�\J��vΐ�ϲ����D��h�j�$
X����"J@�9[Sm6P�3ƦWi�!zĽ���/��hפW��+<B�{�Е���R5�6�0��A�L')չ@��W>�5\S�f�Ev�,QJ�痎�T�\q6謯aGZ6Tzܻ��c��`3F�f��؊CWY��*���03V �+�[WX34���+3F����8�X<�rsuU���І����$K+���;<�*�Uz�hQ�2+�M�w(�!���F�X�X-j�<ՉQ�d]Z�66\h�m���Yɖ��n-�t��V����YD��;��`Y��)2�k
�X��]�av�l#��R���JO,�Gkn�rej����%`-u�nN[i9��;��=5��nh��s��@!7ghge��X䋻eP6�$�a�j'!6]�h�}TV��N�!Ѵ�A����cc����m�I�`��d`
�n����v���h6H5����\g�����w<Z��R��%W��G*�-�\�0��7Q�'=���oR�݉n��^Q�tֵ�d3TW���O'$�6%<��P���� `�pC�8�B)�����799y��%�Sx��6��f�S"�d�3�<��՝B��:������Uh�<�6�!���wBe����6WHinBG��u�v���!�u���͢f���r���cl�NZ�ވ����X�m�e�1�f^mƤ�1R94q%�i�l�{k�<f
� @��[e�!l6�7X|�rn�(���۰ѵe3Zܤ����O�u9���9���q��wn�v�x�Aܛ��n^|l�������d4)e�4&��g-����� {� �����r��A=�� ��z�*�5e+�ZWn�nǞ������{|�`����J�eYƮ��I[x�I;0[��nǀ}ݔ��WW�N��n�o ����x7c��lx{��Ҷ��*�Sv�Wv^ M���<v8`�W*Hz���,tI��F(�V���1�;��1䴕� �뎼C�n9��t��͵t3��='� }Sc�'c���/ �oyM�uV��0�x�w�y�Ol�a�������@?-�����"���	���J4U�v6U�Ӥ��'c��v^��s��� ;^�x�x��T�񻤕� �ݗ�v< ��ǀN�t���cVR�e�v� &�x�M� ������x�G���5K�M���J�ej�A&t3�*,�I���B�kb%��v��՜j�Eݷ�k���7��jݗ�M� �vQx�Z��:t��t�x�\0[������<�9UI�W�m%mնR�T�� �O^ }��[�"?����@��+�(6(ࣽ�;�krO��7$��S���l�P�j��>�� >N�׀w��j���>���իl(�4+�������/ >� �{�e=�,��q��V�t7\;���ٵ�3�y���������>9L�(�ҕ�4�]�����5we�ݑ��6<d�x��T�񻤕� �ݗ���URA��� v�<��\0Ҷ"�)�)]2һw�vG�T���U%��-���J��b,�t��V� }]���\0�v^�s���r�+��'����{����u�Me˙��;�p�>]�x�dx�wc�;���i�H�;Z�m�ڠ�i]*����4f�eM�i�L�d���L�).d�� �we�ݑ�ղ?W>A���߬��7M������ |�޼ �6G�w��un��>�S,@�cBV� }[#�7��un���ǀl֒�Z㻻vS���o�Sfx�5I���ǀV���񴝊�>7t��`[��Ur�w�������'߾�f���c"V(	H-�D"� %bD��Ky痿6ۦ�sf�͕�@�*���h���:Zݔ������u��q(J�vwb.��j�Q�azI|��,򮀍�,Ӈi���qs����]�̊d���3���^{�g38yݡ�ϦR�+cc6m��0f(��U���u��:2q�x[���2[��&�K���	.F��!��M�>�87a���`t�3��i�;b'��4��q*�`sc��f@w�'���R[D	�)r6�
�#�^�>��uvc=
�WT�a�\6Z��ٌ�2B�)q.閕۽ ��< ��G�N�ջ/ �R���Vp��b�o >�����8����O^ N�x��J�ڵut�Ҷ�Ӷ�	�p�:�e��ǀ'���>}��2�LfRl���[rz��y�ղ<v�XdU�L�l�̵�Wp��׀'���'nE�un��=\�+�k�)૪i�q�����s��k��dZ�a/O@�-`l6Mӣl@���u��Zƃ����ߞ;r,�v_�ʮ|���x�i/;��v�"k���w��o>������p��P1B�a���?'W_׀��V��ݔ^:i��>7t��XV� ���ղ<v���>�'�!I��h�ݝ��$��V�������nE�un��;�T�bĕ�.��[o >����w_��T�� �v<{��L�� ��ۺ�31���Ԯg9a�2�b)D2��Z��f
�T�i��s��������o �u� >����84[v6��*�un��;�p��dxݹ����E4�������N p����H+�E)~A;��N�o�6^��r�e�[iZm��l� ��"�:�e��`5���\j�ݔ�WN��>�p�:�e��`ղ<w�Eh��&U�w`�]y��љv��N�M[M��kƎ��ӂ]*mX+� ��[rp��{�߾�0���c�ޚEE"�ʻ�ZWn��\3�j{� ����:�e�#`������ջf v����0�%��`vB��+�����n���}��uI/ �u�~	�!!Z���h�����[l-���+t��ـuI/ ��� J���>�p�>�h�K
C.��m�[H�s���Um�Y����Q��Kh�i��cK��b�l4V�Z��}��� 6�G�}��uI/ �^�,Tիl(�	[f ml� ��� �^���J;�Ʈ���eӶ��0�%��`���	*J1�v�n��I[0�%��`����0��*)�Ո�bI�xݙX��<v8`RK�9���y焁�<���m�X��Q�c�Jp��Vʽ��4X]����%�],M����4i�<�P�/����O$�������OC�i��������Y૥5�`�%�>�#z]v�3��\b��\��>���`48�n�p�f)�0�6�� f04Ԍv��#F���I(��0VlsS�6�w�nNɜF�!�u�1t#I�&��E��X�R�=$lλq11c=�<�$���u,��k�f��_���%˞�X��ڛ�Օ3g)�<y�ca�����c�J�
�������ߞ;0�%�ve`vB��+��`�[v��x�p�:���Mٕ�[#�>�84[um�V�m� �^7fV�U%�W�x����L�˫������w�Mٕ�jڒ�	��uI/�|��ō�(Aa-���g{��p�:���Mٕ�Ԩ������v{�mDy�;��E�!�6��7G#�Bve.�;]5�E����f.��ק �^7fW��W��^���IE^�fk��<] ͽ ��<����$���`$A��ȠfYpP4�Y��\�bI)r���I)���K�!^��.�.�?>t^�ߣ�$���I%ے_�$�tx��gN�+m�Kv���JlyF$����`~|� �y���[�R�F9��I)���K��_�$��1�K�O�� �NNI��u����Yb���������C����lN��I�o$�F��x�q׵j�gL��afV^���}����΋В]�r/�I)���dP��][�*�����Ρ׼�&�?y};����Ē]������Uݣ�(�����
���KIl��/�I)�01-����l%���Eֵ����D��)/�88hHa�(q�u��BS�+	"��i�]l"���1 @���4~��C����L�����d����p��Z��L�>tRl����m�a�k���!����u�~ۢ<#Pa�$ � ��N�BP��5X���Qt���ʡ�	�@�l0�0��`�� D�00`E$`�JH�v��m=��s�9�Ӥ��C�CoA$
��T?|k)U��v���
��:�}M�ƴ�&����`I$d�H~Wi�ڸ�������ȏGt�܁��b����g�߳I?~8]k4�H�&��u��F0���PMIe����b�B�~���	�H���,�!�ӊ�����~W� ~*o�!�@�D����t����@0k�px �hubT"�'rK��칔�$�t����\j��-+t�_|�Sf`bI.ܒ��$���X��fw����[oi�Iw2�3N�km�Ē]�%��IM���$��9�$��:�ހ�0�y	@6���2���pvc�������Nӹ��ݴ6��2v�܍4n��w����C������`l�s���Ko����Il��Ь�ۥm�Ē[��_}�]���`bI-�{��`~�u���l�{���i�R�S�m}�Iz{01$�od��I)�2�$��ӑ}�Iwa�ĭ�[`��@[t�$�od��I)�2�$��ӑ}�K9�^�. @�T)U6��X�[7��*� 08�$���[�������n��r%Qw}�y�y�: ?s�r���g��Ԓ6?Iv�VbI}w�QF��r����+]���a=n	�Cx�8E�����إ�*]����Ē]�9�$��px�K��_�$�v�R� �����;M���'}�o1�$�{%��In��X�K�NE�ޫ�QW��z�i�<].ˎ���}�����X�Kv���K��W�$��QJ���f�.�߷�C������`Ƒ^$���/�K��X+8];t�a���|��y�I����v ~�{�����ݗv�h�����b( �,D �H$	J��v����Ҷ�R�Ѯd�9te��L�׶�S۫�ʼj�̧��p�Y�Pa�o��#1�hb&5�G��sYty <�M�ڛ���|cnXݏj��tc�D��j,J�ҭAOj�ݷ;�q/ckg;*r�ta��+�u��ۣ�b1t�'��5oVy'�<�ѵT:������O67�WpL��e8B�S4ۚ�j�3Y`!��9�Ig���;� Z� �u�<K��7=�B�X����n�q/H2���F8����hԢ���ޤ�����I.��|�[�2�$����}�~���Y���f6M��{%��In��X�K�NE��%�r+��ʻ���OomFi�\�T]�`y��	%ݧ"������o�OIm�z��$���6�l�,à>����};���y<I%��/�^����,I%'�*���x�b�}�_����>�~�~�$�����$�v���Kn�F�P4R۵�ŗl0[�^�taۊ//��܏<]�2l����e
^��W�v��G����w9m�}��wm��ƻ��"!�'�j�;������~���"����߷�.�*qL@LOo2��׽y�m���= ���n��I��'"��Yo��X���9�Xt y�~�����zv߷�����7�C���<���M4ma�c�����}���}����y�: ?�G�� ����M6t�P��7@%��/�Kձ��_$��O�_|�]W�^ NI�O��}��K)[���\\���ܣ����oKe
�x�
.���$�l��K]Y�հv�Ci��RKe�)bI.�nC�K��+Ē_^�|�F��V�ݶ7B�X�K�[���꽊�$�ײ_݀~�u��#<���3
��g9m��}ۛ������r���
4��*Z,�%k-(k`�E* ����RĒ[+r|�QH*FX]���݉�j�$�ײ_�$�v�RĒ]�܇� /���� w�|��n�&�
��I.�̥�$�we}�I#ny<I%��e��Ӟ{R�����l�K�v��*a�*Z	3rR0��̫����c�.Bq�'��V���S^]�,?��{:����߼���/�]�_��$���ū�����FZ1o}�_������T?o=�w��ﺇ@S��ӯ/}�$����!��m�+�n�$�og�v�RĽʻ��Y��/���ߟ�/qk4ͮD�-��Kܽ��RĒ[����$��؞$��G麢%�X$���]	�99�$��׿�}�_7��M��*ʅn�$��v�|�^Z��$�w���� ���� N{��(O}���:�tA�	a��k��W�tse͎�)����m�	��e����3
��������}�>��I.�̥꯮�[����$���*T�\��;g
= �y�s�����ܑZ���KII����$��؞z��.�Ǖ�7q1�B��`������ӯ/}�I'�V���z ?y���� ���|l�Vp�v�m�Ē]��C�H��O���{Ü�� ��k�����[o����s�ɦ��2��{� �߼w@ܜ�I͟�mn�����Ē]�2|�W]��9A������Q&� ��J�:�3�&f�,�lqy���n<��6A�8u�tͲ�v�.D���9v�(��g&�ri��.�5qR8�bpƚ��k3բ�l	 l�߻�S�,�D�X�r��&n� �J���#.���<i�^|��Όv�[���\Km��c�&�#�����O(�o�L�F&-ZG<\��=�������o
����s*MAm�4���NI䓒{'�>C��+q1���5F�XBV�g��:���j�.ܗ0��5!�[�p<[�ﾴ��V-�3�l���~���`ߟ:/@��C���m$���I.�/|��WV��M�u��%�s��ݥ���Im�<�ɕ��W8�l��i1]�aM:HV��� w��r�.ｕ�wo߯ ��v����Qj�N�y?�I\��ߞ����܋�\�R��yz��z�6�;�v�xݓ+ �9\�y|�?��xҭ#h��+&����͹���\Xu]=���c,��ø�{Z��y�rb��Л��l�As;��~�y`�0����W*�A����������Y���E�������]�m�f��0�h`f`Zf�L�fq��˸򅈘�i�,���(LDڏ�jOk|���}�rN~�����9Ď�Z��vL+m;0vy�vL�?s�+�U˹/��Ox��"���;����o�\��w���������ܪ�W8����/b�jk5sYl�ѹ'?g{w$�O�T;�~:'�<�ɕ�okJN�)7�@����b���4�!eud�<R�=��K ���p���NN��F�e�Ք�N�l��w�2��&W��s����� �Y���Ʈ�����0	�2��W?r��f�߲���~XwG�+�H��yz��K��݉[���e`�"��r�@��*��Ȩ�dAj�M
��W�Ng}���'���n�B J�)���t�7n�=U�^��,d�n̬W8���Հ{��^�8*v�[k ���{��'������X��XwD�������ֲ'b����.�3��v1D���a���>�I6�k�.��\��>���' ��2��Ƚ�s� �`=�yE]�N�n�`vL��U$w��,d�wfVz�����^�6:����m�]��;�������ʮW�s�~��e`>��ն������l��e���}���3�$�V�d�����++���W��00T��"bb�bY M*���.��ܻ�w�vz�j�[
��6`�2�ߪ������@�����;�8`��(�$��1�W����ny�v�O�r
�֧J����V�#����y$�#`s[|ev5���~��K�`�?W+���\��{����o��>�����:\έ������rrs�.�?��Xݓ+=\��W=�N�/U��uv�[k �� �ٕ���\�8�w���;����d����郥m������\�+�������6~���}.v�O��@�9�7$￿�n�fj��+n�`vL��*����\�o���t	=O�n���+��ʭ��]�UW�0��g�t�����Bff`��Hk�W��䶜� D"@���h����.���
��l)��[�K��Yp����i
msD��7M����K�B���IB]�0���]���M�@	 8v)@ȱ"2I#�"!4�rY7�6��H�HT
�mc"k�$MB��`vD�$��P�P����B
� �`�%eVXI$���F���!�%4j@��G���~	�A�7Z@�Na��o��!@ۢ��\f�Ye->�s���Nh!���<�KK!	�̇}��UUU�   B�*V*���Zꪠ*�[N    C�]�lWn[7���Lq���K������S�:��ݫ�fW��X&#�D�;�GN�pH��;���}�4=K�bM`L��ͮ���C�r�{\d���=2/%����;t�r<H&�X�Bܳ���;\������n��=z:k�%CYꝽ����9�8f��mq�]u���[$�%�r�m����=YD��E������l:�q�4�π�ntHj�u6���@@�.��a��O����`"�ƶ�-7��u�1�aU!̮M,QN��
�j0�[vҤB�,`P	��31��,�\Pt�άG�QHK�ղ�D�.��d&!AݓG�(���4��u*V#mq��KY�{Y�7�����s�;q��6!R���%ؐ�{b��ـ���(�.�)ck��@Q���-�H���M���L������t؊� W-�T�X�W\��6�d���"Զ�R��]<��;���ɵ�k��4��8�V=9]��r�����K���ձ�$�A��� `.�孞=�-;j&A�.�/baV^]�]�,}���y�Ɏ�������<�g�BO;=�[�kb�^i�#p9*��e�ʆR�t[�u�V7L���4Xań���qRí9w�4�[�g:����e"�fFқ��F��nC	ʴ�J�r��R�9��6m8�.EDt\Җ:���.C�ѫ�Lk�(�6�x���[v�(�zu��H�\
re'e����47e��rEV
.:��u��3eM�d�+�v�c�w���X��]q�)V�(c3`�l�ܪ��ˁX�s�e��̼�m��t�֬�]�gm���Y��¼�6y����.�ͨNw+�мc:�[�t<�J���^��r ��Z�|�r�m�c�[��d�����/2�Q�����<e�3]����fbN<�ssu���%��`�|�MgS$��35fdֵ��>�>SJ�ʠp@o��
?�Wj h�
��?��&*ESt{��P]���]W�Z��xn�/%��"sɁ�d�fh�HQ���z���m�v���t�s���q��f�,	�^��.h����̣[\L� �ԅq岔盪��JSR���Y����h��m��1�3�9��'k�f\1�=��\4��,����v���/gTm�h���e4�ݽ�藳��G��8�c�m�&͋��C�;��j����$��NBI�r}�NI+;�S��a�]IK2Gh�H�˓����}qp<Y��4If�Ĩ�Nrr.:�][i�"���j��^��8`ݙ^�*��A�������iSV���+w�w�N����W.�O~��6~���}{�w?y'����~��Yr5k�g���&V��s����w���^����`�EQ+��K��݂�X�r�l����O^��Ȱ=ʮR�=�`�z�sv��ʹ������O'���_6{+ �ݗ�n�
J);�v.�'��+��.�BTaH��Ⱖd�6��[hI�_�I<R%/&]6f˾��~�w$���ٹ'����l?�*�ı>��fӑ,K������᫒a�4\֮�f�ӑ,K�����!S���X�"2�#*��vF� )	$X1�(���M���Ȗ's���ND�,K��{6��bX�'���ӑ?�(dL�bw���;�h:95e�s:��������{�ٴ�Kı?g���r%��bX��k޻ND�,K�w�6��bX�'������2����N�!y9������iȖ%�b~�z�9ı,N��p�r%�`Aȝ׽��NNB�����~��F�e�m�w\�Ա,K�M{�iȖ%�`�����ӑ,K��;�fӑ,K���ﳮN�!y�^Ow��������R;\�v{pl���=�����qژp��C��i�'$���f�T�l�rwy�D�;�}�iȖ%�b}��iȖ%�b~�wٰ�F
��ı>����'w����/'��>��d�`�n��r%�bX�g{��r(%�bX����m9ı,O�=�ND�,K�w�6����bX�z���&�W32�R�ֳiȖ%�b~�wٴ�Kı?|{�6��cP긡Q0E$K>�m9ı,O���6��bX�'�	�r��&�p��u��r%�g����O���ӑ,K��}��iȖ%�b}�wٴ�K��AK����p�@�����b�L��Uk.g'��H�~��M�$U�}��z%�bX���siȖ%�b~���m9ı-���m=��`��:1%vLd[{q�ss�����'=�	16μTl����>�|�����W&�5��ND�,K���ͧ"X�%����6��bX�'�{��yı,N��p�r%�bX�w�5�CF����f�ֳY��Kı?{��ӐD�,K�ǽ�iȖ%�bw���ӑ,K��>�iȊؖ%�w��JMd�h�kP��m9ı,O���"X�%�߻�ND��,O���6��bX�'�w��r%�bX��e��F�U5�ι;���/Ӓ�@2'����ӑ,K��w�ٴ�Kı?{��ӑ,K�|/D:�� �F�B&J��������G�>AI�~��K�/'�ϩ=��j���ݙ�'w����>ϻ��r%�bX+W>������X�%�����ND�,K�w�6����/!y=������V���ϑ���X�\�����CT+!��uՀe&`��$�6��|:aT������{��7��/�w��r%�bX�}=�ND�,K��C�,K��>�iȖ%�b}�;f�[�&�tfh�ֳiȖ%�b}���m9ကdL�bw����Kı;���m9ı,O����ND�,K�}엚���h�֍d��iȖ%�b}�}�iȖ%�b}�wٴ�K K���{�iȖ%�b~���m9ı,O����e�5�Y��D���ND�,�>ϻ��r%�bX�}�z�9ı,O���"X�+b}���iȖ%�b}����kS$њ��噬�m9ı,O�׽v��bX����~6��X�%���p�r%�bX�g��m9ı,L�|�r�/9)/R{	���UU��+[f�ͷj�� �ڈa����C�ƻe��.+5ϯ+�ë.���<7[��[��' l/!<q�3��=���'�\%:�-��ۺ�:�F��I�[�����ӮMت:�rh�uی���i0�@`v�ic?�p7M�m.56����� BV8��[���>�<�s��^�j+��mq��֟,�c\��ݸ犍tm���Od�ܶ�snţ��.�[`�ѻ�x��DΚPjիR���r�zԕ�,���2����/!y�����6��bX�'�{�6��bX�'��}��Kı/�{��r%�bX��}��u�.�M�rwy�^B�}���i��r&D�;���m9ı,K��kiȖ%�b{����,K���\)t�C5��捧"X�%����ͧ"X�%�~���ӑ, �,O}��6��bX�'�{�6��c�^O}��m���6�i]�'w��b�%��{[ND�,K�x��"X�%�����"X�+b{;�fӑ,K��Н6Zx�P�35�u�m9ı,O}��6��bX�¬S����m?D�,K�=���r%�bX���m9ı,Ow�Y��.���k$�ּYo&��˭�����]N����v���`�X�N��&�9����͗��9��y)䧒���p�r%�bX���ٴ�Kı/�{��<�bX�'���ND�,B�~����c�V[���'w����b{;�fӐ�=]�#��W�2%�{�}��"X�%�����"X�%�����"��C"dK��޾�����l��������;���m9ı,O}��6��`%�b}���iȖ%�b{;�fӑ,K�C��%�RWUa*ۃ'\��B�H؞�Ǹm9ı,O���m9ı,Og}��r%�`-�����ӑ,B�����q�5]E�#.�:���,K��ND�,K�׽v��bX�'�k޻ND�,K���ND�������a|�� �,m�V�M��1O�� ��צ�we���f4�J�4&����I:ف��SY9�̗4m9ı,Ow^��r%�bX�}�z�9ı,OwǸm�Kı>����Kı=�<��ئ\mZA�:���������^��r�r&D�?��p�r%�bX�����"X�%���޻NAE�,K�I:l�x�P�ɚɚ��r%�bX��p�r%�bX�}�p�r%���$HH��"�D7 �T(��*�Ȥb�$@�Dj,X'��!�P)�MD�Ok^��r%�bX����N�!y�^O߽�S��qf��ŝ'"X�(X�}�p�r%�bX����Kı>�^��r%�`"�"{���m9ı,N�O켳�ɫ-��듻�^B���}:��KİE�׽v��bX�'��NND�,K��ND�,K�������P�Ќ�o9�����]��ˀۆ�:��I)jD���P�Jk���u͹S:fj�?D�,K�����9ı,OwǸm9ı,O��m9ı,Ow^��r%�bX��zOd��\։&�$�5v��bX�'���6����bX�}�p�r%�bX����Kı?}�z�9�P��"X���5v�ّ�E�rwy�^B�y�p�r%�bX����KlK����ӑ,K��|{�ӑ,K��w�=���Ӛ��sFӑ,K�=�{�iȖ%�b~�^��r%�bX��p�r%�`i�Кx 	�r'��ND�,K�CޒsY���\ɩK��]�"X�%���{�iȖ%�b{ޞ��Kı>����Kı=�{�iȖ%�b(?M�}q��.�W<�ס�t����qu�$�sZ�Mu���$!�eyܐz u)�J�r��\��,K������6��bX�'�w�6��bX�'��z�ND�,K������^B����}��&-�Y��θr%�bX�w���ı,Ow^��r%�bX���p�r%�bX��׽v����"dK����x\��5��ղkZ�ND�,K�����r%�bX����m9ű,N�^��iȖ%�bw���"X�%���o��Tѣ5�nI����K�,O���6��bX�'{�{Y��Kı;���ӑ,K�����ӑ,KĿ��=��\�kE�Z�\�M�"X�%�����m9ı,����Kı;����Kı?{���r%�bX����|��~z��6��f�W]	��q)��mvQ�#�8����s��\E-'dTպ��9�ݫ��T�*��1m� ��:�:۬�I��'�z�-֛v��f�MJ[�q��nٲ��L�&
��k�Ӄ���9$�8n���v،u�I���9�t�ƌA�n���ͮ2;9��:x��A�5u����l����kq��/ =���]3kG1f�D`k��Ϲ��Pu��!��R�fW,.,�l5�(����׳�^l�y�آ�qZ���]�s�Ql˵�wܝ�B������ι;�bX�'~׽v��bX�'�{~�D�,K�׽��r%�bX�������Nk2e�ND�,K�k޻N@,K���o�iȖ%�bw����ND�,K��m9�2�D�=������H;'\��B��������IȖ%�bw����ND�lK��m9ı,N��z�9ı,O{���V�-]�듻�^B���}siȖ%�bw���"X�%�ߵ�]�"X��(�"}�����K�/'�}>׸��qfV;e�rwy�^'{�p�r%�bX'~׽v��bX�'�k޻ND�,K�׽��r%�o!y>�����Bbl&�k�7hu�Q�].!��.Ҍ.tg/`���+qjr�]����'��/!y���rwxX�%�����ӑ,K��u�k6"X�%����6��bX�'{ٿK�SF��2�&f�ӑ,K���{�i�|�<@��1�[�@a֥�%��na��ĄI1t	�D$#()��r��჈��"dK>�?��ND�,K�����Kı;���N��/!y�y��D¥�n6��r%�bX�w^�fӑ,K�����"X�\��=�]�"X�%�����\��B�������w�j��fu�fk3iȖ%�b}���ӑ,K�����ӑ,K���{�iȖ%��'�׽���Kı;��K�N��f[�6��bX�'~׽v��bX�"��z�9ı,O��{3iȖ%�b}���ӑ,K���I:KI��5f�3����3nT��]]Vǉ�+8�8+�9��B���'re��i]��'"X�%�����ӑ,K������Kı>�}�a��S�L�bX�z���'w����/'�}���a[��Y���r%�bX�t׽v��bX�'��m9ı,O��z�9ı,O���6��� ș����5rɎ�f��蹩��Kı?����m9ı,O��z�9����s	��eM�4z�5,��)/k0?zS�?���}HƖWe�m'ܤ�)͉!m�&s4�Vݒs0����&�sy�B88�8�N�㎙*h�� B U�@�SH���XH�	!����hO�W�bB1�M�Dx�������\B^50�a��І��07xÙ��t�6&�VX��϶���C�r�#	����3z�>%��`f\'Ex���D:= �D���6�.�:��9�*Q��W�w��j�C�0~M�|"dDGN�@� `)T�X��s�w�m9ı,O��ߦӑ,K�����ˁ�9����N�!y�B�y��\9ı,O{���r%�bX�w۾�ND�,K��m9ı,N�ٿA]��jb�rwy�^B�{�^ݧ"X�%�}�z�6��bX�'{�p�r%�bX����Kı>��^䏀�!+��f�m̤b��&��y��gA
�l��]돻�_|8�J��l�sSiȖ%�b}�n��9ı,N����Kı;�{�kȖ%�b~����Kı?x׽.�5�.�ְ�ˬ�r%�bX��}�iȖ%�bw���ӑ,K���o�iȖ%�b}�z�6��bX�'s�-��at�ֳ%���r%�bX����Kı?{���r%���ș����ͧ"X�%��{�iȖ%�bw���3��u���S��]�"X�b~����Kı>�}�ND�,K���6��bX�$	��������z�9ı,O{��/MjfkSZ�kSiȖ%�b}�z�6��bX��{�M�"X�%���޻ND�,K�}�M�"X�%��'�����&�9ݨ-�%�R��Զ�3,N�1qJ&�H��w1��`��6�3u�4Y���9��ı,N����ND�,K�׽v��bX�'���6'"X�%��}�ӮN�!y�^O�{}�f�ȡnu�M�"X�%���޻ND�,K�}�ND�,K��w�iȖ%�b}&x�W�9�r��G*l3�m�:�0V�I����Kı;���iȖ%�b}�n��9����ߦӑ,K��u�]�"X�%�{�=�]e��e�Z�s3Z6��bY��r'}���v��bX�'����Kı;�{�iȖ%�bw�{�ӑ,K���Ozf�5p��3Z�3.�iȖ%�b}���iȖ%�a�������v��X�%���o�m9ı,O��_fӑ,K�O���^G���m�͛l�U�@%;7����g����#���|�O����3�s	��a^9�E�+�n`(�dK�Y��mmr
W����e�n�@H��"����g���"Ф��:��L��y������+O;&�=jq�`�L@6���6ͧ*�Ucv��3���,H(&��M��
�Y�Ӈ������j����WdD�[,_�E(�!�4��� ���%�~sE�4]����׷3O�fzm����`��R\�kR8�zH;�k]c���r~���/!S�k���r%�bX�����r%�bX�ͧ"X�%����M�"X�%��{g��{2gk�n��u���/!y,N���m9 lK��u��m9ı,Ow���r%�bX�������/'����+vZ���N�!xX�'{�g�iȖ%�b{�ߦӑ,�	�2'�����Kı?������/!y�����{��4Y��6N�9ı,Ow���r%�bX����Kı=����K�lN�k޻�����������R�f��*�v��bX�'�׽v��bX�+ｿM�"X�%���o�iȖ%�b{�ߦӑ,K��N˳�3-�If����	�mnm�4�,FFds]���t��wD�R�5�ML]��N�!y�^O~��6��bX�'{=�M�"X�%���~�S�,K�����ӑ,K�{��u��뙋���'w����*w�^��r q~% ��0+��ʠ~r%�bs���ND�,K�k��iȖ%�b{�o�iȖ%�b~����8�̻Z/\��B������^ݧ"X�%��u�]�"X��b{�o�iȖ%�bw���ӑ,K��wž�d��iֳ%���r%�d��}�&��	ｯM� �'�N�I�$�z'���m9ı,O�x��.�V�ɩ��f�ӑ,K���ߦӑ,K��g�ͧ"X�%���~�ND�,K��޻ND�,K��ޒ]c�6커��>^��=<]u�ꭁ���Շ6��5���L�6{^�1�0��j*޹?�%�bX�����ӑ,K��{�M�"X�%��u�]�Ȗ%�b{�o�i������߽����E�,J/\��%�b{�ߦӑ,K�����ӑ,K�����ӑ,K��g�ͧ!!y�^O�{�z��dR
�듸�%�b}�{�iȖ%�b{�{�iȖ;����� ǊH�'u5�]�"X�%����M�"X�����/^�躦����:����ı=����Kı;ٯz�9ı,Ow���r%�`��u�]�"[�^B�{����ڭ�3�'\��Kı;ٯz�9ı,�{�M�"X�%��u�]�"X�%�����ӗ����/'��R��;V-�te�=���M�-�p�Ȕ�2�n1��e� A6���0��u�f��&f�ӑ,K��{�M�"X�%��u�]�"X�%�������@b��dK������ӑ,K�C�~��i��.�����/!y���޻NDı?{^��r%�bX����6��bX�'{��m9ı���=�[ه!v��vN�;���/���]�"X�%���o�iȖ
ؖ'{��m9ı,O��z�9�/!y=��t�|·e���rwy�g�L��O�M�"X�%��{�iȖ%�b}�{�iȖ%��<@��l7Ț���Kı;�����Z35�V\��r%�bX��w��KıA����ӑ,K���{�iȖ%�bw����r%�bX����悚�τB�·0��5��rv�!;����u��8�1��ɽ���'}�F4�,1ڭjm9ı,O��z�9ı,O�׽v��bX�'{5�]��!?DȖ%��{�iȖ%�bw����Z���W	rfY����Kı?{^��r����,Ozk���9ı,O{���ND�,K��޻ND�@9"X�{�>�v�u��6��'w����/zk���9ı,N����r%�bX�w^��r%�bX���z�9ı,�������Al˵�'\��B��9��?�ӑ,K����v��bX�'�k޻ND�,�Ac�=���wy�^B����ƷGX�v���ND�,K��޻ND�,K�������ı,Ozk���9ı,N����r%�bX���7'FD� �@�ʁB�B$E"�U�����Nwo��l[�
�c���	�t6��J9��Pհ�]���҆3Hˮ��l�+�Q�60#q�8�ll��.��5�g�+��gf�y�g�[Ĥ�nrsx)��C���v�:��x6��;����=�zK��p6�kn�f#	���Jl=[�vQ�ng�s��\�����[+u�2��r��������Q�-*�8�Y���Pn�����#�U�(���$-��XIl���d��n���R���n�su�r���P΅��3��×Қ7A�:����������N�9ı,N�k޻ND�,K���6��bX�'�׽v��bX�'��ze�i��.jf�5���Kı;���m9�"X����6��bX�'}����Kı?{^��r%�bX����;���l�)��'w����/'{��m9ı,O��z�9ı,O�׽v��bX�'{=�M�"X�%����{�^��rd�U�rwy�Y!��޻ND�,K���]�"X�%���o�iȖ%�� G"{����r!y�^O<���R.�4��퓮N�ı?{^��r%�bX����6��bX�'{��m9ı,O��z�99�^B�{�ïq,n��q�Qu#�h��v���;���^�*�E�%f�ugc�>�}]2f���35v��bX�'{=�M�"X�%���~�ND�,K��޻���ı>�����r%�bY��}ﮚ&��T֙�rwy�^K���6��߁W��6��D�,M{[��r%�bX�{]��r%�bX����6��bX�%�|e�a0�CN��-֦ӑ,K�����ӑ,K���{�iȖ?�C"dOzk���9ı,O{���ND�,K�C�$�5��Ytjau����Kı?{^��r%�bX��׽v��bX�'{��m9İ��޻ND�,K��o�2�YsS5��]�"X�%���{�iȖ%�a�	{���O�,K����v��bX�'�{~�ND�,K�zK=���kl�������WAbA�C���͙����r�t�����|�N��完�ӑ,K��{�ND�,K��޻ND�,K���]�"X�%����ٴ�Kı>���e��Y5�sT��f��"X�%��u�]� �bX����m9ı,N�k޻ND�,K��m9�,K�뾷Z���uL5sP�Z�ND�,K���M�"X�%����ٴ�K @�A��c�"�#+	1"��D����"n'���ND�,K�k���9ı,Ow���Z.d�3D���M�"X�)2'�����ND�,K����ӑ,K�����ӑ,K�dO����6��bY�^O��}t�4̻\gu���/%�bw�ߦӑ,K���޻ND�,K���M�"X�%����ٴ�B����~l�綁F[.�f;Lv�N���Q�ƥqE�jL��p�,�	�s}�w��~��cjz����������\9ı,O���6��bX�'{5�]�"X�%���~�ND�,K�C�-��T�xE�:���������޽�'!��Tș������ӑ,K������Kı>���Kı=�V��,�e�53Y�jm9ı,N�k޻ND�,K��}v��c��0Dș�����r%�bX�o�m99�^B�{�wk��Y�Ļ'\�ı,K��}v��bX�'�׽v��bX�'�{~�ND�,$D �0�h� Ĉ~v����'�7�]�"X�%��Ǐam�ɭK���f�v��bX�'�׽v��bX�����M��%�b{�_��iȖ%�bw��ӑ,K���K��9eb1��iuջ�5In�#\˃�vuw^�R�xո���v
-	�6	���,K���o�iȖ%�b{�^��r%�bX���QD�,K��{6��bX�'��w�MI�n��Ra2�ӑ,K������ED�,K��}v��bX�'s��m9ı,O���6���S"X�5��ٓ\�Z�ֳ$���r%�bX����v��bX�'s��m9�T,K�{~�ND�,Kޚ��ӑ,KĿ{�c�)���ڎN�;���/ܜ�Y5Ok���6��bX�'���m9ı,Ozk޻ND�,lOw]��r%�bX�z��jfkY���n��ND�,K�{~�ND�,Kޚ��ӑ,K��{�M�"X�%�����ND�,K��X��FKϴ��>�1�*�N
�;����nW$�JA�P H�),��b����Cc�Q�#R
	�q&�!�v�p��"�KF�����	�fl�@����0($�,w�������'  �   9�� o$ �m�  �� 
�����o42�
���n��$�g���5����ιѽ���_.z�B-ͳ��q�<n���9݊�����g�&�:��s,g"bNl��ڂ6�h�:u�cz�X���l�n���TO	���u6m�xj��%�9�s�܌K���YyaƸ���:nD�nc�D��C��n��q����Slgggb7g��O&�V�U�g==L\�J��%q=�B4��:�@6���^\��Cu��6��ݵ������"��],�gXmUa]� t���b��WYi'�*�ET�NUs[v8곫�n\�����st/)�i��Y�h$H��ٶm�f��Z�� ��m��]��*����Nx��k�X'��xpr�ز��w��Ν�(�#�u7���b�c�gx�9.	�(�l����� e�vua�-�J�ҍ%�is�:Vm�zL��M�j��Gn��k�RP'g�=�<�ݹ#&�Z��.y�s�9���6��G�����52�r!�dc%խ�p��ؤ�Xq�L>����r�����x�r�ñ�mi���D���[u���,M͚y����%���CV*�V��\��l����A�A�i���D7i�N��rl�c(-�]s����@V�(����ҙ�����8����+,��V�9�c���q��d�v�= �],rijH��.PZ�9�W@me#HX�*.V�*���t׃���6��Ԃ�h��'Oh��҉�9�iL�N������N��8��qk���M.�ʬ�W�Y�J��2d]���S�n)6J�J�ىq
��
�K��rm���g;j0K�A���SÛ]3�$�v�'p��a��UxU'�F�q��D �y̍�y�#����zcNZ�U��x}�x�#]��n�zy��IۈUܢ�h��-����&@C6�)�g�9$�'G9�)�O� 4!��RPP��	�	υ������@(�P�/\MTڿ��I~�U�N�����u�2�C�r]��<�����$9���cpDq�'/��3�*�@Q+(fݶv�ݩ6ٳ��ў�,��\���v�x�Ɂ��#�5�u��X����hi����HPS�Ӽs��]wo`�e5����ȞF&W�m�O!s�v��T҆Q��	�]�tݣ�O����nu��u���^C������.�J.�s;=绷��[��> wb�����#u�C8A�L�&�TZ-X�����"]q�	�9$2�:��aJf�V���bX�'����ӑ,K��{�M�"X�%������"?�dK������ӑ,K��������%u�.j���]�"X�%���~�ND�,K��{6��bX�'�׽v��bX�'�5�]� ��bX�t��-���kR�3Z֦ӑ,K��{�ͧ"X�%���]�"X�%��M{�iȖ%�b{�ߦӑ,K���߲�kXk&��W5-�k6��bX����]�"X�%��M{�iȖ%�b{�ߦӑ,K�;���iȖ%�b{��~�R�K�&jL2�j�9ı,Ozk޻ND�,K���6��bX�'��޻ND�,K�k޻ND�,K�|Hw�rDn\�i���n�*	�B^�Mm�f��K���O��V��=����]�"X�%���~�ND�,K�u�]�"X�%���]��?DȖ%����N�!y�^CϾ���m�)����r%�bX���z�9O� $I�A�Q���*GJ�%�b{��.ӑ,K���]��r%�bX��w��O�ʙ���?��.�M��d듻�^B����:��Kı;ٮ��9���{�M�"X�%�����ӑ,Kľ��{J���u���/!y���۴�Kı;���iȖ%�b~���K����]�"X�%����NĺS�0����'w����/'�w~�ND�,K?w^��r%�bX���z�9ı,N�k��ND�,K����?�����X�ϋ,����4S�똊�.4e{&�]S���Ӟ�j���fr�9H�#��������_��'>������׫o�|��]R1-�v��>��?W9��8�!s� �?m���ï��@��=��Hl�).3w$�fw�rO��]��0;J�@2H!��������_���ܓ��]���?���n"h-�v�d�߹�$����ߌ}�,�0��, �ʻR�+�ʺm]$ـ}�"�=U��w��!s� ���(��Q�˶�T6�a�Ls�m�˝�����l�%��a���uvn�P��l�:�L���z���oz��p�Us��e�� =�*G��c�![-ݶ���,�_���U]���� �_�� �\�?URF�x/Eи�Zm;.��$���܋��W9Iw��,��}���h��3,2���y$�^�X}~��>�0'kՕ�iR�Us`B	$"F"q[������������0�g��c��M[.�}.E�}�8`��}������T;����1b�n�Ka��Ql��1�����;`�h�M�D�V����8ε����超BV��; �`�p�>��X�r,Wl60����Vݖ�f���*�ʤ���,���}�8`�Y���e]6��l�>��X�r,=�s�K���?�I@]��v��wVݵ�}�"�>�0�`{��.�X�yW�N����l��}�8`�p�>��X�r,s��>�=��;�*��I��*��Қ�O5"���-�tk��=K�ip���mR�9G�c�Ƽ[�Ec1J�sF�J��[�G9z9�.�����γ�=K�Mʙa^ٙή]N��R*=R���qӣjyL�v��U�.:;t��I��3㴝�.��5�B;fY�nPe�h�v�v6���5k��=a�l�A�c)mXKx$/g]3gv	�xyl=��z?��?7f>A,�a��ð/#��p���䧙���
�O��n��4�f3�q��mP���#�}�ذ��_���s�I������m���-�ks2˛l�>��X�r,��8`�p�ܯ�6�}�O�WGTbf�������T>�0��K�p`}�ذ�/l���Z���}�d0��ŀ}�"�%v�c-SWM��vZ-�w\0Uw\��������m"��6,ihb�]̙���,Ð7e9]�������р��S-��Rh�N���� �nE�}�8z�A�?�T���κa�.o ���o'�x�f�M<���;z8`��}5�?W+��~��W���t���7m����w\0��`mȰ��^[V�q��mSE��9\�˞�ߌy�0��X��[r�t�An��[m��\0s���_$����������S�z��cmp.�����S�N+��ݛ0Z�ۛ�mM�n+�tp�7&6O�}�����0�~�>A�G� �J�~mZWV趒�V����~�����=/�X�r,��r���a��,wcc-ݖ�f=���;.E��~�;EB�#�TU@�BF@$@�,D�	�++���Ϫ��/�X�� l�՞cj�h����~��C����[���` ���[&x�=���,�j��t��X�r,�+��T����#�}��o ���@v�X�ģ-n���3��x�I�eBۖg!`�i�O&�Xu�����X�]�BJؚ���'�?�`nE����U|�������^&��q��mSE� ��mȰ���	 ���$�����~��Z�!�N���X�Ix�N�`F)ci�ƛ����=\������x����'�}����Y��#�"v2�Ո@�@�����n�?���v3�avw ｏN��y��O%{����?z�~X�IxSR��c�n�����>82C�Mڞ�K��ȕ�f���/az
V�25KeuV��4��=�צ6�X�I~����������;�X�WM���0ˑ`)%���0�p�ܪ�W�r�����ߨ��ݫ�Гw�j����Jp��s�����<��^ IN��BJؚ���*����I�)%�~�R��޼o�Z���\�Z���ـn��W9ʯ�U������߿^6k���9��⑋ �@��
+%�������M婠1+m�a���L���]I�[E��ϳ�-�R-�^�&�&W2���;ϒ�����R���V���2[pXi�
��|�!�FŎ�<��9��;J�g��-����M�8�n��F�{&r�rێ���Y�s�[)G��g����y�.��]S�,[cً��|�]W �����5ic�,�hb��E�%\�M[a��I�ry;�ϡ~���S\�8��e�]�����B� ����5�5�^n�n:�ݟ.��fl�U>������>^�^6���G� ��Խcn���b�Qv� �I/?r������7nyao��y���y=T�Ȓ�;�o��� �ob�"�^�엀}Rȣ'i��M+E� �ob�"�^�엀M�� vB�5t�l��դ�)���d�v{{�t�g`KF�0�̒Ҙ,&�� �P�k�f�e�9��{sL�r��&��,�a���V��:�޼v{{�x���J�		[�n�	�8gk�#��� 5M^?t(zns/�XW�� �vK�ܮW*�"o�Zƒ�-���h�`�<����|�%�`�vZۜWM�uv�ݶ����|�%�`��s�Uɞ��߯�EtuE�����y����I$�O��7ny`I/ �*�[�g�QM<�6Wd#����z0m��x�r�h��Y�;Ir�����w��
���ag�~���0��,)%��s�[�^���[H8T�q��շ��~���@��{׀uo�x�8`d.�KWc�]6��l�"�^�^U]�}U���8j��2M^���ք$�B�.8������U���en�"�v�ڙ����8\�� HLf~%�.%�\��ٕI�Tٗ4]oR�.ٛ5�Zܩ"�`\&b�f!0�o��;O��4��F403I��hL�?�XCDJБ�)��BbͶ�D��y��kO�lI$0!I�IA���)
J��YJ�$�����U�#a
� F�a�E� �1"
B\(R����d&�il�i	B$%(P��h�Ȓ$)[
�勢
B�l�"�w8V4#`D"Ō`��V-�aaF0C�������&�.I(���)))���$����F��
�) ЂUaL �`�X�9�Ù�6l�R,V$
(B(XZF��! �F��$,�
X�h�4d��5B!$!�$0�B|�?�B���8�� >M��/�a�X��A���?�Y�xu覃�-��68` Qw�7eՎ�I���_��������?���RK�	"�X�[�!+b�m�6�$���z���x�D�(Yz��[8[���V[Jq<U�['_����>$w0���WA�X(����Fm����)%�)%����zx~0B�w�M���e��;{��|��%��=��=<?w\3�9ďz�Iz���ƛ|.��^�� �w\0���M�N6���(�B�+w������7$��צ䝽�sr��TJ1h�`:48�T�hC?_��ܓiJRS���6�ZM]����)%�-��	��X�UUV�(Jx�����nD{O\��g�����z��l�֞r=�W&�v��p�����묺�3�����-��	��Xv�,B��w�7auct$��-��ܮr�=<{+ �s� �Iy���H=�R�:VĨV�i�x��e`�ذ�U\�K����^�� �eDc�/��V�47X��#�X����>RK���s����~�p��_��)��32�ռ����)%�a2��ذ��\�mW%��s�OC��U[1�Qm��q�\2m����)�), �u��K���d�^ޕ�����l���Gf-�n1�nw�#��=����K�{c8���m����o;mӋ�a����R�f����q]N6!�ton�X\�ݻh�Ƚ띷bMXx���hX�����i�g�{k���O<��g��n�ar�۷a�:�v�q9wZ���p�k5�ms��6A����8�s�7'']Q�Kh��f4�;��Xr�]q.<-����3���a�0��I9�C���e�j�|.���߿^6+ ���U������=9��ڻ�l��
�v� �	��n�������U\�~��*���>����
�mVum��_�V�I/�Uĺ��^���X�t�Wc�]���ف��������xW���&�e`��HT�.���.��I&� �I/ �r������W�I�);��I�{�׹�����e0)������̦�V��[���r�{u4��8�-��.�m[w�M���7u� �I���{׀v{�Xһ��e�t����7~�f��Bn\"H@���c�k!R!-T�HX[F�jK�����p8������;��~���ra2�	�ꔇM��ƮـE$��$�=��U%���X���$��)7t�ݴ��v��Wo����=��n���*�������~c�V�E�Hۼl&V���L��S޼�$� �n��J�t�R:wC�k]`3m�F��K�JRk�Q�ช{a�ra�WN�m�����w\0�K�>RK��s���e`�´yZ0���fv^�^7I��n�z��=����n���t��xW���&�;�pS�$VAH1�7��L��,IJ�U�ݗl�����UR���	.y`Kذ?W*��v��^�{Ŭb���պT�l�7ob�=]�_��z��0s��T�<4rr�Ɏ�g:��[��7O�%�1V`�I�#]��jU�~�:�u���sj:��~X�Ix���X��T�ݴ��+k �I/=\H��%�,�{~�F��'�:��eШWn�	 �`��a��w�<��{׀J���N���Ube�l�7ob�>��`)%�}���⪕���0aa�B����,dbV�d�B�[�~��CQԤ,wL�RVRknݚ$!7$H�w�����v?� ��J�wc�E�Uun��>��`����$�w\0/ܟ߯-����c���#�R�h���v�g���c�ΝH�v�0�n9Jt��=��9����^�� ��� ���{$�*��+�.�m[w�n��n���� �I/>�=U�����;���vUұ��y�0��`b���;�Æ4�S��v��6���0��X�Ix�RL�{��/!�M�6����|���n��n���>�}۹&�5 0 ��G��UV-A�m�Uu�r�5� ��`�NT!��W��[���|װ�k�#f�'a���k׶vz��
k�nm�Ylf�t�f�MJ���c�k��)��M����+�9�����ȋ�`��;vDz�l����{<�n�c�<IrF�B�(Ǜ	�
�g�]�	��-�J��l�Ol���7�Z�í�[���l��Εl�U�I��<.q&�����{�ߟwۏ�~s�]�(B:w<�LXvh��sW=hP�L�GGmsX�:�gv��۾����n���>��`)%��B�N��m��2�`�2���X�Ix�����]yZ�eիu�w�<�����0ݜ��'{���,��r���IK��z�	 �`ݙX��,l�-,E��ڶ&���7tp�7�2���X�l� ��Ud������Wn�,lsl��FKu4�)�a�C��;qŸ.[��R�W[拙�L�߾���|����|���n��JZ���E�-��Z7$�s���
S�e���� �ٕ�Iq%�M�6&���>RK�7tp�ܪ��%�{+ �y`�uwn��P���7tp�;�2���X�d�R��m�WM�V&]����+ �^ŀ|�K�7tp�=\�R�EA�Sj�t�&�bN:��K[vrˀM�ٙ��7g�\tZH�	��jWQ.��R����ۿ� �}�w ��� ����$*Ab�Z����V��>RK�7tp�7ve`Kذ�JZX��+��lM+w�n�2�ݛ7;�!�&�3��Z�h(`R��@�MvX�1ZU�+��P,R4 F� � p,��F�Fg���ܓ���nI��ZX�;�˧v�顺�7ve`Kذ���S�SM	[�۲ݷXe�X�Ix�\K �ٕ�{�ҽ4��\X8k*���*��ͳ��	��57>��۷O���4����Eb����>[%��q,��+�9���,z����նQv�]	�x�\K?r�6Oe`�X�r,�+��H�/�&�%t�Ubb�i`'���ذ�UĽ�~0	��, �u*����c,.�`��`�� ��`,�YJ���� ipSp����x����Z����V��'c����&���;/b�&�) �����I�c(e�8�R$2��[�Z�j�چ\N���q�x��ٛMk6K��F���}�����+ 콋�9�����yy&�k�M�]�X�`��`H�ouĳԐO{���E%n�n�wl�$��}#�ٮ%�n�%�%�ڦƛum[0?�K��x�7��,w\0?)=�0	�$��j�m]Zm�f��7\0��N��p�lt�їM���wz^�g��~�������_��C����ٰ�0����s��|E�ȄH�@�]!)���"V���@cH\ٺ�ѫ��C|���6W�ֿ~�KPR�LS$!a�t��bK��3D�/ �1cB�2<�s��9�0����@�p�62怔��ҏ��i�F1#9	�����g7�m}�M!�"bs��q���Cp�҅R	��		�0"B#�&�h71at�b'x6x�01�- ��*�b�� ��AzL�	
�����~`97#!�5 �	v<�?FE�/�|B�x/U"���3dX��`oRl&�%w_��7@8���`˜~B)��ф�o�*�}
}��H�c
HHA�,# M� U)`�)HȒp�y���2���(K��3[)h��o���� m ���ͶUUU�`��P� $ Ӏ
������g���p��R���;���E�
��s�3�m+�ën6�vP�����O3����֎����8��0��2nӅ�m7n��G�n�l���N�'3�����`#b.ڶ V��A1q�LYX�Ыph�+�|�M\��@�P�5RV����k�ikX�����H�\]�4)35*Į;Y����|Ŕ��� �y�U�ؐ�u���n	Z�Hp��͑x� 3q���b�y�v�uu���K����:�n0��nzg6�Շ(��.6af���]�01[����Ӻ��s��4�o�V����W�q��0�g�u����i4���k�;{�#NvZ��85Z�'N�y�:l�]����.%�ic0ٻx�m�
J�@\��vm&J�яr#�fN6ݑ6bُu�h�`�=r�gs���T�z	6�N����������S\s�Gl�d�-�s9fb�e�Qk[F#�Ԫ����Έ�J�MY���]<�=�tZ9W�ԩӇl�:����2��&�Y�[S���u�ܛ��=���T��cqȩ�R[qoimI�[r���H�=�0����0b��S#CZ����ݦ��rr���4��=W[74�	��c*�����!v���`��s��'[,m����x+I�&�Z�4��K(5e����;e�`��P�19�����ɞNe8�-{]�Vtp)�'n��i8ݣY�;&{7e � 
Űs.�i�\����:%k'VBm��`A��qW�Pq��L���2��Nʹ���W<-�p.e�%�'0��B/3*��-�XD"������Ѫ���N�B����s�a�8�݌��0琨`B]���)�1�K�<sV�s	dA�������؀��̖��������ˤ�:I5K�U��k�����Cr���V�@n��,*1b�d�\���h��.�U|���!�PL�j��C�k�:&��|�:/�â�U�H��@����S�!�� !Ӫgfs33���f����Z��flqȨt�'j�l1�jڊO>Xݠ�\n����+�<�ήCM�vrt�M��n9�Z��R��ڃ�칌�i�xnyu��F���b�cOEV�6.Ln��ԽM���*����V�Pr�uGc���v��K���y$�Ţ �'��+BT��f�-c�-U��.��)]�t	����M�(����S/��K]'|��94nBW�c,���ܝ�y��n��4��ef��n�\�x�=�������%t��I�v��7u� ݎ�p���~K ;�V���am��p�'c�ٮ%�M�� ��+��I��t��jـN��\K �{�0�J�U��.��Z�`��X�ذ�ذ?/o���x^���Mr��Z�v��&�ŀ~���_���ouİW9��^��0�;XZ�t���r81qH��T�K:�I�T�=��0���V�ݒ�C��X�p�7��^�r���K�X�q��Li���1[X�p��+���?�T(�Mg��]�9�}۹'��ŀn�8�+��M�ui�`��m�Xe�X�p�%(J��I:le��ݻX�ذ�ذ	��n�˼ �����`+`�Xe�X���x�	��X�ذۤmN۱`=pa�p����۫؎mu��f�-b�2�Z�f쫑f�痵����	��ou�`ob�s�ϐw�<�	=^��v�v�]5V���Y6�,�{;0�Ebh��t�R��"���>�ᄬ�Wj�G*����SD�& D1L��J()3{�]��s�;pIJ0O��E�m17x�*�}3�����E��s�׳׀{��z�m1��t˶`��ou�`w{�����~����Չ�Ѷ;SI/�l���ב_m�ݛ��9��]�̻�`&ں��0�,.���`���v�'M��Wl�"���Us��q#������� ���.�`+cv� �k�;�z��)���<�z��B�����U�N��f;��\0���6� ���4(���rnI�~;�,ٖ�v�]5V���\0�����`��l".�J�����`�C�Z��!�b�N#u\���O�t�;��`֗�Ր�.]7V�]��<�z���`��ou� $����n�N�w�}5�?W=���&�� ��/=I���7t鱱7�v���w\0�8���^��� �]ۺm]Zm��`��`�2�	�p�6��q��'M�V�����X�̬w\0	�p�*����:l�t�.�����Lm��sub��vゞki�`��B�S���7�F8�]a{,6M�-a�m�9C0�[�;B��Y9���l`�v��j^WY��"��H��,�'�n1s�91';fw�4n��e��m���GV�n{58����d���%�1��ל�ɛ�f������Ua��[�jݭ��y�Rʤ\�to�mK0��IӬ��h��Mu��3vwl�ɸD�[ٴW�� ���Mn�vQ�M��eX[f����'c�;��`!*��:N�U�N��u�vk�;���X�̬��W*�6z�v#*�vZ�h.ـ{c�onE�N���;5� ޒ����V�"���X�̬�\0	�p��J:�v�Wm��k �l��;5� �����W*��W��WOj�]8�P�z��8���.���L�Ÿ��vl���QmX�π~�����v�/s���ag��4�݂n�զـN�>q�����6�� �0��B�)�� \����'{�vnI��jҒ�:wBt�Ui�.ـN�ŀN���'u� �� ���.�:��-�X�̬w\0	��N�ŀvBU��t���m:V��;��p�'ob�'d��>ҭ	iDV׭���LΔJ����n�0�8뚍9n�5Ӝh͸�mlv(͓lk�f�8~��N�ŀN���'u� ��QyC"�;H�f;{{����l�V��;�$�$���
��mnI��wf����70��؊b�@��A~<���nwZ�ܓ��*F�(n�66&ݶ�w\0����X���\D��v��.��`w\0	�ذ��߾���ޅ�^�6���+��bѶ��X�)z"̂i��QJ-�1��J���էh�f;{�u� 'v<�� �u]�.�:��-�Xۮ�H&�`}��ooFۦ�w��[at�um[0{#�>�`��`w\0�v�Ytբ��H�o���w�'����I��k�r |Aj=|�I}�ǀvw�����i]n�0	�ذ�\0wc�>�`�96Y���jC!Nl�H׍�Km�D)���b(E'��ey�l��p^�56�����`�ǀ}�p�r���������n�66&ݶ� �������Xݽ� �(-�[e�m���;{�ob�	ݏ ��$t�&ƙi�.ف��s� ����	ݏ ���n�tB���-�Xݽ� 'v<��߻���{�ۺ��Z�;d�Ӻ`�-K��/*���P���g�ދ�tvClb����r�mD&��k��F�Bn��VtJ�E�͙� ��ʅ�ٌΆ���OXv�nx�z1Y����8�uf$��͸k[ǰ;R��:7����W�+5-��XB�)��,1myl	L�J��:X�H+*��p�`�q���vu�����Ԝ�s��L�4BpR�퐚-�d��j���;p/g��Znܬ��#u�À�6�amvw0WZ5e[v�[at�un� ��<��;{��|��s� ��R�MZ�.�E�x��v�,��ŀ�z���J��Rb�]'il�=�<���{�\H��<�� ��(�'�v�Wwv���}�p�	ݏ ���N�ŀI��`�؛�v��	ݏ ���N�ŀ}�ذ	��'R��.��n�ƭ�	%�iE.��먂��g#̷<�:�B2�sC)�6W�|��v�,��ŀ�)DK�ATk�Jl��w���K�琓�5�,�	`Da���A��F()�� �!�M�Oٝ�ܒs��x���) �].��ʲݵ�wny`�ǀ}�p�'ob�6B]�'�m���n���r�/l��;���'ob�>��XvD_�V�˦�v��u� ��� �����I��}�����6�L]�B�h�pG%vfz5≮�P4�sŸ����.{8���N�.��۞X�� �����%JQ�O��Ю��+k �����u� ��� �4)Cv���ۥm� 'v<��R[�s�iM0�!���	��3M�����6C�㔉R&a�'j�R[�# �!r]�L5ie��g��RRXI7Kd�۰�����! �A��q�$� @~�k��$e�9����Ϳ���pk������jI��Sh���J;�B!��Nr�g�$SD4���K���͒)h}����7��ӌ���Zʖ�>Wg>x���?|*+�=�� |��b'�� �'Qq@�����g9�����7�� �%����wE�o ���Eݗ�}�p�	ݏ ��%��&Ʈ��]� ��/ �����u� �UR�������v���Y���M	pg �.���*u�lj�i̷c(�[tl�@p����~0wc�>�{��|��g� ��������cum6`�Ǟ�U$wc�yl��w\0�vQ�tժ��]��}�p�"���>�`�ǀMڕb���q:j�i�`z�ʥ����'ﻯM�'}�nN��(PjQ,�H��"R�V�J�Z+�A����s^��Nx��щ�.�	�݊��w\0r�K�<���.�eh��$��WI+��HgX����q�hEЯ��۹��g�m>�����`��S���^��Nv^�c��.B�'M4�wE�o �u�=�U$yl���?;��$��=)�PZ큰ٽ[}?O^�c���G�y�����Eu.���ʱ�w�}�����v^$%��|V�]1���0�c�;�p�5vK�>�p�>T��XB�
��E E%�Qa%H4q�w>�u�kY���nU���)��^[���/e2웎'p��h���WC�6Â����v+������S����癉h�4F,����r��ų���vH�cf+��������p��PnMj�r��lɈۤ'�x{h^7K3�յ�P��Rq6�<��[��p�X�#&)�%��&�U,�Fe�����m-�6G�?�΅v�cp�I>�<�y�&��πj8ϖ�V�i���%��ń��@W�f+�5@MTԣ��fݦ�Ѻ�d���}�� ��/ ��� 'v<��E�YWGt픮ـN�ŀ}����� l"#�v"�Н��V��ob�	ݏ ���Eݗ�l�
Pݰlt6�]�X�\K��<����/ ���`�\��N���˺m�w\0����ŀvG�ulJ�����}.,����^Sh�c[����R۰���]ӭ��F&.W���ݗ�}�ذ���U�W�;����º���`;V7n��{w�\|+56/@7�}�w[�}���uwe�B]�'�m���m��vG�}�p��ĵl��۞XvK�сt�]1v����]ٞ0[=xݽ� >� �R�U�tpn��+�`]�xݽ� >� ���oOiN�]]�)GGL�,���9�ڭV�;(�t�E�h�*�<�5s8�v%���>��X�dx��Us���5l���h^�����mһ������@m�}�znI�����9�;ۿ*/�������0�Bl��6�'�� ������!�@�	F`�c��G� 颀�������<(%��'m:��4��`{���[{=xv��vG�w��H+�ut郱�����nE�~�����n�� ����?r�t�^�e�`���؜�ۚݏY�VƊ�6/D���ڴ��� a�ƻ9��fU� >����>�\0���܋ ��сt�_Wv���{�����[=xv��vG��*����iWG�"�����܋ >� �u� �DL�v"��I'e�w��s��{3��?~�䟿}����
dG�h��a@R�`�,��5��)lX#� ����H�����z���Q�����#�?UV���g� ��"�;؞�눵��U��0a�v�L1��Xc���)0�4��ц���Zδ���d.�M�����:����r, ��< Лr��]ؚE�0���܋ >� �u� >�WR�����xݹ }��U\��\�]����"��xʒ��|V�]1���X�dx{�Wv^��u�� ��]ZJ����|v����ܪ�\�G=�����`ݑ���9�2��|��Y��C#�=�33Z�Z���2����씧�+��[�q��;�S]۝���"JO8xk��gt���p�L�X{zѲ�n�Y�%<q�ǜ�qW*-����k���x�͡��vyM=q�۱$:�@\fݣ�*\�Y�3��,������]�v�����छ0���Cn9:����i���sa�YXP��fك�`W0�ծ<��(s�����n�!;C=Ĥj�I�ǜ�7U)zӪ�F`�G�EaY��q��x�^*���<��9�3fi��-�*RTP��WG�"��߿��}ۑ`ݑ�9��*�����=#�V�*�hI;�.��>�ȳ��UW��r��}�� ���nǀM��(j�lt[t+V� }��� }��ob�6�]Ӻ-�v�wBm��� }��ob��*�ݞxS޿]vӫ��l��#�>��X��x������B��q
njj	1�r�rX7��oMS�3�!̠\=vF�<=�/O=[i�慼�� }�<�뇫� 6O<z��W��[at���l��G�VmW9��Q�UVr��n���w\3�*���'��V���W�j�wc�ݏ�T�v?��<�ڕiWG豗l��\�%�y�۞X���=��R���{O#�V�*��I��
��>��X��������s���u=KB8X��F:�T]����l�n�'Eۀ��U�]��5�����TQk.]
�k��ߞ�u� ;���wn�����f۩\����}���>��X��y��DT{֫�v[�դһf vO<��v���\�*���r�*��{���p�>Ru.���ʶշ�}�p��c�>�`}��96��=[}�}�7C�-�(̙� }�<�wfx�d��>�`B����c#�Vfڣu[*0�h�
�θ����� 8џF��sȎ��p�Em�w\0���w\0����jU�YWGt6�v� �v<�\����~0�y�w\3�)#���^Rv�[i$�U�o ��� >ݏ ���nǀM���պt[t+v�������'ﻯM�'��'�A��P��/�hlwz�.���^��ӥvһI;o ���ݏ ���`�#��J�
��|j�i�N��k��ڡKh�%��M�Lѹ0�aw\��V�3ؑ�N�WV��.�����{ }6?W+����<���u�����m[xݽ� >��u� 7����x��V7C�k >��u�s�g�ݹ�l��ի/(vR�;V��� ov<��ŀM� �6�ZFU���H�f ov<��ŀM� ���J+>ڪ���r��%M�����S��#$J'�׽�>�HD�7��O�P׸+�����7�%#Kc	"Bk�0sE8����'!�sz%�S$�F�O�]�c~��4x�| K)c&�fu{T
@1�I��1����#��"M���Жyi ��l+�`�2����2&i�L��dH��m0*f5G4�u��M� ]�pHa nO�53�M��}�	e����a>0;J@�zB�~�H���Ѻ��9���﷛~�6�3>���Is���JtO����Ҋ������EX2V8�h �����ޮ�F&�)+(�$�P.��}��1h��K��
Ҙ�3�)Z��:��9�~$%���8aQ�w[SO�|<张 �  
��j����b���p� [N  ����T4�X`A�q�Q�\ч)�1m�A��K�U2=���iю�R��{t��M�ݘ�l��x�E�����M�s���u7$m�8��c��Drsf�3�qr���lHtR3�㓒�IDS/m\ix=,��X!7;��N�b�SY9T��Ir�7��ʇJ�:(i�����8|�5Pc��)mM�m�u�ޡV��Y���R���vpc�%/n�.�v��[.�/8}\�jXlz���6����B�����;��q�i�۲V��.��	[";Ǘ�l���x܎-�n�e&�h�y���+��m�*r���g�.�̴��vZݟ,oQ\p@v觷�rn3���U"pi�X0y�jn1�r��/k�wh��=uj�h��;y����^���'��kq���g<;x3�7
.��{X����Y]�S����i�� !��@�ƋVu�S�S4)0!GXG
J]G���c]�%sV�M;��Q��"�L.�Nݰ�M�m���AL����m�6��Q[�z�u��-�����]+£��kn\�2%��֝R�U�<��̙S^��M�&�ָ��t�m�c+qc�C�Z5��FV5�+#s��lm�q����,��p�ɞڣOd춤M�����Ͳ��u�06��&��UM����g9-�t�8T�³(�h��6����v,��$Y�Qt��	�'�W���{�ۈϳm�ޞ���ԫ�.��:I���[�����а �ʺ���'4�� ��mɘCgeIy^`��C��YV6Fՠ'\\u��p!��a�w.�͙9$7Ε�c*���q��9��{)(�`6�%�mU�:��AW[RVL�4�h��`���N5V��GX�����y���Os�I,b��3�'���V�v&�O=.�e����nU#�g�d��V�P%iUWN��#*�mc@���7<Cl�s��Z��v.�څjf3Z��u�Z�j �S��
��Bo�5^�?�*�f����:��b�����~Oȿ!�;��n��cB�c���k�����r�c���{r��ϞM'k<�+�\�[�e=S�^
�nu��-żc08�'+�,󇉻u��Dcٸ�xL�g�����s��n�4Un-�w5{#T�N#u�@� ��8籗����)�+�����ţ�=n63N�8��F9�N�N�W-u�]�-� ����GR�3,�)A�*G�Ͷ��U�
Yvmb��yBrp�Gxu\\��;:=v5�S=��b(E!�=����~������$:n��o�{oߖ }6<�� ov<l`�6�ӢۡZm`�c�>�`�c�>��Y���g����էJ�v�V����ݏ�ʪ�R]۞X�O<UZ����Z�L��`�c�>��X���?R���E�����պc*�w�}�ذ�����Wv^��(�"cV���N�A�gWj9밳㝖�p:�)f��f��s��kF�8�����ݵ�vG�}�p�:����{�i)Z��b/�+M������J����3'o5�ܓ���\ ��<�W)#|J�ZFU���H�f�g� ���`ݑ�w\0씯);J��"۶+w��r�u�, ��� ����r����^��%�M7J�:-�Wm� ��<���ݗ�}������Y٤��u��Km�v�<�c�ޔ�Bn�B4��\��9竬mp�$�yn.���o ���uwe�v�/UUW����Ͼz��O����ل6��lޭ�c�ܮ$wny`w�x���s���w^��lmr�V�ݹ�vG��^��T*eUJ�3����o� I�x���]6�-ݵ��K��<�� �v<��ŀn��]���E�i��}�p�=UKvy�v� |�޼ �z]��\Bd֚6&̀ݴ\ے����R.�N)s؞',��y7�u�����m�> ݞxݽ� >� ���vmK�NҢ��Cn�o ��៫�H;���;����c�&�%)4�+t���� >� ��~Hݞx�����R�Wn��E�
����3� n�<v8`f��Kt��>sY��$���.�4R�2�ـ�ǀ~������	�����	�'Yn��S%��{!N���� 
b�����5M5F�嶭�v8`ݑ�u� ;ݏ ٱ	,�m�tںV��Wd��\�G�~0w�x�p��H��B��Ո�b�ۼ�?����U\�r�����5o�xt�*�2��4�X�f w�<v8`]��	��wv��'iQm��i�[x�p�?so}��H�`{#�>������9UN�l��]D��[j���&���َ��E|��8S�e�Q͘�i��icECK�k�g�]���S�on1���M�덈b�T�:�m`4٫)
�Ǘp[۞n�J��G6Lb��������b0ñ
��ttY)��t�=�Gy��@��f��]�|?u��x
S�t'cu�k�h�g�w��盤Aɑmܷj�&�q���s����]N�������]�<VЅ�n�إ,6K�>`�!�B͵@#��R���X�3U�98����&� w�<v8`(�-Z8��
�vw ﾽ9��O?�{��<���Wd��Ď��/����v&]�0w�x�p�:�%���w��jV��[j��'u� �엀N����껓��O���FX6�:���ճ �엀N� w�<w_N��^�Ж����6����}��ß�b��upmEf��ɬ�G�r���Ј�b�ۿ���� ;�;�Wd��H*ʺ8Ӥ�V��������M���� ��;�ݕ/쫫���Lj��'u� ݽ��s�{c����	6aj�6�ۧV��f�#�X�?�����{�z�\�36B�r�߾�8��+�����{c�n�ŀEؕ%�#cQ�猭�;v����Ǯґ\�-���M�rE���mڴ�ϖ]�K�p�{׀N��{���U|�����w~4;��\�շ�N���/ �� �����e];hX�+f9߻��;��vn���B#b4�(��� �w��[�~��ٹ'~��*J�)�)]2˻o �� ��x�`z���Iw�� �{�b����:M�jـݏ �� �lx�p{�S�B�xj6�|��̬�].��uՀ�WR\t#�in�lU�<OLi��Ԑ�`�w\0������r�@M�x�=���ۧn�Zo�������UW=���	�� ��J5�V�e���IЛo �� ��x�\0]���KmD'v>
�wJ��s�\���� ��j엁��@P���k}��v��٣Vk2��c����`�%��p�͏ �=��� �	�kcur!��|:��`��n^�$L��LiӞ�ʈ��h�J��}��7���;{4�%IV1�)]2�m�7\0�c�'nE�j엞�RF��-R����:M�]� 7�� ����^7\0	%K�;,Ӥ�L��N܋ �ݗ�M�r�Iw�� �����mӷN�7�M�Wd�n�`I��{��;�;۹'�BY @!�,`�!U`�H���<��Tەm���1E7cNF]�I�z[gj�v�3.ka�C�Q- k�P���;=)�,���8�<5�(���V�:u�UX�kG\,�'W;�e}l�!�8�q1V[�����.��@� c��aU�Lqż���P��;H2<��M�C�n���Y�'lZqf�b�*ے�7Yƌf#���`��g�v�qрD��T�:�~�ry'9������	,s"��X�ŷr���<�`�A�-%x�H6)��A�F��g���sr��¶ށ��� ��x�Ȱ��.��J!;��]�ujـݏ �� }$x�p�URG��K��c��Э��~���� �����6!*�n��]��I7\0�p�'nE�HJ��V1�)_��o ���ʪ�g���߼��{׀rw���t>Pm�b���.�n��pGGGn�pr����V��$ �[�j��]gt�H�g@��避^��ݶ��L�JS'Eۤ�Ӥ��ȷ�b H�Į�8���L�vu���wu�?�s�v~��aj�6�ۧV��� o�ߞ7\0ݧv�X�6e��e���IЛo ���ӆ;r,�w���:�J���@�ں�l�7v�0	ۑ`�G�M�v��	$���ʲ�O'S������Ajz���c��3��e��e�Ahv;��bul�'nE�I7\0ݧf�RYN�݃�wB�k >�<n�`�N�Ȱ	�V1�)_��o ���ӆ*���<?,H�)��	u.J}�ռHR�S��a�$~��9��p��\$#��ht��f�-��Ą	>3��Ki9�s|?|_�~��g��ޢ�Q˩��4���	Hu��dB:6Q��.��Cwf�-��$���vs��B%�0�>�G ��h?T��$�E���tq�%!$�4X��M=aBl"��� �"�4|�� 4�X����#O�qMP��wK�|!��TH��& �`�A0�h"0��t�pB* !�~�
�E	��#C���1Mk� :%70��"�������c/�X6(h<�!����F���9f��f3[�k6;ٴ������h)*1��$b}���3z�iމ$�>@?$�4�%hPhL��+��f���';��l���҆��S��AH?P:T�|�����h@$Q�+�|8(sJH�b"�A�U����+�Ums�x�wc�;�J�R��8Ӥ�E�0=�RJ���׀I�\�+��g����YN�QvГi�ul�"엀I7\0ݮ�p��Y֍����J7��VdguWe��n-�Ib����F����uYL�]c����� �H�	��n�L�W9_ ��z�J'�U��ۤ�	Лo ������"엀Iz��:�J=i'v�
تճ �W���%��G�M�v1(�hv;,�bt�`vK��� �����Tz���A2��� �0 ,0"� s`'5�ٹ'}��%��[�|n軷x���u� �ڙX��X���З��QIݻj�LGl�0�4ex�˙�P��+S%�5[��I����65e+�wm����7v�V����W���x��W��YVq�I�+�`�S+=��$w��, ��n�Ӏ|�zk��a�KV��g ���� �dx�`ݧn��.��M6Qm����%��<H�`ݧ�r,i�e[]�MН	���p�7v�0�Ȱ���6]���B��+�\[�\04Sn�P���`���'�O\��R�#x�[�l��ht<�/N��x㳇���	ER�+�K
��8���#��Ͼ�}�Ǻӗ �S�ۧT��#n��}Չ�pgc*��ǝ��ęEQ��la�.ܒ�X����jȩ�^ݸQ�V6�-қ:k:$8uUܢ��4�g=�����m�'Hn��pf�jS��2��\eiF�I;��V=[	��p���	͵��u�Khn����zt���dˉ2��`�k�pK5��=�� �\� >����(�V�c�\�'V��r, �H��ذݧ��URD���)��`���Wm`}�<I2��W))%?�~��$ N�)�R�;Wv�$�X�ڗ�Ir, �H�Ȓ��YVS��ڶ� ��%�\� >�<I2p���'A�ĳL�lJ��nv`��)�k�B(Y��S��Mvc�����I6��xˑ`�G�l�+ ��%��+,�V�6����� �w��z��+��B�\���D0A:����{7$����nI�rE�M6,��.�&�N��x�2�]�^��X���RݢZN�Ӱ-�1۬Wt��l� }$x��N�%*��wk��Wn��"��� �0�����r���S��`��	5�Ѣټ�1��P�,����lE��¾*4jCb��y�������l��{r��"�$ N�)�R�;Wv�6�,�x�Ȱ�#�;�DB�)�ձ���$���w7$�����p�(�~� � �b��f��krO{>�ܓ��f��t.��j�gp߽����� �{��ܼn��.��M��o��� �H�W��_�r�x]��{=+;��l�ZDU�P̸+��mbF��B&��]�]&9��bƌ;1:���v	��	��`m���	� }$x�}�ֻj�l�7�|�{��;#��� ����J4U����-����vK��� ���{����m��M�1�t�e����	;���ܓ�g��ܚBPI �����[��;�vN���WP�jYwm�u� �r��_�yo�x��x����K�Ў�X�\Bf���:.m�둖�3p�ܮ͜!n�v�n
;� �՜j��)+k�;._� ��/ >�?r����,����ի�]:I�خ���G�I�{��ܼ�*�IOs*�n�e+uBn�����{��ܼ ���	�Ŗ7e��	Лo 콋 �on^����^�{����j������=���{0�#�;/b�>�kxW
+�2��Hة[ ��I�֪ۛ��&`�j�N�d턢ճ�#�Y�9�^�Ou�0t�^9sH]*����b�X9����� ��Wm�a��b���k��6�?__�÷?	��AHѱם��V4���v���d\��g�ɝ�a��ol��)p[����o��&�</-�Y�.�7"F�+�5��vᱍ:s��B��G���v�M*�3�ap6��5�aY�tj���TC���FG��v�7�k.T���δ-m�;8�p<�ȍ#+m�lF����ciSW�NN��m+��� �dxe�X�ۗ�I"��h�t���Jـ� 콋 �{r�{#�$*T�J�e+�X�o 콋 �{r��IE����޼��H2��WM�%m`on^��^��/ 콋 �T��-]e:I��v� ��/ ;��{6����z�,�]���v�L���B���)��-4IPם*W[z��	n�>&�k�U�-���V������ 콋 �{r���޼�/)�.�&�N�=krO�ϻw�m!x!�ؿ�$!X�i�ǘfpTWB�'���׀{o�`�G�}��D�wv�)��i[X�{r��Ȱ�#�;/b�'nRQ���e��i[x��X�dxe�X˫c�$���j�t�񻤮���#�;/b���<{}���%����;i�ؖ��MN�F��U�b�K�K��lN���>�7C)]2˻o�7�<���� �܋ >� !VU�j�ĭ� �kc�7�"��#�;/b�>���j�)�M�N��{r, ��<>��@pbF!�D ����s}��N~>�{*V���)[�I��vG�M�� ;���	ۑ`�DYN�v�[�M��M�� ;���	ۑ`ݝx�O�����h���
Bm����m��u�wTq�mWc8}=u@�\��1�aM4:.��v��;r, ��< ����)(�WI�n�m!շ�N� ��< ���{[��`�:|n�%l��#�	� w����� �*@��Ք��i]���9\�)/I���<v8`;�o*�QH�2�ZY��-if�)J�z�v�Е*ʳ�]6����H��p�:�%�ݏ �A�;�4%f�.<�qҼ�m$tsj�y{r��J-�bv9����4���K���p�:�%�ݏܪ��^��7exʷE�V�V꛶`]��ԐzO< ݯy��� �ݰ����al����	� }Sc�'c���/ �l���wv�)��E�x�8�k�� ����5we�ݏ �ƒ��;,cN�o ���UTrz��z�$�>���$�TU�TU�E_��Z���Ҡ"��"����J����
" ���P �A��B
�AH* �D��F
�A� �AP��H* �DH*
�D�� �F
�D �@
�P`�DV
�H*Q`�E "�EP �D  �@@��*
�
�
�F*�F��������� ����
�
����� �EH
�P"�@
�D`�D��T��T �E*��H*��`�AH*H*X
�*�H*��
� �@��H����
���B
�H��`�B
�H*
�T�� *�� *
�`�A��A����
� �D��
�`�D"�D��A �@`�E
�T��"*B
�F
������A�"���*��H� *����E �Db*H*
�A��
� �DX��*`*��
�"*�*��H���H",`*b*H*
�V�`�E����@
�TH
�@"�D �@H
�TB�
�P"�@`*
�*
�H��� *
�@� ?����(��ʠ"��@EV�*�E_�TU�PU��@EW�E_�TUҠ"��PU���d�Mg�W0Ps[f�A@��̟\��| ��@IM�	���Ev��@Qk[Ě P  � 4 :N��$�E  �P!P�IU�BQ)P��$��H�E)%U  U     P��J�     � �  @@i��%�[��.Yr˽�K����7� �z_}���w��׎�&��YB��������i|�� ��drw��/�|���)}Ͻ�L���_G�7��wy�J� ����+�Z��n{�z�y}�[xh  ��@ 0� � i�k�V�w�o{z�[g6R�k�U+��۔���k���=��w�tv�����*Ź�+��x ��7@������}��}��[��{�����*��m|��wҷ�޽5���zy{�{��v����  �  � �Ͼ�n/�z�p4t@�}� �tpA���{: ��P�hӧ @�   ��s �`h =*����@�{� S���U*�@)� A���� @�  �  (   �RS���� � �Ͼ�o��o4����駽��qg�ܼ��{��yS�>����n;�G��e� r�Mz��>�ޚ�> }z>��O{>�O�7O=�����v�O]���;�o�y�t�6�m���owy�+� ��PPV� �PJ� �[>�����R�n>��a����. �iw���y�z�����qez� }>����]�t�Z�� �o��r��\�ӵ)�}4��׭^l����N���6o�K�-���y3�NM=��7�mx   ���¥H�� �j������i�42���R���j  �'�T�3IQ�� ��J�iR�  �!JH� h�OA?������_�������>�g�is��ePW��_�*�*�EES���*�� ��_�TU���y�bH�@�#�	���̬�<������J@����F���y����[7�Hr46��<XT�##cRT!G�hEl)�5��!i(˩�>��a�h����G�"���u�a�D����˅auG3g3���Æ������{!no#����=��V���.��ۋs����8�C5�\S! ����˥ ��o�E���<o=֏��]P����@�I�Y����w��f�xg7�P��e3Q�4ܭԺ�T�]�{s�j��+-%<�sd�=E�:�b���E��x���/V4�����xk�Xh��F�Hx˚�+$�+�F�'��a��}���_o|	��V��Wm�V��}�݈��!H�N�w&6~���×��	�;5Ēt��hB�,H$HH1(�� c#�L7���ko7�J��0�e9�9���9�VL9�͛xF�/��~bK�F��D���X�*F�)$ �~�5�y��xJf�Y����H��S���4�y�=lZ�!L]n�8o^{��>8
��s���\� @�Q�9���y}6�!�\5��$OC�^���6�Rr]�ė	��=�Ѯ��wFU����Oj{Ի�-W��V�n��m���g�+Q?5�;7�����\ �'.��ٲp0�Hr����H��Z}�2�
l����^3��=;u��\�����SRh�=��E�,���L��WD�y�Շ] ��)�,(А�#`L"d�m�y���?->����b���>+���m��A��W�++8X�ʲǞ��h��?/���˃�4��>����ҫ����\a���\)�)�0�,C Q`Fw��u�<��y���ک��O����J��ߵ��ǲ�q�P�o�f̙��c���JB�C�h7�8��xFh�����/2{�	ta�g�g59�Jx��=	L%�#	0�$���8nk!�e�j)Y������L�󧞴��Z�RB��]ݹ�}"w+���f�|�O����/�S.�t=g��	��y�8�(8�a��s�]��3�o��9��`@�`��Cc��)�f�t`F,6c�!P�H%�&��S"h�l2G��|ٖBy$Yq���K����x�aL��o7��}�[e�]ֵMjk�R;~B7q�3��P$1%J��a��<���o\����,
y�2����6z{vG��D|]W�>�b���1�Օ�ZR�:����y�N�����Nݥ��at�eS�2�ґq4DĮ��~�[(��+� �2a�Jzg�Wv�"'�WW���k\���?:��?;��U�c�^j�^窭���"��=���V�_/���ϡ����٦P��Bdj��0H��F�o��4�kfT�
�H���X4\��\C�H0 �Η"������ؚ��*T��*�_�!R�壺>�_��ur�Z�__wi���qccd! �R�)d�|H^h羞zk���H�Ȕ�0M�j�ٜ�9槷|H�u�}gԙ��jį�W���ެ��|��=	�-aL5�!s[	|���6zpu~_��g�o�;.!�X���_��_����y|U������n��¤+��Fr4�e��mڎ���o�_}���Ӝ�Ɇ��L&_7�Z�`�{Ho4�<�y|�0���5��xr%�e|d�_`C�[�mA`S�#�6���C��ۤ8�����sÌ<�/���a�Q�tB�BɅaI|���l�5sE���]G��5Z\�ӽ�yL3��U���,�bYOz�������w[��J��_��f�|//�Wy��ʍ{���+·r�K��U�:'���z�K�i�+� ����2��'����x6� ��� �m�ߧ5垙���)�����q%+K�a�q#j��kY`B0�p�4F�Au�B뛹�Xq�B1�h�5�Cf͹�k�I�D<�<��Ղ"A��4��B$� 8�ָE�.��J��!j`�B�B"VC�F}��Z�X�6������mb��}�un��Iu���3���>�~����k_p=���8?B%ɭ���e�l>k�a Ͻ"��5��{|f��9�g�\�,~�������V}�6��T������.r��~�Z������;�ً�W��=�q�]b1��a�-�E�k�}0"N�W�;u^��9zƀ�:줨�*��W�U��V�8]�S>�o��׿u�։�.��8A+�1����G"�"D�H�p��D� @��(!��C9�[`J�y��7���C���}+�_�!�řd@�qY�ݴ�S���"���W�)$�B6��,H&��#`\��h�L5�D�+�"���6�)$�Hr,�6{��W�����}�EJ���.B�
/ԏ����Tϖ��?��X�չ�!W�͡&ؙ����KB����O�v�Xh�4]nq��7�%`F�L(�`�\�$849����?O�n�����������s�08bF����9u��Cl�6i�
�ad�Y������z{�ă-��5�J%��ed�g�9�����!='���%T����U��Y��+��z�]���������:��r$y
��{�zï~?�莥s!`�Hm�fR��yB��T�i���=w=�$���^��s�K�����ֵn�,�K-W�A6��՞���sș�[���n쓚������4�4F��B�F#X�bSW V+cs�	����1)c5���\����d"R�������Nk��F�!$����לLv�)�6�յ��X�z�E�q ߊ��O/_��CūF�A��E$! �$)
1"}$,�$�d@xA 2d@"�VF� � !�AbHȤ�P@ �1�@�@�"� � ��	�H�$"�#c� �U��	$a  �H&Ԁъb�H`� bZ���q�� A� ā\X
�10 ���dZF$\��L)-L��H)�5�ĊB5̃LLX)*P(1b�ja�̂d�\�� a�$(8��2��\	(aӉ��04h`I.@��0h��`E���$4E�I�(bi`6&HjH�F��`lp�C8:B%L:���0"b)� �h$d�G :	HH5�f�� �l��2$�2]M����ir3&��b�0����$�� A�ne��g�˜�Yw��ʞy"B����$�"2,˯9䥶6���+G�f{���
N��Z$�4�>a�$
C�$=�D*B�Y�6i�7�ٸ,0�mb��a$	"� xv�4_a���9��vy�����,vA�.��ٙ+�@����[���5w}Y�~Jz�ϊ��כ�5�0���	��#O���4ȑ!/��#�l���0��\�$�xx�S�H���nkO��3āS�\ԑ�uu�a��n��N���,)��ԗ�g��I
��@��a$R1!)Mi6G=�o�!e.�
��r)�RF(n@��HE$!��I� ��,#Bơ�|��6����}��n}���v�a�1��(KB35�.�6���y?�$*Y��yciҼ��G/,��|!�|<����2�p���N�E�L#e�~�a�.��r��B%����\=��F�	�X�4K�ƅ"cL	L n�_���䱌�����b�1TL%��ٽ�ܒ�4��r����)
��1�� P1�VR�!B2A�F�"�EI1c(�P��ȍL���5J����HF�d()���!n�
p�������T	 HX@�4F@��5bD�3Q��Bf�W� �͜X;H�x��
�$-�fL3�
`d����z<5 x�j`h6���! ���5���L�M43N�o+B��~`@	B`0��w��D�|㙩���	�1�䄋�i�H�!d&��&ke��Î��<=f��~�L5�n�Z1#2�*pu5xn,�RQ�%W$����̶F X�H�����dy�\D��H�H�4Ny��JCZ,,����0͛*bfAP$�hi�g��B��r��E�;<�z�#u9K�z���	4�@�c E`�/��g*T�Ԛ߽~�HW��{P���Ͼ�w�?]��_~~��� m� m $ [@    �� l � H      �m�             m�6� �  � �  �llXΌ����Uî7e�q�6.Q3ay�^��-T����k���U�{\�UUUNR�y�oK���3�jڗVհ��YPf���fٶ�t�mm�i:J��@6�A)��U��RCfZ�j�8*�j\�	z@�z�c ���@�<�u�W˭� 6�pҭ����-$S`  )N8l �@�m -�l�dʱ�R�!#m"�א9ɳ6sI���h&*�S�k	�U�ͪ��CC�ɩ�˒n	V*2bk<G/Y�� �k���g�ۮ�w(ιм�@��q�V����ov��:M���=��C�b:���M[X��[�� ��r�-OF�Ÿ�@(�Yx�)v%�"���}Vݵ�2A#����;v�oZ�/;�]�7��A���ڮ��s���\�O���Z�m���c�4k��%Zڜ��\H��@(�d[dR��� �ݧ^��&Im  �V��J��j�'���l� qz�Ž5�M���&��v�p�v �%�sl!n#a�X)�6K�)UH��]#�X�I �B�4�;�4e��3aCkm�V���t�Kx�z�B�r��OmAt�Z����!Q�	V�mmӒ;�A�!ղ���{t��J6��>����0y�8��u�v�p�Y&��j��]۶��vn��-Ep>:JΞ`�3�0�ÞBy�ݠ�Z�D2v�-�]V}�N{l�m3V� s'g�q3n�\v��:[��Ĵs���nx;�U@SOg�Z��R�P��IKu��v�[@d��U*ʪ9�jB�.��-t�W��Y��jq&�Q����
��+:�)ܹ�t�ۖn�Z���b�Z��p��=drc�j�x��/J��f_=ݚ�͵��M[7(�2�����:d\]�Z��-��U�q�lljN��Q˽���]G'[�mI,�骐��Z�J�i� 5	��k��j�C.�	*��4�/P%]Gm�륝�]��S���t�]v<HN��vޜ.�̵F;���&�ؖ�F�[aV�,CT�/5,�.l����L�]&Ԇ��	2w]�m���p�:췻t�ŁN��&��J  A�,�kn�W���7K<��x�����qD�f�8�g0�6��v�Ts:&�K��[��/+�f멶��v��E�][�b|t�7
��X(�MMR� }o�O�l�6H��	1:I �:�u�K�%8�-����8'Y)�k�wӯO�,k@  ���[��,�om+���{#U*�
v�v��ɳli0A�UV�-�iejڪ�F�U7J�R���kl�l�U���}O���.�UU;> �<�5��>�6&HړeS�W��*a���+��UI*�����v���[U��/%�A[��-Bg���1�kn�<��\���P��aa��u�ۤ��˹�s���t���N�b�w[\�v'Qo[N�WL�h��6u  $�p6Y5���[u^�e%��v!�jRP*�<N������(:�@��kӶ����m��ljv�([���mJ�UqhA�-�ljY2��Od�C�79a[�N��v �ڐk���M��]�v[O��m�m�����If�d���d��BNnz�u�R�Z��C-�À  $mV�$�n� �e�fȫk����y�8�y@� SL�� ���빑��t�ll  pm�6���r�� -�dT���q�  -%�k� h�m��6���l5��vZ[Rn�H8�l �`  ݶ���$˅�Qyqsm�`�	t��C�~��   �  	 $�h$���  �2R�UY�L��h+�影�պf9x�h��p p  ��k�� ll6K����� �t�)��W��6�m���\ �I=���ǜ��r�~��}r��.����,'LӔ-ɴtv�c�V���W!�1 p�@)�z��m`-�M.0�UieP%R�:i5��E��Hr@�x/[���0e���[@ Z�6�Y��8==+5sm� -�g��[Ӯ�X*(�����Z���d8{r�UT���6veC��j�ʻ�[��̪�b�
C3�a�U٭��S��k�Zl�s'kX��5Qy�Og��������#�į^�Z���ؗՕ��n]�BA�e�;u�e��� :mW*�m�ђR�n<n��G�ڦ�=��!�4L���9��
��� v�ƃ���Z��ͫ[vDt������6ȳ#��/-��UFK��:f���mMmGͷ�sy���Y�m
��r�UmUg�V�6�����9�` *�uԪ�q�*���  6�m �@T�'�`*���%�X�le���b�  pY���`ٮ� �m�$	6�����M�m�@�� �a�m� p �� �	   [Cm�t����ڐh4N�e��jt@�Q�`j�\�*�l����P[B�m��Ghp��a�   h6����U@Q@
�.�֠#.��ڶ*�y{4��Y�Y�QuTHl8m��lL��tv�\������]���v�.c	����>�[g��R���g]����c$8;e�'䜺�E�c��[q��ڧ˞�,p.�ʹPm�U/-�R��@[@V�L�[��T 屋%�1��n�m�@u��PE�H�۩IA�ug��WU;�;ԮY�*��f�ۻl  [KkI�:��6-��v
���ql�nˇa����u#ŌmU¨�꙽C�O�y��F��1h%����NIą-�(
ʯSj�U����*�R�UT�3�Bc�*[C�Δ6��f��K�mC`h�m�݆Ԯ�[�`I�d�s`���"�R�mUV����vڳ�0n.�B�U��
j��y`�\��'^��I�E��֬\�����:�5� ��!�U�[uj�VU�r .��nBYjlڦ� +��[Ua�1��ql�U@U*��S�մj�c`:������ ��ٶ�Ŵ �� �A�A���ɛv�d�y��hI  �$    ��\�6Zx[�l�_� $'I��f�l�ۆ� ^����`P�ݸ�Z��D���?�@�Æ���UV���[]�I:J�p�m�W*g��!������mN��@�*ٵ��v�N��JF��Es�l�*���6����H���v��JvjU��UZ�jV�]X!%�ڕj��j�%�` � k ��k�Zp�o�|��� �[u�kqm �m:��l 8��V$  my�K[mm��N��m  ^���u5m�4�  	6틢Ԁlm  h�� �� �am�� h  �oP  �`j� $  �l ��ni�g m����)wf��ﾠH5J��m���b�����UJ�J�*�S�+. $[R�L  �Z��\(m�       m��ٶ��� [@p       m�& m�[[��f�  �   -�         m�6�	 �h                �  $                          -��      ��                             ��smml@     m��8$$q!�H~}��|�J��Ѷ�i �h�[BY@� m��m�����km��"ڐ����[� -�'l��״�� I#m���Bi@6�-+�8�f���vݵ�.�lN� m i2dZߎo� -l$           pm�`ld�m�� ��     ��h8���m� ���h�a�l��[R� �`�`�5�� p �am�l ul $[\J��H`*��ҺVUԾ� �hh/[5!4�UP
�H h㎳���pٺl smm�ӁJַ�Z�Ā���8 m�m����&�`6�m6�Y�e�Y@���m6�۴�8� �m��Z���4���6�m[j&M�.�l \$Uu*�t���pg��:��b��Uw*�3B �8�$�83�.�z��N��
�m�m���L���� �v�[I�jMm
U�B�1�U�j����LЖ��`-�nI�n�In�m�"Y@����-]���a��|L��cz��h�IrL��  ��mi6m]��h  �Nb�k� ���m��m  m��  �� � -���!�fM,{j�8�k������宪�B��Sjo<�<��i����n[A�#2�[j���X�[Uu]�M �s�m�'@�`6�V�鱙����w�������gP�P���T��J�E�XA	YD���á bB'�mP	C�x��8�h#4	�`*�<AM(��@�Mz� U4 x�S�>Q��S��G�⇪UW�UX:GJ� hP�bA�+WB��xh<=XCQ�����.�6�zx�x�'�*��B1@6�= =Apt><WѨ��?"|: �Sj)�
��1~@��8�D��s����~>��$"�A'��
|�Ax��i_D|S=I�p=v���)�/_�`	�p���O��Tt��h�a�O��B#T�^�=W� ��鱒�B"����G��G��.�p
"��x��+�)����(x�]"2*	  �@<D��	X/Q�E���OL H20`�p�4��5� 8����@��8�
Tj�U�JQ��	X�k�`�p���! !����ڪ'��Q�A�z�"B�BI&���%��@r�@M�����OOE~/[چY	�eQئ�=�H��"����_ECa�}<$��	X2Fҍ#F[H�����()��C�>@��>�	�@18І@�@��+�}��4��¡��=ڈF!�x;�S��@_|M��ҁ�[R$�40R��DB5X�A+Re�HE
�DP�^�33zֵ� H[xp�n ��Gj�[RTI/�y�q;��Kɢ����;3�����v T�-&F�� Y3�� ��P�-z�xS���^)�k\s�w��v�ч�r�U�t��f�/q��@�l1v�k۶��ƭ��,`�؅�cw��8m�6�|�ïc�'.���+Zƺy�x[�c§;�7=n�'m��go.:�X3�:(F�(^�On]G�grֆ���ʣ9�Z����h�Jn6���Ѱqk1�v��M'EXӶ/V�f�XF�[:A����7-����z��{e�QW�`�:�if��89З�N�간e�g;#�� �����h���n�m����1��v.#�g����e���ln0J1y��(�(m�b���&��iYf��y��Zvݎ2%��;�["�d4ꂊ{b�쫰��p���t�lk�+;�ڪ\jΕ"m(	GX��6��Y,�u��<ur�yn�^���l]sy����W`�v���%#s��rv'T���UJp]tbѫ#-�+UHOU6�L�
�d��+�Cf��g��]tdjW�6��ݭ�WTGB����C+��볞@��r��ܓ��ӵ�x�$��l��h.��m�4)�Y�u�.�<m����F�iZl�N���3+A�]�OB��mp⵹=�S=��Ĩ@trH����/<uU�|Is�wm��L���Ikq2Uvy0�15��!@Pt�̓�k��n���D�pi�Ƚ�I��@�fȺ� d�۳m��  6�   l    ���     ڶ �n�@��
��]mv���k�� W��JV�&M�jU����֨��t� �d�d#T�Y��^��m+�+��c������c�)+��ꭊ$m`�
��;sVS=�=�u[Eg����&9�Vn_q�#4�Wm�q[qPR��Z��nU4�]j�V�$�JfK��5��{�����Sh�OñE� G�@  ���>7��lVD`�?��㗮��{Q�+��2�vۜac��lF�Yk������@jN"��t ��v��c��a,v�(.ZN.:wh˲�9u2`�#.�hg<��!m�؛u��`��]�9���������\�-�[���@������&������!�n�5�	�5� j�m�;d'�!�n�5vx|�4�P�0����uȍ�)�Vx<@6
hGvCr�d̦fKi.[h
&�y�v݌���a�AU�/`��{<�#��^���)P��z��&K���T�5?�y�lv�{7lΦ�{�pt�0&�i��	uJ��eᕙ��&���F�z4��r�9jۣR�
�%C��ww�wq`ٳf[��\����+"'i���`M��u˖���-��#L7����<�N�7	�NM���9#E��܁wm��l�W��b�f�u�]��Z,lg�]�f/߯�~�7�0=�`ztk �w��M:����Wf w����VVRǄIJ�kJz�z�y����i�푦�Ζ���+&e��U�^Ve�=�`{di��I%U����}�L�;�&"TKJ[-X�Z`{��l��lwF��"���݈32�w���:[kd���L��ŀy%�Qw��9+v+)"hS���٩z��*<�p�J�#L�Z65�8`:h�Z��[-����0����7di��9r�
�1U,YX��.���07di��6�K�JrC��^N��vV�ʰ��b�N{�߳s�(ADNA�U�0������y��~��y�ذ�|���A��imX�û0����07di�)˾��R�E�]嬣2�[%�=�`n������O�V��M�ȩ$r@��ŐIˮ{	��$�o�`6��-��iYNḆR*��f[�Ѧ�0=�t���ـ}�w��)U�)l�`l�?�}�%?c��~��F��59��A�
KV�}ݸ�۷r%'��b�;��� �꭛FBT[y�Fe��1����vF�lB���A`p@��L�d�y�'�C�Ċ�ڪ������{���n��?vـ|������t��N)�Ic�kG���|}�D��J%6�@���L6�h�
�9|�:�5t�V'G�vV�ʺ��b�?\�@[��97���T8�f�� �eb�,��Lu�-�ս-������q`ޮ�S��Q%��al�:����L	�`{��l�+'ف����I\��.?�}�`������_�ـ}�w��)C���Հg�)P���3c�5�6(��,�H)�D��! �(`,����D�j�.Y��V虚�L����wFv�lh�p�r�mi0�܀�v:�s�F�OV�;b;m=��s��ι��$�;6@��I�<��8�@.���,lZ��;�5狝�n֒�ځ�N��R���ms��z��q�kl���7Z���ܸv�3m�hi�vm��Pb�������Nm�  T�d[vt*�/A�6�r����$��Ea�b���Y�\���4~��U�J)yl�6u�0�;pQ�gCv�NGR�W6
��2
���K8M�T�#�-�qں���5�ݘ��L	�`H�Q2�YW�32�2ܙ�ב\��fm*ov���yt;t�Z�V��hIf���X�#Lu�-�+�[kb�U��Z������fA��	�1�����/�M��;D�$����� ˼�뼥@g�p�532d��!+����Wo�3���EmM��l���Kj݀N��d��V��\=<��i����k�lP]�*�yKY�%�ؠ=�;�Z�49i+�`��ŝ����송��R��I���L�E:ɒ��f�3+�"���r(fE���m
�b+0�2�gF��:[�d���LEUn��bx�T���._6({݊뼥@{/1`�k&�A����u�f����52���������=�P��d�F7A�,��yz�cEF��������������kkķgf�����Y�c�Ѧ΍0;n�[�d���>�J�Npr�������s�I&��{�k�0����:��鴀7h�̼ʠ/���@[�2(d��gBL$�'f�L���l��R�=���-[bqY��K(ݳ ��v`��ŀ}��X~��0���B�&�-%r���L�`v�t�V�l�o��h��G^�s���ca�.����ڐ�sB�I5��4ƭ��F�3�mΕ�1��`v�\�V�loF��-Np���� ���fy6k�0�}� �{��͞��ny2^[l+�Y���߿[�Ѧ΍0;n�[����գ��Y�~�w��vnI�}�7$�$4S`���B��䓻�������s���`N�0?%;*~�+�~���L�X-��srf�Iϕ��x���ik�p��QVP�o���}`��m�>�`q[��^u��l����06ti�N]Z+ Ӓ�e�`n��K��n��o�`�>��7���%h�n�^Ve�=�`l���륰:�K`l$m
�b+ef^b`l���륰:�KaJ��<����-�ʬ̱U�&m�K`ul���ti�����8��k�H���J4[i��1%%7�=pY>B�ݛn�;t���xw>�j[�����T}�y�@�YY���:εS�lv�v����=+��8�ɺ�.��R(:�WP���ix�C\�5��e�g���\�\������[o���;۰�=��
�ƶ��O�Nِ-�m� �n��:��RM=�q�+��1�2���M]f�M�2�c���~{���(qd�Y�Y�!$�j�&��dr�g�2���`�^͒�u�`��!s!�R����r�l�n�l�=����X��ŀw��� ���kR��u[B�-����oF��]-�+z[����x��G�rT�*�7��,�G܊93�����ͥ@[��y#��̊�^f&m��`uoK`{z4���� |�]C�l#�Kh� ���0o^o��2�iP�Ƞ=��M.�Zw6nk�-sIG^gB͓6y�n��;6�=�]iN^J��hr�W,�?}��@_�)P���fe������"���v�V߷qg9Ļ��r�a`�$
 :@��g��}lT�loF����-�ʬ̳3/���6�KeU{z4�푦����(9U�Z7]�`=����`v�����;��JW���aX�0.��ލ0;di��}r�S�`Is��ׂH�(J�텬��(�e�d�l�Q��L��MRHC��9�V��qJ�e_���ذ�;6`=�����XX��v����;V~����d��}͊כJ����Z�6]Z�B�8G,�Q�f���s�~ٹ���,�!�����a����x��)%���3+�C��R�}�e>53[��,֜@1 ��Ck���/>�4�$ܞ�̐t$$>����ń��l�X4����3B��s�׉�6{w��g�����B�>L4mZsG���oo�|�"֮�y��$:Q�e��#	!���I�8D���Ha�<*�M\���0��
CO!H��YY�:�p���86�p�s�Q�\��%W��Bp���k~�x$�T7��j:	��L�JX�Cx�� @�Aࡀm�����j���8�P�i���p:��|��P��
����3	&M�^]/����د��^�δJ�����;^��wߖ��b�;���F��L�7�y��w�DB�"e�beP��U�;�q��G������6���q|�[A��C�9A(8�+�<*����;<�8&��UQ�q�])u;��un�l��ٳ� �gu�����\_8e�Ҡ���N�9�ħ����bb���׮d�^oR�77�P�ȮI6oCj󅉵h�-��w}� �[������釛��|��y���qH�*Z���Şl�c�L�M��j�'�({̅f�T�K �ha�������;�rN�}����F[j�7��� �������7��X��T�k�묮�l�ص�%�]8�7�+�WU��d����lK�3"EbU��;d���0�;������F�n�[�Ys�Y�W�]b���`v�i��#L	�]-�����>�׬D�Ih崖Z�����6륰6�K`{�4��Ȋ-��U��fe�`v�t���lwF��w�������ʣ#v�緑@k2M������Tz�(
ft��`0�H��!���P�|I���
f94d$z��r��zق^Ʀz�lV�4�BM�&�l�ZK�����mՊ^�7^�5Dv��ܹ�۞��8�ݥ\�t�7 ����ۮ-�no	/b�TUD�d�m-�v��P��	�K>�Sm��m�ܛV��n˗u��m��-�M�K���8  �UUT�aPې�X�z3d9�ˁ�^|��٭]�s)5U�q^�����%�3%nd5�4���@����Z��NhvS#(4M[{N�x�*`�&գ��Y�~��ŀwdi�6륰6�K`E>�V_�h�ϋ�L�`M��l�����:��;�`7Ud�`�}ـ:c��L�`�DK3,�.�.�0�̶��0;z4�푦�}ـ~�ټ�X�Dv��wq`�����|�>lP��h���O���b�e\�%;�sGLr������ʰM
N빧A����tΛ�3��`M��lgL����^�ޟ�`}�y�"�Q�im�`��ٛĹ�ʒL�7���4ٛJ��fR�I�'g�4��#r��X7�`}��ﻸ��{�{�͞�zGײ+jұf`]�7z4�푦���6t�[�(�*��E^|^b`v��=��/"��ה�fI-�s`S=�u�jӓb%	ӵ˃�܌M�l\�ev��Ql��t�cs汶ZA����~�`mN����i��#LV����p��-����ـ~��� �۸��wl�?wP��U,m �N<�`{z4����*b�_ʂ�}HT�l(P`HՕ	)>��{��'�Ww/}������ -��0�����ӣL	��-�ս-�����"(��O�+30�����}2(Y��ͥ@}���L�Ո���i�EtA����lE�ȏ6BJ�M�4ΣEPN�B��qtl�vZ����~���LN�0&�L��ofȬM�GU�$� ��w�{�0&�L�V��[�(��v���������m��`uoK`n�i�.��ݵ�#+��9*�7�ٳ ��߳rNy��7'� D����0	��y�2ke�O�yP,X��f�fc3��`uoK`{z4������e����M[k�ѧ*�G��@�r��p7��1��T�ݨ4 ۋ�7�k��Ax������LN�0;�.S����7Q����-���V�{��RI~Q��s����̥Z�z��d�r��I� ��<����&�ｋ ���X{}Z�V��Q&b%�5��5�^�*켥A̙�(�{��x���S�V�V��� ���T2L˚�{��n���~�Ǡ!��R$!�K�-	���R)DFӸ)�Ֆ�i��7��8�DMu���<F��@���yo:Ѷܺ�Bo�ɇ^�����M��Jm��a;7m8���{ ���Ѻ�C�`ҙ��m��])vlE�p�3�AI\a&�=�O/�k&��R֤')�Uʼ,C:I�T;�ֳ�����v��m�`  l�Vp��J�Ilu����Nm=�ɒ���׶qnntA������jo���4a���d��տ�����h��r"�ήN]�:t�P�s��@^Y��YW����+�t$R!ʂZ�����]����}o�={��b�͙x��HO*��ܾ=	.Q�o=y��Lm��{����JH�Z����p��-+�m�n����o�ܦ7䤟{}�~��{�\���j�x��KQ�TS�ߙ�r���IN��}����w{̚�����)7����ͷ�#؀��-���i�m��߸s���>�w̗��~���s��|��cm����WZ�¨Y(5BY; n�h�ݣE�ĕ��A��U�l���b��{���'	���ھ���޹����sNr�o�}�N��2��~�r�~�B�ݹ,V��Q-��m��柿cky��u)�@n���`a``05�`�ѣRB�s�AJ�h������Sm��������۔y�$�RF��ߔ=+Q�J��)��m���Ln��e���$�S3��R=;����|���:)�A-�6���9'�������l�������[z��{���cm��w��dAti�W�ͷ��bzww~I�rff��qv���PP���^}߯���[�	7f�J��|�7gj�Vڬ�����5�6�x�u-n����������U��kvV~m������m��qLn�Ͻ��EO<�o{�f˻m���]޺3X�J�J~��M܆$��_�r����_|���������u��jJ"u�壖�Yl1����~_�6��ى㿒�
�B�$iE`D�;T	3����9�m�;�y7m��}�i�'�Tv�H�_�6��'�쟓��{���6��w!��.I���/ߛo}����V��Q-������sOߛo˝���~m���ߗ�ͷ��bx�o�]�'P�F1:�C��y��� �=hLs�k���l�x
��u�[>)*��$��P�Z���)�ͷ��;UUzt������mW�t�z��V�c,D���n�cm�����~��?{�bx�o{������n�3�\�6֮�}l�#���;*�����Y��m��y����ɹ�fr;�
ww{���;���b+Tpn�mm�S�߹Ĥ����6߹��&���~��[v<گ��0G0���T����w�"R�J��_�����{��R��o���T�pa*	)��m�7r�o���M}�j��߻��zww{��|���b�r��DM�x��z޵�/^�\���q�[�:��=�sI<]_���ݟ������4�;���7������5#ӻ�߮�䛓&������m����M��~Ge�Gj����v�yqq%$o{���������o��/߼��JH�����il��h���s��ͷ���c~�8���o�/ߛo���<m���dP�Z����j��w�d���e9]ނ����{������5#ӻ�2�Lɦw7�}󻾭i�aD@sYu����Ͻ��9m��_����y�|��߻��9m�g�o&����F��#�'�B�g�)R�3\����k���.�o3+�	pqr�$s�-�\hhN(|��7ʆ�j0�IHB�k�9�!����)
x���}������D"Sh��ɻvK��	pцs0 i�3�*���|�Hnf�K��y��F�mG|�)Y���MF�"ɼT�6&m V�0��.�L�6cc���EbFa��	7"�+�G\���ߤ @	�b���B(A"��X��
E �#��,P�0
D 0!�� �H�����b�E� �H� ��GQ�'��!�A��?lW�!�n�$���އ���(ċ���?_�'B
5�0)��40���mn��&�{0��6�+(��$�q5�&�����o� ������ I		���Q�eW��p�F���e��N�9\�Bn��Ui8u�H�\]�Gm�����n���锰Ӵru͸�n5c�8��.��#i�cb�絫b��t�ݰ�Fٓr�Xض���p�� �<�q#;��n6 $�ã��fŵ�n���C�k7���,k2�m�V�#i�nk���3�;Ov�VԀ�'?�`fEaT���E���ړp�u�0��V���v�9��2�킄�E���Cxۜe��v ��D��q���R��1�[��γ�'�v:0v�T�ݟ;!stiֱ��ƥPs�%�N�=����^8n��W&Z�x����#�#m�;�Oc�Ƅ�F�.۫cn�
�����O���e���%i�ڀ��^@�(�s�2��UUX���8�B�E9����۲9ñ&s�宦 ֶE^H,���s��g���i{F�n7S�Ӈ:K5�VmD:��N�Irjk3Wc���N�˭��n�m�@���+�h��
�ԓ�-`쭲�g 2*s��\������m����ܚ�6�d7b�W�n�κ�������;�� ��R��jn��^^d���u1�#��Nܖ�idʛ����x����!��$:����J�6.%�9@���6)yj��F�-��\j�r8� Thm�,�bv���;;���c��l��P��v:��r��7j�荵����
��꭪�(S����헼��L��H���l��nM�j k5�� � �`  �     �       m�m���vHp�q�殶�]�����IH�� 6� ��j���1�Z��N�
��P�B���~Ār�S]5��P{rpܪ��fk�u1����F�.�a1��*o@ت�[�N�=hF�l�8rm�*�1TuE������ 'r�Rf/\֩(]k!�f52��N���?>6> x��|A`��} O�j�|�<U�꫈�,9���k3	�k4Im��.�dx�-��6�Mn-���+s�7�fc[C6���z&��狀
����WmN7�qd�gy�f�-�j��Y%n����Cu���!�ĝ��έ�����GC�\8� �B�/���.�x`�D�����wn��MmiNLk/��_ۢWvn:��fZ� l�,��n�BX(�t"����A����Uۤ]Z��O����NK�Lљ�`�\\�]���x�H�4��r<�S4�)W�w��p?*sr�K�Bj�2�FG]rU����kz�v�}�߸s���}��uP�e�����m�5y�87c�����}���}��K�&S2��;��������2jG�.$����FG�Ui J�Z�~m��ڂ�����}��37$�3=�5#ӻ��o����m���r�J崖[m���Df��}���H������/�w}d�;�������ڜ'��Z�v�ߛownj]�m���w��-����Sv�~�߸s�����翇��t�̈6�s�]>g�{��d��m�MWr�6�.n��{���b��[%C�Z?Ͷ������m��r��ov��̹2I�����jG�wwΞO.�tə3Z�kZ9�m�}��6l@��)��$`Ȅ`��!()��ս����[o�wm�w��~��s��H�o=��b��X1�f���w�9m�}���woE3;߻Ü���{)����o;�Ȃ2:�Ӓ�ߛ�L�{�j]�m�~�r�o�}�M�~Ț{��}󻾹����T<��$�ėv�~�߸s���Q�{�jr�o{�xs����bx�o�u�j�JV[UnԬ�;D��k(����l6�1��f%��w�l�����w"ǜ��8@�V�_|�o��Sm��|����3&)?2nd���]߻{�����r/��r�J崶[Lm�����~�\\����eݶ�����-�������"�[��A�����K]����m�Y��v߾����p!U^���w]��1�߻���~m��OV7��,�v�S�w�3rL�g�z��;��wT������.r���W]��M[m���s!�j��Lɖ�m_�6��l+m�\In�~_|�~������w�����#���کc�������L���p�1���2�N��r߂�1�ݚ�3$2�Yu�N[m�~�q��v�Om��/%�/����{)�����7�Ȃ87J�e_�6��ى�Ĝ̷���9�m����ݶ߾���E̿3W���p��-+����������m��r�ߒ�9$��ߗ�ͷ�z�Om����>tkS-�\ѫu������W3�߼��woR�33"�̹$��$�!�2vD��X!�R
����
W����`��{i�I+���m�7o)P���2��/ݽJ�>�ɠ1?��RI��T-TrKh)R؜NN/9煲p���T%cdUt����w��g��n��L��̯��݊Te�* �3'Y&o�{��X���1���*�U�f^R�L˙�� /����ޥ@ffE*�qq6w���/ZЪ��-� >��h��TjI��n�Ҡ7siP��-��$IYGm�����ߖ���,w���$������姭�pn�蘕@^f=*����]��^ ��w�� I'ē��cnI[l��r�Y�gխ�Gj�9aXr�3<Ӄ�c��z��s�smݻ@@c�:�;��<;�r��[b�vy���H=z�G���nX��ϛ�pq�뭹�S��ɝJ����/��Z�3�ŻtjD�p23sq�nj�s1̙]^�������T�%WF^{I��m�ݎ�-�m�n��m� N��n,�*��3d��s��)��
{7a�]Tqm&'���8�sT���U�Y\+-r��K�E���b!���P�ڬN�I�uv��6���{׫�KTpn�-��W�����`�ݸe�/ܙ��7�����1�$�;ç�R�2��̚�sw6�������Y�ĸ���{i�Ime�ۀ{��T�cңRdﻛJ�=��@{3 uE�b&^a�U�&|���P������.$����}��#$V��ba�P���I�.I�_wO���ŀww^,{�f��E	X����0¸:u� ^��td�����g��pߞ���Ae�nIe�ڿ }�z���T�c��f��w6���eh<�35f�ֵ�'�{���<Z��'��Y2x6w�@n�Ҡ�2k�32\�� �r�y���2�bU������Tk2N�vh��T�^RL����-	eXI'�o�, ����7{��92\�4v�G���L?4�/���Uf&�ti�;�����Om��6�~�o��(�(�]4z�9�dx9zR��y�hV���&U�;����ݜ6$c���m���ŀo{�������~`}�z����	�)]�Z�X]�R�fL�&L���Ty�4e�,�8������t�[+�;*�;߻�rI�>�[���dHH, �D#�h�^(;N�s�_?f���� �f�Am�nDLL�Ĕ�2fw�����J�˼�T�e��̙Gv����-�䈄DK�<�����I2f[����ܝ(�۷ ���u��P���X�`Da��;N�M��'�\�W:Z�Bܶ��Ws�[�
�ʬ2����;�����ۻ}�$��0��ذ]��e-��u�d"bU~�ǭffgp����ͥ@e�E*�L�32�3�&�d��xt�(%��h���;�f�*.3^���n&�(8�mN�m���{}�`�����=�=��J(L}�
<8�ď�}��=���& �m��j�'t���Ҙ�L`zti������������"�^���G�& ��VG�.$�1@��h���<��o�9��o�/S�DC�J������&��/)k/�73f,��D���m�U$���n��w=����إ@_�p�d̛�Qcl�'�"9.H�3@_oR�2�"�ܢ76x���k�Ȉ�
!DЪ�ʿI����~�L`ztk ��uR�8G\�����v�k?�v~ۛJ�˼�T��9�ko����z�q�u]W�E���<m��mT�n�l^x�__e���eK#��-GX�h�r� �	�\7=��q�����g&��4���a�Onsv�n5[<��C�F{y�]&K6v1Зn3�0�i7@7i���N*���k��9��۪7BS�wl�7�Ѫ�Z�����`��,���9�k�Q��F���+O3�;�Lnf�K�a���K�����+�������"Z��v	Mŵ��9���[˫1��UK��Ո�����'ޭ	��-��Κ켥@e�E-K���(���@q��v���qg�l���*/'J �ٓ_�����b)��l�Հ{w��v��M�w޸��ŀ~գz�t�[hH�ˏݜנ^��w��9�L��Gn�yP��DP����n�R�^ ~�v���o��73b���Ǡ9��5�dQ-*3�3��[�}���	r�y�N���I�'h�T�9,�n��ϋ�O+�-͆�ͷ���Pw�J��Fc�I7��vhb����h��:�X���;�
qr����L���M�ѭ��AБ�a 	)Ī���F�Y�ə��Iz�����=��@e�R�L��W}�KTpn�-	j�=��< �fM�K�3Dv�R�;w�Pj���ZW�)`9^ o۷ ߻���w��q?v���{Gh�ڝ�fh��T�$ۙ�/�����{2h�7g2�:X�!d����"6Љ���&���Պ�{n|���h��~{��}?rs�}��m���n��f���v�$��2nd�/@noR�/���y"�8u���Ҙ�1��ѦI|�.d���r!A�����`�w�z �������IN����;�HW�ꄾ}�d��q_-�n�k۫7����p�^lޤE�$��kf�łBjx�\�>�*yᰜFz[�[٠BBs�d%hFH�dB(ZB�c�)�����Ä�.��+*�`1���!SY�j�P��^�R!Z\Dߓ̵ӈ�zd�F�=4l&���P���#�z@��A�04x>'#H�<U�H���<8
`�������PG@+���/��!�)���Q6�� � ы�>
)�D����Q�A�J~����=پx˼��V) ;%R�4ɒ|�ߕ��J��#1��2����$�
4E
�r���� ��/l����@]�R�97�hBדl�dt��|6ٵʪA5�:�=��4˫r�z^'���N��I�m�&¼�������4�yK�s3/@v�b�7��c��V���� 7�� ��)Py���/������m ���2�H��ٛJ��̥G7&M{�@��@g�:�w����̼ʠ�I>��ʀ�Fk�^d�G̘$�&a!2�e�*�X;�)䈒`�����@}�x��d�sv~/6���ŀs���5��¢��
��sm��jDf�<�y�prٽP���;�r:����=�}&�d�V��G[������w��,{���\���M��;�y��V)"vJ�rf0;z4��#LK�Lt��}�U@�����PF��c,� ��ذ�;�q$������b�5}�A��9DL˼ʠ�ܒh�����/ט���,��,{ʭ$�P�W�y�@s&e�&�����Ԩ�3�0��MP�X�����J�o��w{�;�5� �-�����;�{��ش/7��х^�'p�7F�1y�Y��kd�:w5��
�kn���Ǯx�u�C��unT�	���Pq+�7E��l�� Y��c���H���&��C=)R�l�G�/��n�틎:�Z�&gDv�Lʫ]8� v�]o��Kg6�   �l�-�L����2�k+�!yhm8f�8�w�w~�M�:��0њ�Mh։5�������8���r���[n#TJe�nIUV���W������Q-E%��o��� �����)�N�dWJ��t,�̂fU��J�&w=�����4��,��g�^�RJXYB�*�>��� own\ow}� ��ذ�lm�dk*�e�.���1��Ѧ�a�s��_y���r�j�i)$� ��R�5����|�7^�ˌǠ2���:����'F�)����y�Gh�L�4��R&�����G���7�=D�;<ƒ%|��*�Ǡ2�1��|�y�J����RX�D����X~��1^q��,�����:��C�N���`oO�0'H�w#.�Ř]^R̶ە��v�owI7���`��<��@n�D�)-������@��ذϽt5&��� ����x�����y���i��rS �&0>��,������#FF�)j���r�O�r��n^y[��7#�`�"���L��������:IK+�,���og��{�p��������b�=��p�V��FWk`��΍0'H����*���{9U��d���-�;��,{��
�@)*�����C5��z���\ ]_.�����*�ʰ��T�3�2�&�S3����W��Q��D����X~�׀y.?o����`��Xۼ*���e����Nnf��z,YMי��45�1�ݶ�d\	4���%���y�r�\��^ own߷qPy��2e���Ѽ��О!܉�&I"fh�e*�fgssv�{� 7�� �{�jq�L�-��Հm�R�=�x�jL���ݚ/v����1��-vXX�X\I>�� {��@_�)P|�7��'I�#)P\X�A��n�,� 7�ۀys�w�����b�>ٺ���]ldqG4�Enu�n�%wg�Ź��v|9e�z�N&�e������ȬM�IS��o�7wذ��T��ə|�m�� ,X�^be9
@��T]�*�f\�do= vwM���\̙�(��o1R<��"$������������1�7�Lލ0;�V��R8�v��x\o��� ��Ҡ=��T�fnQ�[�@j�GRܠ������w��{�������I9��krNq�ȚY� [B&!`(�Q(�� �P��k�$D��*�v�P9P��� ���흐����vػH �qɅ�k��q��w�u�y�OO<���Pu��z9���mT8ᱎ�kv��ǩ䛳�5N4�L�x��l���I��ժ:��c���B�Y��9�D���ݸ�g� �Q4m���{�@�Wm��  m��e�vĲ�売۵u۱��i�r�vM^*�������������w�CB�!��;�2+U�|�q.6��x['	���1UmH� ��7��w�������������m�L�&0'H���F��q[m����{;�?ĸ�(������뼥Z��0w �![��Y����\{�� ���X�n�����Ebd���-��{��*�6���A��74E�t��Z���20s�H�0��ŀ~��x���`{�%/*�2�Y�te��v�ά�Iђ˝�b����j�p�}ƞg����Z��~�M���y4��dɛ�zsz���G�gV�Z�#����ܼ\����ƒ_w�_|��� ������S��F�d��������L�wqa�ēzo� }���7�o*%����y�*��@e��k�2��=k�~F;V��D%� �ٺ��q���<I��oF���耮��
���I�1se@똌��U��ij�j��:0�d�E�d,![��Y�������oF���L��?�Vyuʛ�`�ۦ6w��,��|�ݙ��/.������^9i�w��,	�s����R$��dH#$���X�1$H�C����0�o����Gcp%�Z��Ps�'5�{݊���w�@]���q�9e-vA�0�۳ �_{s��;�{��v`�(>�d��pV���鵺^Ԝ�X��=�v6��Z�w��J�沢�m���r�Wl���ŀ}�ƘRK`ml����,W�STb32��bU�fR��h�_������/3)`�hެn���Y	j�:�v`fE�%ɒ���@fwR�>��
�*n�ll$���I�wޘ��Ź'�}��ɜQ$Th��NI��O�M/fH큫����Xe�d<��b��̥@rnd�fwyx~�����5��u�����䨖Ѵ:h�vt$�0܆����V;e��`Y`i:=�^�w#
����U�`n��jIl���}��q~a��b�5w��v7Y%��U��Ȯd�rL�ɢ|�w���۸��q��/V��I]-vA�0�݊�2��I$�w�J���ؠ-{Q��dU9#�;f���{���v�iP|̊I3=������'��Ve�f^&�06�����-������ �WzL�>$򐴩���aA�@��2�(Z@����z���$H��uOfɸ���%�z���D������B�-�����da!��!@	�
R2MaSHI	����6�_���I�	@t}@M�18�=���7th`�=��a)���4Cg��߷x�{�����T��U@i6  HHH�[]�G���-���;X �Nz����v����0c� cvv�K�pl�m۬/�<��u�g,t��<��nnY':��XLV�"��m�VMq�v�V`��ޝ&��#���\�Jr�ix�k�D�Wi�6�'9ݭ����=z)㮫�=m��E봊���������f�m��n:,�kd�N�t�q՛�^u=�hs�K�w<��lP{m"=A�W\��p�n]��ԧ]�wRݭ��t���1۰k��r˼�ۘ�q.1h�b�*��S͡�yY	9��n9������8�dC��Oj�N �*ݳ>ٕ��xD�H ��啴a�^)�˝j�ǁ��k]w��	��粮�sp��q�5��-�	s�Px]���C����)�H;U*��UNˣnin��#F�K��^����]��Ƅ�y⎣�n���q��U�t�wVV�דz��']�:P�i÷Z̛�w=r�V��Z$*Ƅ��#�W\�C�9+{9�i-0o(��U�a �n�r�[[ld m�j������L��ۓ[iڭ�		�n�dwX��䝺��^��Igl`�en�٧O%�[��I��ۚWL�{o`{^�u�k�;���9鸙	�ɓ���Ŕ���.x�W�m��h������XwDQ�q���ne����t��p4ͫ��f��Uq�<�F6-�
{A�;�ն��ivy��`���TF4U��+�{c��m�1�F�ڶ��iPS���^uսۚ��YB��u�v�i0$��S��A���   ��    ��      i66�/NE�x��J�s]m�p���
��lm p0�E���i�m� ��jٚc:5+ Pn�&h<@lT�/�R�k���t���rvL��/R=n�ogn{3�uSn֔--b�6�a��k�LҾ�����l�R�[N�[E�]%��v��+�jk[*�a���PD�`iң��)TS�_�O�lv���>Q�!S�aPN�w~��������^n..
)N�8:��պ5f圢^nݱ��N3��n^��8y88�3�yK m@Br����C8�˰���(�jٽUԾ���;uŷJq��r�CO/g�
�9L�S�­�p�ֹ֚7A^0D�Tݜ��؜8uF�h���[E�ϡn�c�ƹ���  m�
U���=+U�X��o���4��.Mi�ۅ;G����?}u���O��΢8�'U�b��6B�
͗�"��H��N_.%�A�X�n+l����>�� ���0�w�nf^���@^쐠~PJw�yyp"&�[%�;�i��#L�%����Wg.��P�A�"%�C����J���)`{�0�۳ :����T��9ʇy�A��=��ʀ��ؠ<�̊f|�{��5w|#(�n�KUr��wckd�I`n�� � ��-RD�Vͺ��|b�{]v2�z��N�<��Ŵ2�lgj� ����~�l������]���'H�vF��K`r؈�U�h��sY.]k7$�߾ٴ�X�H� S�H�0S��N��P���fMs3����'��<�LLĪٛJ�Ǽȣ�;�{�@nn��?jѽX�n+]���j�����d�y��5$���*٪a�59)�n��In o۷ �������b������h�*�����;D.�|h�\�8�wk�)�ΌqU9ẏn�����KMfkYu%�krN�~�xm9ı,N��xm9ı,K߻�l? �<��,K����m9ı,K��Zɒ�\tYu�iȖ%�bw��i�~T9"X��~�ӑ,KĿ���[ND�,K�w�6���%�b|{��~����-*�/�8���'��u��Kı/}�u��KkhH�"�E^Av���2&}���r%�bX�}���r%�bX�z}�s��Q�L���e���Np�4���v��bX�'����iȖ%�bw��iȖ%�b^���iȖ%�bz{�;��0�s2�f]k[ND�,K�w�6��bX� =����r%�bX��w��r%�bX�����r%�bX�����~6�N�������:�R���.F$n+,v��*]�gS��^��Lֵ�6��bX�'~��6��bX�%���bX�%��(�bX�'~�xm9ı,O:v[ӗR�ֳ5sZ�.�m9ı,K�{�m9ı,K�{�m9ı,O��xm9ı,N��xm9�TȖ'��o�Ś-պ�L�ֶ��bX�%�����r%�bX�����K�T\��?w��m9ı,K���kiȖ%�b|}׼0����ֲ�K��ӑ,K? �����xm9ı,O���ND�,K���[ND�,C�����a��	).���A���~C��z*?���i��'8��O�9i13�:2\Ѵ�Kı;����Kı/~�u��Kı/}�u��Kı;�{�iȖ%�b~�߹O�̒aN<�q�M��r���Sk�IЋZ��+r�-hj�˜�Y�u�RKBZ��Ȗ%�b_���[ND�,K�߻��"X�%�߻�ND�,K���ND�,K��vr�a��ֳZ5u�m9ı,K�~�� �L�b~���6��bX�'���ӑ,KĽ���ӑ,K����w��f����̹�m9ı,N����r%�bX�����r%���b^���iȖ%�b^��u��Kı<�퓭�.]�Y�ֳFӑ,K��w�ӑ,KĽ���iȖ%�b^��u��K����6��bX�'�;-�9�rkW55�[�Z6��bX�%��w[ND�,K�߻��"X�%��{�ND�,K���ND�,K��f���^����T��WE��t�S�\�f{�����:�;m��/<���tg[������㊣'N9��O����nV�<t���K���@�xc���g��r�3�ȷ%���8�6]�*M�Ƴs��w.��Ѹ�]t���VTۋQ�+���6km�!��ͽ�����5��V  m���R��5�F�T�;]ps�mmx�q�����*W+����qo:�3�>������jwG
�V�j\ՠ�/�{\�N-O���ۭ��t�r�>[�pA�k[ObX�%���w�ND�,K���6��bX�'}��6�R)�L�bX��{�[ND�,K�?�au-5��e�u�m9ı,N����r��DȖ'���ӑ,KĿ����r%�bX����iȟ�b�L�b^���kZ�K-��R�Fӑ,K���p�r%�bX��}�m9Ƌ��wI�2Kov�3 L�����rC�3I�$�ؗ�}�m9ı,O;�y��Kı;�{�iȖ%�b}����Kı;��g.i�d�.��ѫ��ӑ,K��w�ND�,K���6��bX�'���ND�,K�ﻭ����&q3���p��-ajn�V�B���3�r�6�;�؆�ݞ	R�J�V��\a����B��ӑ,K����"X�%���w�ӑ,KĽ���a�H�"X�'����ND�,K��~'��.�u��kY�iȖ%�b}����:��SF2&�X�>���r%�bX����v��bX�'}�xm9�$rP�g��#�$v�ilqڳ�"X�%�w����Kı;����r%�bX�����Kı<����Kı<�����f�un��3Z�ӑ,K?!"w_w�m9ı,O�~��iȖ%�by߻�iȖ%�b^��u��Kı:}�gp����ֳY%ֳiȖ%�bw���ӑ,K�|����Kı/~���r%�bX�g�w6��bX�'�v���u�d�]f=��hr�n"��'D�Ƈ+����Z������)�=ӎ@��l��%;�����=�{��{���m9ı,K߾�bX�%�߻��Ȗ%�bw���ӑ,K�j�^�tm7eh����q3��LK߾��c�2%�{�kiȖ%�b~���ND�,K���ND��,��,O�t�%�.MR�Y���m9ı,K߻�[ND�,K���6��c��F0!�������#$ ĄH�O��x{q?y�xm9ı,O;��M�"X�%���I�ن���5�2浴�K�,N����r%�bX�w���r%�bX����m9ı,K��w[ND�,K��;:ۢ�u%ֲ�f��"X�%��~��"X�%�'~�}�ND�,K����ӑ,K����"X�)�_)ѧ�#N#��HG��r7���]<�mÞVN;&�-q��j,���)us��YKWZֳYr�Fӑ,K���o�iȖ%�b_����r%�bX����D�Kı<����Kı<�����J��B��S8�L�g8��}s��(1ș���w�m9ı,Ow��"X�%��~�fӑ,K���]��jZk3Z�a.���"X�%��~�fӑ,K��w�ӑ,K��o�iȖ%�b}����r%�bX�庼[l�T)m3����&q.$�y߻�iȖ%�bw߷ٴ�Kı>�~�m9İ8��� E�@H� `��ٹ�y�fӑ,K���N��K�i0�Y�Mf��"X�%��u�nӑ,K��W����i�Kı?}���ND�,K���ND�,K��͹�Y�Y��Y��5���]�'�
��k�,���y^�&��wd֠�zد<:8��c�w�{��7���������Kı;����r%�bX�w��؏"X�%��u�nӑ,K�����l�E˙��̹��r%�bX����m9ı,O;�xm9ı,N���v��bX�'���ͧ"~Q!�2%�~����]��I���u���Kı=���6��bX�'}�ݻND���2&D�}�ٴ�Kı?}���NDg8���/��#��l��j�/�ű;���r%�bX�g�w6��bX�'}�}�ND�,�Ȟ����"X�%���3�f�uK�D�Z�ND�,K����ӑ,K��!�����%�bX����ND�,K���ݧ"X�%���:D�B @F��嚟�Y�L�f�.[�l7l�-]ZS\F˭Ӳ���ۺ"98����˵�ն�S��6�����y��.Ρ֭�����T�s\���tY�xԖp+{��G,�z��.���Dm�͢�x�bԖ:�\J�������O'd�cn!u�n�{i�{t�[u�s�\�۴�� l�6�:%V�7��sIX�v4��6a�����۬	�.qg]�YpU���_����2�g_6莎m�n9�h���@25w5���=t�Դ�f���.���"X�%������Kı<����Kı;���r%�bX�g�w6��bX�%���Y�d�l�I�5���Kı<����?	��,O�k��ӑ,K��}�ٴ�Kı;����r%�bX�|vNj]KI��֩u�6��bX�'}�ݻND�,K����ӑ,K��o�iȖ%�by߻�iȖ%�bw�N���u�5�[��ND�,K����ӑ,K��o�iȖ%�by߻�iȖ%�bw�}۴�Kı==�;��0�r�f�3.k6��bX�'}�}�ND�,K���ND�,K���ݧ"X�%��{�siȖ%�by����Q�~]��f;[#]W
�B�Gf2)�LVf���9ڠ����˗Z�ND�,K���ND�,K�u�nӑ,K��=����Kı;�����g8���|�'��;]��uu�iȖ%�bw�}۴�>7�U�D��ț�bs;�siȖ%�by����r%�bX�����r'�ʙ���g���Xe�-֮ӑ,K���w�m9ı,N���6��`ؖ'���6��bX�'}�ݻND�,K��vw	�i��k5�]k6��bX�'��}�ND�,K���ND�,K�u�nӑ,K�̉�}�ٴ�Kı/N��5��L��pԆf�6��bX�'���6��bX��E���?M��,K��>���r%�bX�}��m9ı,O��~���j\z����n��������M���S(m 5[TX�z�G}��,�
���Ȗ%�b}����r%�bX��w6��bX�'�w}��<��,K�~��Kı;�����:.��u�֮�56��bX�'��{�NC�Aș�����m9ı,O~��iȖ%�b{����r%�bX����m��.\��K�5�ND�,Kϻ�ͧ"X�%��{�ND���z�����Y��5n	~u��SL����ԇ�i�JRP��&��$��`�;�$�oE�Д)�L��BF�\���L�i�i7L��@ZOY�Cl̄ٮ	���c.2�n�ʉ8��f"�I!C��I��׺4�<�Ma�	j7F�%	14hB�T�xc	�͘�����\��orc3&;��u5bcB� J ��$"E��"I!#$H���ax��5�71��i5
7:j�J��t(&�������8[+��
i 6�'�<P�R���8z<Pu����&�Q!^ $ � ���'�����PSA�f�:X���<ߓiȖ%�by�����Kı/{�z��u2S/�N2s��W��T��bX�'~��M�"X�%��}�siȖ%�by߷ٴ�Kı<��dq?�q���l�8�L�g8���6��bX��X�{�6�D�,K�����Kı<�{�iȖ%�g�^OF��
[dV�D�r .m(s�k�p*��7L��Ӎ�Z8�[�q7ate�jm9ı,O�ﻛND�,K���ͧ"X�%��{�D�,K�~�fӑ,K���]��jZk3Y�fK�fӑ,K��o�i�~�L�b{���ND�,K�w�ӑ,K��>����ı,K���f��d��5����r%�bX�w���Kı>���m9ı,O�ﻛND�,K���ͧ"X�%����d�R�an��[�ND�,R��߷ٴ�Kı>Ͼ�m9ı,O;��6��bX�@��������.���q]�'���m9ı,O=�?ו�֝���q~8���&ql߻�ND�,K���ͧ"X�%��{�ͧ"X�%���o�iȖ%�b~..����7SN;BѲBB�my{JsC�2��f�%y�j�releeU�^����}�gR\�sZ�.k6�D�,K�����Kı<�wٴ�Kı>���m9ı,O�ﻛND�,K����.�ff���f]jm9ı,O;���r"�%�b}����r%�bX�g�w6��bX�'�w�6�����,O~�~���Q�(Ik�ʳ����&q3�}��6��bX�'���ͧ"X�ؖ'�w�6��bX�'��xm9ı,N���t�E�k-�.k56��bY���fӑ,K����p�r%�bX�w���K�V���ٴ�Kı:{�gp����j�Y2]k6��bX�'�w�6��bX�����~��yı,O����ND�,K����ӑ,K����6bdHF�WG�w{�?�&W���CI'���3�{+�R��sYzB�nrpy����H�m�G��wN�wl8����Gf��!����M��. ��q�� .�ݛ�ƥz�[ʻ	���r��j�"�y�h��݇��Z-���٣�p�:۳tn��� ��M����nwn61�݅�`�  ��0�iR5�Y��.˫S�훶oW#�6^H�����w��������6"�,���[�[N�OZ�^&���ګv���߻��۳����٭0��6��bX�'��w�ӑ,K���ٴ�Kı=Ͼ�l?#<��,K����iȖ%�bw���/ai2ۭZK�ND�,K��fӑ,K��>����Kı<�{�iȖ%�by�{�iȟ����22q�gr�Z\"D�12LD��ᓌ�K��fӑ,K����"X�V"{�߸m9ı,N���6��bX�'��'xZ\4f\��K�5�ND�,����"X�%�����"X�%���o�iȖ%�b{�}��r%�bX�߻/\���I��˙�iȖ%�by�{�iȖ%�b��}��6��bX�'���ͧ"X�%��{�ND�,K�'w�kZ�kT�֌޹�kH��{\��tg��3C3"Oc�B�������;]�гw�����oq��}��6��bX�'���ͧ"X�%��{���&D�,O{���"X�%����x�~,ѫ��Y���Kı=Ͼ�m9�tv"XYIdRФP�(�i,C)B��m��S"dK�<��"X�%��~��"X�%���o�iȖ)�L���/DPd��al�/�ı<����Kı<����KK���ٴ�Kı=Ͼ�m9ı,K���u�fK-�Za34m9ĳ�$��s��r%�bX�w��6��bX�'���ͧ"X�
6'�w�6��bX�'�����-��	sSiȖ%�b}����r%�bX~����m<�bX�'��~��Kı<����r%�bX��I-/ݦ2�.H��a�
]��֙MI�^�<�#��&���gf��ͶدF͈�im�������d�>����Kı<�{�iȖ%�by�wٴG�,K���ٴ�Kı<>�;���2��j\���r%�bX�w���Kı<����r%�bX�}��6��bX�%�ﻭ�"	bX�%����3E33R\�[��iȖ%�by�wٴ�Kı>���m9�� �B�@�F��8n&�\���iȖ%�by�{�iȖ%�g�����h�u�l��8�L�b�,O~�}�ND�,K����ӑ,K�����ӑ,K� L��s��r%�bX�w���2f�Ѭ֋t[���r%�bX�߾�bX�������i�Kı=����ND�,K߾�e2�d�'8˓E��H�I�v�y	Q.���|o�����E��sv�=��t��5�&ީy��]�բő,��(��Ӊ�L�q>���p�r%�bX�}��m9ı,O~�}�ND�,K����ӑ,KĽ>��u��l֘e�ND�,Kϻ�ͧ"�bX�����Kı/�}�m9ı,N����r'�*dK�z~�8k	d�nj�\��r%�bX�����"X�%�}���iȖbX�����Kı<����r%�bX�{ޒ^i՘][�f��ZѴ�Kı/�}�m9ı,N����r%�bX�}��m9İ �>�[� 1,��B#KIH���@��--�--%#!pI"@����BĘ匋P>X$`*>�OP���߷|��ND�,K��F�R9-��-�/�8������6��bX����fӑ,K�����"X�%�}���iȖ%�g����?�����c��)��X��ج�8��d�^A�{H��k�.upz\Ib��r�����'�,K�����m9ı,N����r%�bX�߾��`DȖ%����siȖ%�b{��ŸsY.Mh�3ZֳZ��r%�bX�����Kı/�}�m9ı,N���iȖ%�by�wٴ�H,�I߾�ie�2��sI�$�O~��ؒ	"}��i7�;ϻ�ͧ"X�%�߻�NDg8���,^���a-�8�,K����6��bX�'�w}�ND�,K�w�6��bX6%�ﻭ�"X�%�~=��Mk2�n��e�m9ı,O>��6��bX�'~�xm9ı,K��w[ND�,K�w��r%�bX�������'ݲR��Z�U�ݎ��������=��!�6W<�ڽ��֛ayے\����uy����I$S��Gz�^v[�X�J�@)��K|v*�Z���R��sc���z}\�Ή�>8�	:(R�M�f��p5m$:u[��i��Cu����.�ٷ#,���6Lk͉ۥf�f��  � U8�ldꚤ�c�۶3��[;&ƓN�����wQI~K�Rg�?Y2�qʇ-mwn'�ԯN�3ksp�u&N�����c�����}�R�0��X�)�Zq3��L��}��ӑ,Kľ��u��Kı;�{�iȖ%�by�wٴ�Kı>���������mY���g8�����m9ı,N����r%�bX�}��m9ı,N����r'�2%��g�����4\��֭˚�ӑ,K���߸m9ı,O>��6��c�V"~���6��bX�%�����"X�%�|���3E33V浩�3Fӑ,K?*�"{���6��bX�'����iȖ%�b_~���r%�bX�����Fq3��_w�M����7%��i�_�%�bw���ӑ,Kľ��u��Kı;�{�iȖ%�by�wٴ�x��{��������ϨN=\��B�"����ˋ�|���vl���6V��n�\�*]�e���f�Ѭ֋tff�m9ı,K��w[ND�,K�w�6��bX�'�w}�ND�,K�w�6��bX�'O����5%����Heֵ��Kı;�{�i�|
�|/�NDȖ'�y�ͧ"X�%��~��"X�%�}���iȖ%�b_�z�SZ̲۫��sFӑ,K����iȖ%�bw���ӑ,"�2&D�w����Kı?w��ND�,K����Ma,�m�XK��ND�,�	"~���ND�,K����ӑ,K�����"X�%����fӑ,K������N����k5��֍�"X�%�}���iȖ%�a����xm<�bX�'����iȖ%�b{����r%�bX�����<�\�ŻFl;���ێ
��9m�٭��ָs�N͕Ur�:�՝p���"5���,K����p�r%�bX�}��m9ı,O~�}�ND�,K����ӑ,Kľ���f�ff��kS.f��"X�%����fӑı,O~�}�ND�,K����ӑ,K���������&q3���ɸ��8�M�m��gD�,K߾�fӑ,Kľ��u��K�OO���6�O�����IT�YB��LHd�]���!^!�W�*�R�&χ�>@Ȟ��~��"X�%����q~8���&qww����U����M�"X�~BDϻ���r%�bX����ND�,Kϻ�ͧ"X�%���ҙ|2q���e�S���D���]k[ND�,Kϻ�ND�,K��{����Ȗ%�b}����r%�bX���w6��bX�'~��-��Y�d�]{W&�p��Z=���XEA���BMZ�'R�Wk^��`"��������K����iȖ%�b{����r%�bX���w6(��bX�'�w�6��bX�'�O��̚�Y2ۚ��56��bX�'�}�ͧ!��L�b}����r%�bX����ND�,Kϻ�ͧ"~L��,K߿��jaun����f�ӑ,K��;�ٴ�Kı<����K,Kϻ�ͧ"X�%���o�iȖ%�by�l���ԗ.kZ�f\�m9ı,O>�xm9ı,O>��6��bX�'�}�ͧ"X�"��A�3�PCQ�t�4�P�'7��ͧ"X�%�~���f�ff��kS.f��"X�%��w�ӑ,K���ٴ�Kı<�{��r%�bX�}���r%�bX��?�q��'/��*�宑mk�"O7.8�yi�h��j����:sz���W �Z35�iȖ%�b{����r%�bX�g��m9ı,O>�xmyı,O}��6��bX�'�}����4kZ��E�f�ӑ,K��=�siȖ%�by�{�iȖ%�b{����Kı=���m9Kı>=;�z"��T���8�L�g8��{��Kı=����Kı=���m9ı,Os��6��bX�%���W4f�]4˚6��bX�'���6��bX�'�k�ݧ"X�%��{��ӑ,K�T"{�߼6��bX�'{:~��5��ankSS3Fӑ,K���ٴ�Kı=�{��r%�bX�}���r%�bX�����r%�bX�i ���H�B$	3�_c�>�}|�$��Y�>"@��0�>}�����}�7�^.��=�x�K��T�!���u}����r��ɨx�,XF ���Z��)��ߌd�k����LH�fq�3D���e�Y%�׬m6 ��37���Sq�	�$�b� Qp.���$!2c��>K�	�����| 0�YH���/���bMkDa&�呄xI�/�*�&�C$4�L4I��B0��o�����.JK�zR$���!3��@�㶬 A�`F2�R��� ��8�7!�b�:��(��d@g�	�tMPС�������m����mp [�� I		^$�t��]ctf��ۇ���B�@.�pr����g5$�+T�ָ4j�6N2���Y�ӹ�����<0ω�ưq1�˜�y��e���s�:�U7S��umVmU����!��v����.o;wd_[��;��g�u����u�N�dVxv��ݰhm���vpqa�z��:�ӱ��<��È�n�#��a�=NA.�ܾ�N�b�3[3���ʂ���ϨC��!�m�tCm�l�i�4��v�1Ì�:Ӹ$�N�&�vT�uWYNw��i݈�q�r�<컕8����'.���a��c��t�.��رk�ѰX'^(�u���ɬ�:v�H�;bAܤq��ѻZ��6ݗ*4��v!6J��]N����es���as�J�[O+[\�æ�#��,�q�1u�v��a;x�<����p��<�3��ʅ*���b@�H�\�{sփ:���=`���\mV�.3��h�
y�rh{)ut%����BY���ڜ�H�hj�j�A�YE"�)MN��e�l��s�Q��'��r2��zճ[P�׮�Bp�O��Kk�q��qU�6眜�W�x��c�� D�[sR���K�T�<׳�6�c:V�2�w);�B[�nvS=A6_=$���6]��x)�͵P�/ex��竲�Ӳ�ͺ*�v�U�u�nl�G9�V���n�g��lq�c���ff��v]�ڀ�4�j��{M�!-Հ@�-�k�ڪڀE6�z��պ�<!5R�;�^3���PZju� �v� ְ ��  m�m�    ڶ       P�iN�����WP
�\���'����m����EjU���ReU�:Y:����h2�y�\��msdhd�'M��5���S��8Dg���Y��{��e���.y#<t�Ό��c��*Ⱥ�tq��1U]�qc �.�^SKu�5Ԡ��5�k��f��Z՗^hG�\]��>��'�^/����^z(��
�Qt�����L0<@�~��z���v�@����ЁGZ��q:��OE�&5�஍�y뛶\�.�qm�a�q��ٰ���ൎ�tI�u�mƜ�]���[mI�-���ʗmp�p[lf:���n�a#����������;e蕎����p���7<u��m��Y���],�㞴�]�Qh�R���:*U    v�Y4��$f]N�n廧Kd�#�C<�SXf�:����~����]�����{}�Y�&�n��	JI�g�M��$�G5<]����d�%��pWl>z{A�f�5����%�bX�g{��r%�bX�}���r%�bX�����(�bX�'�}�ͧ"X�%��{m��f��sZֳ2�iȖ%�by�{�iȖ%�b{�{�iȖ%�b{����r%�bX���m9ı/��뙫&fj��h˙�iȖ%�b{�{�iȖ%�b{����r%�bX���m9ı,O>�xm9ı,O=�Kp�ȇ�N����3*�|2q����e��qLr%�bX�g���ND�,Kϻ�ND�,�<����Kı>���3�h�h�4\�jm9ı,Os߻�ND�,K�G�����%�bX�����"X�%���o�iȖ%�b~�����ܸx}����u[8��ٳ�#����ۗ!�TfV&��������?絀�d�2]k6�D�,K����iȖ%�by�{�iȖ%�b{����~y"X�'��fӑ,KĿ�:~���0���5u�iȖ%�by�{�i�x����z�s�D�%������r%�bX�g~��ND�,K���6���%�b|}��9��-&[��fh�r%�bX�}��v��bX�'���ͧ"X�%����6��bX�'���6��bX�%��t��ԓZ�kY�sWiȖ%�b{����r%�bX��{�iȖ%�by�{�iȖ%��'��{v��bX�'����l�Ir�5�kYsY��Kı<����Kı<����Kı=�_v�9ı,Os߻�ND�,K��н��'���	�tr	��ь�rG$�����r�un�j����!�^�����,l�Y�Ȗ%�b{���6��bX�'�k�ݧ"X�%��{�sa�D�DȖ%��~��Kı=����2�2�E�Y���֍�"X�%�����iȖ%�b{����r%�bX�}���r%�bX�{���r(X�%���-�̽2h�Ժ4\���r%�bX��w6��bX�'�w�6��c���dz0#@1R1 0 �J�zb��UD�;<��O�ϸm9ı,N�_v�9ı,N���jZf�f�.��ND�,��"{�߼6��bX�'�~��iȖ%�b{����r%�`~B(dO��fӑ,KĿ�:~���0�YsN�]h�r%�bX�{��S/�N$�y�@]�k�^e* �����Sbt��	.��,�3�)c��E��Q�q���mQ`qvk�;���������x�K����})��#_�}��{ {��9�Wm��V����Z��2N�^�*׻J��d�rI������J;-��W�o}�X�qQ̙;����f� {1>4D�C��e�3/�#L�!l��L>>_�ǡ���C{���'�}��2�2�"�^^a����$-��})��Ѧ�q`o]�clnR��-n���ӑ��똌��EU�r1�\FΨ�1�c��
�%&�Ӻ���ŀ~�w�?0������y����aU��)��Ѧ�F���[v�S�\�@r�\K��	�a�Z`��@^wR�>^G2I���f�w�J��v�*Kh��AY*�??���>�w^���Tܢ�ʀ3��<4'�%�fd&d�ދǠ93]���׻J���xE �$�s��y��Y"$VV�|���LZ�K�.'��b:7���bq�/';���9�)���{K��[@G;n�����X�&�]V����+Ip����Z��M��Y���2N�f�'M�6�ܖnk���۱נ��m�(�'w6N5�T�ݬ�h�&ќ�U���<��L�m�  ٶ+Ż	�Rژ�[�6�"�ni*dt�NA�7L�j9s����J��B�H�mx{H:�7^�LF��t�S�Ge�j�9[�ͱuy��e�V�7��Ll�0=[ж�;� >�y%a,�Yym� ���,��(z/���R�L����xP�%�6���ڰ�}��?�7��b�>ｋ �tn�=P��XT�)�Ҙ�`{di�������xEQ�iTn׀}�w��}���>}�����6-���D�����Y#%Ms���cnC{��e�k:OT�q4�כ*m8�-R!��!e_����,ս`n�J�_/PwO�0"�~C�1U&[��fhܓ��~��5L��$`��,B$ ������jk��X�=s�0&���`��nr)@��h[I�}��ﻸ������,���0������9s2��`n�i�푦�z�ݾ� >�y%a,����V���X������s�07z4��&*2���cEu���k�����Ѥ�g5U6S=��U�I�6�f���:f�]�����[v�Sw�Ll�07�U��ET�ҦII�}����g{�ŀ}�{���&��7DQ�V�v�޼�@}��TJ��I2�g-�&�fc#��ʭ��~�n����<�=�����K#��xJ�X�'�}�� ړ�l��Lލ09w(���UuWxff&�z�ݾ������n���gv�$d�:էNeծΙH��O2���0���۷H���ߞ�}���>�R����ܤ�{7� ���X�q`�{��;����YUrڥu�W�{ה��S4A{��>n�P�Y<�2l;��J��Z[D� ���ŀ~}ҭ��})��Ѧ�EUj��b0yy�fU���4\�����@{ה�'���X���!�D�9�}�`w�YI�*�-*c���u���T�̥@|��x�92O���)S0�k�.ߟ��o��3�f�{]�j"g�T	ŵ㥻��ww��۵���ӰQ`n��T�̥@|�x��$ɾp��נi�ԕ���%�*�?}�� ��Ķ�����O�}�Q!�;3���(��L���ݾ����i��q`�ֆ�KX�M�$r`};)�����#L?%򭸧�`N�~w��U\�9e�����ŀ~�w��wf�Ӻ�����i���'9x�p����UI�	�T]���ݱ����p��ۂl����r v�w�{��.��W�#��~�շ�_Oo[�l�K�/�L�Z89ٹ�+0�/<�9ȩƣd{M�ћ��f��1�WE�1�)dy����js���(A�kn��Ǜ��v�� m�5�x����YT��<9м�X�N|�b!�S�t�h:������{�#�K�;757c��X�����qٺ�½J�Q�n�Ԫ�]6��Vd�ʚ��K/�|w�ŀ~}]ـ}��?���f���*�;w�%;��f&�WK`n�J`{z4�����Z�H�AU*���K0��׀~���&Q�Ԩ|[�@b�0D�VVau�Y����i�푦�WK`}�� ߍ[IdcvYlD�U�~�e*��\�ޏ��@}��T�$���<�j�p݆����3�ȯN�-���tę���ad�ܕ��]�WnKc^f&�WK`n�J`{z4���� ���oT��4ݲG� ���yR��BSeJR� E"��Qk���>�M���<�ۋ �wذ��6g�l���J�eU��XY^��b�?}��%ē>���;پx���ISRZ�m��q�����T�q�@{�x�����Ѹ�o)St��� ���f�Ӳ��`{di����b���̡eU#�n���Y��ҘY�\gr��ٲs[A��U�ub�$us����#�T���:Y������`{di���K`E�Ԃ0���.�(*�)��Ѧ�F�����u�ĸ�y{�Ե�۶�j��J�={����2(�2j�c�+t3ta1̔i x��ClKAH54���.�9Jb�NQ���@���y.��.�A�2�Fh�3|���9�0��$����Dԁ@�aA3d�K&\q�X��@���i�<I���,$a��RcQ���B@��NNM��\�pe�v ��A00dc����	9�E+Øq��s�%dP����֐1��X��Y$�mi$x�~ <AO�A=T���ʂE1X��8��*�Q�Oh�� ����>}���R�_E�%*���΍0;�Q�6�T-� ���f�Ӻ���Ł�%�?��~X����)J�i�d��yl��LwF��`z�t��;��?J�CT-Qъ���8ɺRn��y��m�1�ݝ5�6�gF�-q2Kr�,VW���ŀ~�w������s�@ݞ�x��AISRZ�m���#O�$���S��;�~���Lotn(�J�m�Kj�?>������̓;��iP��T��D>(����`q%�����>�����[��� �X�
W�I b.4P�A��T'�������������;n��q`I$�+��/o���^M��"wqd�0��ݺ�#&Q�M���2[7
�7h�4u	5�Ϧ��^��7��s�8�;����0=]	lw�0;�4��9D<V�6ܢ-� �����9Ŀ�% foM��J��ٔ��$�wj�}QJ�M�$r�`{��~�����8����`>���;�[��YUr�,V�3|�N���߿4��l%�ޘ�;��)*jK]-�-� ���,��-��c��٠3/)P	3,HH�L�¶YF�C �B����P`�SJQ�$i@㗮���j��N�Z���v�r�p��En{>�y��ݷ]���հ���ϩ-�y��̌�s��m��Dѝ�Z��|��
K�����l;���\�k���j�ڐ�S&�Fn��y�)����<�ʹ��az�9չ��[�Q����S�Q��u��s�Yb%YZ�  F�J��X����t��_=Nۊ�䪎حnV�_�RI%8�����>?\�(��b���Fּ*��'���Z�*����)z,�:�i�1@:���`�1�'F��`n�n�PU7%U��� ����7{���`J�K`E�©]feV8���2���)Q��^�ؠ����V�WnT媖J�?ĸ���0?W~?[ ��	:4��9DSY�M�(�Kj�5�������_�{��X�q`n�uhY�ZX�j&\��������k]cnU؋�,�])؉�����J�M�$r�`�wn��ŀ~�w�8��}��o�_K-eU�t���krO����@���~O�I37̙rT�_���zlP�y4���IS����Rڰ�n��5��E�$̓�w�4�m*�^���a�&ePjd�(�����4�0=�4���.��ŋe�,��lw�0&�i�푦�]-�?����\��˹���̉��	��H�t�N��d�&�Ú�Vz��7�?m}���Y�<���m*�fR�1��#��7�{���^���9\���U�~�2�k$��潬ؠ�٠3ה�Y�e�D��CҙBww��Lʠ9�oEI'�{��8�� D @�D� HH�E�$	1$!&��|��I/�������ߚ`!r*+�8��8���8�}��������X��v`ޫ��YUr�-�Y�3ה�d�{�/�׵��^M��;�x�e.��&��]%����rC�����x�k�T�icvyL�����q�Ų�̬��7�~i�+T��7zcwF��wF�8�C��붬_�vg�$ܢ3zh��T�̥\�3;�x7c��U�*tjY������X�F���u��eU+���!�f�[����*��k2(%/?���:�#IQ���(�L\ �#b��"�툸�� �\�9��UK���ӫikq�W-�2���J���ջ ]����K ?|��UR��T��! ;I+v3�F\�d�6�Mx�Rv��Kͭ��=���}���m�!�ڿ���L ����7wq`��ŀ���7"n�#�� 7zct�0=�4�����Jʙ,eU��[\� ��ŀ~�w��f�#��tPf��e�
"�����o/3�#L	QIlw�0�_|�~���`w|7 ̅�v;]vՀkՙ���37��wwR�>�e* �����>����o��+�fڮ*WDj��U�d�P�����r�|���k�z!ɏv���8\e�۞v"N�m�68��:YV���,d�T��ŉt��s��5v��;��yK�X�d����	���݅�̡��J�M�ct�c�����'���yҗK���cO��@m� �`�$�g Ҥ�tuL�sX4U���:Lrآ��۬���n�w?�I��fy��������F^�U�٦u`���ƨ�0p�
����El��������y��?*�r��ӽ��:}���M[L�$$�3@ffR�L�o̚ ��@s������ۀ�մ���+��j`{di�*)-�n���4��9j+P�n��Հkջ0ﻷ ��Ł���}�� =�/!�Kpn�.�f[ ��	:4����T]-�ޠ��ȂP��H�h��R[!8�Δt�;b�F�GJ�v-�n�[ 6�j�5��WXfe^cN�0=�4��K��ޠ;���;������KhYmX�Z~\�Jо���V'-�{zcN�?�s��g���H3!j�R�j�=�n� {דG3��m*׻J���<��
����,����}��������X����������+mF�T����`{di�%�-�n�����]�ט�)mR���E�	`���Z<��4�� ���n��7}�~���0Z/*�0�������t���5~a��P;ӫP�Z��v�d�����{{�`{di��|�P~�/!�GY#v��v� �w� ���â�fHԁ$j��_	}i|�/���&�&�������E��eU��[\� ����?}�� ����d�s34Ff����(�N�"],�e�`��ŀ-�{����\w�� �F�T7l����)�e+�{s=�gCv��#�j6)��J��P��b�.P첕�Vݏ�0ﻷ ����?}�� ��d&�
�����`�y5�ɓ���J���Ҡ/!�"��6yj�<¶�n)x!�p{}� ��4��u���L`���/*��2 �*��$��ߕ���בD�� ��?�!��xnC��Z���&۷�%�`��� ����ti�푦�@Iy�j��x8ᛪ��/4�,�1p+*�M�q�J�uKZC�2��H�����7/)P{2��̹������@^���2���,�Y�n�q`��ŀwc����v`ov
LMIk��,���fR�/!�"�L�oy�@n�Ҡ>��d�2��e+���v`?���'F��`oqYv\Ut�컪̬�������`{di��륰�s|�4�i�$��gڦf�y��x{s���Ӛ�#ু�e�Ԝ�n��D�%��r��ϯ�$�>h��6)�HB_=�hw<��LYR�!`S�usU0 �3��~fkq�7�]@"�ӯv�l��GN�F�XJR҅v������k������Ka����7��F�����	q@SYB�UJ�b������WWU���S�B��L�H�*�$ H��H�d!�!�@*�-F��B!Zח�#��2��f.�R��7���&Ќ~[�fe�l�2 @���\|v.vظ�� ����$�?ImjG �� �Ą�		)-�t�E�6ɻ�`�+Gl��m�&�۔v{TJ��MU�QhS��d�xm�-�f�d��8��#�|�w\�\�*�[��$�2�J��}e$�Ķ���X�FV�Z�6��ƶ����l�Ǚ\���Z��Nʷc�ص�Ϙ��snt@f��i�ƴ�E�V.��]�܆I��ӫ�����p<z��s�!u�1۪����zk�w&�T�9!��"�;��p�jX댝���a��1��i���u��t��M��5Ǝ��.-�B�רDQ���[(��B���`���sƺ��:���V(�� AÅ����	;'���^�����r8�2)vX�:��7�\��gUj6T��YW}U���yIvڧؑd�j��*s�X.v·;��]�U½g��˶z��9T�=�T㐳��a�Ս�\f��W
��s��]��X&y&m��+Kq`ջ��t<�/6�4vu��z:�\=vj��v��Yqa��ncqE����2�J�Z�]@BV I٪�.j��A��;iiX-��BF���9�Ϧk]s�Ɗd�sv�������b7Y���Rq��+��>���vۍ�Y礜��U��
�^nVi���Ȝ���k{Q�Gm�pѴ�x�4�V����'��8nl�q)��w��β�Z;WIiQ�=��-�[r�q<к"�v6�='�I�v]�L��r��Olq3k/fMlAK��V�R�[R���[ Z�:�ɣ�����ѷZ�l�d�9��`M�`� 5�m   m�    ��     �>�6�Ic�Z��u�@*�^�W����t���Ѥc��eA����n���l*��d�����5ͱ�����B�dM�6j�4�88yWi��<Y+rZ:�2뵻��u�uۙ!�Y�]��J�͈�f2��v�5,X��4�vح�� �]t5�z<���;��m��I�x��vh B#�R����A �4�#�Ah?��P~(8���Q����"(l ��GХ���35��5�2˫�Ƚ/i�	�d�)��s���M�]�-[y_rHv��s��/]/m�gjy��N��h)�t\�a��4l�b��g�ݖ9���KJ�t�\���!3��Bl'6�p�+���<6.���W=�r"�mԗ.���۷iy^�h�Vu�۰<�p��i��_UR�UU@��n�ڷV���%�u��H�dX{c��g��Fʣ�W��9߰��t��@���){���o��.s=�nۇ����5�4k�[vE�Nl�ۉZ(ڍ�/ vπ���X�q`��� ��ݘ�WuJJ�D�HV�j�>�e*�s66({͊2�k;��W�1Z��v�-� �G�����Q�&fN�y��^�* ��X��J�*�.��-���-��Ѧ�F��}ـ~��v2�%�K,�Y�w��*W�w��p��@y�y����V������I�XV8l�s�a^e.kin��j�%r��V���lT]��l�0&�t����oF��R�d-C��i-X�vgx�����K�+_c.��`{z4�������6o�Y ��j򨥲7,�:���w�Ll�0&�t�\��*�]U����0<��}�`w�ŀo��f�\O���yo����J�h���#L	�]-���-��Ѧɂ�O<���V�X��4�yE��X� �`ݎJ&�1�%�I�t�<�m�K`moK`v�k��7�~i�}�/�l���d�;f���3˜�f�}� ���0�>��.6}���u��%�K,�Y�owذ�m�%��9ذ�>�t|
���y5�ܓ�߻��y�{�15%���rZ��m� �������oF��Q,T��1�����t���N��`{fA��3��^4�b��j���	=�.��u��l���+U]����J�&���:��fe����ޖ�����2K;� ��4֊6�rV&ـw��,��g���}�o����0��ꔕ��\��U�~�n��v`?�� ���XWz���R�/,-�����f�oy�@_�)Pb����C3/�:���0�B�=M�87,�BـmoK`v�i����-���_͋��nV9���8x{�
x�W��wM4��ve���i8.��1��eKL9lލ0=� �����6���7c�I�����KV��g�ĸ���?[���`v�i���YC�1�0�H�(�Ƞ<���5&fd��y����� ޚٰq�jB�,�6���;z4��̃�Ζ����R0�����PVe�;z4��̃����>wf���:��`�[9�6M��κ71l�\I��{p�nݰ���ێ�g9�:��y����7n������<#ۥz��b�b�j�Ɩ���_2H��լ��v���"��WA��qKhl���vß[�!z��\�]¡;s뵣���.��݄d��m�סxM)��nl�  �`�_���t��`�mci<5Ju�vwg�V��K/�i.��Z�d�6�V)R���pFL����=��ɕ2�l���j�O������JJ�D�Eo*���� ����6���;z4��ܢ��+����"bJ��+�fN�����J����3�6n��&�������`v�i����K`{���*��H�er�ﻸ��m� ���&��O���n���b!-p��]�&�d��큵�-��������ʩ��B�`Eu{*���d��ܝ�f���	�:�T��:3�4���R�.�`z_K������Ll�0魛3����� ��ݙ�d�M�e�T��m*6�
�Ȋ.WJ�f
̶��Ll�a�$�ޛ�0�� }�uJJ�DʻY�x�ِ`z_K������� ��V��
Y%�d���;�Pə+�͏���Ҡ>�N�ӏ-���6���bfM��v��9��]Mk�]s�dMpt��.�z�^:�x�g V[kz[�Ѧ�d?%��/P~럲���uCܪ�d��W,�?}�ŀ~ِ`M��l��l���m
�2�ɐx��@}�(�^LQ�0���mNS�֙"�(�]!�y���~��ŀ}լ��YTv؜$�6��`moK`{�4���������l�pĜ��Wm�����?w���dnL��Q��W��Ue���`�T����C��J4�Ui\�{u@��9xՁB���il�?w�� ���0�n��0���`�{�RV�%r+xYV��g�\I�ݞ��_w� ���,���1[P��X�-��&ܙl��lwF�ِ`˾��v6�ܪ6�ˉq'����>߻�rNy����W� +ǟ#�Ng��ـoMN�o*�Y#���0����=� ��re�6���?|��/�U��?�t<K���!%<g���Kd���x���KTf�g��(�3�]�h�[b�߳���re�6���=�`{yk"��\Q�bp���7l�>wf���X��I$��/6yG$3��fe�^e����0=� ��sl�5umF���Ҧ�m�?w�� ��8P�̘��ffw�͚ �[�$���\��U�~�n��7l���wF��Iy��B _�!!�!8���?u�Ej��㊗�x(c2�����Rkf����F��q˰m���i�����&p)�䛶"r��˓x����jv��H/�O��������9�wVœ1g���5]��)��o6�s[i%:uٓ����/-\qEan����S��m�n�)c=�j�m�  m���T�V��<����l���1��� �]�Ѯ| !��{熦h�Au�.[�]d�b1ur2-��u6�r�4q6��ķQ6��ٮݚV�)l�+e?���l�����Ѧ�drU�UVx����`�1�����2	��-����y��Id���-�?}�ŀ~�n��;6`�wnս�����Dʠ�I�{ZPq��@���k$��}�`wW�J��	)�o��m�n��oF�ِ`R���$2i��A�/m�&�3����b�Hr��j*���q����Eu�.)���z^��i���Xz�z��v"K���D�34��|̔�a��D��8!�@���k�'>ϳ������l>������J9YeX���0&�\����`rޔKP��X�-��7�ٳ >��p����?}�L �Wy���m����f[ ��ލ0=� ��}2�wlc��y�tP��8x]�T�k�<�ܧعsRf]��xW[�i�ɋ�멕:�����Ll�0&�L����w��))k���Հ~�n��nˀ�1������Qj�w�wYyh�"J �fD��y4f�j.�N�,�H�3�e��N��Jpm��<�=�MCl�,Xl���n�<�ڹ�֦��p�Ի9�[Oo���������i��&ba �OJ�;�9i><~�����fk���#����o�7��+	�����l��a��C~�	35,d��5�y�U�ao�x�����}���o!5�KB�ry�'�A��b3I��g��!)G��kC�M���c�|�ݨ2��o�=M7���pI��lԺ�8T�a|%��|פ&�"bE�(����	C��ƍ#�U�G +�ba�#��<���Ji�g������>�F'�2���"$�p����H^���r���H�7�<+81 `�����q��i>P���@0�}_�ڃ�SHW`��Ds�z!�(�wdC�W�Лx;�CC�#ꇩ�_|�S��od!A�ڷ�]�2�fbh5���f��fҠ>�N��s��w}.��y�b������poF�ِ`z^07o�06����;�宔�I��]�F��*-4^9�m0�� ���e�:��n'��0=�a�&�d�/�ҿ|��6O�05w|є�����`��.�Ӳ��0=� �r��+�Te]�^#*��})����Ӳl���k��Ul�H��p����?or�J�_�|��B�H�ԭbI0����~�W�;��>;�̻�e�Y�w����`d�`�1����X�ė������)yi+lWmB�Mvy���W�gU�V��B�8�&�Z2(;+��b$r��=�z\ ��ۀ}w���o�=�:P�8j��QLZ��\ ��۞K�M�n�����7�fys��^^��Ktd�MۀN��`zti��.�oL`�𕸈덕U���}�� �g�& n��oF���!��0�ϲ�����.��L`v�i�푦�$��q$q-Y����"���|�J�^�Φu���m�q�]���i���Q�2���;�wmg�s�w��.��������m� N��]t�뀀ۆ]��=���r�wPd��l���dMsی����x˜R��_m���y�j�M�{p]7Z��1���[�m�  6Ͳ-Ǚ���L�ș����4��|6i�*�����n�s��g�!����r��h	��Ѧ�!qkR��b�T��Sm�f	�uk���7e]��}�yw���1��Ѧ�F��7d�?wX�&�cM�]�ۀw��Ll�0=�Ilw�?���F����4))Uv�$�`w�ŀ~�7f�I���\��ŀ~�Md�x��b!-Lu�[ ���0=�4����eHKme� >��p��ŀ~�w��ݘZ�����u�vk=k���6�^0�����=�'�qs�i��8�|t�e��X��$*hv��wwذ�n�`{�K���E"�/*�VX��Ll�<���*�䪩$��VX��_�T�;A�=�?[ ���0[ґ�XaW�e�����K`�1��Ѧ�n, [���R���r^XK0ﻷ ����#Lu�[�(���س.�V^Vefc{�Ll�0=�Il~����q'��q�Wj��v�J�㥝�+	�n�谜6Jդg7�Kv��ajW��\))U��$�~��ذ݆�������q`���9:�vX�KV�����L`oti�푦Ȩ%ӂ� r��f }�v��w��uC$��UJ
�EU?w{�O=����\,N�IMy�ލ0=�4��}2��L`u�V�[���+E�`��ŀy{�/���~��F�&D�V��V��g�y��zᬳ����Jۓ��7j�5�Ѧ�KZ-t!G/,-�`�{��7zc��Ll�0ܫ���UWuw���`�1��F�ٻf���T�Uj�7ev�n��`{di���`�1�Г�����e�Z��n��>ٻ& }�v�VDcG�)��EqG���պ���;,!-X�r��ޘ�ޑ��F�����+;�����+ֹ#�=�=�˥�8@���9��8	��(�:�.��˄�ݰ�A/1��l���T�̥���p��،�W����%�,�?}�� �^R�=�y@c��+RI��Q>���Mn"!�QY*�?��ذ�nɇ��I�>���ذ���E��(������}.����=�4��Ѧ �uw��M:����[& o�ۀ}����y��dfDPt��l���2HbАc�V {��p�.��ɠs:tni{m@z4���c��Gس��v&���CrYď<a;s�zN ����mv��vk�,9[�XL>��[POlNp����k�Vu�%2�+�s��ʛ�C��&qج�eS�rVܖt���SY']9rJ�<��v��3	��m��n�l��`� UH�:�YT��������ܢ����iݬ�MZ��� ʀ�E��<35��)y�i�)݆�wV�%y�4�E5��mvi+�;RFo]\�U��~��Ƙ�`l�.�oL`t$���w�*��˫�LN�06\�l��0?ww&Ϟ��^G]r;,$v�����v���F��`{�YWI���2�*�.�oL`{�i�������[V�,R�VZ9f��)P�����͈�1��(�y݀�m<s:θڹ���8�ړĝV��U�1��9(I�����}�'i�z��gغ��w6���(|���8e�Ҡ�x��t!G/,%�`l;�<�sP'�SU��,N�QR�D�B@EX�PL���s>�L�Ѧ�`ܻ��Q��˼i�&(ȼz��J���w6�{l`�5:��Ti�hK+�;��,gF�,�l	/�0=�Ю��Uyyuy��'F�,��_J`wH�����FI$�Z�U[%�rH�׉U�l�����b&�%U`��B�җ~e���DH찑ڿ�Cޘ�����ŀw{�����ƱP$�Z�l�:����4��Ѧ�$�(�)J���w�fyl�`t���H� @�IC@X�;Om�w��>~�L���N�"!�_,�`ލ06Y%�:�K`wH�hR� 2^Y�`l7f׽ـw����w���/<�	lq�Un��x��W2�{uA\%!q��u[�GUӭ4/a��sʜM�I	/,-������;��Xw�� �a�0�N��V���$��N�06Y%�	�1����1
EUN[c��~���>�n� ߻� �wq`�jz��뭖�8�T�fO�/���4�e*�����(PZ���0�C	$HЕ�� �W�����y�A�@��Jݳ 7���;��L	�`N����Q�V��1Q#������Z^������������^4�-MЮ�Pr���ŀoה��|��o�5�6({�OK��a�rYV�wqg�;���y�}0���<٬]��� ���V�O?����-��#L	�`ܻ��'�D�ļ������3{�P��XϾ����5;�*�Q�����0�2����o����ؐ-����TU�ڨ���U����U@_� ����W�J�
��QP?��� *X
�D��@R"�
�H
�DX
�E
�H��E *V� *�H
�X
� *��B�
���D"*`*`*`*��A��@D��@@��@X��D��B�
��*��*"�",��H����D *`��X�� *Q��EF�(�V���AQ"��Q *D��D(� 
� *","���D ��b*`*� *�"�
��"�"�",`*�,��"�H��@H", ��@AB(� PF�AH",(� ��@R���Db�����D�,� �E�@_�� *��TU��U@^ 
��U UҨ��@_� ����PW�  *�  *��1AY&SYc�+	��Y�pP��3'� at�@lT��  � ���� �JPIT*�� (HP(�T��HT
T �@�(* * ��
	E%  �R�   �@I U��
��J�`     h 
(*1 ����.c{N]��`׼< ���kq���}<] Yo���f�� 1�z{��}��9��{�n[�.a��X�}��G�>�w w����t��{��> �|�� 

( �0 ��O�+�ݶ�A�8�� 
#
�u�q�!ܰ:qt�@='���� 3�F�� �����W�s^l�e=nm(��L�@����76��r������@��14 }{�o���nͯ3U_p ��S,*cCʬ�P{� c�d�4��;� wW�E�ث� O{����/]�q�/g>����E�'�ru�q�������{�x9>��U   ���4��F6�ʹe͙��,f��X }7>�R�,��� h�7�(��Ҕ����Ҕ��Х)����Ҏ&����t�� ��JR�Y@�3��J)O@�K,�)F�Δ�.�:R�w3��v==(��� {� 
�
P(
�` =�R���)Jb4�����[�����������/^-�|���E4��=��� ��-�x��>�� ��$���}����o���G��r>�{�{=����  ��JM�)UC#��j	�R�! F"x�T��   "{J�e%M   ����)��R�  �F�ԤRh4MMi����������R�w�;��>���I$�k�ow�� 
��@T�E W�J 
��P U`*�~Ͽ��z�C�t���B��dHI#��i�ٯ%�oF��d$"��,@D�҇�������P�@���d�,����d0"�$R!$
F����@#��0��B4t0��j@�"I#�ԓ��AbI �bH���c$�]@ ��F0�"D��B�T�&P�$	 `�đKv7,��ܻ�P��ie�n��@�4o��a��j@�q�D$�Y "Ae��H�A�H2&l6�h6I#"B�(i�$@�{��4�6�!�J���7�5��v���E">/��J��d��90����P6ʐc
ʡ���X�$*4�i�Hi�Ad��$�I��-�oPѾ66zm6P��7A54��5,a�H!�	����@D�,�S�Ep#�@V�+l�MLz�J����J��K�k����Aca_"�+J�&��a$`��B!�����k� �"D � �nŃ$X�db0"@�Q�գ$�1-�M2�)���mцjU&�A���A��u%)0��bA�AQ^:�V��,�$�T��(J�$&���������m=�Ս�h#u��g'8�C� ��XB��9���rC�1)M:7�	�pऊ>	 A�F�fBBK�S�C9!���E�9|k�os{�]*t
%
��N���|P��΁�ĕ$#�I�j2q�`�5�ተ�I-��2��H� �� hc�(�Z�
�JB��fM��cC,�C���MӅ%	M�9=u�o��sfl^h�o"�T��5��(ǩ��(j'-��,˷��҃�va[�F%��7f�Y%<2#B#	!�WT�m��B�D�'�Cm �B^�頉7r2O!O�efV�L$ߦ8����B����H7Fi��Y
�cL� �OK��taa��e�Av�]�	(!R榍��˫`٨xc��=c]3lo��
@)B��I)&�^�0b@�$ZB@�N�z�xK�СK�/ǔȠ*T�H�-Rn&��;���P���� Y�l���M���&D��<%�
1��Q>r��wE�2�s�z�V%IHda
-�&�S%"w,�{��J�N%����"D1���.��(b��  �HR"XQ��$w� f͍X�%eV�X,c ��,X:cM�j�Ć� $�b�H P!	�tAd1�0$d"$X�XR!��4djŋ"�SD�Ņt;#b�$�`F#R5�`HR@��I$A��bB) � :M��&I �R6Bą星xm"H�Q��P����F�F$B*�I"�aA�
$X&��hh��(�Cl�!�"Z&�5��*H��5吾�5�u�֔�	,bP*B�B��	t
�^Jԥ�&$$/��w���{W�]��vq%�+:���JYQb�0�~?����$א<���!*fsn���F�f�)�s|n�6p��MF$��vp��TАbE���# �,�R!Si
���a�:0���,jiٵ`SF�񅍘6{���
�|��D٠ф����S����q�40#,m)M����6q�V,�/�;��p�%M'A��S[�\��{�2�����t��3V�q�
M����l)�	�SI�m3����{1� �q����*��F��k��p��# ��"ń�ȋ���	�a�a �a��(jCk��$xq�RBHD"1�6D�BFp�$
D�R�C�Ą�0�]�a/�+�^c%)�#�����ە�dD/@��(�##X�-��5b�j�㲧��6�D��0%u9���h��TE��vP)��	yX����M�.N�[��xzS���uM�,�|�3���t�����D�V͚*bÞWa$d���s}T�6���#*\��.֨��b���H���Btg�&��0���I�u��z[1[�H��SB��S�7E�~��߭�Q�xs�Iv;(�RJ�4+ār�7r=x{-e�O'��t[-U��Nc1��A��S�My��Y+�C�KR�!�]b�<f�aYwJ��nk�y�5��/)���u��{������]ı�0�+�+RV�XR6A`XU�!#��*���H:�M&�"&���I���!+L%4���1�K�CI��rI ��vnX%�#D�-�:dT#u�C�	u�x��2f���3�])� �����=ᆒ���-�$DƐ�ٹ;v��$�6�-NmLME2T��[���V�EKՎ�*թ(0�-�Ij�mBB��\ʡC@p	$^L:[J�(�(s`{�b^�#-�c	��R��Y��(̹DE��T�P<�]N5JF�d�L�P�B�[녱[��/0��ޭP���c�|6��6�)&�0�$6q�$`F��,I
F��h�%��m$	�bI�H�B�'=�'�ʐE������t�0��8HEhF�+���ђ�ă&���_XB�U���LhTġ(r��)�pb��|с��@��"�XaX�
�jJ�F��FD		 @Ml�!��BI"؅A�I@�M��	����x�,}���&yK!�� v�Q7��
Ɓ�R�)�^J�Jbp�KT�E[�3�;O�A��S[!a������)��}%�|$�p�b�F�tZ�G���V�Lb��iޤc$H@�6B��hZx�xl[j�L߼"�ڠpݡ�j�6�ִr�x�ޘRHĺa7�%��4������ m��#`$bՑ�B�����sz4��]}|ӿ���6U��}bT�w�q��Խ
V4?Mg���H�K)13D K�����y�1
i�F�b]��徭��)Nf[�1"�R�l�
:�u�
BD��7�ۭn9 ���e}=��`��"��@�B�e�a�dQ�r(DBM�0`Ո��"A� �	s�� ��H�P�JA,�Զ�Z�)�V8b0p��ַ��7�
�(A��癇���mx�Im�0��J�4h!��)�"M�nnj��8$pM��(D��g�w�;HP�/�$�Z����"m�/ ���"��S<۽��� h��cJ�d���H�C,�6U�˜�%4�(j44o��8kn�ńc#'֙
L�nW�֩$����l>�\I$6!
��Zk<��[\6����%4�4�^Z�����aXU�Tȶ���j.d�2�B�^�@�<���x�S4���)�J�1B�x��lhJ�ը�^p��B�-R�"�� B�)c-5�%�����I�uXGP�#2�z���p-����l��4l�`f�̄IXl�H���A�Bۆ�O5�ʱ(��*���!!&A���T�*F&�sS�3�KM��ֵBh�a�H�
{�cRĈKl�T��REؼ�WUfΧ��M��g	NF���5��,ĕ�ڐjhٳ���l��l`]�ى�$���xJh�Fm%�P�
�:�]H:�}ǎ���#$�	^��@���\i^�K3<�H`�9J��8��"�����m��X�oٚ�.��
E��.a=)�MrB�<��)iَVB&��sF�sG	����A�th��,/>!MK$��X(R��&�%(1��BQ�&�\za�14l��o��8 ky���ۄ'�rGW�y��Q4��&�z<89/7>s,ن��!R!ao�� E��@l����#j����T�� 5d�P��4��z$	EY
�@8r��{��U�/P�e8M�d�ŭ��B$�#�1\�R�5��Q	 @�Ȓ 0�	X0���
@���ЈB�(�Iau��H7N�0����,	!J���U�lƚ7���~� 6���           �m 6ض�       �[F�Y�;�7:�HaA�V���m�U�����sM�!v�l�Yȼ��P�:l��/mFC� ��	�����NjZ�ƀB�Plֶ�[�T�0��c����=)*��᷁Ŏ��鹌vѽ�b�a�WIjK8қ�ַM+$��Y{2�'�U��жtֻm����o��	��0 m��m�4�m�d�\�-"��r�T�����k�I��w`G�5m@U_}��r��� 琗�0fٳgm�h�`-��Q�Y���mͶ{(��d��զ-�F۲��m��P�#� <�˽X�AU]b�xD3pMO(�U �8�]6�[`�d���c�I�c�J�pAW�2�q@���*ʲE�/-�]�m���:j��-��ݜ��`M���� �m'f�����m�el8 5�P�hm� ۤ�J��,T[-�U��VQ��Ueٍ$�hm-^� [@���[%m��$q%�u�-(6֯N�Zl��I -�����ֱm  	9!  �� -��ۀ4P7���6؃*�Z�-�g[��̫��:��,1�"����*D��e UUul�;E,���p-M@  ^�m�<��,�ݫl�2pl�@6���� �m�km��pj�� �%۵�6���q"��>���� ��` �m��uV�Ѷ��,�-����	���UJ�܂�P�� G �m �m:��am k]xb��Q�+�*�*�k�[M�,���6`LB*�j�nW�<���*�T�-uSʕ`�Z��=ev��?w���8���ژn1U+%�\��f�^��m��[�l( �FA��m��ɴ��ēJ�jk5�kX^��a��m�:�Zv�	(�.��ۀ]h�i"M�Vv�������sU@:@��.���jBj�u�d��m/n�#��`v���wm�n�n�$9n��u�v{N����q��*��&��n��j4��{v���ݜ�[F���m�8�96�^���k�V�[Y��]�m�s��  �j�  H&�ۖ��-�mZf�� $��6�ݶ��r�5V  �E�R��m�h[G ���TnXv$:@�� 7El  6� �	������p����+.ˢUz�W*�p��m��;d0pv[V�m����� ��`�i��m6Ͱ ����� � �}h 6]n 6�mٶ� �( z�-�` $[\����b@?h������ �oH�̫UT�
�T��-J�C�bFH��%ٱm�7m�j�`�`   �� m&�n]6 z�]Wh��6�rM� zޮ �CH�UT�UR�J�J;`q �`� :EKʻ/UpJ��7UT�J��A�l�@���WUS���%Bj^W)�d& ���  �� 6��7 �ͻ`�E�m�� �M�  6�      浶�   m��ۚM� �t�   �{98��%�#-UUJ�P5� �ƶő��J�Y4��b7HN��W/-V˶ͮs�
�PN���ꪧE�&Tf������t���Y$��oU\�PeG*�]�K���︉�a�j5p�i��jڏ[�m�R�
�V�7��V�;<�uT�GD�R��֜�n�  ��w[��$�8m���r�����@6ۀj��Zm��s���t@��M�L�:Nku�z�Ic�`�
�V�h!�b�!�fěl��(%�m����e�I$��Y^d��-&����o���j�{]�_+�!J��c]t(m5�
��������7��e�'HJ��m����g�5�M�m�i��մ��Y3VU�]"^��"ǛB�6�m��Bn�:�;�e��UI�x�İT��J��96ȹ�q
�j����7��y^	ԛq@�H��n,�͜:�n�U^��f�N7K$Ivě �kp��m^�r��Iz�,����q�TQU�E�,��hIn�m�� ��ID��u��p�[�ݶH��%��u�f���@�ʬʁm�n�`� rGHmm�����B�:8q��*�)	�ir�m���,�T��+��KR��v�h
P�[d-*U�5T��ª�UP �\��K)�	���[m��2Iv��[�m�,�� 6�h  ��l� m� ls� [Z/ �m��!#��3_�>m���m���v HӶ�m� B�YA��6��	f�7T���Ip�lQ!m��pm���պK;d�M�8v쾮H�J �t������#�6�m-��.�6�i�[%\�ӡ �*�*�Uҹ�Z�� ��l�@�b�$�k�6�4�j�xB퍶�S���Y[PŒ�TƮ�V�v��
�W��bR�2�sʵU�]Uls�uI����kZL�-�;7)5��2-�{��9sŞ0��8R&�OC�,8�9���A=�`��+��l��467T�<��nC�Iw nn���kP��2�l=+<f�T��r����3�L� HMW]Utvq�i7i9�db@�m�bnڶ;v�h��U��<)]T��q�h���V�u+��������RnF�kh�m5�(,$�09�[\s�h�z����ۭ��V�� W��~(j���B��d�8��2첦�i�T�hB�3E��ļ�JzV�vU���u�J� )Ki��� ��l$I��m�"H�I��� 4�+l鲔t���)�Z�6� ��v�Q�z�6��m� 6��rT�M-֨   ��f]{[�m��[��k��  �m����v8	���'m����k�m'P�N��h 6ؗ��HmkZt   H@ n��  ��  l ړ�ڶ�-�h    n�-�6�  6�M�eꑶ�*� mM]�b�N�kf��K/2鈓��` z��`���k��eh� �h��$���  -�[A��ڶж����  @ H   ��ͱ�Q� � Hm� m�v݄��|���i�iK�kmC[F�tKV�UJ�ʵJ�ё�u[;T�Ys5m�ҩ�    9�Ŵ  ������׭��.�^�@��]�IX3p
��?/ʶԫ[uV֠$���sl��m  m $6�m���ٶ��` m �mm���-�m��  Clհ�$ [�6��-� p^�[v� 6��B���k �\m6�m �6�6�� v�f�-�{i$    @ ���m ѭm� �aIk��^@j�8P%�@T����U����H ۅm����9�� om�m��� m���Ҫ��Ԫ��[���n�v��n�e���j�
���u�m�` 	$��f�@{j��m��i��&�^ m]m��}�΄��@7m�ꀶ��yz��OR�����7C8i{8f�*���
U��V��J���;@�g�ཫeݔFG\�`*c�n�"v�vs��m���4�^u���	68����mY �`�-\�Ssn�a#l���p:��3h_5m*�54�ۅ���jڽ"1�=�p�0� V���[v3��V�}0+��T쵲ѶK;���N���*��h{.�*��X
�UYZ�&H0R�%�if��$���� �HM'\2�sJ��m��iJZvm��ʵTjiP<Ҳ�f 
-�ˮ� H��@�j�K�S��x��.�ꪨ9�I�[�h �e��-���C����|�h B@��R�� �qJ�UU 6�$[4�'`ڻa�l H� m��� [@ mְ  6� ��� �`�m�m�e���n�B��} �[D��R*�UJ�J�q�� �7i���� �m�e��           ���n�m�4SZ���� �H
�`�����U4��`j����Ij�*UU5 īU!JU!5Uh�$  /�	�U*���h	Z�-U//O��u��X��� �m\sF��'���7i6�K(��#V��t����v`�r���k��wb���
��v��Ij����vj�v�Dn�ɔi��Sm��y$5^�h��z��J�K҂@:�٬Ν�N�6ʀ�Y�*�2�3�����h�H�Xd��� 9 �t�mΎ��*�UR�V1Q*H���k�6� HYA����+X�A�ڪ��l/\F���-ln�D����Q�/�w��q:UTJJ�P�x&����Č�M���U�֛- ��h[��Ir�n�[��-�/AbI*�k<ٜR
R�K)�%�P�e����P	/��N�m���:�v�iX-�K��	4[h [dmٴ���[k6��`E [)� �`��e�Z�mh�}h��Ia�6����mKC$�MTj�5�h�h�-WT�pS�Z�\@����/�k{���*������8O�A*���v��!���/(!��Lh/ʨ���D��1D�,P�ȉ���1�S�q҉�lA(	� @��&����
 ���ػPҎ5�����D�" ��lOC�]�DS�1�=U���0Sࢂx�z�S�4徚T0X�áO
 �<Sb�>@P�N �A�>LN(	��< |�U<0CR�O��TJ�M ;��DN
����"������v�G���������	��E\A!��iA� R EUN��x(��E��D����#�L�@ء��Fx
��T��	�Cj���1U
	��>���mpT=����+��~��� �T<�1��H�"���P��B D��a1�1!	��=_ ���B:��X�Q�!P�P���Lb'Ț`'�*�a(")�Q�}x�y�0A8����|��Ep��*@c0C�v����T�`���8�M!�T%`��?� ���E! �)���{w��������;/�PR�PRp5UVS۰�G^
��&�-9���S���wf��m�u��GA��3Hlf2hT��R`Z�����ɽ��.Ξ̥ܶ݉m�Fs��rndW�q�-�2u���X�p��a�s[6�$ h���+k����a�E ��4�݈3J�$\���H��)]\��a�V˨|rc��9k�7Wek5��:�fv�k�����j�l��yma�6��͜p<�gOc��	�nWvu�ͮ63u�;��U/;+]�.� ���gB�Ui� �'�1��eؠ�,�����m�#v��-k7$�8��i��-kv��J%�WD���gl��	j��U"�-UUW*Ԯ�NR�<��s�9�ۭ�Ll�;q7VM�Q���u��]�2�욧wY��`��i1�a��G=��`pûl	���h�v�-c�.[��rO@��%�G>��1�����h��� dVD:7Blt֩L�,R�D���9��.�nwZ@�!R�6��tWpJ��\.^ɵ,�g����/+%��<�$�5��<k4[V�cԮ6�gd���$�2;p�v�0�]c���)�mY��r��ۧN݀EwZ�-;g�D���-hx�cqm:���S�C�I#��k�lx;.���ۧ�P6��%Uʲ�UtPF�lm\��V*��T�D���T�gI궈�q,l颪U1��"Ϋ�,\ҩ��f� 6ͱԭ�N��2[I��c�LEP5�ͺ�m�\�Ye�u���2`��\#�ӡ�ݼ������Gs��0[\��b���=����x��۬��ڮ�Nn�ه=�7VW��@�0�:i�+�n7�
nUy�V-����%����6-��6�]'d3�!U@mm��]�ͳ�ף�̽%�7�%�B�F:�׶l��[�yF�hI7l���+��|t&N�w��!�cv6�v��:�^^A����d�+���ɗ���L��� ���M�݆�j����m�����hCZ�8������=�A_@�Q6�� ,Q�Nny����=t���%h���;[Y��ӕ��%��C���Pvˮ�0#i�;�����h�q� �H��ҽ'C�;hz�8ЕO�t��u�nM=�Z��';<j��瓦�k#g�]���tm�8=�K�e�v�*֣g�l����419�5d�Am�d��sɹ�\�^p`SK�E
��<�V�5rd��9˭�|�n�sf�7�����{�����s�
d^��9y8 U��s�r����2��*8Ȼ�����:���U��(nm��i/@g��E��o���pWj�9&��f��&�{{����Z޶hm��CQ8�8�p�=z�hW�hz٠w�S@>�T��d��L�ܙ�}_U����Қ���s�<��j"qhu�@�t���n��}V��CxW���	$C��1<��b�y���h{#�x+ �NV؊�Pܝ��'b�G4���@�t���n��}V�w[4��Q<q��$��G��Ϳٵ|4W@%�C@��_�Q���?�Z�h��/���nY$l$Wr,Ϳu����9*��������s@����xH�dMŠ��{�4��hW�hR��7�E�w�S@��Z��Z�{� �K�\>�y%۹!%��m�E\�5b	a�cY턼=�k�"�\1i'W<P"��<��E#�ƣ��~���}_U�^v���M �=Re�6H�d����>��h��@��S@��[�7�u�r���q�ǀv�s�<��Ŕ��m&�M4�o��ݞ�9ov�%�,iD)��t��yڴ��Z�j�=Ϩ�n&���2G�hs��ՠ}�)�[�����nbfX�g��38W��i�lҷ۷��R�@�Z��\�ؤQ��h4�ڃNO��w��/;V���M �l�;è�G�)�&ț�@��[��č�g��06�׀j~餅�6�	�p�<���0}ݘu&�u�<���hm����G
54����N�X��y������qa��!��;���$��'�,��hɐiɠ}_U�^v����0���uR�ޮ��\RZ�r�uaN�v2�h���.ŲjƝ��ٌGCp����5 '2&�D���~4�Jh+��ϐ{󿖁s���JE$Yh�{�4������Jhϩj&�"B�!4������Jh��/���N"%.XG.^U?�7���� ���L�z���Q\��&l�8��ދ������w�`{�z,���F&�)m�h��$aV`@5d@b�I�)�`�5D�)��������Fƈ�,���I��]�z&���Mf�)zv�m�`�fu�ֻ-��zf���\�3ɓY�6�U����nw+�oF�K�C�
HR%ڍ���RQy:���޹p���q��79�C��ui )��m����A_�����0�/�(�%U����\�Z[��:�jy ��gh�]l�mr���b#%����s&�zs�c���0�C��؉k ��wwS��jr3�E#
n�H���x;	:P���|ۚ�gP݋�:�H�X�ȱLp�/z�Ɓ�^��}V��}V����Lo$��Q��x�ݼ��l�׼������f��8K�B(ѓ$QǠ}_U�w�U�w�S@�^�@���RD��Q�@�>�@�t���^��}V���X��H�$ФZ{�4��Ϳu���u���KV���2��j^{l�u�g��U�7�*f�;�5F
�<lՈX����������<��^���_x�}��ޮ�b���,	#�/ �o�yK<U�
���p�^�r�j�i�A7=q`wmq`y^�@���xE1�(��;Ϫ�;�)�|�W�}_U�v/qIn�ӊ�$xJ�ﻜ`�o^�ߵh��hm����I%�����������v�}��F�~N��U)R�Vp�yiEٲL[��cu�^1�B�2�3/5���I��QǠ}_U�w�U�w�S@�^�@�ĕqD��Q�@�>�ff$^��y~����}V�v{�	F5"uEDLU������k�5�Suʴ��hϨ�n$�L�,��@�^�@���@�>�@�t��}�Vbq(�H��@���@�>�@�t���^���.m4�SPQ�峹�X9*�'\v���^���f���W�)��:RDG!�	��qh��h���Y�}_U�r=�j,m�x�8I��f�ԛݽ0�{� ����:�*l��w�Z��H���� ?v��>���;Ϫ�;�)�S��cP$lɐ�ɠ}_U�w�U�w�SAQOb��@�RI�����o@��J����D� '��}V��3/]�|����>���/eQ���M��m��MF�x�`} �.f����������nzn�9(kh\Q����t��}z���������1F�w	5$%� <�vgUU&��{� ���w�S@��+1H�J5$$rhW�h��hwJh^����,�c�Fb�G��}V��t���빠}Ϫ�9�51bn,S$�@��S@����>��h��h��-��%���|�Փa;G�5-Rֹ�Ij�����h<��jB��H������n2l˶�p�� |�;U�9ˠRÛg��;�\s�V�m��P�,���� ���s�v�,�*8ꗗ���yv�2�S��ѫI���e�fJ�i*�`�]�ۣm������g�.vnm��W��un�Գ��Scm��=hۓVc9�绻��{�ǻ����?�]�n�A�J;X�游p��Y�qү2�۷�C6Jb�T3���91(8�}����>��h��hwJh��&X�"�2H���}V��}V��t���빠u�X�N4�Q�@�>�@��S@����>��hg���cR' DؤZ{�4�]���������JĮH4Թp�<�w�UU�������@�t�����U	�D�Ĕ9�T���m�x���ɝ�Œ[.U.[�,�^zfbq(��$�I���Zy�Z���rU^0��ذ��gK�Z%إ�TT�X���%B���	5"��) �@��.(^�Ɓ�t���}V���q��q��$Z{�4�JhW�h��hԯP�7��F�����M�Қy�Z{�4�p�*���1Ȝ4�Jh��h��<�f�R�I*݃}e��r[r�r�=�l$v� 1�Ƅ�l�F8��7P���f�M6(8�N4�Qi��/;�h�Jh^��>����u�Q�����r<���3�%I��l� ��8�;Ϫ�ٙ�����A���bőȓ���u|Xޮ,ŭ7��<�,j��II�����E<��3I��A��x0�M��!�#�]�M�y�z��H�P�1����ec47�Į��=x���j�@P���5�h�[�f�_�^D�DJ"1�� � ш�j���F�4 ���6�����4noAJ�@�i�A)(��;� �M�H$0�4)RFh6u!��b��U�6qѰČ-l%������tT���
`!�&�_�MC�x"z��EJ�<C�Xov<Q���_<*5T��!o��<�$�Ϸ���ef)�F�d�'y�Z��4�Jh��*�Ǆl��AHh��=�)�}zS@����o�{�ߟ����a+�[�fl��ft�2u L�s��fw1�ܽw��sQ�Y��Ƣ����|[?ץ4��h��=ԯP�7$������sg������ ��L��hݟ�P$lɒD�z����Қ��4�Jh�m'Q(�4�nmq`f�q`{������_	��">����'�:Y�}��$����+j��ܶ�� ��L�ꤽ��|����=���{��M'�Ln<SKK#I�R���;Z0)���2�[�f�V?����"o�9 �dr$������>�S@�t���Қ�YX�$ځ�H�4��h��=�)�}zS@��QT�<��$a!�w�S@�t����M�*:����N���0��ǀ~�a��������/{ܺ��7$D�.��S�ۜ`�R^�����÷������2I���*(�`� "F(���)"��C���[a���]n�:#��5�˓�sk�<��6�P�����T���M[���η�a�Xk���d@]��jg��@�dX�hRT��)�v��wH�B��䢼��n	GJ�];.��]��7nF����\�b*# �K�bv �e�q�j�ų��pT����#���ܛD1r�u�4�V����å����x��ͺ�n5�,�i�hjX�W�4�|���˻^\��\��$�%�������f��۳B���y}[5���ԲA�p$c�b��w���g���K���0<T�v�oA�r��n2��پ�� �vq��ݳ����hg��I�x���J8h�\X�>k��WŇ�q���`t{ϭ[�r�M]���9Sg�����q�K���0<�{��`���+��mJ�Gp�������.�Ϗ�0���4~��r�EMY$��q�f8�=hg`����hޔ����7�t�	jJ���S ���)�Қ��4��O��UU��ӌY�\�e�iʚ&��3v��o��Kn����,t� ���L�M��.�e���܉�r�����4é��g��� ��&T8�F̘�N�e4�Jh��>�)�^�Y\XԘ�j"8h��=�)�}zS@��� �KV��h�� �+�#:��5��9�úkh!(�h�/+lEH;L�8⺓�,i��C�:���>�)�}�S@�t����W�8� X܉8h^��>�)�w�S@�t��}�V1��!��9���YM�Қ|����ͥ��mQ���`fmq`f�tS��L �4�Jh��>�)�}�S@�{�8�ŉ��Lpr�k���K>����WŁ��Ł�k�߿�߿���Z)���v&գV ��(v����-���H�s\q@�f٣U�H�p�~��}�S@�t����M ��,tB��&I���YM�Қ��4�Jh�W5&&�D@n{�4��>�)�}l����1�Ɯ1�C@�t�������mq`�oɶ�0����y�6��|�kxۉ��BƤ���mq`{���76��76��>I5����\�̪��i�9.�L�(��g�l����?�tj!ˮr�%�<Ҝ�3�'����h��;�)�}zS@���A�G�F������M�$^��{����Қ��(�S&��1��h��>�)�}zS@�t��s���	 ��6�����M�Қ{�4�Jh�	2��(�2d�8h^��;�)�w�S@����p_��$D�j�$=�̒K��N��ut;����m�;k��0ۉbA�bGrO^҇^�O��U{mΐM�Z�I�8w�����Қ����u�L�ڴ��bN��8��2A�Ukj�������mX�����OnyD��N��i6�I�e��8�&�]�Q�� �t�4]�C-Z������u�l�;e�C]/&U㛮zU�v��r)$�w�UrJ���_�]��RWVl�<���]�c�piv-�@�<ܐ�	���D���LrW����ݏ_Қ{�4�Jϐ{����_ٲ��i�wn��=���?����ߺ|`��� ���L��_��j��.�m7 �4~��}zS@�t����M�,��p�
A�8�����M�Қ{�4<�\���E���������,ͮ,�[�>���=�S@��m��ӏ����XH]v�ѽO'3��Bb��`(�%W4i�{�ܽ���I1bl����>��Ɓ��M�YNT��7ݜ`�N�$���)˷.�k�Ƶ1�y��CHc�4�6�v�6�i%;�Vo}j����9*K�*���oc,�lq݊)#�`��������I/��+�ޟ�t��5n���"�vFB���U>���8�7}�`u*����0^�,�wM[�+q�q`�{4�>J�|�}��|~��|`�������I.�.�{V�scvι19�1t�&x�k7�ji��$+��'r3�rK<�<v]�w%�M�rp�v�0?l� �����}�����5p��AY����i�*�I����8�7vi�&���Eq���]TX}�֬ͮ,��k�m$6$�"��BBj�ԕW�>�O�}�|`����YN샖)w(�
��|� �����`s���`�N�$����j8h�M�YM�w4{�4*p��H��2H�LdQc]��ݽb�):�3u�v�Ҿ�%/S2�Ѻ� �&̙$N޲���h�J~��wN0]Ѿv�r"9r�-�0��W-�2n�|X}��`{:��7z�n�Q[�+q�q`�{4�7vi�ԾW~��� ��ŀ~�Z��K�\M�r4X�\X�,��Vn�� s`@�]�m�`F,���-P�P�I=irK/նX�v:�D' ���w��i�}J����ߗ�?_��h�M˰\�n�$�#rF���V���	��F-UR�%�'G�i�7.s,	���$��m��{�4ݚ|����ߺ|`-��K"iݐr�.��=���9$�gwN0ݳ�wwr���9n��H�Gw#N]�p�;�q�y�f�r��U�]�Nŀ{��0��Y�8��RGp�������W������}� ��٦ʒ�*�W��y�|��7��\��n�n���>T�%�R���|~ﾟ��i�5��_�P�0H�@"ihx�R��a�t�%��6f��u��J�! a�h�������15O^C�7V��q��@��4�'-% z��q�Us��C�M���cˢ��x)!$��"Ej�`�����@��ܡ��X%40�`B-7��u<��!"����2!``��D �+ĀH�", p���B0 �ā� H D`s�n�M��q��EB��Xӹ]�k=�k=���x�󌐐$I�(x�Ă@"H�$Rb��1�F8 �4�%�m
u��кH�BH$!$!"�"�1�|�6:MkD#"Hj���d!������m�`�L#��$2X@&���si1��0�sa�6a9Sn"H�c!#4��` O|֭���a���ۭΚٙ#�	3�&2��
Z��t�k7=����u�v�eDp��U]F�<�[q�Z�q�l����ˎ��~��U�E��;�l�S�>�$ފw[�J\�\���)�g��������Z���Zx5�S+m�mB��N�m��$ ����vm�2W��OjRs*=f�v��4�G��v]�ۂ�@6��+)�]A�V����^L�u ��S�n��怊uڃ%�p]+[�p&`f_1��B��*Q,G3��ObE�ʩ�YE�c�5��],諥@�{�����@��*H�� 6�$�/@խ�rT�j�m�����lll Z�Z�u��˻Hf1mh�U�Y6��u;�H�Vˍ�2��ѫT�H�mq�]����.�gcX����9�2�tU���l��9*�Y3[|\������v<ͧn';�CƠcqل�!V7f�*plk��}�ui��]�PWu���Bl�)	�X�L��m;UU��~�����l��;*���7h8˭�+t9�s:]qp��k��;G�k��`MF-����'�ێ��9K��fm.M�NP�閖�WZ�qw=s°.�#�hnʨ5��^s"��6׶��kl2����6ջ\��*0���`-��[pm��ט�U�̑=GA"�ʵK��][�T��� \�V+)��яHդY�ҭV�h��~�}��إ�U��RS��ҩ��ڲu0�Mv�g�'�����9��!K<-�������lgE�@#�r/b�u�ol[)���u��c������Zr��>�>�o7�ElC�d���(�Z�65X.݉L���=�Kȩ�6j��3�F��@疗gfwNy�e;r;F���������J@�fQ�mR�R�;e��ڱW��j��l�'a�	� ��6�#5v�-�e�Ͷ�6(���c���XZN��ݼ�87.<�4��U�ԙ�b�S�	�����<�䑍\�W#�J�J�J�[Kԕv�D�p<T4�F}Q>"����4/��rs|޶k{�ֳ7Zy��'~�}��xVS��':�<j-��v���펵��g�q����ֱ��TL�c,a�)6x����Ē��=xĳ:׀��^{Ev����m̦[g��S���(����{�n���|l��l#nKl�T�gW52�2���)�Y�Z�1��S۞�7c����7g6ZC����9Z�::i\�\��pm�� w#�����s�����rO�S�IM��l�u"������mY�"����: ��\�y����k�玹rA7�o��|`�4�<��N�wwb�5��ӻD�%��rB���3�]����߻���t���Uc�G2'p�<��LwwUT��}���ӌ�e�y�'�w4{�4l������v{�H�68�fF�h�Jh̵Jhz�h��}��_��?��� ���ݨrru<\8]l.�[���[tG=	@�X+��S��CmG�)�}�)�[n��t��u�eQ%fL��޲��}I��J�X��g�Z�>ݮ,ޮ3��l���m9"n�B�� ����=�����vS@��S@������ɍ8cQ(�h�Jh�M�YL}��,_��;��\M�$.�[e4�Jh۹�w�S@���ᔴTi3��I�[@.�z��3��GJJJ�Q"�qf��K�c�9���`{���;��X�\|�ג}U�`z��~�����!2D�[n��t� �٦��gU$�j�N$��.ʨ)IS4�ޯ����5bi,I3?�E�|h[w4���I��n\0:�S��� ��8�7wq`x��� Z�U#@�lɒD�}�2��r��ץ4l����uD�a4M����ͲM��x��MY:V��qq�XNm]s�G�'p)��[}������{�4l����M�v7�Ɯ1��s4�Jhl����M�����D�D�ıG����h^��:۹�w�S@뎪��#�"p���&���o���%��fI��TQAIТ�  A����M*#�M��w��r�g�86Y�.��(K���~���o���}��~m��}�x�f�4��o}^��-X+�[�fzVK��f㌖��ێwb���u���Za�Vn����������Ξ�����m��`cm�wsO<m�}�N�K˶��w��o^��$���p��n\m���i�|�)#>��1��}��/<m��s9RWv����Ka-�R�y�m���������>��������{ݜy�i\���f)&&� 7	�$���}�I^���$�ݧ�$�zRjI+���v�5�����6����������������;gm���/<m���淲F�:���5h�9vX8+���WC�^I���u� �&-�]�/[ؠ�n�e��ts�S�DX�Vx:���@tA��e%�z��:.�g���'Xv�u`�\�fd��<�mq�N9;:K�ٌ���XK:s9�n,�pas�휩�$�����!5K�d��'�9�k�����jWu��?���?n�oH�����z�� �&Ԗ~��K*����m��=�8<NκI��뫥��܏i��3�)Df������5�X�7+��m� ���獶o�I������*J�~��of6��S�]��ԸՑ���l�f�9*J�����y�m��`cm�wsO<m��,d�A��#�Ԓ]m�>�$�]�Խ��;����/JMI%󸸤�$��xᑹ�|�W��jI.�i��$^���K�����%˕�E�+	-ˁ�����<��$�s��m�����䒽wCRI_q����$N9"s�D�e���g���k<�urj�B@�㈸kM�.��%X��9-��`��.���m������w|^x�{��R�W�}ٜy�m�NMd�]��m�@����{��/<J����P����fI��y������7٤ϩ$����7���MEn����g�$���t5$��i��$^���J�~ϾI.���l�I26������w4���7٤��{��/<m�}�灍�����\ �rՑ���l�e&�����Z����%z���>�$�ǿ��G��UefvrYz��o<�+V烘x�)md�n3ƛ�IT��}�.��p�	p�6�����o}����{��r�߭�v�&6���zq�eح\!rx�{��}�JH��}�x�g�>&6�����:����\����9D�r�e������[l���7��Ą?:V��~�@?+��9���Ӝ����d�m��r[.�K.]��|�U���cm���<����m�UU�T���|y�m���e�j�D��"�w	���w4����T�{���}ݜy�m���cm��煐x� �bi�����a]Nb��Of���D�I�i�n�ԃ��96��\�1�(�}�I^���$��O�I"���*^]����^x�{Ӱ���%ˊ]��.�cm���<�%IeI�8��o���y�mﻘ�U]�}�s�p�j���獶v�&6����y�꫻�����}ݜy�m��45����d%�co�+�����o��m��i獿�E�$3bxz�~]��>�7�����#�l���.�����w01���ךy�m���cm����6�ԕR?w�?]��'-��T9f�5�$M�V���{*^kM�ոY�.k���s}�2V)״�����o�Ϗ<m�}�Lm������ҽwCRI.�U ��a�7�M�}�L�����6�of6����y��UR�I}�ˎ�"r�"�w	������獷��`c|�����獶}��cm��"�pV���獾�����1�߽�Ǟ6پ�&6�����6߶]M�G$#x��Ԓ^�i��%ԩ����{��/<m��sm�'J�6���-SԪH%M)�""d�!��Ο
�t0��Z�"y�/:�BQ�mvd�\; �΁���ۦth���7e�PV�cy���!㛛��Iw]|ٮ��eD.h˵djtM�W�w/5�N�BR�z6M�o7�����h�!K*v^t�H6\�*-��Ns+F���*-��Y��>�/N�g<��[�U�R��Ѯ{i�q�/XN�n(���[p�l���ww������]$�-;t����+�a{L��w�m�?h7Gs��Zx������Dq�\E�;[l�m����o}���.�~�gx�m�89����d%�cm�}��y�+�}���o����l�f�RI}�T�S"�ن8A��|�W��cm�۹��>I]��8��ow��獷�~�nA�d�Kr�co�]���x�gl�cm�}��y�o��/�*�w߿6�}�,�F�r;b�.\<���i1��$�{�/ߛo��m���<���K�wo��ng������qs7vpB�m�Wi'���M�R��]�\�k������w��o}�����sO��~���8��o}��v[�+������~��&x�!>�"&�����R0T>:���s���r������~����Ϊ���;n�\��ڹrˁ�����<��٤���_%RN��y�m��c�cm�ٯZ�A��I����H�RjI.�~ϾAz���䪟������Ⅴ�d%ɀ{��,�W{��^�t� 7wf���er�S��ZF��m4s`���ܒ-�	�:YE�9��zo��o�]��p��^��<X�٦ n�Ϫ��%�K��w�b�9=�\�ے�-�s4[)��4�w4����ىw2Α�N9`�� ��� ���2l��}`����0�0���md�7��|�����+,�µ(W�a�����iU�]U0<�6^	�4 ��� �C��)$��`2$e]��|"��a�R�1M!��<6�G�e���рHHy�w�l淬��5�� D4�V��@ � �,�a 4��q�:��v�е)D��<b��(�<�A()��>D1QUجN�8�� *x!�	���@!�*�z�����}������\M)0q�d�������߾�֯ۚ�����@���˰�;��ӗ羽ŀr��{ݜx���ﻸ��*�]��F�w%��;��j:�{i�x�[�u�A�4S�<)X�Ղ��������k�9�+�Ͷ����7v`����_*�K�����X�_��dp#L�qp�7v`��� ��^��?n�3�%TٯY��(ZQ����&�݋ ��^���_RJ������~��y�M$�5wm
���9U$�n��`�N0�ݘV�UE^����ї.2����Ȱ۳L�R��x�v,�}{� �W���o��p�6��RnQ�r�OQ��bA�����ݮ��u��#^�e����_|g}Ո�������� ���X���*��u�<�w�2�Eȋ��(r`���=��,v�^ y��:����/�Q�dLN��֯ۚ�ׇ$���wL���n�wwrI.�;�܋�UJ��>���}��7ws4����-uV�(
bpmŠn��>UIR��%��}�~���,v���UN?c
V!B�
���tD�*h�W]�k��w��\+��,`3E�ztٟY��R�n!�G�W�Év�y�:����Ln$b�ءuJ�\u�tPZ��V�z΍ur�\��Ǌ�[������n�U�&�lY�V����M-�+Ů�(�	)K�[M�Hs�+!9�R���|Y�X��u��r��TvѲ��eԛg���aR����n��bʃ�1&�����z�5����1@M	2�?�W�8���[q��y�P�1��ŘrV\���u��&JsE�g~=�q�_���7r�"!�������w4]�@>�f��b�2,m�1���>���ISgu�< ��� ��ŝUI�Y���$mZ�$��Ȱ��x���:�&���`�_b��e��n���q��ݘ��,���,UI�N���������d�4��-�s@�/ݯ�^�}� 7���=�\�NKRUb����^փ�ۮ�=[Of.@�mpp�j�۳�f惥��[�%���lu��=�`���I�@ww֬����H�)iݶ�X�{�"���0!�����7rs��o ���,�Ow��v�G�:w&f��=��`n�Z���Q�}j�ϧ�x��~�\P��w��&��*�߼�㾵`z7b��J#�z��#��$��pĤ��u��>�ՠ�f���s@�jƶ ndi<RI���'�����6�M��5{uk�ۭ��AXh�}�Y�L"���仄��?u�< ����=�w%^0���, ��X�Wp�1��@/������u��=ou�R�پ�Xe�G"�wdP�r`�{�I9���2b��#�  �r�	�*��~�sz���{���I>�u���'!�5��}N�����{��'����7��.��H���'v�"�?m��$�����ذ��s@�p�$�P��7��j̗b�ўx���O)���8��� Z��%�Iz2b�_���Z}�h��hS���/�W������>g�T����Wɀ{��,�T����,޾��v`V.�$dX�Xc�(�hS���ׇU*l�w��݋ �~�F\�d��v�"�ꤓ��s��z`��j�P����i$�8޵`�� �q8� +�ǀ�ݘR[��/ �����=]�@떤�odMG"�b��Rq5���8m�<I;<��s`E�!�XNm]s��nUNIl���.ȡn����X�빠z�V�_u��u��S#�W-�q`i��ϒ���ٿ_�< �{�{��,�TټwawwrE%�q;�93@�����f��n��:�h��n�j'��p���:�7��Lw���,�U|����� ���>r�җp�qܘ����>�K��/ ����}�o$�xDE@(4(��"���6)�3�J���<�Rv�kV�A����[t����2�V��;ێ�����+l㠲�^$�铞ٙP�9�2(�=t���4�\�wZ.�;��n��H��уf��@n�)��;r�K=3q���$�ӻb�]�U����@1v��M{�5(���l�7tY�b�$^`ې��6��'����.�̶��)���k�s��m������I�E5�Tj�U���=`�n1=����-���c�ط�3c�:�V.�ef��w��>�jtv]�6�f~�~�����h�Y�w[��T~�F\�e��]�n�ou��U%�+���w}�,��n,�y���/� b�'�_���;���;Ի���h�T��H�9&A�&��ow� �x�X�ׁ��+�����z/�ƦE!�5��w�w4Wj��f��n�Q늉F'�F8��d�'=:���1�73C�SLQ�0�����7?��.��HIq[NIe����������wqR_W�~;�X�?������QD��Xf�ZM�cM�i5�T���X�7q`��^rl����#�WPw#.;� ��ŀy����7�_s��z`m��c�F�bj����>���`��< �}ف�=����xe�.�w-[�nE�~��xʩ>��x�v,�7q`�{n��rGs������9�`j%m8[��U*n��I��J7�=��.�X̸�R8�r�� �ޘu���빠z�V�ު��%#�r]�B�ɀ{��,�l���,޾��f��H�u��ƦE!�5��<�׸d�ϵ��'ሐ i�Z�[ �T��{��}�{�I=�}�o.�\�4�v܋���8���`����I��}��=�����dqӸ�n��v`R[��/ �����e4r�U��)2&܍�0mxj�� Y��:��-p�;7�n��u�����s��S�܌��O ��ŀy��ŀz�M ��hV.�$dX6b�Qŀy��ş$�UJ�߾�����=�ws@���DN2I"��%&hzS@7����Ԫ�������ŀ{��6�,���˸`rT����`�زIϽ�Xd�] 
�4�Z�"}UID�߳L���y#w.+���L��q`U/�T�����/�w�>0z٠\�g2��Q��!&F�F2
u�u΍����<1���n��NMK����2)pjL�>�^�ץ4����UU���X�܇���%��v�ŀ{��3�I}T�*�vw�L��`o�x��M�ׯ���n8��p�p���{��,>J�U$��޼X��0v�W��B�	܌��L�%T����`�z�`����J�7��0��,��`������>�^���V��V����䔡6��K%Z)��D �x$>yP�'�dRR��HŌ��(r#��lMȕ4TaxF�(��)G��H�l 4�E�����3Bat�+%�萴���	u��Gf��0a7BB$�����ļ�*"���`BLJ�4�V�$I ����B��P���AP#�b�ֶ;D�R� ��ow�^��c��!@*�M�E&�UUlp=�s`n������Q�Pn���O�b��!�.�[��*Fu��r���[��j
^Ț�9�w(��N��r.�{�Z:�%A�,���FFx�0�%�#IIų�U�KH츬Ŵ��ٲ�mm�Yx�\��(���aZW���֫5V�t��8���N�8�7Z��aMl'HX�=�pֳ�nG6�5��b�	G]	���=�9k ��0�����Zh�$MH: �\�HC�٬��6�]�Rڅls�P!j�vV�Uzv�f�"�+m��u��  v�m��ݛ6�/F����7,�P+��U�Z�  H��֐s�*e�5�A˭�u͊�m�6{a���3[6��T�6��i�$#���N��*�f�g f�gr����g�j6�cG ��Q+��Uv�;&yVcEK���{c���S�.��z�d�a������	S��g=+;�9�P5��g�0� (�d&]��8,�� �m=*���肜
���*6v��a+N&wnJܑ�Җ+g15N���̔���FH��`x��66y�h͸��ی�5���@�����z��t�lr�4v�6%H؍�٭Qt�g��%���)�E�lh���;v���iY&�TUmʼ��+*�=��"��q����XX�\�4�1�]�p�Vq㐊�q���'�rCr�GR�[���8���Ԭ�٧y��PBW���.��m5�<:G3e�I�Mt�О*�Pي��rӕ��ms���$=�d��wbc�q�[n�Ʊm���k��b$����#7�u��fz��<q��Ny4Eq�\5܏�1�����-71hހ�5J����uώ,��mm��X� 9��lm�{;jZe���
Ưl6��4l�θ�=V݉���1S�)�ק�̄����
|��0����.Rv���Iх\f��7%���v����ڎGI���3�t��"OG��W{�M"l�(q�?'`|�������x��"�H��"�Q~����v�Χs�d��
���gc����jԸ����d�DK'�]f�Np���m
V/S�S��S=@;�\�GF�`<���[�8�У@<��9���8�n���gl,Y�MFӕ�۷VW�w�Y$�h��m�6m�٢ZGt��b�_`6�����/n�۞z+�;s�e�ۖ�v�Na��{4k6��[5����]������wv�S�}��d�X2�rk�N%V��7��ꂴ[v�Z�.h�������}�	Zgvmw�m��{� o�� �}�]^0��׋ �cqqFc�'�^�hz�h^��ߺ�=ߟ���"�wdP�r`�}� �}�ŀ{�� �wf�����wr;�wp�"�����ŀo^���v`u'����7��c�$rI#�6�s4������]�����m�����&됙�Nڒx�f쯪�l::E��|�w���un�x�O*���o��Cq�Nˎ������{��,��o���Z^�Q��<�'&���}�G���@
���4��C&���?u�< �wf���֤�4�Ю
]ŀy����=��xrM��� ��ŀj�ёې��Ł��R{ӹ�ot�=��X$�v�����0댲�+�ǀ���9R[��/ ��׋ �ou����n�\eݚ��"��.�ꋫ��ě��=`KS��0Szn���Gk�v����o����,��o����%_U~�>ﾘڻ�ۻ���Yˋ �}{�>J��6o_s���`��,��l�;��ԑ�$�;www�}� 7���UeU%��V$� I��T4��I�`���D�Z�=�S�`n޽�Q��-�e�wp��I���`߿nh^�����*�H0���\w&����9*���/��ot� /��,�'�F4���jB��S�NŔ�<	4n�f�tU*���G7)u��ȱ'�c�F�h^�����볒�^0��ŀr~���q�,.�ǀ{���I$�w�� ��ŀy��ן%J�;�Xî2�$�9#������,;�IR�����>�����n�["C�"l&A�&�m��ף�d�}���#�Q� �R��>���&ܪ!�v#� z!�R�������0�}��V�\��B��9�ף�@�ڴ�٠[n��IU/ڻ��I��r�"��E�z[��9էr�Y'-/+�t�R��[���}�����o�F�8�4�n/��?��h��@�����ŠuuV�(%#_�m8�}ݙ�UT�UIR�>��`����]�@��j$q0��"D�ɠ[n,��lxuUR�����ot�<��:�6�ᑹ����k�h��0:�T�v�� ����ㄉ8�q���h�f�o]� ��u`[p�~M&��{�HUT�DUv���m���ӝ±�0��� y��'�H]h�N@�k�ݰ��	�즊�vIё2�M��YH�:}K����V0j��u4�6�QO�[��s�ah+���.�ų�gkm�8�3��W#�%Ӟ�d(�G�m���pVU4s����Xv���6��.�Wm{nǭ���;�m�i�yg* ����՞���[����������X����_�bʚU5Zj�s��KS��c�:ƫ��nM�/�2�1/M�a9���1�m�����`ﻋ <�v��I*_%U�þ�����Z�m�Dܻ"��ɀ{��,��UM��޹�o^���vgRJ��R�>��b���Q�"dMI�����4����$z� ��s@����m�b1!�J��g��������7׳ ��V�(%#_�M8��٠~������> ��M��[�&$ӭ$祩�2�5�ɳ���n&w"R��=sZ�n���2DH���G�!���:�����f�ߺ�I$�������{��w�K#Eؚ�(�, �}{3UR�+�e�� <��0w�ş*�UU��{�6��p�;��r`��� 7���=�w }yY�Z�+�cq��8�Z��ϩ$����� ��X���`����h�$���LcNM޻�����^�W���;�h��@�Twq�$R�#W]�˺+ud;x�9+�4�¨]�*�s�u�sE˚&t%w�m����0��^ o���UIxû{�wQ��ܹ�v�ݹ0��^}T��ý�v�, �}{3�J��$������r[��r��x����7}�X}T�A#*U���\P,����I9淞���Ip�B	l�ܘUU$�v�� ?v���������~�l�rYWb�pQ�X���`*��]�y���Lw�ŀo��[��w�w�U/Dʽ�wLv�s�m;��V厙˻z�Fl'����=S�$��ߟ����lo�ـn���*UT�`~�}0��0댲�]ڹ#��{�>��I��{ {��`�����$�g��[2パD�Sԓ@�����^Vh��@/����uF4�QI"dMI��3�*M���`׼�n����HJ��ٟ�+���/����̐��6Ԛ��� �|��%o�O�}�}� <�^�҆(�5X��N8�K"jF�\7lv����T��r� 9g.��3�%�d�H��bj,�����V����&��׼�{��-6�2Z�R;� �޵`펫�w��;;��I���Uv{���9,�bjࣸ�߹�0��^6w�� ��ŀj���w-�RK.[����%O�o< �{�������*M��}0�q;n�r;� 7���9UU*������� {�?���{��'��Di �M};��j.!�:HxL[Z3�D�nm�k�D+��Y��O]�����kdPbi�ƨܬ!l����
G-
�㱻]x�qhl���$���Y,�{u��gD��
��.V��݅3���u�ժ]pYpS������@U͠z]3R���NJ�,���J=���{!�i��γD<�!�yԩT�]ZF�3ʽ����YN��ȷ!�oa����w�{���|
��&��]C֌���ظ�1��9�N���3�ں�#;r��,W@��F��o���, �}{0��_�W���`���,�n8��mGnE�o�f|�gu�< �{����ϩSf�܁�%�p��6Ԛ���Z}l�-빠^VhyrePQ���c���_[4�w y������� ���d����	�)&�o]� ���k���@���H��1��Ġ�2
�ɏU��m��m� �+\�j��{�|������"s> ������h�f�o]���T�G&I�Q�o$�}�~����R�_TD6<����y0ݽ� <�v�|�*�M���d��܊9ǀ�� ��qa�U$����u�<���.89i�1�94z�hު���h������R����v��%۷n89#jݹ y����J�t�~ w�� ��qh.Q4�"�,�R8��"!�5�L=ga�k4;�2�ѕ�\?~��ѝ�����}�_�$����jݹ?���< ����7}�_�T�`~��L��]���˺,W.�ǀ�ݙ�*�l��ŀ�_Lv�ՠU�j$ia�P�"rh��Г�{~�O@�SPd�m�D��%#Ye	e%H�et��d
�b ��;�22������6$�Kn�%B�
@�,HE���������@h@��/�M)��.�j����R��.����i���bHq63Z�8�p`P ��A��m4D4`͗���GF��M2����0��<������)�j0�Hlb;��N���N��$�������"F�,���v>Q�08��54"p��!Y@4���)�6��Xy��O��#PC #�!��@�D�Q�x�����Q� 4��4����L�ŀn�U���UB&D��Gq`|��T��߹�0������h���./uK$$$�#j5&��~��>J�|�%�߾��}�}� <�]���ZikrE$��cx��+�z�Ԭ���R�,���v�v�[�۞�Gl1��HӄR'�W�z�w4���ٔ��׼�}���ȣwn+��^o]� ��@��Z^�����ċ�lM6�PRD���� ��M��hzנ[�s@�[���F�p���&U*}�y���w�Ł�W�?��.�
	���f��� |U�2Ƥ���N-�Z�}�X���`����RIwsO�"6��ZY�ۨ������Re� gWlY-ѻ!�xm�u�R������w���i]k�q�����s@>���-}V�W�z�c^�##V�
;� <�^�ꪦ���x?{� ��qg�M���HH�]��r���������䪛��Š�9�u���5c�R'��*T������X���0>IU>��w�����6���q����?͵�}5�>�{�:7�lI:z�$�;���Uךv���PG=i���e�s�uҰ��k\j6-�u�v��QF{Ǝ�J��8	��yM� (ĸ���O�Z��<�l�u����`ru����yzX����n����,OS��Z�(;	R��ۈm6�x����3�e���Ct�F��,R�pch�>��J�J��Xm��:�sq�g��S���^W����޹���t�܇&ַ�'8qg)yhɦ���œ7zR��L1�gw����O}�С�rT
ݹ����v�׀k�v�������?~�ZH�r8�E���k����zՀ{�����I���M9����ϥ�%�W.�ǀw�Lw�Ňԓg�޹�w^��5�[��[d 쑗Ɂ�IRO�{ŀ�z���Zz٠}�Yőf<pȜX���0IUUR�����n��w�m���~ߒ��L������@C��vF�ު�`�U�֔�����Z�Qěj8�k�
�נ[�s���߯�4�/�B�EmE�ŠU��f���ꭄ 
�W��%Y�M�X��\�7}�`~ݵ�r�.��n����, �}ۘu$��o�g=������ۅ��HڶMR�v�Ձ۵Łѽ�a�M�o���7��o��w.Zq���0�٦�%׽���v, �}ۘ��]ܒ7\��*m��y�=�����Y�@����⹝ȕ����`GRQ>̫o�{�x��ŀo�s��*^0����v~��1�B6�Lq8��w4��s �}�`�ݼ�I���֝"p�*h�*��3��j�����*b�M������= ���^�,NbI�Իr���T�w8�9�u��ݘ�*J��z��-�c�9qId��w�{�����>���}�MX�\Xw���/�sWS+D,�`���@��ppmk���9��۩�u'��w�=��Ѝ�����߿~�����Қ]k�;��bm(L���	ɠ}z�3�Tٻ����^ o�ٟRI&�㺛�.��˖�ww$0ݜ`�ݼ>I&���`�{!������r\��c�������@���h{���(&+0���<F����x�.�H��F�5#�0n��I/ݽ�<�g����;w��ع夭k�m]:�Yz��l�͹6q���{*�&�.���n��5W�ϻ������;{��_�������>{�6��;w�Gr��������7;�K��i�2|��6�ƛi����~Z�� �����>�@���[���M�LN- �۳ ���Y�o��I$���x��퉴�"qı�94���������ՁM�$׷Ar�R��<ܻt���ɰ�dv���[sZ{"�WX�2�ym���=�k�sÖjv���v6�6�TH�n���F��ږ�ӝ�j�uv�b�'V�r8�jк�e�3Jdy^l��Е>�ˉ۝�읭u��r�a,t��B[�HA�C��q�AY$m�:"m%��U&m}�D�ѝ���vmTKk�)^֞��#nc����qƷn�]�|<Z���trK�t�OFhv�XF���*�I�X0-%���j��p̦�˸��Zq�$��;���]�@��s@�[��
w:� �qM8��ՠw���;��4m��:�%M��[�$M�ƀe�x�݋ ���Y�ԒM�׼���x�jS���f�L.�7��'Q?
��~��X�}��=��x��i�k�귶�n5Q����Vנw���޵nhּN�0�� �F�c=p�=%�;B�.�.zƫ����z����{�����I�R5�ڒ'��*����;�S@�Z�4W�h[^k���P��][��$�������x>)�tD�'~�-�󿖁�����6���ˍ�e�0n�X�u��UU&��u��N0tݬ�#�n�ȜrH��䪾J��~�������=��L�ۯ ^\�d�ܑM8�Vנ�W�*�߼��o�<X��i�y逸,U�@���u��D9.���wW���9�&��Ĥ�+�mH��j�7m[��3�۽e4��s@��M���V�,�26Z�N���^,ꪤ��l�@����@�YM�v5[��&�J51J�������鲒z��N���H ��CH��U��UrI%�*����w��ŀo���r[�ݹ#�w�*{}�x�Ӎ�]F��YM�kŲ)���+�ܼ��`�R��R�������@�mz����)#jI��1�ګud;r���pAV� �a����.{.�njM�&(H�X��4�u�e4^��U%K��ӌx�X]��܊Zqː� ��f��l��׀{�N0w��g*�l�|Ԉ�\���n�����a򪤛�w���zq�o�6�$Ƒ�!�&�z�e4��$�Ϸ��>?,�(B�d���� ?�����d��ڷ�;��r˦b�C@��4z�hu�@�����r�\xI1���ܒ,�������.x��[���!E� z�F�/i�gf[cL��U1J��������3:����%��y��;M�c�ܸ����p�*�^��YM����=�)��331#���FȜn&
9�$��;�OƁ}�nh���*�^��wJ�I�H��j컆�J��w�� �ޜ`���*O�{8�7�����H�n�K4z�h��@����}�Y�fp���H�b Њ�\Qkd�� �#
'�1By��4;�h�� ���I��L���
|A�&��x	�$�u��������}��"�j�M��'��HH�&Y(n��+�Rꋮy��HHm�k>v+�B�$�����TW�#4�
`�'�V$@@ַ���{��a������ܳL���j���[&�	9iH[�\[��Su�9$dr�q��A<h�T�9r2h�jT����A�k@vDьx���]._F�����*�]\�$bv4�҉=,죌��c4.��2��(mM<�闗k��X��!K����b �Tk���.֜��(�]�')�4����k�=�+��jΈ<g��=1��G\u��1{k�O�A���[G&�b�s��c��;n�c<�f^n��Ct��e��f49�ȻO!d�qk֋����iY��U\�l��� �K%�r�Acd�]@B�����m���M��z2������IjP�]6m� 6�m���w\QN����iiK�VIs��hN��G �!dM	j�Ҏ9ʹ��^��������t�k�ڮz��OeюN8��<q�Í�r�Z�ֺ�7Y{�֜�ʹ'�q��'�9��oj��t�9䔃�.j���ݍ=���GI���	s,��U*��΍���W��`�p(c��ݱ�X�����gv��n��ui�;p�$�D����-cWV�8��#sź�-�N4��t쪪��۴chͥa!5�n��.��V��I�����&:.x�YuUH@���u���	�Y%��Y\�J&�	�y����6-�vqau��H*8]�����[�t�e��$;g[)�5�����^��e���
[61UK̭R��#lb�H҆�CA��:��,Rq�m�\O �:�,,��V�*g���9΅�l�t.;qώts�`�=�<u��ʜqڷ�q�9��KF��α���gn�u\˙܎q��ӻy��;�aQR,���v�J�J�Rq�.mZMSmv5�� ��c\�x�n�R&5F��cW�@HhϤL����$�F���2��sщne7k��������p�L{^�z݌F�����G�My�JĚ�4Z�Mw)�(,�W&&	Ex�V�&���{�=@�x ��Fn?"z)�8) ����J��4
��B+��x$�ڷ�bi*���3SSU$�Q34�U�d3�:q=	�Qɵ�70����!h��yC�g�]���c�η&�hLܬ�I��K-��tK@�eM����Yqn�X�k�h2�ʲ�T��鍝)m�i$�ȓ;x�Nkԅ�v��NG��ӣ[Y��4�QJt��+s�E�����)ga+[\��6h���t���ƹ��
vJw��Ac2nM�l�L;�.�.���u�&7M��DZ�\�MED��$�Q����ܽ���ʧdg&�r�\Y�sI��L$�I�,�&��{��@�����׋��T�����}�}�D��`9�b�@����}�nh�h���M����D���pD��?u��4z�h��@����W�m\��.6���>~����}� ��f�R������;M�c��qK�$v܏ �ou�{�g��<X�׺������ݿy7񀚖�d�[�u�2��Ƹ��d4�&��n�t7dlWJ�����7�3q<Q��������/���޲�R�K�����vs�n�r\�������O���(�*��P6w<Ϸ��?{{� ��f��%M��r��AȤQ&♠w~���h���/�����VI�BG?��$�4�ՠ~��L{�U$��������Ek ���=�)�_u[��e4}ݘԩu��RZ���rⶥ�Yɧnz�M�������۶� ���9a��XU���y������"$��>����?o�M �l�;�S@�݃�c�d�R	���Jh�f�޲��U���&��{�$���$w.��� �Ϸ�ɞ+�|R��4B��B�*�HD�n����>�d���4�kFȜn&�d�4���+߳���x�����$�T��ﾘ�z|�۸9%��Բ�X��^,9��������Kı;�s��,K�����'"X�%�Ӥ�wW��-ݺ��E1��k�Yz���4;��{J��+e�[W3�����}�3%u,]�����K���gf'"X�%�߻����bX�'���0?
Ț�bX�����)xRe&Re/����N�"�����bX�'~�vbr��&�X������bX�'�����Kı=��ىȭ�bX��s��oe��ka.�19ı,O��xbr%�bX������c���j'߻��'"X�%�������Kı<�}���m�.�Hod޶br%�bX������bX�'��;19ı,N�����K�� �*��� �"o�s��I��I���t/�W"n�9n,ND�,K������bX�'~�vbr%�bX�{����Kı;�ݼ2��&Re&R��5�e��H�HIq6��b6��ԭtI���[)`6kn-㨌\7nz�y��M��)6�����{��7����;19ı,O}�xbr%�bX�����Ȗ%�b{�s��,K���u�.K��;NZ���<��I��I�{�{��,K��v���Kı=��ىȖ%�bw����? D
����K���w ܒ]�Բ�YK�,K���^��bX�'��;19��CQ5�w����Kı>��YK)2�)o���%܊G�n���Kı=�}���Kı;��ۉȖ%�b{�{��,K�DQ=����'"X�%��]��{����r5�w��ND�,KϷ��ND�,K�1��߼1<�bX�'�v��Ȗ%�b{��ۉȖ%�bq?i!%E!T��}�����Ir����Y�v�V�R^?��|e�R�/mp��jɷW�7n�	q��)�(�%D�宕#Y�&�@�t����;uq�u��ɭ��C�dF��N��bKbRwyN9œ�K�n.2�G=�[tb�C۝L����%2/�M�A��ю��m
�[GNU����[v�[��;t�؋�l+��V<�C��Eu��v�sVm�N��ۮt�v����dZl�;^�O>h�	���9(�9�n8��c ����(�ZA�Em0.(&������L��_}��,ND�,K�~�ىȖ%�b{��ۊ�"X�%����n'"X�%�����M8�D�*�TҶ�5P5Y�ىȖ%�b{��ۉȖ%�by��ۉȖ%�b{�s��?����R����m\������e/
L��N'�o��Ȗ%�by��ۉȖ*X�'��;19ı,O=��f'"X�Re/yox���r��R��LKϷ��ND�,K�{����bX�'��s��,K�w��ND��)2���~[�.K�Ӗ��]�)xRq,K�{����bX�'��s��,K����f'"X�%�����NDe&Re/��|w�Q�;�
Gr�cʧ]7ZꇰZv�]C�ؽq�鍆�hc*������\q�Բ�R�Re&Re/w�|br%�bX������Kı<��ق'"X�%����ND�,K�����r܊G��K)2�){�gf'!� ;�O>TШ��O"X�����Kı=�����Kı<�띘��bX�'u�ڇw-��(�7.K)2�)~���D�,K�{����b�bX�{���ND�,K�w��ND�,K�N�/�m0.(';�)xRe&Re/}����Kı<�띘��bX�'�ｸ��bX�'�o����bX�'��:T��.ƤD��^�I��K��\���KİT=�}���Kı<�}���Kı=��ىȖ%�w������~�᪙9��rу6 !�Q��S�Ӻ�jM�jj\�K�N���ك�䷸K�[��ND�,K�w��ND�,KϷ��ND�,K�{����bX�'��s��,K�����f���k{�ֵn�q9ı,O>�{q9[ı=��ىȖ%�by��;19ı,O}�{q9ı,O~�u�w��;��Z�A�yK)2�){�gK�,K��߮vbr%��m@:����x ���qT��%��7����bX�'~�vbr%�bX�}�[�kr8��n+R˸e/
L�ĩ$�_�����Kı=�}���Kı<��ىȖ%�b{�s��,K��{;^;���#��re/
L��L�ﳹ�r%�bX�}����Kı=��ىȖ%�by�׼��Kı>�^�M�!3
�X6o]��E����"]���V'ng�1��XW��w�����Hm�f�m��'�,K�������Kı=��ىȖ%�by�׼��Kı<�{�br%�bX�zw�k��d�ٸ]��ks�,K��ﳳ��A�$O=��i�I����!"�'=ݔ���UK�J�L��8�(\VF������'"X�%��ݿ��Ȗ%�by�����Kı<��ىȖ%�e-��2��&Re&R��B��$R\�4Kw�ND�,��T5����X��bX�'����'"X�%���gf'"X�D����������^�I��K�[�1�$n)qܰ޷�ND�,Kϻ����bX�'�}����bX�'��s��,K�����&Re&R�Zn�Er����i�m7h��gY1��Wk�[�VB�Y������g�h�rG]Ym������,O��;19ı,O=��f'"X�%�����,K����f'"X���^�c}w$q˹dV��p�^�Jı<�띘��bX�'��{�ND�,Kϻ����bX�'�}�������L���/e�.�R2Y�)xR�,K�w��'"X�%�����ND�,K���ND�,K�~�ىȦRe&R�ݱt�q˸
)IyK�,K����f'"X�%���gf'"X�%��\���K���]�u��)2�)2��Ws/�m0�d�"��Kı>�����Kı<�띘��bX�'��{�ND�,Kϻ�,��I��I������I���p�v�R`6��������
�d���k(�z������ݻrY<�髜�c��n3��tI���@p�{I��z�y�z�8��v㝭[��Ó����y��DD�Fp�dŹ�m� �̸od2\����?o�x	 h�H�
��e&V��S��. �� Y���k�Cu���F��}�dJs��vwV�����B��W]6M�ww>�s���w���9���5LZ��WEN.\a���@�G[��;N:�Ux����U*&���!U"��kF�j�k;�?LND�,K�w��'"X�%�����Ț�bX��s���K��K��V��RHK�"Z�e/
L�ı/��w�Ȗ%�by�{��,K��ﳳ�,K��߮vbr%��I���;�RF�ܴK�)xRbX�'�w�19ı,O��;19��]D�O~����,Kľ��锼)2�)2���o˒˗$d�����ND�,K���ND�,K�~�ىȖ%�by�����Kı<��Ŕ�)2�)2���7�Kd��Ȯ\ַ19ı,O=��f'"X�%��Q���~��O"X�%��~�Ȗ%�b}��ىȖ%�by�ܺ-��a�2뭗v�v��r"�3����2�Ҳ��-C�y��d��#2WQ�Co��Ȗ%�by�����Kı<���Ȗ%�b}��ىȖ%�by��;1<)2�)2�^���]�QHK�9ı,O>�xbr6�=$O�!X$%�b�@A:!�P8�*�'�,M{��br%�bX�}۝���bX�%���9�&�j%����~![dd�8B�YK)2�)w{��'"X�%��\���K�D�K��߷�Ȗ%�b{�߸br%�b2���ָ���X�ڑC)xRe&P�by��;19ı,K�{��r%�bX�}����Kı>�����K)2�)u������rX���)xRq,K���x��bX�'�w�19ı,O��;19ı,O=��f'"�oq����������`MRnc7eô��m�*�i�N�(�c��J2<�C��w{�֙c�Hܖ�m�R��L��_���'"X�%��~��ND�,K�~�ىȖ%�b}��ۉȖ%�b{�zߗ%�.B@Q]�"�^�I��K��;19ı,O=��f'"X�%����n'"X�%����N@D�,JR���%����%�ᔼ)2�)X�{���ND�,K�w��ND��o����"�J��F�`{��b�o�t�Ѡ�H15�f���ʎ�15��l��-�Ox�D5 �P�U�sTCet� �tB
�p�֔� Mh�acc!6�Ȱ�NJ��L�ۈA ��9�"i
Ut1� �St!:������Y]Jh5"h��Fl&�Br��������+/�����m2%eaP��t]7e�Mo�]�T�&1kd$!��M[#<S��Ah����j|
���4�Q ؁�z	��� �*���~
b �D��ؙ��919ı,O��vbxRe&Re.�9xݻ�-�$L�Gp��Kı;��ۉȖ%�by�{��,K���gf'"X� �'��s���I��I��f؟D�phV�[{���Kı<��ىȖ%�bwﳳ�,K��߮vbr%�bX��}���Kı?(���֮��~��od2 z��.��k\S�X��x�wg����i��ԍ��f��ms�e����oq���?w��br%�bX�{���ND�,K�ｸ��'�5ı=���19)2�)2���7u����n��C)x%�bX��~��'!�R:���'�����Kı=���19ı,N��q��)2�)2�_���ڒA�b$����9ı,N����r%�bX�}����KlK�}����bX�%�K)2�){�w�9�9n]�{���bY�`j'�����,K�����Ȗ%�b_=��x��bX0BlB*������O=)}~���^�I��K�}���Y.�.٭Mks�,K���gf'"X�%��k߻oȖ%�b~��\ND���������@�o�?T��),BVϱvV:6@V���l"�Ln|q�L6����b���BN�}��D�,K��׻��Kı;��ۉȖ%�by�s��,K���gf'�&Re&R�㗍۹pr8� �㘜�bX�'}�{q9�,K�w;19ı,N��vbr%�bX����S�?
��j%��ﺇ�m���!�[ջ���Kı?w�~���bX�'~�;19���MD��sS�,K����~���bX�'};�5��M��&�浹�Ȗ%�X������Kı;���'"X�%��w��ND�,K�w;19ı,N�[���f�$UU׆�j�k��%��İ��G������%�bX���?LND�,K�}����bX�'���DH�S< �cA�% !	0@<�!Ӓ]�z�˽���s@nU���nK�1�s�OYã�8H-B^݄�e���ɷ/8��h��l"�K�^��Mq��;q�m��-c���a�(�oI�J]c[b�Wn6����������\�����ї�2jx�YS��*�mm��[$�g��x���Ϯ�󘍵ӎ9A�Ω���j�岳�]�,�ٶyG�n�ܬ��+?{��{�Ͻ�߾�}���,f��t�/:)#�5�[vΧK��tF��%�0��U+��uD���vWtj�;�����{��"~��\ND�,K�w;19ı,N��vb<�bX�'}�����K�2���� H]�-�m��&Re'~�vbr%�bX������Kı;���'"X�%��w��ND�,��_�޷��w!pWd�e/
L��X������Kı;���'"X�bw����,K����ND�L��]݀��Ӹ���dV�K���D��y��Ȗ%�b~��\ND�,K�w�19ı,N��vb�)2�)2�w�n�˃�Ɯn�K19ı,N����r%�bX=���Ȗ%�bwﳳ�,K��v�e/
L��L��o1_�2Ӗ2��������u���Bv*!��*bp�	-�\Y����D��Erۑ�/
L��L����Ȗ%�bwﳳ�,K��v���O"j%�b~��\ND�,S)}��~![aƈB�YK)1,N��vbr�0W��D�K^����,K�����,K����ND�,K�����a�����M�s�,K��v���Kı;��ۉȖ?���j'�����,K�����Ȗ%�bw^�i�H��d��R��L��$R�?}��\ND�,K�~�Ȗ%�bw_}�br%�bX������bX�������qKr�r<��I��I����ND�,K�����,K��v���Kı;��ۉȖ%�ow�����@�0P�,񁶗u ��=�����'�f0�ۢu�":c�.vﻣ5�hʨ�Jd��mxj�j������D�,N��oND�,K�ｸ�Y�MD�,O����'"X�%����#��l��wrȝܼ��I��I���������Q5����~���bX�'�����,Kľ����?05�L���/��pwi���)xRbX�'~����,K����ND���N�p:L<��K�߹�ND�,K���xbr%�bX�w��Cz�	#B�rۑ�/
L�ϨJ�_w�~YKȖ%�b_�w��9ı,N��oND�,K�w��ND�,K����nB\�!�e/
L��L����r%�bX=�����bX�'�ｸ��bX�'~�xbr%�bX��C�w����kg���������k��8���zs�Ʋqr{u�\h��*�0s������w��<�bX�'�����Kı>�}���Kı;�{��,K����2��&Re&R��x�2\E݊Y�˫��,K�������$D�K�~�Ȗ%�b_�w��9ı,N��oND�,K�}{�K��{�[��ޭ����Kı;�{��,K���gf'"X�%��~��Ȗ%�b}��ۉȖ%�bx{�u�kzޤ��
+��YK)3����w���bX�'�����Kı>�}���K��S����`� 	X��t�B�	!�J' v��ȗ����,S)2�{عڎ�q\v��p�^��%��~��Ȗ%�a��������%�bX����ND�,K�������I��K�!����we�G$�ŜNM��e�r"5���b�gW����nX�C�r��8�#�^R�Re&Re'�����Kı;�{��,K���gf'"X�%��~��Ȗ%�b}��Y�%���ܓ)xRe&Re.����bX�'��;19ı,N��oND�,K��{�ND�,K��̿�w!#RIR��L��^��ىȖ%�bw�xbr%������{�����Kı?w��br%�JL���݂뉑ӵr"He/
L��X������bX�%���x��bX�'~��19ı,O{�vbr%��L�׻ı���Q��YK(�,O��vbr%�bX~����'�,K���s���Kı;�ݼ19ı,Ms�#,'�O�O���.�l	���-$�avm�αN�עnJ3�I����km�Sk�΋s�6�LaF�s�*
^�'v�1�Яe=���n:G�<H�L��(��bh�cO�EAOO.w5�b�Y�7n,��*2"��vQ��� L��b�L�Uٴ��yk�Y�^2v�ܱ��W6N9Wm	��.s�0� j�M���\��vl͕\ݏE��g��_��}����5�����+��n�-�Y`���)�����F-��P��8�Ն��&ߞ���7���ￜ19ı,O{�vbr%�bX������D�K��߳��^�I��K����v�H��$X��bX�'��;19ı,N��oND�,K�{����bX�'~��YK)2�)wvp�G%�w.�d���'"X�%�߾��Ȗ%�b}�s��,K��w�'"X�%��~�2��&Re&R�w���.���owf'"X�%�����ND�,K�����bX�'��;19ı,N�y����&Re&Rޝ�)"	#�˻��'"X�%��~�ND�,K������bX�'{�oND�,K}��)xRe&Re.�o���Ȥr�m�8�{!,���Tt�X��qZeQ�Vܺ�3@<�nݒ�OVb��w�{��7���{�vbr%�bX����\ND�,K�{����bX�'}��19ı,W_kv�&GN�ȉ!��)2�)2����'!��ۑ2%��;�br%�bX���xbr%�bX�����xR�RV�YI�����X�q�����r%�bX����br%�bX������K �,O{�vbr%�bX���[�^�I��K�_yc��e����r%�g��~���19ı,O�w?LND�,K��;��Ȗ%�b���2��&Re&R��o_��ܒ�(������Kı=��ىȖ%�bw�guq9ı,O��y�Ȗ%�bw߻��,K��/��sW�ٺoz��8��odv�b;:�T�ޔ�.c[�X���Q/��=��F�6���oq��%���s��'"X�%����19ı,N��x`q6	"{߻��$�w��<NZ�wb��ܷ��*AK�۱2'bX�'}��19ı,O{�vbr%�bX����\NE�,K��Ф��8���rL��I��I����'"X�%��~��ND��!�R*�F@U<x��ș߳����bX�'{�vbr%�bX���l���.9R��L��^��K�,K��~���r%�bX�{����K���5����Ȗ%�e/��n�}q24�W-C)xRe&Rq;߳����bX������1<�bX�'���'"X�%��~��ND�.��v��Q����櫷����S��W;"N���\2eb�Y�{7�r�Ft��7f�.���Ȗ%�b}�s��,K��w�'"X�%��~��ND�,K��;��Ȗ%�bw�y�w�u0MQ%LEM׆�j�k�Ｍ�	ؖ%��~��ND�,K��;��Ȗ%�b}�s��?���b{����;wr��v(��e/
L��L��v|br%�bX����\ND�,K�{����bX�'}��19ı,N����Gr㻒�d��2��&Re&R���\ND�,K�{����bX�'}�;19İ?(x
Ŋ����">#����5��<���bX�R�����\P��ܷ��)2�)8�{����Kı;���Ȗ%�b{߳��,K��~���r%�b�������KvBf��Z�yzQ�-�&�"�D�V�Հ+t�wM�"$ѭ��[���bX�'}��19ı,O{�vbr%�bX����\ND�,K�{����bX�'};�5�V�[������br%�bX������Kı;߳����bX�'��;19ı,N��xbr%�bX�׽�R��7K�5�{���Kı;߳����bX�'��;19ı,O=�;19ı,O{�vbr%�bX�k��57�D̊��"�b���@�v�׆X�%��gf'"X�%��~��ND�,K������Kı=�ӼԻڪ�&���"��k�P5P5�]�[^ı,O{�vbr%�bX�w��'"X�%�����ND�,K��Q�(j9f�F+�w��u�1�2��h
�j��]11|J� E�=�m 0�4�R��d.qe4l��?
�(W{�"��n��MSAo�'� �}�9���3E���kȐ HH�JB��@��Ml����$C�7DH�E�A� 6@�A�����LB2ԁ	HU�`h�$+!4��!L.�bx�G�Å
�0�jcu�JWJ�@��"�Ig��n��FIr�MS`m)'�Vצ�E9���:G!���1�8�������M�.j�q��N�\BgLRʰMNI@�i(��͖�l�B���»�d���8���\���8�;nJfcc�Ɨ�vU���]<��îk^���A�J����)T��:�bj��l/��Kss�뫨;ss�-O���`ڝ�5�=�Qg�;#r�j8�.�H[��,7;0X����!N$��6�6Ӳ�n�#S8l��մ��yB�঺��y��sI깴9"dk�f#v��d&8�䁷��USkh���u�j$A��e��T����UjU�Y]5k �l6�Em��J�s�8�j��.��n��M���t�wLuS�����h��ۈ�
�7�����.tl�uVܓ���g\��s���{���w��p�t,mƐ�quru����{ s�!��NL6W�<�����9y��\U���]X���P�(���dK�� �F�-� ��C<�Sm��4��ƻ,��h��P�d�pl���$�E�<m�#��&v�ëQָ�6�s��ؙ��#.v�݄��ӳ��n��s׭��C��q/��RKf�-�X�ۧE��$lԤ[!�˭�8:X��a�R�m�m�6�(�d�j�V�<�7.�]#[�ةJ�搥j*�M�Bn���m�D�֚�U2e6���s�Ɔ�S��8�VV��h�
�l+A���lf��C9鬳�$�Gl��R��l�+�}����WD�pc.8��݊'�9��g��<���v�a1�M�mA��0a�t�%�_K�sۄ�׷���*�8�.�q�{�#�-96y���mHJ�%� n����\. ��&����f��WW@)���7mt��÷Y�.T6�>�US?Y]�K%n�qܮ�n.

Nu;�q�r�^!R6ڊ76M��vܹէ[n�e��lG9�-��uPR���WO5!��S5�]�ַ����A�1@4*B(qF�E ����h%_t��	�t��x�x�R�z����EMTI*)HE7l��Ɛn�4�C�MN��M��u�Ga��ƸN.)���-=V����%��S��`�X5@�����n�M��[�G!�`oc�c�a��}|�l�iյ�Yݻ+��#�Z�^�n�on����wH�H
�*�v[�W4ҵ���� ���87n�^A^v��vR�[J��]̖����۰��ƅ�|��������7;�.������bq��M%�s9��z�zݦs�mز����N����˗%آ�;����&Re&R���2�"X�%��~���r%�bX�{����Kı<�����Kı;��n�K�q��n2X�K)2�)~�η�Ȗ%�b}�s��,K��߳��,K���gf'"U5�������R\-�%�w-�/
L��L���?LND�,K�~��ND�����Q5�����,K���s��'"YI��KzwX��$�E%�p�^�K��߳��,K���gf'"X�%��~���r%�bX�{����FRe&R�Ws��F�ツ.ᔼ(�,K������bX��B>��?j�yı,N��?LND�,K�~�2��&Re&R��n۾v��i˒���n��ӓ:6昖|Z��
<LAnfy�2�Jkn��2Kڭ�������ow��;��Ȗ%�b}�s��,K��߳��,K���gf'"X�%��}��VK���FH9-�/
L��LO��vbr
18`J��:"dK>�rbr%�bX���ىȖ%�by߳�����@�MD�>�����Ke�+�n\2��&Re&R�{>���bX�'��;19ı,O;�wW�,K����f'"X�%��o_��ܹr]�+��2��&Re&R��;19ı,O;�wW�,K����f'"X��f�{�y�br%�bR��}�;�]ˎ�Kq��p�^�I��O;�wW�,K����f'"X�%��gf'"X�%��~��ND�,x������v��l6)c8 ����v]��3��.٥���cS%��g��.��������q9ı,O��vbr%�bX�{�vbr%�bX������Kı<���\ND�,K�ｚ���n7E%�p�^�I��K��y�/��&�X�~�~���bX�'����q9ı,O��vbr'�U5���������˃�.ᔼ)2�)2������Kı<���\ND�擠��TJ����P����H�D��g�Ȗ%�by�����Kı/�Y�.��v��D��^�I��K�nu�ND�,K�{����bX�'����ND�,K������bX�'���K,�wd�r[�^�I��K}����Kİ��}�;��yı,O�w?LND�,K������Kĳ����~��lWJ����L;L�y�;���X�t�jF��z�j���qT.+޵w��ND�,K����'"X�%��~��ND�,K������K�@�o��mxj�j�C��D��MMT�57u��r%�bX�{����?(�Q5���s��'"X�%������,Kľ{�w�Ȗ%�bw���joZ�ܖ�!nᔼ)2�)2����yKȖ%�b{��ىȖ%�b_=����Kı<��ىȖ%�bx{�Yx6��[V8[�o)xRe&|�!+)n�?LND�,}����O=��2LT,I�(m5朝���w��UH����54�u�޲�ץk@��SM����Ј�\�1-i-��ʗ5�-��EwrS�2�#
�Xn��+x�0ݶ��v��@��S@���h�Jh��4�Y���8'i�89��m�����#��ƀ{��}�)�|�e�ds	�(��"�b�����=��gͤ�j���h�g�x��$��Hc���{��>���>�+Z�Қ��k�9��Ȝ�޲�ץj�����=��`|��Hm�I.�A}ɷ��'2	�[���;��o5��#V�#�=��5u���b],�'>��g�.�Xer�=X�]�]�3��jl�,�v���6�{y����شm[9l�/\)����4�ύ�_tQ�Z۫�k�N�8�l�6�2�7mѩ��v�=@l�����Ӹ-�z1��d��dܝ���U�ĸs�N��K*�N�n(԰ӭ]�R�Ww{%5��Z��9_���&�nn}����vM��*�
�h�l G^|`H�����L3�H�F���k@��S@��)�}�)�}���k�p��Ӎh�Jh{�4?l� �}�o>M����Ȝ��H�p�=�~4�e4�Jց�t��}��=� ���n޲�ݵ�f�4�7���3���N(��H()�ҵ�{�)�}��>���;��V�jLR'0NH�2I�;����[p��t\f6�0�:�0�/a��B�q���A)#Z�Қ��M�YM�ҵ�[��)$M�CmG�mqr�?6�Z��ޫ,ͮ��36��>�uod�E#����4�e4�J֟�����{��h�Sdq51��Dp�>�+Z�Қ��M�YM��_�X��1A��=��>�Jhz�h^������x���������OP�֬��Q)���p�`J$Wb�і&�����Ƭ�H{6��=�\X��4���WŁ�g��'�J< ��}�)�}zV�{�4�Қ�J�W?�1<�(�*�ݵ�f�m%�%�1�(n���^�ږ�Ԗ��Յ���q`z;����	H)�=��>��<��L��O�vu��oc�.�r�j8hwJhz�h[+Z��������~v>	�n�m]]�2<;�k�*m�]mz�4��n9��jM��e�>�Ɯ4�e4�����O� ���wt�vK��W%��[�`nͷ���7z�,��Ł�̹"*bL��Ӎh�JhwJhz�h[u�����"� �#Q�C��7�o��`{��K	��Q �	$��b�"E���!�])�� ��~�$�x}��XD���i�@��S@�۬�=�`~�i�rI$��Ng\��q]�q'L�ݮì�V�h�ǝF7N##㮲�u����L29����D��>߯�f��t����S@��S@�^�b#�6��I�h�Jh{�4�e4�]f�nu�'m
CmG��M�YM�n�@��S@�=R�"r7$a����������=��>�Jh�Sdq52H�Dp�>�u�f��k���Ł���V�!
R�h�F|eD�D�3U2�58�����_q����m��v$[n��c;v�7^�O�,�\۲���h�B�@�������S��l9��j,��s(aa��{h�icb$�ӗ1�knpq��\byc=x�j��<�㳭�n|Gbݝ@x�.�!�ծYCc���.4 U���/V���=�%�c�NޖN��i���={f	��d����	�''7b���B+Nn����m(m.B��Y5133Ъ*��3#�6�$�o\�j���g�f��L���7�ܽ�ı�%�-F�%���� �}�X޲�^�������ɀ<���}z�hz�hz�4{�4�$�#n(�Rf�����׮�@��S@�����T2�����D��0>������� �}�X�?��~4
�_�b#�4�2'!�{�)�}z�hz�h��h/�/�n��𓦙]Qb�m3����t'a�z�N^(a-��
p�'b�2�o������ ߺq�wtd�8�>�rWdRI��R�MTU+�����M$�&��7�4��~�.�;k���oZ�;�����52H�Dp�-��=��>�w4�e4�u�5�)�2%RC@��S@����>���-��=Ϩ��"r`$j8h^��޲��v�Қ��QL�$�q���<�[�5g����#t�1�<6����:�/"�6��H�Qd��L�>���-��=��>�w4���('��J
C@���@��S@����>���9^�b#�6����=��>��>��_T*^��UI�HC�M��Z��q[� ���J2+ ����
���t�4���++C�h`������͌`�HP�4?.�HF?:.ͥ01o���ѱxG|��!
	,#sN�$K�K���|�-tT�~Q�=<ָ0#�#� mӆ��(�Bx`]!�ѭK�I�{O�O>H-Y�ŬXp
��i�� �"���J�&��I �8x�E��8���CG�fMKC`i�dؘ�;�ڞx�����'�AR�_F%ГF	�C�3�O 1��v�Aڔ�}OTM �F��1���z�U !�$(��E�\���Cj�Ҏ����jSiCi�����E�q`fw]����r��+�n\0>�UO�ox���� ��rT�R~����{�����I�&9��}�)�[�a�{�)�}z�h�AdVc��6L���q��u:�^-�ϵ<�8�r�-��ҌQ��(����d��#qi�@���@��S@����I/~���w��m�$�n]�TX�\X��V����z迒p�v���-��E�#��wb�<�e4m�h�Jh�j�0�9�䃑��>���-�a�{�)��3?�N���B���tw 6@@�jR#A��FR�]
K��$%�@ m=Xr���$���\�PRc����m���M�n�����|����I����u�6���)�յ��t��Z�-�2!�ر��e�N � �"r�Қ��hz�h۰�:�u$�p�Rh�=�֬gWwu�`fmq6�l���vH�ܵn��K� ��N0m�h�Jh^���T�$Ȋ��4z�4{�4�S@��S@���P��G2%RC@��)`v�q`{6��=��E���c�w��~?f�v�C,I���AO�u��S�Z�����V�lq�x�z^+��4%����SKp�����q��^Ѽ�I;��[�P�'F祉��y7BTj���t��w=s�&6�v�
t�y�vܛm�K��������Ȩ�g�L,��n6st��`�7&��|m�ێ�s�4q�l4����FM��;�T5�k�1��zػr��{���w��}�3$7MC�۷4t���v���c%�~���^d��,��+t�Q�V%e�m�䄎�������t�����>�Jh�j�2)&8�2�@��)�}z�4�Қ�)��P���F��4�]����S@�e4�u�G�����ddNC@��)�^�������a�u�u�$�I�c�q�@�e4�u�׮�@��)�yx�d&(�$��#I� ��UƘצ�<O�m�mn�۶Q�aF��JRu�f��(�L�n�����a�}��/YM��6Is$m�D��I9��f�p�=�� �Mfo�����h:��j�I&D���>�Jh�S@>�Y�}�v��m���`�BG�ڴ�u�޷a�}��;�j1=�	$�x��@>�Y�}�v��M��x�K��iwnƹܴ��r�B�08�L�slQ���
�O��mgYc�S#t�m�x���i�����~4�Қs�h��4
�u��	6A���h{�4�j���h�S@���q(�1���h��4������uH	bAN�-Q1AM�I<ο�۵�`yf��U
f��lɑ��@>�Y�z�M�t���e4�*ے$�Hۈ�NM��h�����7zq���f�\���_b�M��Xض��a睰��:�+��V���:���{.�znع�J�B�m��ץ4�)��@�����&�H�p0y!#���e4��h�S@������Q��I&H�H93@;�f��e4�Jh��h�2��xI�#MG&�z�h^��/�}�I�p!�T�G�T.fff{�~٠y�!��l�nC@����z�� �u��)�z���t�j�(��U%&9�� �u�WMM֝��^�n�V3QNl,ng3��z�� �u��)�}zS@�=QvE��(ٓ#���@��Zץ4��hlU�$I�q��L}�׀y��0��ov, �w�s��5�jI1��Zץ4��h{��/;V������"n$$p�/[���@��Zץ0Ԫ�J�٬r\�d�ۗB��^��^-������e�zfrQoZNY%6�:GI�s�P[����	�����]Q++p:$��\4�\��7k�7D����$:�;l�=���)�G/�q S�`�T�i:��}v~�nz��S�K�<����a����P:`X��k�=nu��M��1m�U�u�֎3M�+�;"z�l�Y##o(VA�k�f6E�����_AE�����[rɗWWZ��KCF49ڴn�\��F��WF7�\s�@:@Z��uŘK�L�k۪\u9�������^v��Қ�w4�(es ���@��Z��M��������D89���F�$Z�Қ�w4�[4�ՠ[��<&8(�6���z�h׬�/;V���M��W\��Q�&F7 ����j�;�)�^���bU��i	�kV}�e#��8�a�-&��v� =�.�خnӭ�l=[-Ҥh��o�4�=��� �vi�*���oL��P�4廒&�d�`��i���J�%�qς� H!�K!�R*.� �J
��Ͼ>�4�u�@�e4����)p0Y$Q�@�e4�[4�S@��S@��+1��d�<Y&6�z٠wYM��M��hv:��Cc�1F��;�����M׮�}�f�|v)[��18��I!�8��6�f�PZ����t^3��e㛻Յ�6���c0���$pr�Қ�]� ����e4[G�xFD�����z����l�;�S@��S@�=R�d�2UL��Jf�X���ޮ,�iS=AJ
� �������d��>��(�H	̉��4�)�{�)�z۹�}�)�vu�q�I&4�#���t���n������e0����+�[v���Z�KmF���ƒ�I��jjT��h��1� �ѮV���x���CW!.�wb�<��L�vi�{�)�_e����2H�,��4�e4�)�{�)�z۹�}��2�xI�$�'��h�Jh��hz�h���I�#�!��M7���֬gW-���2� �xU��7�$�}h��#j5mG����YM��h�JhZekZ�
9"s�5�մ>l"ь�ֹ�1j���;NogLAf�G6cId�<l��ɓ�4�e4�4�?~�iԼa�wb�7oGk�;�;�w�vi�M������ŀy�f�ʒM�����Z��%� ��?���޲�u��=ϩ�<R%2$,r�@��s@��S@;���Қ�YY�őd����4gW�Ӟﾬz~(nm��
��� _� _�P Uj���D _� U�@U� ��/��)E�A`�Q�T"E�$Q�DX!P�Q"DX(AbE`�E��(��Ab�E�Q �`,Q*Ab+E�E�)E�)E�E��E��Q �DX�E�E�E�AP�AcE�DYE�DXDXBEdEDYE�E c T$QDYT$QPG�� 
��( *�� ��@U� 
� W�( *��@U�
 
��( *��@U�� _ _�����)��H7o����8,����������0�� *
� h ��2�@b�� S�k��Q� 9}!�    4Tꚅ)P (V�	J��!T �@UP� 2�*25��SP^�{� @)<�KlP �p=<�F�};���۔U�ݽ��ݎ��7��)���>@�{;�����m�nϽ��r����SN��wc�vM�G�� � �Ǘ��-�.ϾãG�z��}���:=����n�݁�:�8��|�u����y�J�x:�܃�F������f�ѝ������pzw�|
 �5x& ����#��Ó݁oNl���>M���2*�;`7g_}P��aː7��E^��n�Gv[�p\�غ�G!�u�w�
(��   ����_!�k�]n��s��:2�u����Q�`gu
�V��=�w�%�}����;�����>��{۽��8�׃lY���A���� �h��tm�]���:n�{:���v {0 �� ��\ �� y } �>������*�ݏ�� oX ��ޏS����ݝ9��;�     P  4�0��J=�d`�`i��OǪ�Lj�b       =��JI�Q@C@ �� S�j�b�U?T�       RRBb����&A�yG�y!�i��MB��ԁ�i� �����W�����	��z~l����ף�����JE;���TQN���E���L*E7H��_��o�v?ѯ��E+�R)�i�:��S�K�[���W�|����O�������+�U����{����www{�7wwwwwwwwwwgJKwww4�m0�wwwww}�{������������n��7wwwwwww�������3wwwwwwwwwwwwwowV��ݝ�׻���bŋf�tn���ݗ���㻻��/wwv�w[m����ѻ�}��{ۻ�������w������fm{����~$$�'Y$'P � !�'��Ty�yЏx){���=���{���^�/x��x+��{�]�.�'l�=�����{������{�{�x+��|h^00'�0^�{�{�y�=�^�K��ު{������By�Chy�y�Q�BpO8ƫބ{�Qy�{�z�zl���h/z��^�Oxު�z��UN�9����@Hu�	���az��"j��?�X|w��~�����sI�⯤|����J��N��,�V�^��2�hփD���h54�&�M�d��2PjK��QU��YE���2�V]oa2Cz��2CsV�P��!f�jKkWh��d�
4s+���]O���EI�6ڜ-be��&M.M��V5zԼ��/-�b��6(ʬ/��n5y��.��W�4jh��<���oD�ְ�,�f���[Z5ɡ������(����������)�0bU��\��5UT
�@�Yrz����Q �b�����w:H�z@"b�0�n��M�_����׹���f�G�2T*���(h�D�AL0��A��ӑ
�5�����CH��sB�*�����*�W��W�Ճ/��)0�����ZP4��R�D�(`*(ʱ�x�Jjok�Y\çw�S���N��0-����R͛��r�v��Mk��ܠi����J���0�	�@�$HK�0h�n,Y���qu��4t��h1#&ᔨ���ӭ�%�)�U%�k8�4!E�A�j����+��Ś`T���Vl�5�櫭;쾍&t�/5ؔ\J@����S��%N�h�B���40`s8��t�N�\��W����o3�V���䪼Љ�
+E�EPnZ�1"Q��n�5"���e�T5�K�v�Q�U��9EQiK�U�u.��E��mvT�O�@��,?9�oEJ(�3G9�j0,��z�ʽ���E	BSrtP��a(�`1[#���m���8.
��Q�e���5f%A�@h³�ֶ2�s6ѩI��N��GѫcE�eoU\�S�j�&�Z2�&c����Ʒ;��6�*%T2����D��n0�׷ww��4X�`�5��-���D��3	f*�F� +��f��m��_O!dj���E".��'��ŧ�y�1rҺN6��s��\ͳ�@`�b ,I[��s�(FD�l��*]˻0J��h�R���8l6.N14j^j�E�Ӊ������7efW�Fd9�h�����f��R��Ki����`���\�N�9��MZִ^�]�3��͘TX"0(N������ $D���W��҉����b�r�%CX�Z��x�yy��jwDA4���f�z��
zl7�*���Ό.D��Լ�#9ǖX�0��U�a�Ws�"�X���Ѵ�Ы��o�ֹ��@�)R����x��*i��a��5�zPt�9�
�T�`0CJ!*5}��kG]t��N��q&&R��.¤�c@��Uwf�)��E[3�噭n}^�b��
t����6W��5�D��
gbJ/Qy���]��羚\&iv3k�5��kF7�0��F
J.iw�tCF��H�H�Ȭ�� ��`0+{Y�<΀�N��w8�wN7͆U��
+n���3Mf���$Ѣ2�Z�kW�oon�/�4Y�����K�Y[�;��f�f��E�fMCG%ަ����F���^P�F��wW�n�6S�6�)#~��� ��`B��w�	W�y�<�!�^�2,�L��H�5U7w4i㙚j�H�]�`�*�X�(�-�����FV�©���ꎯt�p�YL�}�
�Rfc&E<�8/*�O-��^��/vZ�F�5R�/!Ux`ݗn�P�o,0�fĢРeCF͚�*:�A���E�J�fA���/�.Q����5��gE��Rɨ�MA
/bp��T�%��Y؝U~7�W��f�X6O��1��D	���e	�L��A*
2���$I���X��7N�Y2b�����fd��Б9W4ka�9�t5�|�x�{�r4X4f����_4%F���ɋuI�щ��y=@����kGz��aE*Į�I;��e�ˈR�����%�[�*��7b5BC4s|q�+S%�(�h�H$(��/%���J2A%E�Hu�ݖ`��]$��!Q(�B
�B�*���
��MR��BD�hU�D��H�5��6��g�E)§�(�Y���Z�13�9<��@5t(����YU��$*D
Q�ͱ��d�w9��]���xN�N�Z�w�uz�3��њ4r\��jl`�w��w\��cE���C�캣Y�l��Z`��+*W
-�%�mz�ݞicc�^$�kʠ���r�~��
�Sѭg���l����/1K*nh�q��5ʺ���-Zrc�r��lj��u]�ȶ�e1���7U�܆L��еy%hV Ȥ��YL�LB�f�͐J�Y&I	"E���A��eKֳ}��;9;:h��Hs],���0���@��$�qݏ ���R2G��V) (dN1��GT�6wC۾z<*����+{�����LB��*Ptge#E��й]��J�W*�^*d}�s���eoa�E��@��Z�u���hB��U��U���kg������B$	��t6d_��2*��4D��l�Z^hFN��se�lb0
,�u4؀f�{gf/4H0�j�;Q�0@b��P�2@�/Zm�~����]mb�� &UП1g%,H��#@x�-eN�D���ic�Q�����L�v��F����{���atX5fA#��x��:+]���*��-�ڮ^*`aPEB�ʹ7����%p�cL�����v�](����|���
�G�W��*U��h�NoON�Y���U�l�g{֍�+���n�Y̻MY|X��^��kw�w{Եޘ�c(��Z0���s7�ԃ�DT�E�R��ի�0aխ���e��q�4e��ic�O�8�ƭgYk���F0(�d�ɛ)�7�F6�,�,K0����P��jC�`$J�z6g7�Q�p���JӾw97 ���o6s���E�:۪��٤¤� C��bUUh-�B]�D�u6�e8��6[�<:yL��y5��݀�ƑI�#�W&�4��+��$�aGK�Y+bq*!`)�c�on�w��G��gy9�瞚ρ�;n]H闷�[v�&�JNƴ8G��'�;e���5l1�z�U]��I���o��ܢ���?�O�|Ѱ�Bpu��N�I����~�^_��>� m���h8 ��V�    h    m  m          臠                                                                            �A�                                                                             }��                  �l���%�m&Ű-M���M.�J��('G��Ul��(  k�[�M�m���j���i�#����ΘM��b�(�P�;`$� � �A\.'��Bl\�Yӳk/F�0�m��ڀ4T�!L7+�誃6�z�-F��ۜR7\*��er�
�JT��7lAi�]����"I#i��v��'_}]|�̫u*�UA�� ۶ZV�������[,���J��m2N�֌�I�k���@�R�ݶm�$�m�n�		��6���E��%����a�m#seU�d��UU[J� ݶ�6��m��H5�y���f��l�M� �O��B	U2<�u:9�m���-��ڷF�8 �b�� t��ٙz셽�\ӵ.Āն�! M�KoK��sgj� ����;s�#ϰE�[�vұpZC�]��k������a@�톨�ѶϕIN8��A�Wu
��h=�����I�kH��۞ێ��NѲ��k�VC���UTy��AN���C��c���6�7/�L�\�a�RA�Đ@5Z����l���}��eD%�H@h
�`-�@uT�[�2��mU�br=(�Hq,�%Wiu,
��9de���U�x��9�kn�� h��V���@nU�6�+ڿ����vP@j�Wv�g�@nC���#q��)s��
�H��s��k�r�l�-����`�B��v�ny�uu�;� ��60��-se�l��K���wl�4}�N�﵆Z�ݒg��ů�M����Ь� H��l!�t:�Nt�-�$��^��m�z���Iל �F�m]��-�0�a�E4U�Y�Ͷ�V魗Y�l8[P���ݓ`j�3��Tmڕk�*�P��I�m��ڥ��ŵrz�؃�$��-�9:ʶ�{m�J��i�q���A�7I��4�l�UUD��@�%�}�����[����(^�VxH�N�^�!:^�LJ�J�Qƭ��ZGv��l�T�UT��}O�t�&����-Vڄ;
�]J��FR�Y�p/Oku�s�j^�{4�5 ���u%cu��vn{6����xu�n����ST�����eU�Єpl������ 7=��j��<5R��!LR���F�ԭ��#m�a��mÇm�[@�	zS�m���  m�m�-�nٲ�m  l/m���UBK��� u�CA�H@��m� ŶF�mk#M��hm�� �m�` � �9,M\�ZP�V1�KK�Q�2�UWC���@�V����
�U�,�U�,v��614����m�m��[,�v� 8�m�lH �km�m�� 8�h��uJ��U���U[h�r�`� 6�  �ઐ���i�!K.�h�  ���H��;m����z������m�v�l6�m� I��z���m�ն�m 9�m�5�Ŵ�m�ڶi6(< �m�-n�6gZ� =6����B�X[�� � ��7]uꎹ�t��m���)rjۇ`�}���e>^��[UKn��w[� ��o`yꪫ���*��K�0$b���k�{f��$�m��h�ۮky'>�jj�
�n��jv%�V���r��������m����U7j�FA��y�-U��vyD��k�\võ���te�v�Yxۋ����� ƭ�dD�Ue;,�U꫃����p	f�m�m�6�:ye^�-�hеTl�Nh�t˯K�D�*Z�����e�{e�V��YlӵvId��8]Y&2��;&��]DUT ��1R�meI���j�5��J��Ą�f�t�m�0���]z�[XQ�QD�J�Y��kM�U"\�֩yӺ"d^q��nM�:J\vBY��'`�ڣ��c�U��S[n���n�΋9:�Y������p�譸#i������lXqfq��1�a����rھO���ls�,�a���8]��Zf�&�f�V:Vf�-����ᝦ��6�]5c�%+'�K�F�_�Ȗ�k6v�,�B�Y��a�`����m)/$U��!�`vN^8��<hE��r�A���
IRM]��a� m�(��P�Nܰ�r��l�mE ���d��ôѰuR� �ʵuJ���mU,�(����,ң��[��q�f7:펎*6玢[	���wj{[
ʫ�i�.aL!�v�Uwm��U�Ç,�$;jڔY���j�VZ���$�U��Z�`�6�m    �l�F�z��%�Z�4S�*Ŋ8�h�Um�W-аp���K-�E�yI�V,͌<����RkhI�l  �m�Ἂݢ]�bB5�� �lX�`�iV�sr�y]��ڒ'�����Qێ�Nm�݀I��Q*d����媠-��m�Y��Z���;qSծ6�J����ƶ����v�el�:ru5�v��*�&J�
<u��Y������N����-. �Iv�u�ڻmi�a'kՍ���mN��KdͶ@q�m����,کT�c��d�M���u6 s��_(�%q�x*��ꫢ�A��4��b疮����}P� Ҩb�aV����Uiv[��w-@�vw�0����oZ�
�:�ˏܯU��[�J��-饋*�3M.+عkv�V�ܵ�u�t�eHԄ�J�A�d-y�]�V��[W6��@ �T�m���@as-V�P�q���g�՗�ni �S�E�$kx��88�lU(��[n�*�W3̗ɸm�m��s� UU*ʡPU �0��vyVX�e�H��uVª���|_UJ�n��E�T�H�L\��ur���.��U[uR�� ��Άצ*m?/v�=����'�����R�_\�Y�]?[���#�88p�8c�8c�8.1�j��-pYe�b��qb�����eŗbq�d��������yÜdec<�1�q��u����l�Д��KBR��;pln7nǎ ��ǀ���q��(� �=��G�#��3���q��8�xc�yc<1�c<�1��1�G�8�#�g��22���.�������5�Y'���Խ�_��~������Qh�F��y�6�1����I���ާs��|%�=K����fZ���Tu&GA���=F���N󺝅�rJv�0wnԹ]�#M#�.'T켫j]�]Lzq�Nz^k��	oGT�����;GU��S� �'�Ү���̧�>*OGK����D�qN�r��Wa���d���G�|bv�'~��H�j�Κ����eރ��
wy�>�CA�<�T�N�*;��it.Jzi�zU�t�G����ȴ,^}W.O���薢�x�^G��4r%�OG�^j��|*z���8�Q�9Zks��s��rm9.[Q8SQx�����G�U�#h:��]����^���d�\3�����VACP9�C���އ�=��xN��ٵe�f�q��5�)ړT]��W{R��&j�CԯI.��_�zk��nsN,��͕�<��+�9�� ֍eQ����e����
���^��jt�橆z_�>a�>��
E5���;�C��SAL
J�?j���1��e�c��]Y�N.�lΔ�ʮHT�6���ӗ`Z
��S*,��6���*R�TTH(L޵�[� � ���              l              ��  �d�k�	5��&��s8^ԕ�m������\�E�1 �����0ۇ��g'Hy�J��]!�i�K�<��1b]��ZYZ��CX��S@4�(<!1Qs��R������ӛ�Vӳ�,�����ŭn�����1Gks[Y�0c�A�F: n��H�������n��zۅPݸ�ܔ��eM۶�v�r�ݮ#p(05�E��ƕ�+p=��h�֍!��u;�D�aƚ��SJWPK�aT4���;VU�8ej�����0���� [���d��3�86j52��E�V�vd�qa��5������ζ��ԁ�j��VP&�Klaj [m.�;�r��s�'W�7@ҠR� 8̇��"��պN�.�g����l��G<qC��k�sۓ%&r�
����W<��7#G[&;'my�8�X�{C:x���ts�r�>2k���q�Si�DI5k\�S�	8e���֒[��ۖ2Ԫq�GOR��g���Lt�^��X77aCutE��U�\:�q��;����݈�"d��2`z��p!\4c�s`x"�uU2�9g�A�
����@2��A�gk���%-�JneJO�0 t >P� 񧀾u{�$1/+ڌ�ҧ��������;)��;��ϙ�O�}��m�� m� m��f�ۭ�r���d�����U� ��n�ؽ�F�4]dݱ�VYJ�#��!�jH80۷�] Vs=E�Nу��f�q#I�f4���[��sr�s�<ɱ�.鮀֠T&��.�ڣF6�rO;����޻�Ux{���ʼ�r��@2)퓓'?���U1]���4� EWs��'YbfZ�%8��_:b��Ǻ�я�5�i�jhi̘����q��z�]��HL&����=��35>1UXN�ࠤ)U�z��f�c���\{7m��r-��L�]s��Pˤ9�Q�R�e��v���MT��<�O�g*�X�޸�d�-�(L����D>*4l��XC��!�:sZ�wϲw�B�n�A�2Q�6X�^1����0َ}�6��JAɗB�88��`��ݗ��2��h�m7�BόUn��y��?{=�Un�jL���J,t�]uہ�"ղ�Pc�&�nFY�����{��آ�FaiĄĦ̑}��]��BϮx �^��[���t���y�n6���EkU&��uK�;μ��q�X�Bd��e7�����1�qys8�\�&S�i�w�X�޸��:{���UY��Y�ttG`m��Nh�tG�su�n��Ɩ��)�gv�//WZ|ck|&�r�J�F��k� ��a7 Ww���!��2Z,4[e�m�g�p�����s���e%.YT4��~�f�5�'�O�Tnd�	���ϽG��Q�&�^n��q�hY����m�B`���v8��v��aN1pq��bg\�ƍ��Oޞz�9�L�{��z�O!2K@�Sq��d���{o\^\�Z��-9
p�]����B�n�L�a��� 9�ޡz��{��6a=�E�A ��T/s\v�1��Wu��DC�*y)m��l     ���Tu*�LB�:�Z̑;66ܗ�s��͜�m�����m�@Ll���b�`��,�9��('Iؐd�tnҍm�ŋ+�.ݣ:���ɈͬL�`=�q���\.Uyl�8��Ѳ��L����Nr�rt����tQ^���zR�<u��`f+B�dx3EJ�)�f�,��n1�qᛣ[�2�H�8z "�1�����/$`ƜHl&�fޱ�`g�>1����%�)șT/s\g�X�f=[n=��L��l��g��2lǻ��u� D/$�sm��������.�s�!#Q���h����`��8I^w�=��_��Dm����R�0��s�`v'��X�+�ʸ�� o�"<��|����h�$�SB�5�^�g�&�n�t`�\�Җ��: A��l��=����e%.e�i'?]�=��&�X�黖�m��Yg��ݓ0�$�i��k�֨V̳;7h��,Y�s�}���x⽥>0����)�!J�{��P��v�{�'P�%��M�f�W2E�! 8L��0����{w�Ʈ�����;�c�z�P����R�%3&'ۧhV^8��,��j�U��m����=����?vW���s�	���U�+�f�F�w<�ߞu�,צ+wm�˒������_ 1]�Ǻ�ǆv�l2���sH��w�=��+7X���q!��1~�c�x��%*|��D����yxVdI2�B�5�D_cl��<G��6�;<NҘ����/7 �7H��ƚ�FRH�t���n+5ɲ=�=��3�8��)MCNK��=��
�B�n�MJ0�F=��{-a��Bόk�i�(Je���+5>0�m�퓌�!��-$�P��v��޸����b �:���m�     H����[�Q>0q:o3�����;1[j4���z�Z�v��j�lЍ��s*�yy�kkRg��9:����x����� ��H��պ�D����n�-��v�$�qu��w"��9�b�X�A5VX[6v�R�rI�x�s�w�j��Ԙ���j����h)m8""�l��0�W��(L�S���~�q�a��B�E�i��L�Ƿu�e��Bό:�$7	��*��k��_@����q�p�Bd��e7�(Y������KJ�������SvǶƸ�ԍ]�V�m��nL�r���O](��"�u�JL��L�%&jPA�J1{�ǲ��f� 1��\�f�)��P�I�ׄ�&�Q�P��f:e���ϫ�rCJZr�V�|an����5��E3%�ӆ���޸��=r.�N$&F+wX�^8��,�� �""����v�C���
�y���'*��it�Sh����w=���+u0�mǽ�u	�Z-9n+5p�l��wc����D6�u.*R2�E:���s9�?�J�������T[�QTU[k��d`�Q�t*}�������?�� ��&��|��u=��Ԧ0=��j=G�x=\��L��tӻ�Ιw�G2��XM�澐�>�m��H�D>8N���;�(��a' �H�Z��X�V����Oow�����_;�w�P�ԃ<�h���� ��hK���D`^G�˒"(ꐾ�:6	��Yr2�� �H*���}��H�@2��]�f�ks~�F2���!����eOf�WQ��i�~����qO3Ի���ʻGȏ�8���x�lNN;lͧp��ʏ�Qw4�%��/U]��_w ����y�>������R�"
s߶\f^8�j�� 1Y��١Jd �I舁UM�}�pq��<h��4��6�l6�3,F��L��k��mG^-��A�L��w��Y��C��\X��͆R)�sC�~�c��ڏo/�\��Ӊ	�ы��b�1�]�xхU�D��)�*��s��{�>7|����ɗK���P>gK���4 . @�ߗ���bu	�Z-�n+?!��v���������m�s���]Ek��C*�z�e�Yu�uؼMk�k�tq���O��Ǿ�qY�?M�i�AC	LɎ��y�Ⳑ�N(�vhR�%I��]����,ѰEn�b���J���-0+7���8�{�v8�v�a�R)�sCM��\�]��d�~��@�M���4FD��J�0�B��
��>�ym5[�     U��d�4�4�V� �"�ŗ)�n���V�1,�XT�Gd=��n�F�3ٵa�4�؍�b�$���l$ta�N�,���G�b�z�di���I�_�[l�p��3qEq�⺷W��&:9��d(�Rb�}�w������}~*�u�4�xx�Gm�6�<�Y)��2�N�7��4a~��x}��B��!Y2a�h�!2
Dʡ}�\Vo1�Y�wc���<�˙�KnS�=��d�wc��8���\T�e4U8A.��}�B��&MZ�5( ��_w1��7��}�h�z���UY�i�
�v���e��P���b6Sn����A �Z>��:������ \�}����^>�ɗu�Yy5��3� 0(��b��,O��+� ��s2�L�sC�~�xo�\{y
�a�91�ퟨ�ڊ��7f�?{��	�Pr&U���P�F���g9km��NC
��(2�Y9z�K#Ǥ[�e�)���
8X������<>0����v89�KJ���d�6a������*��6�A�f=��{3o�3�&-2/\�f^��2�����5ϿY�擙�q�̖$%��}��J��L��wkG���2\4��-8�rh�D[�B��j+�9>!��ʫt��fk.�9J9�D����M[+������a�T�e͏��~�c�}��G�����Ӊ�Da��b�u�Y�Y���D��)șJ���{W���ӸX���8�Vb�fM��g(3��|�p>�vHg�k�_�����ub��T/�LVf1�qY���̕��Y��(eɢ,�)�0�K�ш��n[k�Y��Jd��c���ߐw"�\�nH9��{w_� G��1����������)jZqY�;�a���1ǳtk2�Mʙ���ح�q�  ���Ӊ2J`{�X��{���?@d�	N$8����5��UUUP    ��Y��̷P���Y<���ru�X�q���r�;�{;Ԛ�.:���d>-�;GS�h����q�s�P��2m�--��'G�<���E��Nj�l����|��ָ��F��un3�m΅���-Ӝ��NNt�Uf�tj����$��89�Z��1јu�6�`L��k����?��E}�1�����%��rCq���
�����Ը�AI��{fK#��ʡ}��=�mZ�d6��@o��f�q��*�{�C		a&�{w\g�rn�ݕ��۝�WK�)%F�Y�kx��k^Q�U��~}��]���N��}�g�wc���Ѭ0�E-M��!�9�a���
+:]�9D*]	r\!�I�íoz9���3ܺ A�H�iĄR���c@v��U�<$&ANDʡ�"wuv�!��
"  }�q��Es�%��r�n�1� @� ����C����3���n"v^�M/@��8��X���-��?����O��"4<3'��{��e��  ��B�s�$0�R�hD| ���@v|�Ԍ�#���5$%������g�~���~@$ ? ��9_P_��4�t�.LJZ������z@��xH���o{�0�)�SC�@���ME�k��B�}2��i�T�:-dJ�l�M�s�X���?����o��,
3{���}����>��p��9*�ws�y�m��[��Q\�hL�ۖ���XO�>�'����}�3�3?�Fe�4: �,�o.��k���vy�q'ĺ��t�'�=���
�ߙ�$�S'��c��ޢ/~C= } {�%m��js,�r
з/�~�|}�)��/�B�\�dhe:T��a�*����+5q�d~�	n���<>d�iKR��,.z@�p�=ݏ@n�a�RRY�d�uv�  ��c�'���vӉD����� '���3{����}��Ow%��?�/�����߾����	 {�����>v�����?��b����m���k( 1^�99d$��N��%x�����Nse�|�W���CA����	$��Q��1�M��tMh�������fN�.9h���q^E�$`]��D��e��th�\��!,��M�:��[+bK�Ӗ#�uul�D$�9#��F��㓶_u��+��%�kV%���Ss��Dv�A ����p*MF0�������0:���Р�y(��vM�����3q"�<U�Ŋ��vYINJI,!�ve�m��m����                           ��       �ˤj�wGe���w2�	�g����mۨ�R^Nќ�kZ^�<�sgg)�f
�h�;#"�]�q�O&�]u%`�5HXŧOv�]�� Y���\^�l>gnO>[=����C��n�nY�u����P��W]4�Ť�<�kZ��aI�*N�</+X�+.����Ӵ�*n�`8���v�VU�mj:��͎���.�����q����/	b��X�6��E��5�kA�]��H3m��VnV]�C%�mp���6���R4�*���m����52��R��c)���=� �)�Jʄ<#δᐞ��
� xLI*��A�Lu}�������k��v� �y7WF�Gqv������������`��jz��	^K8��m�:�;=gi�z�V��tŞ�r���V�i571���b-���ݬ�+`�3�r��c��jq]#�ŵd嚲2��y�&.�--����ژ		CK]d2ۂ6�cac6� g,��Z�j΍�`-��lq���7iW�
�@9|�ˍ�[,\S�ى+x#Fnru����V=_#ű�\���\���ӚjU�dn����Y�T���[Ԅ!˧f����?�?���UUTUUQEQEQEH*�*����������*�������l��^��}*}���ʟub���.�}ǅUץ"� ��'�#��tH2h�t�˺��     �ͥ6l�nS�;�'t��%�&q�%����iT�,!�u� A�u���]4�[q�'nY#6x(��ثlr�ېG3̫�6�c$sqq@u>��[vv1T`	�l�!��(���y����Tk
�8�q]�w~=':��I����Ufdu�ֱɹ���ozF�J����æB�!$ʦ��i�q]��c=#���쨀"�o���ə�҂H����� D���3�\_�\ A��1��RHa v�1���>� x���F܆G�@��Ձ�h�X��� ��D��B�c  wcNd�iKRӌ�.$DFyB>�����<���~��q���*/E]%�݇�e�ŮLM����DKlS2�Neȟ���͡��_�� ��!푺ӉD�S��z��@���g&�s��ዚ�p���I���Ϸ�N����?��!C�s�~(�A	ɕ�}���o�"\���.���$��r��  v�
������ 3�f���2��SP쑄� z�(_v�#o���k[m��L�2�h���j�0h���]x��'&����XH�
@��M�덾� F��s���CE�r���|  ��X}3>��TbǧF�5u��x���|��!dԒ|����qy��a�RR̹����DF|���v}��ŏw>L���iĢX)���� �fTe��5��mʃ-<t�Fh(&αUٚ��rIrΥ�!3m���}�����G `we^�W0D��NS���� � �vM
�Ǳ ��;̡)�����  ��X���\@3��,$K	L�~��D	߾�1���=��ק_5N8p׊N��*���:��w/�P�@�	5B�~���� v}C�o'_�ߞ����UU�2�4���ւ��S�ղ��j2�s�""r�9R�Zq��;�×ݾ @��n�j/{�0�))r����� |D	��_�s��˄  �$b��"XRX��Cٺ�@���d�������!9�T2 @����ȓ� ����`�`�.SjS��C�6" {X���}�8�D	 ��$��>���m��`     �(\�l��HԵYl�[�"\��pa��͵�=��3�!l0�*����&��
�H�u�i[�]&�h,�m�J�m�i)�p��A�y;k�ۥ�3��*���V�̳W��FIg&5�rʣ.�2�o���H�MC5��`ئ컷c.��-�ų���/b���������Ì�Xk���fc���8	��=���,$K� {ﴱW��/Pw#�uu��CEE:��35p�@����Ӄ�s-0� ��A��QywP��ڏoh�e%-&懶@�@{�a��f|���8�m��mSP��)	o#���,\��7,�raPH5I�D�S3�=>��(����=�h�!2NRJ�����	��l<@?I6{_�r�{���!���a_�2f\��8��sH���=�u�7 n�����C��
�c
������U�c-ʕ%�) =}�C����h��g���y���:��������Rʨώ����T�K,�@�k����f��G@D�vW�ӣC�m)IǷ�� ������k��z �I�ߏ0�)6�e��{��|���<]�/m�Sd[B�������<B� �}����*�Z��"X)�� @��1��a{��@ �����$&A	�ʡ��\p�  =��d��ݔ8ݬm��I�a�dBP`frr��U[#�H������,(9��:��>��'_}�p" @�}ݴ����$�li�л��BA�w�7������� jH����Ne"XH��+>����b� �~L�H]��T�XI�/��=����� �䟤�@;�~�}^<a�ʖ�m����rV���+�� f�ߧ檇�O���!Vu0���G].����,�rp�N��R-�e͌�I���+�� �r��8H�����O�A��F����� � D�_a�HL�	��Q�}�_} O�@��k���J��$�Ӕƀ��+&�;Ǳ�z�V����eP���2���\{y�XL��\�'Ͷ�m�     5[�f�<-W;a�ыv�<��mY�3�V��r⡀ᦻ�ڛpbSRk[�����Uҙ�u��&�Xh��U���7��}�n��l�'K]C�<�]���u[���\�̫5�t��I���I%�9��v�W7=�%���6'\�鸱̝j���}?��_���M�R��f�*�a�����k]g�fP�bST=ݯ�m�f�@�v;<zthaÔD���q��qY ��>�������⸰�E3.hz"�Y��w`a�" t ��Zw$%��D�S"��P#ٻQ�����m��L�S	�H��g��������t�,�H�!7"CS2Un��A܎ Moc�����*S��]��# �ܫ�����櫛a�˧\�n�]�ݧ]�v]�G�)��s�{1��ݪ{?%�!)ٗ��՘_�� oﺣ;���\�%��@��ky�x�5�O��^I�ZV�feI�D��ڢO��U}�"MOX�D��m�ە	�傑�V�Sј$K]�rew
'k�3s��9:�gQ��k����T
��O��� �@ț��$�����E9���'ڡjn�kw*�>�o�� B*s����D�)��I;?},�w�:�g��ب������VҕV�����JY�%�>h*Tkŉ�f͠l�,&�Q��l9{��@���̮%@d����l�
���޴F�D����j�ohy��� o{�2Tw5�J���q��h����#K�{�͘��nLg�O1��T��ꞩ;S��Wj�P�S�����x<��~{OP�$�\H�Uސ��l%́'!6I� Nַ�1^b��L�,:$&A%&�sD�	�t����u�����P:���ް���{s��$��'<�I����s�/�`8��5"r�2M�8�bƮ�YrK.]D��NCk�TR�a��I�A}j�$绷ߢ="�=�6I����.T�D)$�ˎԓy�j��w9�N�
��=�g�L�h� ��ĩ���w9��@: 	v/�����t�1�s�\��I}��b�單��9گ�~�����@�}�D��g�|Xe"�j]{D� ǆ�7ݦ���͒D@�s;���mj�-t�GC/�ӶDGZ "��y����5��yv�:����=���MM�﨓��� 
�v�"Mڳ�Bd��(�ɜ��};�L��҉>�e�&O���`��*S�N�6I�Q�&o�H>�ڢN^O%E!)�2�'�D,I�Ge�kﲨ���d��5���I-"$�'5id�� ��{��.�_{��]כW��~�I��y>;����      4ҹywK��r�lv�Q�i%���d�Etl]�Z��z��t����(G��3bij�	XY�I��e$�����iFC]gtcN��A'u܁׮:��0f�s6�5�#Fꍩ�9z�DxQ���wm	\D��kU��F^V_�'�@�	,�H�{ʪ��d�'���_������nu�1���`�y��s�uzN���&X)��ޙ9�U���d�N�I�+9ROON�8r�̴��gs�Q��2}:Q&�ad��ʭ�d��+����-��&�$�ɣQ3��$��d���,N$0Җh�s٪�>�ڢN�6OI
w~q^r��Qx�yM]i]���i^��ΧRO�fQ%�Z�$��m��O��M�v�=48��ٖΫ5�qX�9�6�鄵.���'s�$��,�sB�RO�������ޛ���1�һ�7g���n.��R��6�C�	�Ϋ?Q����TI��͒s��2*CRQET����O��TxDL��d�I�D�Jʹ.L�,$�M���2�oy�I�$�&��d���p�I�N�ٽ�d�N�I�VY&��������sm��a'&��v�͜LE��r[��R���ɺ�+^�����I�,,�]�[=$��y"NjJ��X!�[2s�I�n�v���>�*� L�Z�̦�)K*Y�M�uQ'١��{h�J����O)�/�k�d��a�|/�	X���nS�M�͒jp�M{Xd���wo�����QHJE�)Q'ӥG@ה(���$�s`w���*�鑖�8�-�]cu�i��(���ڻ`�׍��l�ʒZFMo5�zgٻTI���I>$7k���r�ߩ��,�1˚W}�]'7���J���}|�$����Ç*\�N�9����N�X�3}B�>�ڢNI�+K�S-K�z@�\Q&��1]}�u���"��'H���s�c$�!��8�\��ɢNg0�< @������u|0��Ҫ�
�^�����{V�M�7R���#���K�N�8���.�d���N^�I��� �_0�>���&ZR�o9���#� /9��9_0�5��U�� G��䨤%"�Iԓ���&f��2O��j����I�-�L�&YFM� N��d�f�Q'/�T��@"��~��l���bKC=&f���jI� _u||I��>��d��|�<]�q���(�՗y�|��3��u��u��      �e7��˧A۴Yu�&�{�f�l�B��#1c��U:6'�N�]7o	�9�p#��	���6�'��ù���U����7O\]Z���/$�hq�G'=�$�{U؋s�^�6���E�q�y��Cd��W�I�y��$���}*�5٩�I.E�--�\�Y�V��M��ݯ��_���BA6����L��҉>�a�k�&����⸰�FS2��''��� 4w�I���O�3��V��7�j��#)0D�D���;RO�v���͒jp�O��y�.
E��h��}��'ӹ��>�(��@,����Ϟ��.W/@y��~�����y��B}�κ���ꪮ�vujk�Yzn�9�G����(s/���F��1۰?_�w���vW�@�Nw͒oWd6��S&��z��@Y:OBvB�sz����}L��Ү��,+$�e	a���>����7�?���\Y&��I��ڎ�4���~>�7�S$�vejz�2r&��z�h{���bld�z_������������ߐ�ΕWc:��x��lnz�pძ�2��B�'	,gĜ�a�j�*�ٽ�d�L�D����T�)0��8=$�wUx	����S�}|�v"d�^�+�i����+�}�����������H��&a�352�/h_:De��2�;�>�'ӓ��*R�H��TO�mp(��XY&����y͒j�d6��FMo̲O@��x�{͓����?I9�ϊ���E��ҭ��t��+f�[TȜ2:ޟ8�wXKt����?}��t�=P:�WL�Od��=<��Æ��-:$��@H��D���C$���n�'w��e"SR�]nt�O��z���	_}�D��$�ŉ�EKY�v	��R�j��{zW�>�}_��!�h#$�����I���������[�h��k�I��"� o}����s��W�Od��|y��UUٱ��Gg;�$��뜪�G�����P�[Kw���\���t�����}?d�@*I�v�w6yS		A�]�&��*D 7;��7��TH>ϛ�DL�bѬ�ZFAI��I�̪?@��7�6	>�(�z�բɔ!���g� N}�ޢNq���>�(�" k�����ǎ՚����Zw|0���I>�گL��������A��I$RR�ZP��mwC���)9����F���H#�a�٢uѡ�F�SC�xKdJ�*ʺ���XL4�F"3+��*DfUSp��r�1��\�9຺�SFG�ɚ�1�tE!���^",�a:&bsaAh�AQ�"3m1d^Ô�� ��Y�� �UU�`m�Am                                    ���S���V�wI���u�i�<��y��'�W=�;.�����P&Ik�̡z{[sʤOFRq�.m
�:ہ�kv�1�'ݢ��mg���g�fBM$ljƵ�zw>�qn]��g�5��Fq�S@�/$u��pvp^�G�+7k�{���0뗰Eð�뀚�4Z{7�����$��H��ti�i��H�ڶ4��E#�v''�n4Q[8�[��TT��Rz����sY�p�.��y�c�(��D�8l���f�mJ�[�)*���e-�8A�����|����
Y"Z�6��*�&[)�W.ۋ����@�Λi��c���ڦ�)�&b�]ʜr���ϟG1�꣰�V˃��B5�C�<;��\��'m�5�n�5�u�q	bw����g���J�%�;���6��)2(��Za�t�y��RCM�P��IksR�j�ks���	���(@+]�����kB������4<��2���"R��c&:W��ѭ՘��th\[p�)�A&�,Q��.�N�X� �[W8�(\��9Ӷz�{@]4�6�h	]4�h�'K saZ�=�Y���\��ۢK �ǯ��<�>����1�p�������qe�XY��㳳�d�̳�'�=�$=�E�(��u}h�x	�+Ĵ�^.�.�⇋��j�*��<�j�<��k��      :m�a�;l���r<�t��qۉ�Y��ӵŃ{.[g
 Zޟ=��v�Ӏѯc\�����.̶�7����_ 'C��4\�$�=95XHUyU�is���ًڢѴk	�g/M2�0�{�w��j����O1��୭Q.����8x�������?o����jS����(�Sw,�]�_�>��ħ��jg9\�$T�D�D���d���Us&�$��_ >�H�,:ʗ&���I3�}��I���&�
$���I��pV�2T�2��#��u2MΕs&��&�O���I���L$&B4�����I�̖I�v�r��Mz̼m��L AM@Q�c�7c+�+3�t���Jc,/��gIj�;��Ւ^eQٝ�l��҉7ޛX�368kU�;W�}���	���HA�%�Z���1^�ͫ��\�T�����.ë���}��[���o���@�j�'/���)�j]z�I�XY&����'w��}�j��"���h����O��x��ު$��D��u6۪l��%
;Pv�^ġүU��ֺ̮��p��O��k�$��d�������Nj��J��PW���e?�{�?�" 	�s�}k��5��U��'wg�L$
D�[�O+��T���4 � �F�+���=��D�bѬ�ҙFLQ:""s_I�n��nNsg�noe�O\�̠�2�n�j��1oU}:`:�| w��n�Uv&L�6 �ͧ��-�aܙ�T�4�q6�A��us���C����w�|n ��'��U�w8�2�	�r�s�`�&O�ad�wmQ&��dޡ�S����D��Œj�*���9�S$ז�I��|̴AH4�'� 7���%��G�n�Uj'ҁ�Q����Ke�a�ݵ���ԇ݀t#�SD��
����e:$換$��D����5��D���p�sm��e�����&՚7Q��w+�伹t�I���J�ѴԎ6���D���5��T`��l�q x��l�̚$�-/� 	��ݪ$��d��(�z���d�[4OM�w����l�f�J$��I��.&PjZtI���58y�>�œB .}ݷd�gw�0�	̹tI��!�}k$�vUo>��Ӯs�9'?����EUUUP    ��%W�,g��Y����Y힤�l�Ǜ�6���l�ui�8���/Yt6]�@����u�p.�>¶�g��Zs$��@ƺ,u���	��%9��hB1�Ĝ��s����h$��h]��c]߮�}�g������m����[V����N�[@��7�%���_�Oj��>�ڢM�?�G�#ț�(���>E�[I�4rf����f�{�d��k���  H��pW��&e:$�|�'|��q7?I�wo�I��zjd�Bf�؉�Ҝ��,,���$�sd�����ad�L��Œhf��NoK`w}0u��;eWE��V��G�����%�4�<<����a(4Yl�fN}��D��l�S�b��\T�<�B�K��@��I����": " \EQS�{|��'��U���=��l��f\�$��Q&���M}��nNkd��1bp�R�Ӛ��O�}��?y����=v��^jj�@}}��|3{��M�I��I>>�m��7t�0M�:�Ӟɴ���i���p������x:��M�I��	��\h
�}ݵD��'��($Z)Q'ӥ|	�ֳf��9uQ'7�����\9�\�Hɣ非�Y'ǟ^���3E�m{\��i�3���+8q�Bٳ|N�r�~-�jx�I�M����,�~������I�oU}:Q?O��Y'��B�K����o9�O�yieL��I�vMQ'���} 㶎4��z�K��l[.\��سlb��m�ͨ��NBR�s�(�^Ve�>����fU�W�$ޡ�S����h�����L�f�Q'���$�t����5��-�	����M�uQ=9�LЁ L�t�\��I������U`�Uy�� ���b��v�]��q{s�!PE�## �T���}�$�h�J�AI���ҽ2~����M��Ulɜߪ�;�ֶ�m��N��b��/V�vK�95m�[ch�h:뎀���Y&�2��y��I��D�ޜS��(6C�D�wmQ&�[$���I��艓���k%��Rm�&s~�$��Gb"&}|�$��j��'s�ː�L˗D�&��>�a�k�+}'� ���w��_K����D���'��/{��;�6I���{��ba�i�)$��p�$�ē�Rk��U]�T    �-J�YË;�i窅��ݵ^�:�`�m]-�9v��}�U�w
�\.��83��i�*�0"�g�R�*	a]����/��
�����!�`��Nwe$1d�5J�l�9W*vל �j0�3�������K#9�;ݪ����v���I�];NrI�5��6
՚[\��76sS�?�����7�$���ԛ\�T���h���M)n�9���'ӥ}k��5ݕ������?%�RKnS�雞�d��mI���ɼ��>ţYE�@�*Q�I��&�2��y��L�>ZQ$���d��D�wmQ&�[$��D����>�n�gjۚ�ۘ�i�M\�-c�Ҹ)�%9���-A�i���ϪI��D�Z�d��v���gpr�*Jf\�$� �l2!G�Dg|��I;۵D��o�ɽZV˄���D���4I�ݪ>��ߪ�;h"K�>*[�M̳D����Iħz����?A^WŒk}��-8�s2��9��? �'־R����$��}�`�l�[�fI�͈9+A���.x��q��W����J[)Y'�Ak��T�}��@�w�l��Z5��e�R(�ٯ�D��ڠ?y��z`<��|�Ȗ�&g`y�v��c5��@����I0G�$�R�ZSK��6B��~�HO��.��ϝ���L<^Ϊ�,�ژ ��nD�輎A("�
�Y	����7��kTЗ�#Q�e��o�w|��ٳvrIbf��Q���mTJ@p���\��'��Ư�p!���ֵ��2^ި����IC i�%�KՍa�-`�Lm�nle�iZ�baƂ�0)*A��H���*��>��c�\Z˖�����n���F�v�5����w,��|W�_)R}c�,�fٷ֓��ξ������Jx�
�]�zB���8@ɞ!�%�����w�+��rD�KN��x����y�a}1u$��mQ$�\�R��r��$�ۆI�"��Q=#'������d��wi��H��c��������c�iі%�Q���Lכ��t��'יTI���$������⥸A&��D��ꯀ������{D�Z��dؾ����L�3)�'7�$�D���4I��$�`�HL�YR����+�_\W}�ivI8�L�
��4BQ����oǱ�)��n�+�ߋ$��*�7���D��"�Ս��	��]S�lp�OHU���"�gNrq�_��>���l��}�Q&�kd���^ZY'gl,e�(52�o5��3;�"O�qd�u�W��2N��s	J���.�=� I�+,�$�kd�Ň��B�P�xNk���sw�E�����1;�"Mz�-�	9M#D����I?o}_zI���$�+-_�)J�L)���R���t��o>��ֶ�    � :4e��l�˶o:�l�%	��݌<�d0�,BP��il��Z-
�e+n�i�B%v��3p˹�+�LT��Y�K����\��۔�����png&���]�՗�9�=q�GL[��Ј�;�Z�3܄�Iԓu�UUvlfums66��o*#dz{rg�N�cC_gSn��s�mM��=�@���^\~>�'>ߪ�=�'��4�ReD����5k$����d��脎j�̢�Z*Ew��,�뼪<"����N�9$���9J��)�'�N}�z�9��'wړB"�uI����"e�[��9��5$�a��x�d�u��@w9<���U�at�%��-˷�v�'=M9���k̆��%.eˢN��L��}}�� G��ߛ$ರ����D�����Qq�#�1*�or~	ͻ��Q';�d��%�qSa�	4�$��j�;��� L栉.���&�z���L�
):'舟���sV��5�œ�7������y)2&� ʕD��'��D�'��TI���7��i��l&$2kQ���`U"�`t��XM0��v�E"�B����Ƌ$ׯ*�;����I;�"I��S��, �4I��U޶I�A^��L�����$L��i:$�s�sPFDA`253|�q]s��iW���R�IȖ蓶�$�VY&��TO� �z�̛��.%"Ô(��\Y'�^o�I���7�"My{���m�eM�*v8�h��>�|Fz ƶf!��!��͜��	��}�$�l�x��M^��7z��i���N�;��&�Iu�K�k۵]2w4L�&D�fRTI�As^L2M{������r�d6
��Q'׬2Mz򨓹���+�`�D�v��, �.�t�K�%VK�
�@�%PYUDc[�-W}����@��(���$�kd��%��@�NN�}��Uڤ�Q-��m����9�u�0.�1b޲͖������ߔ;��:��?��Ͼ��$�.bT��Ȗ�v�$���I��Uw5�2lNRfJC33齖I���;y-�w� I�-%[�I���'���x�=�TI� �.k��kV�2�$� �tI���9���id�n�T��y�w�o�����      �Zv�+K:VKL&_e�c���n�[<��8�N5WR�j8���Þ���|b�:��:7!�s�j�"�I�:뜄���8�k������d�Z{,��N�v����z(A��E�e�f�v���'S���^�UV(�q��a	6�ux"�r�Z*�a�-�`����݁�`VY'ٹTO=�L��Z5�����$��I�fUw5�NyI;se\4P!�[=�';��I=��'<�$�\Y''l%��*M'D�D=�L����K�Œk�*�',j�%JJY�[�N���\�rO�r�����M�sm����E�:l���XGP�nx��Z�u��3u}kK$��*�s[$�D�KIV�մ8�c�y�{Z����c��oT=����؁�~����=��ߩ�v�G�D�y|$��mQ&��&h�	�iQ'mI����o�v���͒{��k)��eH�'q`,��̪$���z`w�*�赺�	�mO��֞�c����-�ݎB���m�x�q�)�}��t���y���ZY'uM��9"eS��9�TI� �>��2O�r����5k	J�.Y�Ҿ�����n��L���9&X�ȅP�I`K!�}��ZWߵ�M�XqˉH��
'�D�>!�owj�9�$�D�R�U�2��r���ݪ$��d��	̟%��v|u%��W��u�cey^�\^����;ax���9��ѭ�m�n�I� �>���&������'�2&�-5]2{_ "R����oﲨ��k} L�ZѬ�fP!���$�s��̪?DL���'mI=��VR�J[�(�>���u]�s�,���m!V*�IBԀx\�a�$9���v��wZ�2�(4�s�j�;h"Mטd���t}o���ʪŗF.+��Y��QuQ
*���KƮ��������u�݁��`ݱ�쮈����l�pjӮ\JEÔ*�N��T(�{�TI���9�DL���V8.+s��}��t�z�yޘ�X��k�&T9,�)�?	�=L���$�s�����ĝݑ<��4��v�D�ד��׆�;��&EF�`�I$�D
KJAK�B�� �{� ��L���������ܷ�kl�Ƴs��u���*!k��� M�#�Fj�B�E���#ݓ�E+�$,�*HkbG����"D�	��0b��Y�#CW
�3/��2�.sB�Ӛ�&����pu��.I��jA��FT��g���/Y[�Y��)���uy='�iu^��h�6�,���* ă"T�99*,"	cTK��d�vB� ��D0���\܁���Lr���h�3[���ggx�n�'D`���s��w���BQ�*1���J�m
C̅���̪��b��XHBB�u�� ���UTp��                                   9�#A�LR�:���F���J�X�wl��r�۟]�<QIt�t��r9&u����R�A�$�T<N���:ԒϞnkv�1c�+�vb�|��ճ��SGNև� �'vL��6j�a�����cG>Θ������<���<�c�Ė��źnkp�5H�lݤ��&��<m��A����1ڼ$��O$��u3���G#�6ǚ��v]�lqty����]�#��%v�Y�OEλ��X�t�9j�A�y�J#N7��V�J�.�]Vé@b��� ���{�;1� ���U�ǜ۴�s��  �d5��! l����Z9�&S��;Q�:�i ԸW��v���յ&W�nq�6آ��uH3h��.�G$T�;c)��v��F�1m�;�D�� #��v6���4K�zGq:^���x��:�o���|�FN �[���v�����nU�eZv�ks4*��J+Olny**�
�kq '8���=�n�6����m�<��gn[d��7qgl���ۃ�5���&�Nb�ZN�+��i*���x�E�Y����{e�5	� ��i+�1�)�3v]s�n�
���T��hU׈��kmv��NI��M9�Fs���x�
Os���N/Q=��QԪxiai+�x�v���\ !h��3��m��m�    :v�r��;;[B��0�Y�Q۳����:6�:�E�m����ۯl�CӐn��Y�*��۴��;��E�(Ѥj�#XW ��#����5����,Kp� =;�aCeF�vm����9$�%���UU�h#��a,s,�L�8�ZG`M`��.,��L��)��Յ�}��D���T���$��°2�$2�I��$�kd�䠉.��I��	`rD�4�w46I� �.���I7ݵD��;�FJ�S!7D��%Ҳ���*�;��&�,8�Ĥ�B�>���~ ^��Ğ�l��AtE�7ߊ��M[�Yĝ���8�ٗ�i�<�7-��kC��';������k�9&���O���U\�q�ҿw�֞��!$����Yj�w��;�i^��W�h�����D�.��I�ܪ$�kd�����fP-�2(��ZY&�2�����kU2~�'�h��RZ,�S�M�u�{y�Mb��p,������m��"�+��fu��l���s�2�%5�"��R���I���5�"K�ǢT���$����2T�Ȗ��A]+,�[�TI���61`8�ĤYjM}kK$�3*���$9��H)!@d�Y�oي�PD�K	V��2��4O����{y�:�L�z��@����۸�Rz���2O�It��MweQ'"sV��m�enР�@�'Jla�Av!
���{��8��>��A7�"K�e�k�(ԓ���k�2�ʔjdQ'ִ��&roV�{O4�� }������"�߾�u�����J$חI���4d�������W����_�Z��P� ~���eN��m*JdKtI�A]+,�~��]�� ��y⪷M��i�j˺�ؼ˻MK�"M�5i�3����[���ވy�TI���I;h"Myq8�L�.\�D���$�kd�����ƾ��G3�	�n7#v^�}��w��'ܷ�����D�̑<��4%JMQ'uIt��O��TO@����> F�CL�@�T�$�I��w�$��d��%�V&m*      ��fI$̭��A�M@G-]�HЧmMÌ{`%Ԗ�7�/GZn��Q5�ebiQ��ڻg�/kmUvT(!�^����	R�nͮ.nJ�'����r�c��k�1���ৌ��7��h�۬�˒��1���j�6̚��j� ћ6���q��D��Xg��m��TI���9�"K���rvĬL�A�ӢN�I�A]-,��n��N����50�W�>�L�� w��u��I��`��nP�O�id�{2�����wu�I�/m��2�s4I�ݪ$��d��e�k�K$� 	��m��V�,�6��c��ו�<sN�[#a+Z���kr=~	=��&�It��M{v���2D�&evX���]�ˣ� 0H#$	�Ij{yw����i_wٍ�sw�L�R��GޒsI���{��'5I.�բ��K-�$�^�I�ء��o����ߒ�"4ZW:$�kd��'�ύ}}�D�`+9�P��1�jQ��c.���M/W9N@�J����R��j�9�"K�e�kۦ�����hb�qˉH�ТO�id��eQ'7[$� �>���q2��r�}{�D��l��Ώ�9RܜRS��۞�a��2 u���q�Muz�}P:�I�-,�^ݪ$�,��DȚ��sPD�R��5�ڢNn�I��/m��S�kp���AJv�E��f[0�h�&���@ykK$׳*�9��&��I�KV����[4I���`�;�oD�:Q''l]�!4�G=ﾨ����ވ��^��dn-*QR���N��^XY&��TO�  ."N�$�Հ�PE̩&�>���kٕD��l���'�"|��~=�[�ٮ��/R���{|�}At'0k��mN&Q�.Y�&󺨓���o� C�k˲h�x���Cjd�)�'٭�oD�KK��^�5D�̑:��4��Nj��?W�$��U{5�vrލ2��̊$�,,�^̪73�[$� �'nmXNfP,2�I���w5�M���}j�}y���~v�      T�Ɯ���z��t9U�j�hsr�`��;뱎7h��¸@���H�혐�E���W����b�J�f1΀5���=u]��Uq�P�I�샓f�#���Wm�tǈٸa�\����6�-�rrFu쓜�K��v���2��C��;��4�s����Uqe�Bi��|�>P7�"K���D@��M��UOh���JT�rtI�P�.��I�n�w7j�65`:�ĤZ��j��T��=D��l�x�$�ZM�(�r�'�&��I��~�L��@���Ɖ5�@{���7�%���5�ڢnLٝ��H$m�"��t.�Y��j�����&�Z�2�e�,�Û��pQ%Ҳ�5�ڢN�I�,e$Kj�Ю�~s7 YI
*Q;��$2����Ҿ��l���~�����@���4I��$�kg�g5I�.,���%`d�l���_w�d��%���M{憎',n��R�$KtI�ZY&��I�ޚ�N�I�>����bcj\�ԅS;6�h@\�� ̀�=�U��\J	�B�>͗�O�v����d��%��m��F\�`�'׻TI���7�"K���D���$�P��D��l�ye����'뻻�m
Ki�P<2ڍ�2���9O^{u�s�Ѿ�ChnӸX�2������� ��0c��d\�VF	�J7�7C�Bo�*1�̫��@��V��TB<�TÇ"�G�6K�Er�m(���u�%�ʔ\��2�q¥��4B~��Kޏ5u=OuQê��ω>*�j<��]J�p���H�ڶ���0��Wmh�-��C��B�8b�ݕ$lGo8�^�e3)ڙ4=s�����B�R��m�	���XME��tΓiӛ.�cdR'7#��mgnY�;YI��sx����#�\�c���2B&KT>�_���+���{���v0�R�2%���M̏���1ת(_X8�Ġ����v�3|�����D��HJ�&�u)Òr��r�.�KO��x�lo���n�%6b�q�����ߐ}_�g*�3#v��b345��ĉzf�J�p�t\�r�aC��R�75G�u:b���x؝FAa���Ҿ�׋�M��(}�����5�̤Km�B�x�k׏b �j��Tz�+	��}M��|��(���Len	X!e���׈:�1^�tMN���_�u2�d��y�'o��Y�       ��ε׵�,�&��<�����T�7�����D7�\��0��Cq�b�we�b
��c���;k�	L��|�ōɮ��s[H��E���OY��җ���,/-�vz�{�(:�h�#q�Z�kY��$���w{�UX��k��q̈́^��EP�X^��BbKeHM��)�-�o �l�޽�A�k��9q($Ԫ����6�G�Pu:M��&RI�1��c/�y�Q�LW�Ğ
�B�C@���7�f����c�pN# �9Qy�}^Xc��,u�u��*��P�]�3l�Sk�Нؘݎ�ݘ�p��9z���-������6�}^rG�qb%ɱ�2����jÄ��J ֡!���qY�N�}�%h`�(6Z����_��?�����)J2��� ������:�E��qˉ('$�C�:b����(���>��mʆ�M�"���p�e�M9�l&�d��$̙L^��L�^�1������C�%șT:�p��+�^�{vpO# ��iʌ�Aߔv�Y�L����3Vͷ����1 Z��=�Tf_!���H$��D������ÿ��V�, XM��u����P}���}���	�5J;Z��p=.��fn2j��)�u���.P4�)ws�7�^j��5�٨���&R,�n+5p���Yh_s쒞� H�Πuˉ)R�}�
�c�Q��N�m8I�"S�Oһ�߰��\�?YsU@��D?H1���\�.;4������T	 )��^�p(rY
U�Q��]?�u�߾�x~�z����`��+[r�n^� a�]��X����(�-�-9Q��;��w1����چ2���%K��ɘ�^1�1E{PۛV�, Xl����c=�} |"�|�����	X�RT'.P����!����ٿ1���[&L�D�	����DG�7��?w߰����Iܐ��J���*|��}^��ڀ      t�e6�K���/�p��6ڋ��ɠt�zi�^�#m����AIԍ�I��<1�������.�DRD�Ͱڜk֥� �ɢj��͂@�؎�'#nv%�6��.M�q��D�d�b�M8����r_9%�=*��K�b��N;7h"�س�:�^]�l(�-ˉH�Z�����{� � �_!^�'p�2e0:� ~�=�����@W�ğ��%��R���+؃� 7׬W�N�diʏ^�c}��.��p��y�k)�H\��b�x������s�w~UVfd�fSE���}������6���A_PK"Ki��X�b���+�G}�%k%I@���z��� ���U�/׏�" �;[&L���-��J����_�u�=�7	�T>�k/5��!� _!^�'p�32S�9��(��������I�g�z���h֦s��4���חa4玓=-�ڎh7`�ҷw>��P;�G���6�
�����-9Q^�F� 3ײ�����CYL�@��P�Ҁ~�� �5%(&�_gnk��ܮ_-\,p0�
>sy��Q^�cb ��/�=p�̕%Br�P��G��X��z��X'��*�y��8��l�фd�idn���%k��[Bm.=z����kX�b�=�7
T��.��p����c�HQ^ཱྀޟ�Ɯ$̹R�vo1��{�{>1^�t 2�i���@���7�Y�V���.2H!�B>�(y�b��O diʋ� �|c}z�v�G��w[m���e���`U1�t�%��9��a�&R�̥&QsC�8b�x�� }$^|��:� X@�۔c�ϓ�Q��όen	��)�J���+�P{> m^��Ӎ�&XI�Q��όm^���{pn�-Jt=��2�&X�b���� '�wwv���I",��h�r���:8��8Ӫ�vO��&�����=�3���$5[�������a��;5x��h͕���fV��n�;�����/�:���WWP��������C��&��Ȍ�+xN�<�ATG���0�6D�U�N��]�M��Č���D�1�x�Ӡ�o"H	aV	v(�C*B�h.l����.��-�
��.���XƩ������(���      �`�                             u�]γ[���A����h|���W]^�s���X@M�2A�I�pU����l��0���Ƞi8�tW.p�*n�[:��lSU��
¦���hb٣����MC2���X�0��],-]��q ��[���v�-���eR-�q����N�G��u��H���=q�c��������[m�I�*#���)�tF��ml� �1�+�]�*i՟.з[����:�>�����5�@Ӵ�c��`�]��K^�����FYdm#lk֕U5�L����c�'��t��:6Cn׶��� 'T����<*H\J��Y	��
 2�]�.&]��;�ӭki�s��D5��m�
pem�^��7g��T�DZ��M����ղ9����#͋�i�pAƎ�q�eIV�\L�%�V+,ٝ;��wIi.f xgR2�M1M��T�}�h1ql$��L�t(��n���*�y��X���t�=i_\9y�xe�;VR&�n�jU8۶|3�U�88�7,q]��&y­����mƸ�ز��ۭ��M�Z�9��"����B۝gS��yժ9f��7FxEp�k2�@�*x�h�!����e�-�n��rrM�O��rz��;��ؾIG�N�a�3���h:������������k{��ڀ      H-,_&�k?5���p���@�m<�˹�{�ѺW�%�[jeV��s*�wx̆�L�U�w31�8�2�FjK��4J��wLs98���sHk�nt�A�v��C�ڱl��Ͳ��I:M�;f�~מ��@�-�e��u-V&�CcY�4�����^"��i�je�(��c=8b��{>0��$�PҔ��m��P�|IW�����<��,"�i����|F�����~�1�Ĥ
%��N��c}�+m��ar�o�K�P��{>1��X�m��2ԍ5Ff:
A�GP�G��
��Tg���~��Y���ٹ��w��g`�����"[�v_I* Y�A$�nx,;fJ�lo�/��}��p�I�/��?^?�Q{�M�mK��l�>�wP���C� ���*�I�(32�IP��)ߞi��w�~�Τ;/�*�L&��zq�ե5ee[�i�ь��v��0��~���w�~��@�^���CYlJ@�3.��d� =��u�:�h��]̢�K`�:Nw��{���eT�Dc���	��z��������BPM�uꌼA���u��l2�r%8��c��a��~��w���~�x����uZ�ښK��:��cFXsje�Iۅ*K�t6��W�Q���A��6ԸA���W�_�Q٨>�u�'��reȔ�}��75�����X�Bip�/(������'=x� ���~�i �P2M�O��a �����>�0�����8�R��� ���솒����
Aa�}pĂ����|�n��y���74ۨ�b4��f# �RlFc^cn8a�V肐Ro�|�4�R�)�����������&�h�Ne	A4R�1 ��������X}$��_n�AH,5�߲H)�{0i�/�� ���\1 �5��VCl)��	Ja���!�����,��Gt}�.����Ci!���)��}��AH}�������!���ܺ�f[Y�Z ����VCI!��0��X}��d�۾8AH,;؄�<����ޖ����    �6��Gkdb26�LyͩUY;t�-� �E���W���=�t%s��nқ���tl��v�&� ���lPu�oP�`w%YwJ*�j��m��]M�`��1O\��bޫVu�;��p<ۤۦ�%�!1���9�7	��;�Ufdv�"�z�"��CV��.����,h�n��q�M���r���圃 ���pĂ��w�,��[�솒
C}�_YT�-�ʽR����!
H{���
Aa�~���AH~�s$>�BUXp'�_��®�ƳP�AH~��� ���솒
C�=�h��X}��R����Sc�^U� ���d4�R�s)����
�I���)��~���,�2��Ci!��}�R�߲H)r�� ��>�CI<�w��� ���6[n���qr�S*e٣8�v�jz���/(��R���!��)����$���a ��ߺ>̗WNUf�������$��5;!�I��=Y2
C�{0��Xk�7H,��=���fX�c�
Aa���I!�w0��� �L;��H)ܾ�AH,7�|�����]ޡ�����fRu��
C���Rs�H)}�_YUuY�^U�AH,;��Y>�	*}�y�
Aa��8Db׍����g�[m�Ы��f'�7e�v�ؘݗ��aL9v�D�j��>�~1!�o�R��i �s����"JH,=���
C�����.8e�[�
A��;��Ci��;�AH,9߮�Rn�u��������eY����!��� ������ -UY��O�0���%���/��
Aa�s��� �~�����/(��Y����!��.���Xo�}��AC�#'�}� �=���d���j��M���ߜ ��}��AH}��Rw�$�8<�Y���oV�'�r�D�1�2��q�����[�N+}���Ý�솒
C��a ��~�bAH}����|��lƫn�����d�� e$��H)ܾ�AH,7�߲H)��t��U-�5yW�
Aa�}dĂ����|���i �>�s,4v����0���m��6�/�!�g߫D�þ��CI!�w0����X��!�z4���p�AHk���o*�p�ƭ� ��}�CI!�w0��,9߮�R��XAH,?I�~�����tE�q�uܮ��\�N�>|eQ� ���t�5��
C�߳)�;�d4�R�~��Rw�d4�R~�����-Ĭ�R��$��}� ���d4�Rwل?HITAa�߼?fK���Ci!����
Aa�w�CI!��� ���H,��=���f]feh��,9�}��AH{�� �w�$?n��ע
Aa�{��M���&e�H,�=� ��
a]��
CU��)&���CI ��0_�@N@:���/kh     xzN�Rٶ船-<�CC�7�.�-�up:<>#[��9^�@.�F�L;F�S��u��6�L FIG�R���-˭��/��fF�4v��xT���g5�U�:�����vrkO=�z��c�{�����������+Z�l�5κ�9�ˤ9�ă5��Z˲�ʥ����aL�ý�\1 �7�fR�̆�!�}�AH,;��g��*�n����;�a �7��!���}�fRw�$�ݾ�ʺ\3
2� ���d4�R�)�;��
C[�0��X}��W�*��2��Ci!��� ���R�ل��|�솒
A��=�5U����
Aa�}p�AHk}� ���d4�Rw��@���rN���>U[��u��a�ѺU�3��/UݤM��-�R��ׄ�� Ez���� ��~�c �5���e^K3*�4AH,9߾�i>>���܁�B�`q!�}� ���$��VR�/�ٍ]�V^������fR��높
Cu�VY���ׄ�A���J�ʥ�r�D�����M0�
d7\�a ����CI���� ��~���e�Yw�ld�+�Մ�Ý�H)��a�Xs�\1 �>�+;�������W]OOh	��L��.m][��l�^���&�D1� ��~�!����|fY�;��
CU��)����zܢ��[k5����0��Xs��bAHj��a ��>�!���{ϟ�UXbff�,:W=�CI!��5SO���]ݷr�R��$"�Y���@��DM{ρ>.A����F�	s'�����"Q
g �;a"��8MwÐ~K��^]�2w�׬`n���D���`�<m�h��!)�T�6fsz&� N9듞�'n�8plj�p�ҫ5x�I䐨.o~硰���N$C�����VI�b��ŭX��,��1�$�HP=A3F�_�l �����5,�@��	��#Va�4����X��w!,w�I�T�;	 �3���ؘ���w^��t�W*�䦻��ͶO%=@�=*x����^U>T�
�z�d����
Aa��x}�.�����Ci!���H)���^CI���� �?� 4���pĂ��/����R𪼧D�0�~2H<��fY�;��
C[��9r']�����"����!c��ݫ�pN�bD�6�h楷A��q�;u��9r}���@�Xs��CI!�_���JH,;���i�R{�YT�n^U肐Xw߮�R���
Aa�}������>�2 ���̶%���1�w���q�$��!���~ｭR��$��}�6e].�X肐Xs�}��AH{�� ��
a]������(�-&D��A�~l��1� ��t���*�2��Ci!��fCl) ��}pĂ��/�)��߫!����I{������Vin�ķ�t�*CE-tv�r�l�)yj1aUX`���
A�C��7$��|p��Xo��`~�� �?{��
Aa�߼?fK��*��M��;����2�w�$��}� ���$�ͷ��e䡼.�Rw�H,1���a ��~�c �5��� ��=���ĪĻ�Ci!��� ���R���0��×��$A�:W�U.Z��f�)�|}pĂ���R��H)���
Aa�$.zI]Y">y�|����{P      	3V̱�����{*ݱl�R�ZMr��mKN���C٭�����:���&�k�ۆ�	q۵��rfy�v��vy�u��>K��E'��t`�y^!����pkF�<q��S��I9��I�rI;�/}��3�[͉�� �zm�i�%"��Cf`�n6�,�C%��OI���w� ���}��AH}�fR���G�9)9>�>&����S�'"Ý���i�R�)����
C[��!�
����|W��e�mf�������� ��}p��Jd7��� ��?~�i ����0j��3/D�����`�R���
Aa���CI!�}�AH,4w&UӕY�m �9��0��Xk�����
H}�,��}��!�_Ǻ ,㗮˓��bK�;v\ƽ<��=��7�b�1�8{>�a4�R�)����
C[���R���ً�Cw�m �{��8l��H֓�K���8f6��N��P��|0�
a�e�!���R���i �s�}eR�n^U�$}�n�)!��� ���d4�Rw�a ���{¬�ʪ�Ci!���a�F�}��A����AH,>���$C��{��WK�eV: ���d4�Y!��0��X}�\1 �5�~� �� �?~��33Le�b��TjP��0��S���������C��0����� ���d��|p��Xk|�4�Ry��0j�L��R���!�_,��{��$�����B)������ɗtVy���
C��&H)���d4���z���TPYOB��BH��8����ֈ)�z�!�Yιy(�
��R
Aa�{�CI!���� ���\1 �7˾URo���G.���6�R{ﵢ
AO�O߿\4�P�����������'D�?Y�_���UX�LV�9,��/79[f��N6m�f�i]-jΧ N@����R��0��Xo}��AH}�{Z ������v��֡� �;����[�H)��kD���}p�Hk���fU�u�e-c�
Aa�}�d4�RｭR��\1 �7�������nQeٔ�jH)���� ���\1 �7����Q�H.�rMm�o>�i �y��0j��2�4AH,>��H,����\ ����$����� ����~�ߪ��J�(��	�e���-���2B��^z�KUyE��q �=��� ���솒
C�}�h?B	) ����H)v����KE�R��R��솒
C����
Aa߾�bAHo��~�*�,7߼?��F�,ʽCi!��ߵ�
Aa߾�`�R���
Aa�}�CI �+�*�.9yY� ���$��|p��Xk�}��@��v�@$@&���s)���$�}~p��Xk��CI!�}�h��Xw��X|���C�TI/'9��p9�;�k]������    �ݴY�c�1��l��XY�rjJ��i���F���LBTCS6�l�KW����F��k8�I���b��)P��\C7��[��-�:�4GQ���\�(ˎ��F���lQx5�p�v
̦�ˢ��XzHp����+wڪ����)mG�:�N�6�P�Ό"��ݛ����Z�Bm�X�X{����AH{���AH,;��$��|p��X}ϼW��,�2��P�AH}�ֈ)�~���R���
Aa���CI!�~��̍Ud�2�D�ÿ}�CI!��\ ��>�i �>ｭR���ٓ.겫+P�AHw��)���d4�Rw�ֈ)�}��
C|��r�Qxe�cZ!I�;��$���� �ﾸbAHo��	r'S�?}�� ���#:�N��V��:������v�U���]^���$>��kD�þ�ጂ��/�C�) ����CI �+�*�-���� �ﾸc��g�gd�]�"1�P *2�:@�����N�3[^c���5��ӖU����6�^j��D�2�={�e�8��(��[�q!��-P��qy�>�ǫu�79����ޙ̰\`l�����VmGm0�lXZ�Q���=ҏ�1^����,m���2�\г�1^�co1�o5T�YiĄ���ǯu���x���c�@�L�i��{S7�/JP�rT77\^j}����8��<��-��D^r7s��6�psysm��k�)��bM�eû��"h\8�!�k>wf+׌u�?�f���)%��Y�_sy����1��'rH9-P��qy��z|cպ�����3-[L|{������aޠ@�Lu��"Y�4j.]8���iQ��=�=70kp�r�Jr�U������ݗ���7m��H�іч*D���ŵ�9�WQN9�08�a!�Ӊ	�)�"O���^c����/'z�С�R��ٺ�@#��z�������&Ia����z��z���޸�ɜ[.P�	��p�����k�}CD�Cޜ��i	%�s,��s�" ����Q��?������UU	"���i*I�?o�:\���?��"J��U�������a�64v�$���Th���2����b�=*��3)GT��V�Vh�v����KZE�T�x�u):�\���J�d�6�����\�b��5�eQ�8ܤ�63V����eGƧL�Q�(�UE.� ��%O�+�o?����o
�������Q�r�)���ߜ��Ϝ���������H����eG�a�~��O�f��(��xK����GP�Wr�o���
�^���	_��#v�������������򊢨�*���Ȩ�*����*����*�EQTUEQTU$�8x���|���
F�>1����y���!zu���y����<>>TR)����?�?�_�������'ߢS��)?�u.?w�������/k�M�NO��G�5*�_��_���|��G�
��y�~�×�~{޸��گ�~��?Uu�����������k�����������o���qͫW���_��L���Eɶ�f�ڨmIfh�6[#d6��d�m
�؅���9)9j-�m�M�m+`����� �&j��M�Lԛ*6F�[%6%�ShKa&ʩ�F�-�6�h�V�j[&�մl&al&bT6�&�S5E�SdL�m+2�Ű�[Jf�bl��0[I��I��d�!��1�Zed��mV�ڑ��K4��5�KYLɭ3�i��m1�������f��2&d�fP֩f���mn�8���)�VjM���Z¶�[D�Y6/��j�f�������Y�3A�͚ٚk1�flf�mci�fkV�ʙ�4-�Kh�2�ղ��fJ�P��UR��F�Ҩ��Q�!��IK�{�I�������0�c���	�����T�$�8_҅u���_���>w���������<��7�t��;��������H���p����A������?M�ϳ��˵_��?�߳���]��}��~ߖ�+��g�v��H�����V>�?g�~e��~Ϸ���}����&��AE?-�HR)����,�w~�?Ss�������e����������)�o�ٞ�������V�J���������߹׏?ܡ[�(��jU?ׇ�x=N�~�uw_����x
E;p����*�`�S����?�3��*%{�g�������N���u�N��_��������9�ﶇ�9?o�?��`�S���ޣ��~��"��+�s�_��_���}>O��O��}S�<N��t��_�������1���_���=x�I�O]��Ο��)��}_7{���;������ߣ�����|J>5*���w_����n����O��a�H���c������8?
������}�K��ó�;��w�>9_g��?~�7R�l��ױ���]��BA�\ȴ