BZh91AY&SY�4���_�pp��b� ����af? �
  $   J@ 	 �  � 
     >�h _�(�� ( %D��QJ �QT@ J���	(�� ��D $@UB�(PT�
%G    `    @�14 s�N����m|�ŕӗ*X �,�u.mJd�vܚS 
X�g�g�  �q�$N��@���6�J����&� �M\�4��J7TgjWM��   �@
P{�Um\�|�y{�6��w��/uf����/s�{���w��o�-�fܻ��w� gU{sn�r�� ;��^�w�j�  �u�[֗.{s�n����U� ;�,�UX�u[��-ǹK� 8�  �  �` '�}ŹK�]7�.��#� ܩbݫ9n՗7\��t�\ ==�K��;��\�^��6��ۀ ��m˺isj���)�˞�\���qn��,���]9wj�� �� 
   D  >z��;��͗T�ݵ�y���� m�nN��Z�wO,�mŕ, �-qn��ܻ� 7O/v�wyokj� ;rӗv�nv�/W�xչ��y����ڗ����i嫛�y�7�V� �P  �  *� 4��P���{���כK��w{j}� ����->����O&������p rW-٭ͥ� e��}��x��� ������uv������n N�&[�ܷ��Zr���ǹS�      ���F��UJ@�  ���P&ʥR� &�@ ��S��R��      =��Hڊ)�  �� D�	&ʔ�� �   R%HA15=&S�d�=C4���~�؟"~������W����ۇ���:��u��U}_� ���UUO���X�
���b *���,QUu���@U]���AUo���/����'!?�t��1,̢L��a��2�s�-?�6Z�_ڜ;��h#�u����*���=އIBS��XH) (L�%)Ԇ�B�)t�N`QQ��:�R��-!�rLc!)6���\s``&�P`�b�lnw@��NA��%	�N�@a��Pf.:�0�-��4A���X�l��k ��AS��	��`h�A���*9QrP�M!���2��9uۅ&n�#Q��vkHk��w����W�����qA��[��������Edk��Xtxp7AY��tH`@@k,ܚ���o͜�F���ݵ��I�faC����ӀNhՖ�Q�]o����.�8�
��خ+%ЪQ�8���y)\��`����9�]p����J�KBjj5��=59��N$w��2"�����Ǝ���]l���ry�Hft;A�����re��z�ѐd8������ԙf7zz�mλ���ﾎ����;1���Y��ރ3a:$��3X�wû���s\:N��:��3N#58�����kX�u!�kXhtjX����vt��u��Ӓc�T=<���(KPo.s-]o'V�v�hd=C���sX�#2�f�Ck ё��R��a��8K�	̓�ѽ��R�`jq�C�F�5�a���sq��aNEι�5�v�fh۠΃X�nY��e�f�����yq0%9�r�1�����:�6�a��0�гy��Hʢ�B	Ԋ�+-�S8QN�|2]_Q~}�WDU�N���TR��i�d`!�3�!��)X�M)�`��dc�K��"1��D4��޹u�Q��ל�F�o�7�0�j04�����:����:�Z�-gG�Z�^��"��:˷�g|�,d��	�:H��o�r3~i�I�[;��k�!���,x;��䦙rl���P�%A3�bT��uQ�2]Fc��kA�O ���II�λ���^A��V�.�Rn�Z����f��Ĺ8�j0��3ak@h�o�|�f�ε��##x�|��FX飑��c�NK�X���F��:t��;7&��MA���2��ڐQ�oY=��	X�A��BW���p�f	Ar��g{�ֺ�8�gi����;����Nd��4V�35�z|\��P�,ћ��Ը�8:�8b����BP�ε2d% by�P���M[����-BS�6A�@F��=Iy�7�sYÉ��z<�F��X��k0�W!+|�e9f��;�I��9`�=�k�A�tC����.�L<5kY����N�m՜R�Բ��ϻ.OE:v�#����W�r.�B/��2�W�)V6�0Ѣb
��0a�3�}]�u�;��:��'ں���UÔ��8�w���^��)r���Q*�x⩎bbd;NcT3�g[띝a��P\�}���4h�m	CJ'&	�3����s���]�pԔtDFBP����Ms���f�tU�oy�k'��[�7߽ٜC:{H�2���j�\����z�\<���w��341�0c1q�[6C��l���M�9�%c��X�3R�`�r0)�Mâ2� �b5j��i'Z�{���p�acQ��Q���O�+���C���N**Ep�o�.�֠�Nk5�s��˓��㑌�`㱆�����]˅���5��������(՚ �P`�DBPh��0p��LL�,{�¯;3Gy��`Ų;��E:󨺌��l�w�nIQDh��3��ќ= *��1��f�=y����o��j�������Pi7�|�:v�@u.98��n�������f��f�:�.����ְp��9����4�$kA��Gf��1g(��]��}��N	²��ʬE���Ӌ��P�
T0/�ڦ�\�j����49`Pd:�[�޺Д�NI�du4��Z���Z�K�͐m�%	�L�I�Y	Bj6K�5���J��)����0yj͚�癿z��Y�������($ �� �<���M='G7�h۬4tM�F:�
5��g.�fgn�)
n�SP]L�ꔦ��lU��O}ԝi�㓣|��o�k�.8�e&�f���0l�C�a����9F�:���&�49	F����[v��5����;�M�̐�YAX������F�;�Fu�es��Ө�4��r�c��2��S�7�f�c�ui ��9�L�
��n�P��!��4}B|�e���p��58�ٽa�6��m�`ᓆc�f�2<z���3�S��jN�6d%���J��0r1l����K��δa$f`�
%WCD�L���рd1��2�*CYdI��5VDYo0��A0ӄ0J�H����+�qVX�I���\�\���<2��j��Ԙ�� �Hg$�g]I;� ��L��kǸ�cjBn�A�蓚͘5a��l�Q�g�h��j�rr'F!��1Gpa:�����`m�0��sA�h��N,A�20 �p20��{,�'Hu� ����
4N=F'9щo�Ӯ��=y�����-9Qa��F�,"2mE��f8m5��# �Y:Lz�q�hJyѸ1���cY�5�8i�jc��Cs���d%��K105��� ��Q�VW/�}O�ݺq.+�#(���~Rʶ|鳀_e�;�����y�]���.��֎�X��:H�3i��S9kZ!���L3+gE�\��;~�®"���l�q&�Or��h��]�?8�s���V�����T�4rݳ]W6s9��E�l(30ѱ��tkoAcL�cA�,H2���!��A��2r�#Kf���[�$r4�&C!����$�$�9M;j͖�Y�	u�\��z.�S�`b��C$�<�:$�2ō�͖��#3!�e=��\ga�:�\��YӃOD���mѦ3�6���G00rqr0���޻xvo�G�έ�i�$L�!�"���7��@���U�i��3m�{=9�il��J21'�Y�㑉���6�I�)�*NUNy�o�;K����Q�34s�ӨrL�$;�%.�$���麂u��G)�s��Cӭ���M�5	BP�Bw�%L�:�Y�r{�o͜�=6w�m�e�蓐�&1�pz�
��HCN��IT�F=7Z�)5Ō"��)�v���fη��#�c��ӥ�4j��3V����o�<�a��˚���9��9Ga���hd%.VI��d�5c��'r��Y�8ڃCBP�J�+�ò<f�q�ގ�vy��s:�3�c98���[LL��)�$	{3(d�f�;��g�8��M5ٸ�Nˮc��J2H�,m�F�1NA%3y&1��,ԇ!2�ݘ�xxo�j��ճ]lͤ�Gz�F�r8�D�P`l�Ȥ�'s���Ç{��^w�����=5bEn0�2��C-�F@e�8=XJ�"��I�Ō�)�p�̘���%۽�4�����e�5j-BX	F�`�%:!)v���D��'��L�BQ�1@a����!;�N��Q���ܙ�h�G��Ӱ�:'y�J7Dhի{Kre>��	@o��f��Z�uk�k^�۸�::�g}A�cQ�:�	BV�ޥ�-''Q���l�x���s��=��XL��HD�8Ҏ��a�R�bYj4��r2Lc/XrF`��Xi(�3A���-A�h�9�(rC:��FN��	Bn��){7��0����BR�<�LYib섬%�3�{�b2[��z1*�dEhՆ�C��\l�kfs'��c�hц���2�l#F��h���f����ӣF8F�e����g�� �K=���BX��6up���xa%����@e�t:�'���F;ML�kQ���h ֧p�f�ǾrL�����p�ê<v��f.��:\� ��[������&���;�a��w�5�G|y��]��z�,���i;�.�='{���!�q*���\8�I�u�Y_�O���E���۷l�w����7��NF�V9�-&�'
s����#V.ø �U\J���󫢊�B*T��B�o��5�:��:`��F��0ӷwN��µ=$di�� 32�8R�I�=�o3#���љ���'��۷m��z�<s�mс�8:�l��zth��i�h�soA��;i��&��Y�kK�ۖ���S�)BQ��](W�u|��(�j2�!��JNDd �u9.)��h�#,&s30-o�:�͞O���2MDn�1�J�e&���9�C�����f�#����4Y:ͻ�:-!�e:�!+L���w	BW5��ӿ3�[���(ܹ	���A���D��y� 2�4j�n��ѳvum���hլ2��,:-0�X�70��გtNF��C��9�����P7	HfXÐ{Ue�nLL��
�j��s����9������.��$�I$��k� H    [tQ���  ���   ݶt���V;;n��K/&I-��� -���$9ͮ��$�|�R��a�n��(��j!v㝕YV�gʇ�_w���O-�jڐ�f�8�M\)1�L��_[ymOmU��AB��� �+�6���� H��\*��(�*�d�+�s����d�ڮ��l;i6������Hٵ� 8I,��e���WU��g+r���n�d���,���UZ6 *���e%��� �  l�s,�
�^j�+�`�4�Ut��UU+j��:��U�\CTT��[W,J����H�6��v��%�$��@hgHbڶ�(UU@UuP&«*�r�e��F+<�Gn����	vp�`�햅�  ky� l�q'[&�vݛv	@  k�m�� 6�;m��pZv���� [u��/�o��m� p2 �U��ٶ ֳm�ejU����yj�V��&�M���M���5� $�  �6غl� 9�Vm�m��˦�m,M�.9����YGI�vղYVгE�ko�Z�`` �l �f�lp�Ͷ8m�a��m"$Tm�'4i��݆� lֻ�fa����i �6�  ඒv, m��l �b�-��l-�6�N�X�(�� ��d�-��l��%��X6�l  �֟m�(��S�j�&�UmUP [�9oM-�z��J�6�[Kl,��Z@���m�� m&�:�$�����V�k��^@�ڹ�h��P2TUJ�UX��Wrr�Um6
%�{tK%'G:��*�m\�K�mtS`����`mm�$�� mi$��'b�6�g���NL��N$��l�5�dٓ3<�;M���{U�[p$A�l�  /ZP�%�$�5�rD\.aN���n��4Y����Wf�`��U�W*@�%��E�� ԫ ;T	����h(�ܷ[�.�!!�m���9mh�rt � �`-��:BG-� ���ꪬ$-�TY�]ŞL&�Uպ��o0H�[�5�� ��` �sZ�Z�kh����+�*Ձ�kP�Ķ�j��k�
�lhT�)A�ӨНEV�*�1;+U`�;��J�UU 5�5��h�k�+[���*�5Q�]2�σ��YV�x�V�S$��6�&�6��u���P�m��a 6�`6�tn� m��lڥڝlU���Ů�e@��,փ[Z�/ש�u��p6ِ��l�m�qm si6=o{��W@RC�v��Hn(6� ���V�h6݀ ֶ��Cl�Ԡ �#���3
κW4�Q�[��e��� 6�m�    �l'M���u��m�m�!&�t���x6�$�H ۶ ZlX`��k4Q�rl2	6�-R����P�r�l�Ut �qz�d��j���Š@h�l -u��v�����\ �  8ٶ-��$�Cjٶ���	@ ���nm&m���k���m�^P��mq�@	 ����%�)�@[J��lm�݄��e�o� �$2�UR�T�������⇘bv�yZ�V��uH�<I;��'Xٻ[�O@�m��q�j�r �	�q��Y�jc' ��9Uj���媮��Uk�@2J��֏����"�誀�ݰ��ʭ���2KZx%We2�uU�z��Mm H H �8�'U��󗪪Biy�$	U�Z�� g�һ��_Z�9`���u9�i*niWm�HR���fE� צ���k���l[%��M��ppk������n�r��ld�m��p�����ճ�~'�����h  v��  �l��`�R�6�[E� R�D��I��� 4W �f�� �  i�Ɗ��p:@ �b�G	 ��.�V�6Sf�p[C"�o�����6��ŲP $$Z�{l(��ε�  �pkX2 R��m�*��(<8+�Z*�R�U��� �m�M�,�Bu^���vav�d�6u��"O���o��/K*�U*���UJ�VU�]R� < gV�Ϋz�"G��k�6��xb����W�8�n�]���$ �2�ii&u����*����m�^<�����d��/iv�k�v�I\'-2�j^�m���U��jN��Ԡ[Z��%��G��Z��mm�H	5�U�H:N�0$�����GV�˭[�m�%��Vm�M+n��Ę���Jl�3��ڇ]uŭ&Z���`*U���m+դ[� r�ŵ%��M1��@U������R�  }��-6kZ��� -1n���ٖ�p�-�-v��Γ^��`��5��lふl��[�t���{`��mM�w�`�j��Ӵ�:�,����حB�[�"�2 m�[@$m� �ol2�W*ԫW[)-J�i3��lڶ	�1��[\�9�$Zi� u�Ah 		k�ר�vHkn� �[vٵnĒI���'@/Z -�q%������k����u!Oھ�vZ�^��` ^�RX`6��k�G5����I�lH��Ո=�Byݗ���[U*�T���m�Uʻ�V݆  �cl���m���mw]6v����A���p	j@pvC}�m�Ay`*��P%G��UR��`� �m��i5�˷��Căm����UT 	�j�VUU��m@�H% �`t�TJ�6t�6݀M�$��ڴ�  ��\,5��e���6ݶ���m� [m� ��#uݛgm����C;` �km��`�p����z���VH n��^�\H����  ���a��u����ݳl��hH l�� �^l�˷l-�m� m��m���6��n����`�^g��Hà�@���J[���Q��Ym � �C���� �		e�ݶ &�q�ն 8 $  	�� 	mm�-�� l�� H���vZ��G*�AØV�NݦY[�*�UU�\�*�n�9j��/5�� n����]6A&�6���$���#�6ؐ@ 	m�	� � �8�6�ܐmI �Y*�(Ѫej�
��U�ڋjE�4���l	 ��� L�	�3V�J�$.Ƞ;e   ��A'�t�=i�[v�Ԃ�P
l-E+<�n���`F�I �H�  6��8�ж�    �bGN�[dpm� ���m�z��   -�m� ! =� m�gAm��i8p���� 	�  	 m�h��[u��f�cs8[[l�m[!�m��� �`�-�n�2�Iz�MU��^Ԡtgk�h���]�VT�L &�pV4�P�`���퀐���9�q#�jK�����$��٤��`pm�2�  $m�  m��M�[Ki6��� ;Z��H-�mmnkp  6�[@~�x -�m  �� R�j�eZU�+���A��8[@�� l��`�b�඀   �6�-��nm٤׭�0�-����P i-bČ,K��E����.M�i�9I:��P	��Ŵ ��o;�iͶ 88m��֛lH����z��I�,�Ӎ���J�捚Kn�  ۦ�\ Ӏ i,�P�Y�
�mTHI��2����)ݴK#��IK@6�rF�[�8�UU@olbG2��ځ��m�Gti��sft�Ғp/Tb�]�tʻ[UuG�` ݶj�4��m_>h�ց�ͳlt�ݴ�d�Im  �[d�i��m��EJ�Ir�2���� @۴�    kY���Hp  m��m� �f��h ��A�� �n�Hl� ڶ  �`p   m� ��Ŵ �� �mm� ϠŢ��e�BҵV�U   � �@h v��m  ���k��  ��]t�:MSe�֎�َ����[Aɑl�j ~�`�a�l��-��H�`5���@�i; �] � 6�8m��H�� !ZRq'ʰUUr�ls�� �@��*�@R��%^���W2��J��U/,�2�0  $   ��*����j�T��m�8!' ��Zpm�/ku�%�� e�m�6�H���]WA'pmT�~<s�jB�`HN���ռ����v�n�n�l   ѭ��pn­UT����kavn��C6�� ���G  8�p		 �$s[#m�[m���+��3U@UUR�1giXr�U�@WP
���6�"l�E�u�l������8��V�E��%k[k ��-��&�H�P  [@ �$�dV�����淼޷o4Z�R�
���W}��1����?���_��"����?����B��!^��	Tz�4*��_؂
8��x�U[�B�x u������	:?��l���X/�@��P�H���)vS�=*��;P��׀(ly�z�� �F�z�T"Vd�&U�:*�x2��"#ત��;@�x�����U� '����N��
@��t�h:<B@ P�x�j��BK�@U�}@N	ؾ� �8'�
/G�A��
pP@x������"b(��vih@���"�/���<������}�Te�Te��"���S�����������h���Q�=�AWa�}$�"����v�QU�h�Ą$2b�8ؘ#�+$�M$�	 0H��)PRH��5%%a!4Q��.1�b`�D� ���؈mp{š�����A�T6s�B'H*���	��"�u�
 bL�E{TҚA��P@U_�?�������?��.(K#�@� c)110�L��^�{w�?�?����򦓊����M�j�[t�{MO-�L��Cb��m[�oT�&:��4�d{";-u�5<��me�vnsy��{;�s`�Z^v�:r�	5�D�'2�3���Ci�%g��3:���Q���b�� V�$�kF�MIΒ�V�����k�!��m\�/CÃ)X�շi+��&��t�.����mV�]a�z^=ZJ�6���[`W8���t�!d�HV籨7ZcJv�v�=g�h�tX��UU^1q���v�e^�Վ��`���N;rq������mj�eҹ�*��]R.�吚�̕0�21[;*�L�$j�[FKa�s:GgH�Hcr��n2v;Z� �x��g/�K+���j\v�k��� U�gF�HL:�պM:-���M��\��ⴋ�TlR�l��eW�`��t��Yg�FJ:B%C�ڳ3c
�C�oO�����7*�����1i�5.SV�b�BM�L�Q+=ܙ�mmg	�Mt���(r��:NV�V �&��S��;�[�j
X�ѵ��=�-���+n�e��:X�2R*����Eڠx���Ү�ԥT��8�(��g+���+�Z�̄��E�6����RZ7`�E0\���М(T�$��k@9�۰!-Z�Ȇ�9e�vC�;D�QI�{Sl�v���lx8٨j��iܹˍ
�Q�G�R��'�NnQ�k��إm*��qFg@[S��N������G��d�r�`mnJ݌v�8�۶��"$[ti���kYH&�"Je�8����j:ه��VQ���l��㮎�9�ۮy�lѥދ'�Y)�4z�[%��'f�[
�2�N�ȐP�)�,)M\:��@�(�l ڷj�"�ˬ�m��I�Ҩ��Ѱ��٩��U��`�K����ڣhD:[d��Gd,`�\WPQZ�%ʄ��n1=�)�h�f�]����I8���[���ո��n�Z���^�'+�	�%VRM�������t�t ; OP�P��_�پ�{Sj8������j�<ٲ-�0��ef��-�ݭ�.�1E��J�S���7A�\��a���j��ۦ�#"�^�]'7HG]n�[.*�7�^%�d��x#^�{sҖ�k������v����9���Ir�Ϋ0v��;<����0S�֓,g��-�0����cj�fpZÞ��r��1OcM���0�\�2�od�݃i�c��e:�	t�de_����������\q�6����n{���ό����N�Ea��A��N�e��{�ИX��w��+���`uz�U���(P���/r��IN �ܫ �+F o
�IEJi��,�����c�>�L,>�K�x��K�V��T����r�ܭ ���u%8��L�CX&�n��>�L,>�K�<�`b�����P��t�r%JS��!Ύ�X�Ӧ��:2][F��gv��8wg�u�٠�(*T�B�3�d�>��V/�����0�{n��$���Ȣ�t��ú�Ȋ��":ps�u�/���,�e/s$$��TH9!`b��X�Z0{���h�:,���mSn!��>�L/y\�r��l�=�4�ڮW�f�啢֨��iB�TUـܯ �+F �ܫ �+F���L��*�RNTe:�!����eس�m%Nz�[��ꭞkxBr ��x��q�T�5wx�Z0>�X�Z0{����.5@�EHӅ���c�>�`�+�=�юd�*A�,���#Z-�z�^{���U�~{�@bL$� ��"9�{�nU����]�Z��1EB�ʒHX��,��������0���m�x㑥J9RKܭ*�8�Z0�+�:c��h�U�����x�G�9�k�<�5g�������OOf����U��5l�r�ܭ˕��h�:,��#I�m�I$V�Ʌ�A��,f�,c�+�ՂJR4�Clwf r�x�Z0q)�s�rv� ��ʖ:(��*���X{&����]����^ 	Ԡ(׾{�Aܯ�� ���#N�����a`�d�>�L,���"��Bt�u�Oh�Gj�xs�m�u�v.��Mv�Y��L`\;��6�c@�)A��m�E`}�X.W�{�� �\� �qRt��&	��.���\� �+FʹN�S��/y$�<q�ڨԕ���za�r�S���y;f &���Q=�.HD((ܐ�=�ج�� �{%���a`z�2�8��q��9$V�V�Ħ���� J�NQ��;��a߼V88�l��;��׎�v�Î
�b� �)����s{#l�r�*�g�:��8�pt t���ʯ+\k1S���<�EB�P��r$��{]'+j@6��;[��Fm���<s��'>�v�jru�W<&"얺w,�.l�\��@ݞS�p:6.3�a�ݜ�K�� ���[����;T*e'fQ�N����R�A[o){/����{����{�[]�n���Ie����~'�>��]�l�WI�b+�ӹ�q�+qnz�Gj�*��m��V�*�8�Z0���,tQQJU)�%$�>�L/�U)�� �� �+���S �]�՘U�pr�`I^�S�i!,���(E7MH�5{6��ӼܭU�p�N�WSeA0U��ݘ �W�{�� J��ݓy\�y�ؔ�	�C�)�o,�s��<��"��.�9kR]v�r<�.M��NH�*�8G$�͚X��X{&��,�e/s$$��Q(Ԑ�=���s�Ѣ� E�7Y��ە^���Ʌ�8����G�n"G,�9;f %��r�`	u� ��Rƨ��dj�lr��R[����;f �r�ܭ�PA72L���V�*�8�Z0.W`b���
N�R6�ED �*�X�u�=;���M�κ�;2��`�Wupf�����\�pE�MY�%\� �+F %��{&q��gr�StԊ���0��^�V�J�Xw�'+��t*���3=����0��\�ʤbɎ���1X��'Om�Pp�]��h��U�{�)��^�K��	$"JHX������f{%���a`{ï2�TۍDG$WB�x���{��^:�<�h�� 57/V��tl��dLN1������1Xg�X{&,�;��ƨ��dj�l�s�	r�ܭ�ʰu%8���,tQR1T�������0�1g���Jp.W���O�0A%�\i��Ş�`}瘬3�,9˪�TB$/����ەvw��u����$UAWu�{�)�}������ Ş�`}���N�p�uM�B�<�<h��y3'n^{cӵ��I��l��5�=�:T�E`��`}�X��������Btc��JN�,���J�X�Z0.W�z%D���!�AI{���a`��`}�X�̸HМ��CrG`}�h��U�{�� R�V��Ss0JQJ�&��,Y�v�W*�^ͽ:��v�Ʌ�|�9�Y_z�!���{�v�쳝���m8������n3��T����ɑ�v(˸�"V�ݚ(3�[u�ܤ
db��b�ew����Ճ�e��b�ј�-���}�����!h��ۣp��rr��wC��m:6y%1�!&��Q[m�n��58B�S�B2l��4���
��Kbçj�-��v�ն��pݕ���\��������*�%BP���W
�N�W�Q��$��V�܊rι���t���b�a����«A����ܧ�EH�R�I)��饁��V R�VȎG�0A&I]�՘��#�)O�.Y�H�! ��
�n	"�
���JS�K�G�R>Iv]{�H�<J:Dt���������������f.^{ԓ�$m�P�K���w{�G�R��.Y�5?)"�`��n��@����zx&�Nм�x��;(lݗ����j�St�$��$������,����]}�xs�Ͻ� ��i�6ܺ��1v
m�	<*{�H a3K�BA!C)B�H���V���I���&�6 ��F��p��5���~{ÿ<���Q)E*4�d�r�=�_{���]}嘹��b�T�U)�����cÞ��˯��/3�u�+Յ5E��EHӇ=ｙ�J~Ĺd{�#����&S�������EM�e�vB�[Y;7���#�Ε�R�Sc�v��ur�=�_{��{.��$z��(":JT�C���u}�#�����e`�"
�jf��\��n����[�=�_O�w�S�e:���A%�i��d��HR�)�j23F�ͱ�G�LW{|mtJnw�2".�6:y�'�h�R�h&CG�: ��%,	TJL�d�%D����L���Z�L;���j�!�	d���*h�"��1����̢#tBSD��I.��7����d4z�78�M"p	s��:sL NX�"A/Z����("�RQ��X��P*

���J`�(J��%�P�3HҖ��49!�1-�^Yj��]�BC�mNŕ=s��]�Hm�7��p��f�" `�<�!I��%-*:M�? ;�;�P=�T��ä�|UAPյ� 6���*��� 	�����┥'_{�uΜ�9^����!$�B)I�*� )=�<��R������)JRu�����R�|���qJR���>� RN1����uΜ�9^͚_9D�*��_y���)O=�\R��V|���9�r�)ң[\BC[|��v�]�n|�Y���b��9M99mN&����:�_{���q�1�k��A���m�v�������R��߷��)JO{�=�J/S"��A�i�sJP��%qVffo|�)O=�\E�)=�<��R������)JR|wy����	ZS�~���e̍���5��R���}��Y�!{؄��c�"D/c�;�!+M��N�x�j�7�hz���~���):��~��)Jy����$�'�e1E�p�W$@�L� 0��JO�ϻ���R����Y�Y�0�[���|R���]�����(N�Pq}�����{�����G�݀q�x�����bK1�Ƕ �w3֛q�4�c���+Ы�Ʈp�}��z�|�v��k{�o|Ҕ�����)JR{�y���)O=��qiJN��߸=JR�qm,��I$I qI�(9�V|����P�<���)JN��߸=JR�{�����  2R�����o+5�,�����fs[懩J����)I��~���QPiO=�\R�����ߵ\��Ps��dU�$JQJQ6���P):��~��)Jy���┥'�����R��~��R������4aެ6k337�R������)JQ�C�3߿h{��=���p?!.L ���ި�!B�z�w���Us��3\��]\݂C �tp��Y�qu&�N9���M�&(�v䰶�1ո�*볣nv�s'Px=9�G;a���9]m��ݞ���<���(�ۇ]1�*2m�W	"ԩ�ia�����nر�L�4u����<܁f��i�ps��.lq�\�6��`�ѥ\�:1��/�&��n��wDv�Ok��;^����-���۔דW;M��������Nxa�wj��bB���rm�����Rn'�\�:�����瞮?]��{l��H��{��'�g�~��)Jy���┥'_y��JȄ���� �A
�4J�Y��֭�|懩JS�~��)JN���E�":�=�A�}>�J,IPs��SB�Z�t��Q�I�(9�}�pz��=�^��R��Q��>�={J,�A��i؄!6䜒]r�Ku���Z��=JR'�k߳�R����{���JS߽���JN��߸=J9^��g62I"Iq_9A�Pr���ߴ=JP�_�}���);����D �X��!B^a��y%�.|:�a���*��N�V�;&#ΐi���3���{����6+p4����{�JR������)I��{��JSߵ���E)JO{�=�Cԥ)�־ϭnѳ7�3yk5��8�)I��{���8
�H�l�C�������g�)>�>��R���k߳�~T rR�������0���6k337�R��ߵ��┥'���~��CH�@�䧿k߳�R�����pz��=�>�5�Y����[�)B��y����)O~׿g�):��~��)I	F:�=�A�����N�x�Uf��`�)J{���8�)H^����)O~׿g�)<��{�R���W��;��d�3��u]vy���u��i����U��a;��di�w{�����g�TR��s�؄!|��TY�!c��R��{���R���}�qJ�(9_�U�s��Bt��T@�H9;\�R����~�"�R��{���JSߵ���)JN��߸=@�Jx��z�!$�$��ȯ���(9^�<�\��P)������|�_h$~;;A�)>��;��)Jy���8�)C�o�b!I8�r����9�
�s5�����������)O�k���(������*,�A�)�+�.)��N�[��R��}��pz��}�^��R�B��c�D �X��!B[��������Ob;uARWn��Gnbر�X�ޞw�oW!ڧa��iE�?}��#�n�����ܥ)��~��R����5��=JB����A
���D �X��Z;#Yf��R����5��=Gℤ�O_4�B���{�D �X��W���v�@�m*�ԡ�R��s����{��)JRu�����F���}�qJR��|׿`�)Jze�g�}�ތޝս�{��)I׿{��JSߵ���)JO=�^��ԥ��`|�  m����)JN��ܳFgٽku���k{��)J{���8�)@y����)O~�\R���߽��ԥ/~���c~���U�N�:�Q�+��)�v�
���:�'p{d^:{?w����U���խoy�)JO=�^��ԥ)��o�R��}��p�JS�~����������q�F�Z�t�(9������� ��JN�~���ԥ)�߷�┥'���~��IeD�=ƴ��ԥD��_9A�Pr���t�)Jw���┊�'���~��R���w��)JO{�����#y���5�R��������)I��߰z��<�^��R������R���G�Lh�;#Z�kw�)=��{�R���߳�R��}��pz��;���|�9AʕUϾ��L��*H�n":NzG�V	���j���r}��;-��ۨ��䌉���K�Sɽ�bA���P��z�ܥ�ea�tJg�s`w��U�%�͍ٶ�+�3���AѺ�p<Ѥ�Z�уF��M�q��iܛ�ћ[n��<%�6��˺Zl�,��F	Bܳ��ڇ��]r�����3qf	�WFKs��/.�ze��r�m�iƭ��ߊ������gZ�xf�m�v�Ŵa�ӫ��u�5m'b��Ϸɲ2f�0<��6�;���ܡ�)v7.o���u)Jw��}�R���߽��ԥ)߿o�R��{���JS̽���5��ztoV��{��)I׿{��JS�~���)=�<��R������)J+�f!:KTmQ)�]s�9A�W�����)I�y��hz��<���qJT����D �Y�MK�������R+[��)I�y��hz��<���qJR�����R��~���)JP�{�o!J�')��n�Ӝ��+ٓK�(9����R��~���)JRy�}��9Ӝ��(��Z��R�QH8��D���6���r���.��P�e�zu����^sr;}ѯ���F��l޳5���qJR�����R��~���)JRy�}��^�)O=׿g�);��߲ֈ��V+{�o�ԥ)߿o�x i|T�T��6( q��)I�3���)Jw��8�)I�~}��@iO~�O�4E��dkZ�n┥'}�����R���{�qJ@F�����R��~����(9�WsF6�V���ܻ�uΊP"��߳�R��w��pz��;���qJPi;�>��R���{fѨq(��2Tr+�(9�W��ۮt�
T�߷��)JO;Ͻ�Cԥ)�<�|�9A��VQ�4�H��#��t�m��S�rc.�9p:�Ι�0-�n�#ɍڌ���{��I񇏵'khf����{ݷ{��I$y�t�B��ӯiE�"���Q�)<��~��)J{믌�u���[̭���R��w�{�����J{����R�����~��)Jw�����PW=_fl�Iԡ9N8���uΜ��{����)I�{����V4�}��)JR{�~����JyY�գ����&��_9AU��{�ϸ=JR������)I�y��hz��<�^��R���_~�Z"7�Xl��5�R��~���)JRy�}���)��s؄!{珪,�A���N�$ꗞsH���Kv'�c���ҍ��j.vn�9L�շ=n���[uەqJR����~��)Jy��8�)J��TY�!}���B��=3&UJ��k6Yַ�s��)O=׿g ��L ��׽QdB��ӱ"B�����)Jy��|_e��oN��ٽoy�)JO;�߸=JR������)Iߞk�z��<�^��R���ܳF}oz��[��{��=JR������)Iߞk�z��<�^����d$����8~�� ���$�w�y�\�)O��u���-kf�eh���R����Sr�Ȅ	-J �o�v!B^���z��;�_}�R�����ܫ����ۖ6��t�x޼��x��zy�57N^(���][�ݺT�J�8��UΜ�9^����)>�Ͼ��)Jw��8�)����t�(9���Qԧ##I����R��y��pz�A	JS�u���)JO��_}�ԥ)����r���jiҢ��%#�\��Ps��=�┥'�y����V���w��)J�����Ȅ	���*B'���UU\�)K�`�?{�~��R���~��R����>��ԥ#�o�R��y�#T�[R�Sc�v��9�r��uZ���H?{����)O~����)>��}�R����μ���5�4#���_�ߞ����X8���[$͏b`k}�(JմRӬԆ��e�Q�FX�,Ӿ�L�A ���_���RUr�����V��~��tۦ�t�(�0e�v۹;v�+����2�0hluҡ9��l��Ҙ����7d��1oQ��������<:��c;������6ָ�)-��B��m\k@a�/Z��Hf8e]�w0\��R��^��e��_��p-ӕ7
];r�J��n4�6�-��W`(��M�Fݢ]��Ó��9Vm:6We���`Y�]�
�{gaIN�y4��8c�ŶĵA�xs��Q�],�6ھ�<m}�p��9��S�
e�Ռ]+z'���0\����g`xP�#gr&�N�CPz�`�*���յ�"���lF�ҕu��l�+�v��� �X ��;f�mu�����of��ɹc���N6�; ��0h,�.Uyڜ���������q��5{'���f�T�+UFR�ۙ�v�0�[(�g�%	)j+�UM��3������s�� l�mFę�[��ٍ�9ٓ58:^݆��)��za���y�-��P�=��E�G>5�$X�C����Sm6gǷ]E���qJ�l�����6&��K;;*���U��/nL�0%�x�$��;j��U�/�8�N�sPlU@��A��*���[��f������};F���"��7�vʖhW�L!�kv*��▛*��h� �Pl��r���s]m(u���H<�7Yj@V����[ M�d>�kk	��\��4�vD�Jm�ȶ�J�qj�U۩�t�d��3cǷ�gfPz�w.���wN���d2+,�.�]�nڰ�J��O*����z٪�*�K�� B�E"��v[���i�k�L����z1��:�F�V�v������yl(�
fK#M@#l�F��Ti��j�tܫU��fm����I8n��\���phԯ�����t���9�eޤ۩�n�N�@Y^���P���g�Uv�MF5&��{B�Ur�d�2��A�X���]��������U��30�����u���~S���h�b�Р="��z��E�? ��ֺ�e��ћ��j��u�ѣ��ݺ-K�.[n�:6���c0��U�Q5���Iػ��ݺ�G:�7O(s;
-I��lU�"��/S6�nx#Q�������ٸH8�=��$�����`�AX$n!�.s%�7&�9%;v��/kk�8�ջl�u�5l�����lV�������p�܍�mTl%ptc�;t�?�}��������B�'�4\�K��9����g6��`�q���'qF���u�}=���A<�u����m�v���u�TY�!{؄!?z��D �+��U��+�jē�I�G,����R��߷��?�9)I��u��R���k��┥'�y���)k39�!�Cr�:���+}�`�)Jy��8�)I��}��JZ�l���r����f�J��Bq��'4=JR�{���)JR}�}��R�{؄!?K�J,�A��RrF�JGM8�r����n{v�9�B�>3�"B~���Y�!{)��Br����Ǳ�%I�6����*jn`�Q�ۮ���9�S��%!����ׄG��%JG.�Ӝ��l���=�}�MΥr�v�1P�]�q
j��r�������;�!����Z4}V���I�ډ���`�rJ���uSpIEm�V�ʛ��otN�`o�澀z�KQ�"Qӥ*Tn+�otNـ>��h~�����;�K����G��@�l���=�}��U�������m-M!Ӧ1H����O��۝̹)��Pv��g�/7e���S�gHp�鱹N���?n���z�?y�Ԓ�C�N�<oy�*x�$��U�ѕyZ*np����� |�5��$f���Ҁ�)H�i�V��۰=����BJR�JÙ\wV����~^�U4�	�$8��+�a��"'�N��Y�V����S�7}#`A1�E�U5f��U�{�)�s{�=�4�=_�2��)"%S�+p�(� ����Y���\qc�L�]�vQ�1���L]U�IEnfV�ʛ��7�'4�7�ۯ�z�kij$J:u� }����0��ցʛ��sIѤ��#�rw�{6i`}�ۯ�*np���	(xD�UWd�VW9à���Ձ��?y������G�GP�ZP >eQWʮqo�e�o�����2!8��Ee^V�ʛ� �ﾏ�sy�rv���u�Ɗ���*�2T��""&sAm�ꞳϞ���r�2g�]��4y��������;JR8�i�����z�f��O(�IX�nz��J���J��u{�rv̏�" :iցʛ�3�݊"#	�J싈SU5à|뛭�78@�����`�I�ڥZ�`�m�����{��Ͻ�ށ�٥���f���X�f��GN��(���3�n���=���v�e7��L2��!,0�E) &bϾ�����7���Z��Q�:����ӱi�ƹ�r*��$��Cײ�d8l�5�,N7/5˷�A��+nַ=m*���m�Ju�������x4��[�������\-�s��5���Û������e� �ӱ��_F�.	�٥d��;�iZ�t��z������`��N������C��\0D�'��ՂD���RF�cj�7RpU���L��k�����{��?o�l+�]�9��ש�7���;���c�	d�;O1(�
�|j�	~��|gE�:T@�	�}߶~,��u�c�K���n��fa[e'M��pT:UV`tӭ�78\���� 3ٯe:r����;��@�=�`f{^��� �h��"b¢�n�f���p���9;f ��u�r�����aM��J��%#��͚X��V����u�=盻�9�y�XN�{b����C�lrnON'�
+��/luќ�G+z3���Ow;�i޽'K޳�:ꚳ }M:�9Ss�5��h�� �
��U��H���v�-�wvs��*盻��3�|��ԡ)��~��%:��G`n�����4��Γu�	�x�IP2�ɂ��ɮr�6!K��:���X<|�jJ	x�n�ִފiU\U�QJj�t�&�@N�ɽ�V���Ϫ��u��.����W��Z9��c��x�3P姃ty	��Di����sBisl�����x��3�����H�����ݫ?�PJqH�r'%��������)r�G��tm7�`��(�
��t�)J�#���4�>י����W6�I5,)!) #CH4���P�߽�|��=n��$N�"Q���Mp�%
:�u`��g���j�����N��~B��ү�r�)����@3se�r���ɼ�V�Βu�>r�l�������.�/C��Ϥ���Q�ؠI����؅!N�s�q�nї[1���:*�m��otճ �G�}��`� ti�$��7&�ʮPk�u`d�u�3�n�aLB�^��4���p�&
����;�7��-:��"���ܚXnk�Q�N6��征���@ϱ��1��;�D	�P$�-$�D��Հ�Y,����\�]L�\�� ���5l�;��:��������*�B�t��H�R7	J[2on9�c�M
su���7���S��n)Qw�}��{�J �8������3�3W@Ź����ͻ�l�:@�Gc�SU5à{��:|
Zu�w�{�&����<��,*�V�\S"�U7�̀�^�@�ͻ��A��K�ٚ��[OP�#�Q�nf�"#���5l�9�Nt<�`n�`:4�Ң5�rw�f�������6�:|ۻ�$�`��p9\��y����ʒ�R�┇Vi��H&#8�d���6�WM�J�.�+��[�O����8qkS�ٗdر
[�{e��A�74[��/GP�z6�0���L�Es�8z��[u��uDb�,a^n������ke�y�n�����n�k&��e�jϔŭ<�b�h7X�w�I���N�aca6�E\�l���X���l�n�0�P-�Z�>�����?i�~�.�p��Y�פ�p>��']��l�/>!
^�����,X�ww_Z���nH�TINHX����t[���w{\��@�ɥ�f�u�4�M�$W�́���a(>m��"!D} ��N���o���ʮ$n���:��S�F��9,�ݻq��<���1��@~�
mֺT�A(	�@�ɥ��l�] Ǐ�S���X�I�J;B���0�ӝKN�|��	�f�^�r��4��PIȪ$$�FIM�OVk�{F9g�-��̉58�G#a]�:spU;y: �w�sM�`	�z��(u���QӨ����nn���
�L�����s`��6����GJ��r	�ށ��K7&��nl�3sw�sI��67$I*$�%��m΀&���{�&��ݚ�2GI��R��@3se��n�znM,{f��f�.FA��q��շ'S��zێS�<O)F��t�˥:�:V.���F����S�N)ND�����zj�`j۝ M;��)���Q16QtH\��`j۝ M;�&��
dպH�@D���)����=����W�{��'F'�`�QvCT)☇�&���+���3�j�qF��Q�()GH��#'k81 G�aG���$Ѫ5#��G�V��L-m ��P��	҃Ry�h�&H$���(D�u�K�n�Iae��h*^��ރl�e�ax�l� k�hm� ���=�OGl��h<�H  �P�^��C��1��P�DWB�t�
�ś���=�K�jP�U��H��}�:Ӽrot�ـy�ntkQ�"QӨ����{7{�+=�K�ɺ�������>��)�J����~���ni7�Fׅ�y3�D�����y7Q��R��Y#�Dj9q���Xj��@9�y�� �7�L�Qwe�݄�V]ݘ���@9�x�ot�_9T��z�#���n)"�k�x���wf�DB�o4���K2���N�8�i9�ª���{ҽ���r�~��}uJ�=*�����f�r�U4�]*Pdb�w�g�i`DGɥl�i� �7���]�	pUrc�m��f{F�F/;Jju��qy���ځ�5_{��=�t�ݎ�z�Ö�4���;�����ـkL*"��d�AW�h4� O��s�`	���>�r0�������.n� O��s�`D�ӝ�s]����h�GJ��r*NN�
���`�ӝ�������eÉ��	$���}隺9���`o��v��΁	B�(����F�y<$<E�=I\���l�����4���t�,Q�x��s�َ�Q��	��-A7U�r�����/$��ţ������
�f�ps������t�:��]���I�]yk��8ł틋�7Y��-��mg�K7.�	x���V�=^����%f�W��뇌��[��e���Á���`,۴��+������۾�`a�����w{��w���w��R�{v�f�u�H�1
��QÔ���9z�������"��A������m�?��+ o��Γ����@rṊ��ԧ�&�q����@�^j�7}3W@���`na�N�ҥQ��&���:�=�s���yOg�o���bd��(T_%�'��隺y�|��Γ�X�a��&j�d������rw�?4�@�Rs�5֜�	�o~��Ms�A਻s��g�f�p�m���^�'�l��0�F�<O<P37u�?4�@�Rs�5֜��N�׼F�:TF��R�w�}皮��ʣ��G��C�P.�����:����v�����*V�u$$�*m�`5֜��N����Np��;��F'qH+��K�5@7���@�{=��.��Ou��R�R4�JK���@�Rs�>v���;�?DGw����~����9ԣF�S�s�{�'[]k�a�p�u�범�D8�z�]?�o��G�x㦣�N_�{�V�&j��͗T�ot��d}pD��\���:����otu'9�	�&%�N�)�n�����͖�{��s�(�hB!a�Ze�I��	d��H	E�Q
�$�!D.�}��=ٜnl�֣I(��ujI`n{w��<�`>v��|{��c����.���bf�tu'8C�I΀{���}�]UЉ�,��2Ѐ���O�9��ũ-�g��sǝ�F�b��������p����i��d�v��uU�[�yZs��� ~M���{�9����)��n)r�@>�l�Up�7vެs�(W!���l�7eW�R�R1Ĝ�����y�s�F�&j��͖�4�]*U�BmU��}�� |�9�rw�����(��>݁��] D���)S5����:�}��N�����Npr�cn�����m��r�Ba=��LεB��ݞ���V�M�prۣw����}���uE^fN�����7��'?�6C�v�M��B�4��r�.R9��9]����1'���@�|{6z��@��C9�J�dr*JN���}�5t��V�����T�iԎ)#&�qX~IN��ٰS���n�6���o̀}����7CL���Z����[���{i����9�)�!D%��&�峒�66'������:)U6��:vY�͠؋/gQ�noWp�y�kv1G28��m�a`Z�R�o=���8�׬	��r���2�:�S��1jW��^�v��hU٭�g+ӹ��n(�V���O0K���U	�Ι�gz]�v�#k�Z���z:��sj��v�	;=,B\���x��;�sA�ћ��׍@!Ӕ�l=v�c�����x����=Қx��Q��ѧ��s!m�%�B�������Н��Upv�dc��ٺ�]�."���?y����'8�i΀���s5SN��U�Bm9ށ���`>V��
y:��{�8_9�PL���5s�4�9��u�?&�@�y����k���)�ݮ��ٵ�?6�@�� iZs�8aLU�uP]��� ���Γ��i΀g�e��Z����b�9J��r\n�h�f���G1ا��v�s8^�\�5y�.]�ԣ�Dj9Rw�|�5�왫���~��W!�^݁���5R�+��r�SU5\����ݥ�DJ����{A�w΁�noz�s]���f�r(ƜQ�!=�f�3���<wf�3�׵�=�{�@�{ZR�4���iG��s��r���݁��>x��IB���{=�j���*F����@�^j�?r������)���7v	DFc�N�Z�:	�'O�|�x36y����t��t���8+�'�k�>{n�k�`c����h�9�&�@�� MI1.�uWw%���U��Ns�6�@�y����ޝ(6�kijDt�:$�rzy�vα�M�؅""T$�*3����@��V׼F�:#Q��)˰�
(��ǳ�3^�K=X�g�w���:2�TN9#&�q��΁�B�Np���=-:�=/�<��N1k���s��6�y�G��Z��9v�3���n�q�㊮S���]��?8���ٰ3Վz�7v��֨���r�������JP�R�R1�V�{݄�BJON�����{6z��u%&���o�J�Q��&7;�<�o�`o�f�5DD$�I)S���v��ˤ*�T��I�a\�}�5t��V�}�U���_ t $"i@5�h4��@��{ε�3�}ߙ*Z��䈍T��n�@�<�`~�W9ž{��m=�����6��:��*�S5�����Y�<��onFwi��[�,a��`�ø̍7X!-����T}���?���y�s�>V���9�6;���n��L��B���y��U$~͛�tǿ���f�{��3x��Ĩ�rF*M��?'o���9��{�y�s�)MFՂ�I�S��k�g�j�7���@�^j�7�3W@�rmP�R��cJU� ���Γ���@]I� �z�A�8}��L�I2$A�KѤ6�SD��� �vm�$$��ܰ���$�������M�mJ
��\������Û8f�R��@j������2�n<)	�3ޮO�e�0�!`c
ht99�L�����9�����		j$�!�X����j����O:�f�c) �,���:8�d%8���RE4HM$6�]�#iލE
n	�
����`@��Bv�8���1�ޕ���it!� %8�AX,�������������������R���C�3m�R�a0��%��lyj�/+p�Że�l8pBt���M3����\��NN��$�i�F��8�:�7`�L蘷`A/4ܗ����E���)�l���酵�����D�hd7Z���J+h�� �m�_l�D�U��l۞��䲖�9We� ��^K�v�&�Y�N��,#��W�@��6���gv^FWXܝV�˙�|PlU$k�=n��m����&��E�Lj��w;��H^�ۧTFԷ+,�v�sۨt�͝�k;u�ghpl<�m��b�V�)EJP�6�k�.����m������%��^U��u��Ӭ�nG���$�j�̈1c����ָy���t���'XH!�K`r�lG\=4��9��bM'Vh�i��]A���Y�*J�[6�k9J�qR�js�f.U��;@�r�!�� h7nGL�m��ɖ5�p/m�9�3�qu����]Y�^�Q�F��
ʯ\�@i��7f�p�t�a�v��
|�W��	t��c�N��c`�RѺ'ls�rc6���+�9�����{�eT֋U�4;Rݰ<� �$�40m]� �c������+��5'S��@�U۟n�o@%��/G@�N`��"���UJ�5�e������.�OK���*�U���p��v�mb�.9��Ҥ�F�6!sA5 In3�c�ܛi�yU� s�yb�e�qv�8��z�:�Y9�ݔML6�*�7$��NƮ`%`�]� ��|��@N��P�ܜ��ۛ�$ku1���n˳ĵv��%^��o��BH�;,:�o����ܒ%W+J�(G:�j�ʭj�����J� v�J��v�<��s�ut�ڪA)4[�3���)V2�%��:ۉ�M�\�5@��[+�yg����+q�O"�UA��%j5ú��i�'�tgz��@dxL��k[7��Vk5�fe��s��*�����D��xv���k� �"����@��E4�����&c�q��4`��T�cY��9@�/bl��nݮQ��n�u��'6݌F�����k��ې��;N�x�q]dx���gX�Jʛm,�׭�.8d�m�ѻ;��6�:��K�S�p���;h2ñ=u�^�\ur �f�vCy}q��q3�k��e�"��F;V.��l��Ϛ��;Z8��Ɠ�4�'v�����휛����&���{����ww�~��o�/�	qW
�N�d�{q�u�hx���i�*�\�f��kq�#�S��:F��No@�n�7�3W@�<�`oٻށ��Ե�P�%R��N;�X�u'8�otKN��DDL���*K�?6�IB��'l��+~�����`��hR���X]EE�wws�?&�@��� |�3@]I����hأ�Q27
N����BIn7z|�{=��݀x�*������n�{[<kͥ�'�I��
���!K��<pc�u�j�K5:y�g����X��=��ޤ��C�Og�9z��X)�#�D��:y��8�U[EI��=-:�%��<����.fn&�����{�y�s�>K�y{u���6��B��b��Wy�8�X�u'8\��9�PNL�\T���� ��f�Γ��7ށ�{��ϨŻ)7i�QTUc�5��gu��t���'�-ːiͪp=�t�*c�9r$�Qԝ�]��U��f�zy�}�5t��֛�:�$�I��{�.�� |�9�9�s�lwѱGN�dn*��纬�L�Ң:R�P(�c���w`{'-qs�9##�r+�ɚ���>���?r�����X��� ��8�I;�@�I� �7��np��hw~~w���R�ur�������o��<c�����nB�:V.���W�|=�D�rO+�`n����nzy�e��X�nn���N�Q��&7;�3�u_򫜥&�}��ͧ���w`<�] D����D�V�L��=�5Y��\�8��n��+vz��$ˇU\G�*���`y�9����3���1�i	���w��9��]�֖����:���q��{�5I� ڴ�@s�� ����tM����a�s�������^!�շ�B�3uۭ�yq�-����D���c��ZT���Nt<�`�{�'��#�H������ɚ�������sv�\BJ"g}��`k���2q���Q��J宁�ۮ����z��V�L��76-):*"S�F4���b�����ݞ��s�|�t�-���S�$�*�v��=TD-�׳�9�]������(P�P�(���]8��k��"m��9K6�`'��M)-]p!��m�t[uB��YM7��.�}zNU�B�y���,�M�¡�h�ar�r�Ð�y�.�I֎[�U\��ӽ��quE�q�(isׇ����Yb.�lb+��:;@%����޺0�W($^�MT�+���e2b�p<��XXƢ�ث���8���l�*�h�K����3�m���z>���X��#��|�l�e�;��u&�Y�P^g%r� �ȒDn��DT��$���&j�y���{���'8��2��UpTYqw���9�� ~i��'8^��������-��5:u��?w��t�9�����Np<�`�	��І�6���?b�7=3W�W9�W�?,�����w�fӬ[R�$dt�N��ӝ������O7XG����~m�"V����ǭ�˛cpI�}]q������/	a{��ml?`be�}|h<�`�=�:y���NtN�JI� 7�dR;~����ꪦ�>�]�s�O���ɸ�gt�H�ʛ�I��������ӝ��� ��݁�s.�"Q��A5��j�y׳�t�߫ ~i������#���.Ru
�����/n�k��9_noz��]���zt�\��%��6�QGya�v6\�ݎ���NN+��uk�N�[i�c%ȪD�8��:�#M��7���ށ��u�&�3@��u�8������.���s�`z}��7�e����؅	\������7�:������dl������XO���i1�\IG)���`b�� -�N(�p����|����{�t�u�&�3@�w,���ª��.n� M��O'Xmc4��]���*�5�T�mD�u%&2�\�[m����νvN�z���a*�T8&��^
�<d�35Uw�O'Xm=����@��݁��s.�"Q��A5����k���d�V� M��O'X�2�mR��h�Fv΁���3w7��ٮ��ܽ:ִ��5:uG5\������u�1��,-(��UWC���;^�mt�&F�Iv���@Ԟ�>'7k�cx���ߟ��L�1�RY
)�A s��]�]�ۧ���0p ���Ƌ�m�E�4�u�U�`	��4�n��{�t�u�b�� -��q�Fܺ�^�v6��<�`	��4'rȘ���j��.n� M��O'Xm=��ۮ���f���T��m�އ�X����u�K��롪"���������$3늘	��6��O7Xo��7]�$����"=>����=�7;j����(s�t��`5�Z��; ���`ص���qZ��ѝ�<;�Z�DN2���3�Ϣ���P���WU�B�V9V��'k�A�=�N��;�\W,%�p���UҖ�\�m���j�@'k�u흺�H����&�Y�<��ri�<���f�A� �dnD���i̲Omvn24U��Z86�f�F��-h�P���f��˭���z�I�����{e��3p*���[����6�㘢84�T�q4B�	=g@չ��M��O7Xmc4������������i���� �X��ۮ����h�GJ�dr*RN�/k�6��O7Xm=���..�\�FF������@���3w7��ۮ�Ż�@ڐqI�F���:y��i���� �X�:�`��'2���1<�Ztg:w;V�6]"a�#Upv�q���n���z�l1Nu7u�&�����6��O7X�+V�t(�Ji&ܝ�^�w�Ϲʯ��oq���`	��@�/�˨&��fn� M�f���� �ot/n�۩!m1jq4B�	;g@��u�&�����4��rJ�T�9J�.T�r��c�b����`o��K���cd��%M!�L�SX��y,o1�k;���[�\!ر���'9|&�����	*��Ȓ�w�y{u��m�@��� |��8�.�j�躢����O'X���n���FԄ�H�m;��y{5�y�u�����<��Хi����:پ;ր�b$�e�nk��v2v��z<Z��1|*�%��J4H���9݆ᦋE�h������0̤��<8\^�0��Ĥ$��`��	�F � $�Y	� 
�|Fa"���� ��h��
v��*���E�:N�?���g}��U׿�s��Z<�N�D⒑���foz��� ��3@��� ��R��Tu32M��<�`��4���,��܊���P��J8*p(�����J^{:V���t�.c���w;��� ��c���fn� ~O��� �'�/n�7�F���h�Fv΀{�� |������<f��\I*SauQqQeU]��{�wSs�?'����,�x6�$t�&I ���ަ�?����7·b$�" ����}*	��c����}N�ڐnI##d�Ȭ�6��<�`�{�wSs�t��["��j\Z�î���۶̹�5`�V����k�r�Zv���	G��ܥ(���I�6���<���$�@�� ~O�(e'QQ	'���v�3{Ӂ���`wsz���뿑$�OxF���ʐ⩙�n�@R�~��<f�<�`�{�}�Z�� T����R;~ͽ:��������T��Vn�@{�I�R�f�J�"�.�����Ot�n��6���G(u��j�S����+���X+�:�Z�$�9���\��P��ؤrɸ{i�9�(��v2<��U;O#��O8`��6�{aܩƻk�iL�ɹ�9\���V����+˶��v8n�Isxs,͍t��E�$��M��6j��)��l�-k�	d()��;v�1����nE��z�i��7mmڐ�&�+�]z�:���t�n������ǻ��`��坞�t�kۋ�����N�n̥0��Y�v�;����r�(��X��Jpcq��ٽ�<�`��4�n���e�HAu7T]���<�`��4�n����NPn�-$rG#d�����������
""fb5��|Nn�@;���!"�P�Fӻ:�<�����۠wSs�?'��1[����.*긃�\������ԔDBY�ݛ|�������`wk4�n�T�F��r"��nqHk;�ӱ�<'7h��V��v��ήdwݦ��B�b����V��zt���$�@�̒�	��.&`��O@c�-�Q�^�*�GTE���� �i��M� �I#���4\TYAw�hsw�>I��M� ��3@6�Ec4jn�86���f��*��p��������˺���.�����;����{����oz*��Mҡꑺ���t@|�upd�쫶��61˶�l���'��3i��U���Qw5w8�oc@;���Ot/n� ��[Ii)pn�6�΀w7xi=�:y��56�4�N��M�R�JI`{ٛށ���eUr�,��� ��a�k;�n����,����Р�$�&�<�`��ƀw7xsOt(5#] +iT�����ۻ����,��<�`�j��\\�\XEMTtu�a�!���ٺ�u�u<pܙ�r�g�GI���B#j�n�:�G'k���=�=�:y��;��4Ù�T0���⬪�����O7X�x� �ݖ�yF�4#dRN�/n�y�����ܓ��6�誫��������y�f�w7xrOt=H!,���=��r���[B����87��:�n�����/n��ݽ:�V��RC��$�w�8�V�}x���ۉ�p๱�7$�:V.������(SA)�Ԩ9'@���ށ���`o7���� ]��QPL��u32M��<�`ͽ� �n��ꈏ�1hh�)�S�>�ݵ`b���[�t��X���.�uUaqd]\��hsw�w$�@��� �o��IV3dT�u)��%��foz���@�7�X��:��(��%IQ\�����EZ��TH��m@bum�z��:yQ���l��k�vw]$t�]F}Og�����v熕{g�r0q��Q�o:��h�\�q���
���\j8����I��[����A嵸�3����Y�Gg��m2��J4�s�ۋ��2t/+\��e������0d�<�1�P*���%HL,c��b:*�c���mk������v�
�����Y�;���M������9��J�ػ8�v8�I�����l����2ٌ�v�pB��9ў֣AQ1F��{�b��`w۷�@=��`{ٛށ���l�M�$r:r'#�7��hsw�w$�@���?}D�g�~���"��&�΀f~�,{���P�rsv�ۛ�,fqҕ¤8��Wɞs�J"^c߬�ݮ�7�X��,��KV�t
�Q��Rw�zy��57���� ���DG�*���?��$im#`8���ɲ���מ���j��6���S�68�ݴ������u�y���� �n�I=�:y��7�IYZۄD*8�l���V�u\�������c���u�/�/�2jJ��8�ԧn+����^�vlL��{���[��>���*Arh�T����<�`��h���/�����,��@�鶉R�jH�l����׌�;���9$�@��� \��󽝁 ��g���>5�r�1�;��\��!���z��/�����\q�N�l������� �����Sx�1[�T�H���$���foz��]��ݽ:��U���KZ�N�TJ4�JK�=>n��}e�!Dt���!F�)�R�D�0�P�)JQȅ���:�����t�	���n� M�s��� �ot^�v|jHZ�Z�B�e��{���5=�߾'7k�c|nl<♩d.���:��wnz����팘�V����ԉb�n���9�W�n�b�����m�m��=-��v��sw�(H�����R9;�<����>�+�M������5n�vn���}�F-r�jH�l����6���`	��@��� 3�-B[�Q��]���5��w`}-��s�N"�ḿ��㤩�)�9B��`f��z�w]���utY��e�Z�c4�8�N�C�ɋ����h6]׮���Z���e
)P�Rv��M���*�F�IIށ���`f��Z�N��{�6919�����5D(�����8��6��K�v|jI-��:�#U�-t׺�6�ٰ�(�����w{��49V�I)%R���Vn���j��`f��Xj�J'w����s� �4O*n��t-��v���s�&�ݫ��u �0KI5BPLФ!(��2���Z~�>���`}�7�֑4��M�wҸ�"bH��F-���}�'�鳩����5�|m$��1
  :xA2�0�!0K�hIu6��ai�kN��h�� �h&b ����)*e"	%��(�E4:#(:<�A܅	W������)2
i��R�ړ �#xs�����`X���c&�ܰDA,��Jj���uh��h
D`���6Bht�X��Z��%C�K�z`E�@�=��%H�"H& �����I�X%=Y0$�Mu��5������Z��8�U��v��9R:�y�����J{���X@�����i��ڌzKnܠҳnI��ݪ�����-���TD�]ivɲɕj�֩vUxf�n�)�$��On����-,�Ӓ^�g��@A,���X�NT�[l���O���ly���i��ە
x�Q3���]������0��'����n�!+���n���)l�����c���V�ɬj(u��Hi��ָ�6^����y�اZ�����]�ZV_@+˻��ᕝ#�.^�zZ�ȃ+Q�D�ʁ%��W@Þ�,��q��[UT�a�rvG��[
o'6t����9g�D4��"N$��vg-�,�!�me�i�˹6�:#�����]�-(�Wg���k���m,
���*���ł�j�nwTcdݦt5Ѳ��D��GO�g9�(�v$�-���W�g[ ۳m�S���� 6�Ȇ�]V7�N��
cJY�k����fm�����	�c)h�r��k��-���
����ek���:Lnź���i�n-�o`�YJZ�q��W!�4Ofɲ�;u��f��d�]�ǚ�[*d�WJs��GP�V_X���ֆX�Uv��J���<sn����,F��M�*���κ9�-J����x%e��\+8!eq��l���gԃR�d��t�L��$��"=�6Z�r��i��s�ݩ�x�"'&�R�m<1���$����HR�Z��q�U ��!{��Q�2��Z�Н�Jegn��Vzݭ1�,��rj3�b�c!=�
���Av5�ho]T���3���4p�sYd��{*�����cj���nQ�Y�թ��v���]\���ާ6Ga�v�.��\m���6�2�BC��2j��lҴ��.��锎��i*4[����DP�jR���vl���ݩ��T���y�Y3�O,�Hl5ԫ[Og�+rd^�������u�/0 �0Q�V:�]E�
):��u<�u���̪��p�� �	��ڝ�õTOP1|�v�/�<�qQ��D5��a���v���h�D�\vN�����"�%��	t��ʝqt�z�κ�m�dv\r$�.��O=v٣d�Y㝇�]�=<9Z+p �F�,�z9;v{5���\�-"�
Fwc�;#�u�J�Ξ���K����5�Q�%`�5���Ğ�q�\�R��v�t�p�n�U�=U�R�٪�A	�-p�eܶ���kl6ɤ�ztw}��w2|Fy�6�����3�=�.�h確��;/7e�/�N�60�e6ԑ��#r?�g�7W@�{������+���ߝ�o�~B_�"E���N��78m���� ��3@Lɮ�
����"�=��ށ�w]���S?=��`n�����.�e �F�IIށ�w]��ݽ:��V�������S.�bs�@���57���� ���n��NjHsv��z��GE�6�]�°Bb]nͼL�
/ax�ݻh\���'R_���a�nz�1݀�Z�Qr=��`�����$��J���X���r��W#脡EP��@����t��/xH�TLQ����u���Ӡn��`{37�}��[)��F��X��t���{�|�X���-�JG;%�G,��5X����N�M�4��AD�䨛���C���f:p���lc.H@Z�����<l\J��	-��R�c�7V�3{��� ��3@n��{��R2�&�b�fbf�t-:�7��h�s�{ٛޜ�`V%��/�����>��n��LP�"�D(���c���v��6���N�U#S�t?r��wx�z�����]J�>��5��JIT�*'���7�V��ͽ:��V�m�Г��4�z����<[ηm����O��P1<1��\a�NqO���r��J,�����D�_@չ�����h�s�{�{�4�G9aUww6r��*����Y{��7i�������5�*���[Q(��,��@n���'���`�c4�Mh)@�N1��+����[��U�{Ϯ��eVUzECi��ϲ��g�Z��R�IG;�5nk�3�c4�9�9�{�{��:�.���X�]-�+Ǎ��-+�dc��|V����仝�bBTRJ: ��䤁H��j��s�/r{h[u�{��drS�8�r�s�/���n{��D���n�����`w}3W@6�EelDpIT�*)s�/r{�9m���9��� P�6�$h(�(ԒN�[���j��uX��{�7�ť���$DSWw�k�Ntt��ܞ���`\��[[Mo)%:
�I"ElS77��6���^1��c�J�;�v��&��=v�,�m�s��X�wi�VKj}�8�!�����@Oh�p��2���T�OC��u�v��p\cN�c�%�k+ӝ�
4c6�h͔���v֙I���m�=vj�n�q�m5k����7m�7Y�ܛv�F�;=6gVZ��?᏾���Ps`�DK�h�.:�:,ݣQ�K������MU��&h6���Ŏn�st�x�㩬u5��l�cU��6.�D�����̞~�ߧ ^��@��� �֜��f�������{7���u�-�����+��d�0��[SH*�bn@���:[�X���@�� ^��@�:��'늚*�}i΁�I� ���$���9��拊��������78�'� �w�oޙ���z��R��!�T����Wu��-s�k��WK�2�c�\��fJ��&�R"8$�S�R+~�oz��,��5~��{���X��~��#ADiF����f>v��p�Q?{�����?��ށ��-�q�(IJ	�,��6l�7=6L���oy�/؆�j2E;%��v���U��{7� �͖�隺�)�&)�nP��Xܞ�I� �֜�t��И���(�q��^+N-Yݸ�,C��FX�Z�)ڦ��Օ�&�=#�0qk�� I;��ӝΛ�����X��Qn�䤩I%����]�{� ~��@N�x̎JuQqQu1j�|��:nz��ݔ�
!B�	$���%H@������Q���W@>�QY[U)�)��s{�	'x��@<ۼ�D��E(�"�Iހff�}隺���~��z˞��V���)���[qN��{
];�)=O4)Cmv�8x�,N\[C�"qȡ"M�`f�^� �we��7� �w�o(r�軛�6�� �n�dM<����Z0�c�
n���7(�I,g�{����K�m� �*���\�M��]����oy���,��:��w��T�|(��rST������h�w�7��$��BSL������� ��.4���l��u٠9^�:�����[.3/\��q_�������{�	'xic4�9++b#�J�HI`n�w� �͖�e���vX���iH�4�RI{�	'xic4ͻ���@q�
OQR(F��rX~��*��۽�t�~�x|��I��������ªʙ��@<ۼ�ot$� o2����9�W+�RѺWIE*%m�ۚ�=6���s���iV�.3=���7Gm;vz�`�;�Z�j3�����ӡ�Xdct��k�kQOW^@nԪ�����XM�蹮��]v��:��g�z��H��gQg�!z��.*�r⣱��Wm"p�ed�%���ۭ4Y,6�h.ɕ��^�+
/l���;UYr����!\��Jsy���t�cvvx�wC��������� v�`2�6\��[���ŏ��X���82��3l�+V�ɥ`
N�S�ܢ9$�7���@33e�߳���>�=����ҝ&�p�O$�� I;���6� o���2y��m@����S�s�wt��|�B���Ƿ`��@��̒9)�.P]L\�{��y�x|��I� ��zt�5��JIT�(�;7��@N���h��`�	>R�	�)�9 ػ9��a	�ݸyq��\]Ҳٌ�v�'oP�΍m�q%U��m��� M,f��m� �7��VD֢8�P�m�`f�^����.�G9��/�	)PB���vJ��t�c�2�́�eIl��r���wk�|�u����	Rs�>�Nt��+鸫���n�� ~��@J���Zs�zwu�^+��h�'#H#���5X��9�>��t���TF���N�l�S֑��tl�,����q=��1��rW)�&'H�T�$�
�䦔R.��2���=-������� ��2H�wUau1qW���z[u�?r{�%I�~��] ��Ef���t�J#��{���=:�*D+�D��G�C�� ����C�2i@���(u �B��ɐR[܎B��w�z]��&���[�M1!L�m�Ff)a�+����`�B!�3^a�o �@�����.h�Y"hG�)����!K�h�' � 9������ �`8RH$'���@����� �CI�ID�`BT��
 @�EP�S��WJ�!I$:��d�,ǸJ$��L����J �ք==XPSg�v*�ڀ����| ;⊾(/j(�&�BeIx?f{���:����`n��QATLQ�R9ށ�y��?u�:��X�'���w7vI#DqX��j�-�v������Vm{hT*��A#�:PeG
��j�۞Y��=�n^�=S3qr��|'B.N�}�r��4��t��~�ozy�Q!��=�[�좊�O���'�WX�'��Np��@��� ^9�kU'J)AA$�@�<�`oޙ�`|������11ʝ�v�\U3��'�p�P�}�{6��g�?���=^��?�z�Ϸ�g*���Aú������*�Λ�>Otǚ��e��3Ւ�̓c�T �S��۞�v�g� ���8�^�s�.�ʳ5'X�v�Wmp�")�T��n�IQH��f��f<����<��#�@��ɋ�&�j�\�2��u%2k��,mn�@<���)#�f¿IJ2H� ۊ��������s�RQ3�׷`7Og�}�IvL��e�U5�h��`�=�<�`n{/N���mP��0�r����{�%I� �,f��m�?.�j���+eJ��TeGB��d���1W+��ECm����u��m�J��f���)���;k�=��÷N�=T9�ö|��i�;���5ۚ�s� f��9[x�.ƺw�[��tT�p�jҫס�ָ��Z�q�6F]��]7d�[�;]Y�C�W����rµf��ڇ�z�,,cL�6Z����$�[�{[s${F{tn��yѹ�ص��������𝱾j�v�91p�����p���{=�-pA�
�J�/(]�K�R8x�	��9��n�@o3��>��t��ށ�a���Zh*SJ)���zh��`�{�%I��� ��T\\]L\M��z[u�'�'8ne��>E��%I*6��)#��UD��߬���~β��[u�	�j�
�b�9�@�y����^�廮���ozkU�Z�hhm�mR�Uv���q��Eܓ<��d��;/�n��_��`uGFI#DqX��Ӡ|�u�	�{�%I��PGeM^�^Q�S]�`}-��b"!BĊP�$�|�;�5n�7}��@�ն�CAF9C���=��� o�3@��� �I�K�4�����r�6!(�M�t�}���[u��;�>Xd�u;5!2]�`	��h��`	�{�)K]��}����S\"R�@��nII�k���f���x%�ְ�j��h8SE�/Y.۶��a�R�J���`}-����9��".C����tRȭ�J�TmӄRG`k�;�P�S#����>�`}-���D.$n�Q�EQ1F��w�j������}u|>/�B, �`� �a�!*�
�A�ъ<�9ԯ�]������nT5�Q�GMF�����X��۬�Ot):�>�ѩ-��:�X�]4�΁���`k��@R���X�󲾙�d�QU��R�w0���b�[8��crl�J锧��y��T���P�J��(rH��f��)I� �,f��m���K��$��ʙG9˰2swRP��7q�Kӻ���;��<���씅�S'9��������릥	L��۰���;��i�q�U�l�-�v�݁���1�
�Q�c�+�A��ڕ#n�"�;37{�1fm`m���۬c�"��&���E[���vuy����lux�6lz�(;�/bS�qF{$�`�"�
�b�8��@ř���[{��XI��<�X��n����������k�z[u�6��JZ���jKj1λ�7WM;��|�u��wfIL�ok�n���/��Ъ0�r�$������Y����Ӡ|�u��4��Sb!9T);�2st��w��zwv�o�I'� �&�&J�"K#)(�`����o{��i�;�-�n�Ӭ�ܽHn{l�g4.:�[l�����;�r:7��V��z��P�[�y��%��%DMh�5�����c�/&�8���kJ�ݐ'vx�uِ3e9H`�]v�;=��[Ip��*6�j�L���u�9�t��t�ZMv2v��[B��L�MX�`����v��fg5�Yz���@de#ʮ�x���ƀټ�Yt����s�Uڪ��Wd�u�F�D�8���/;U���v�s��խp���仜�.8�% D:*SH�>���������+ջ�`n���
#�-�t^d�V��4\T]L\�{���m� �Ot):�7w/N򪪀��j+v�Gl���`��@R��������
>1�QATLQ����5����@�n�7w7���D�$�$t�q��]`���6� m����`o��{�!߁����n蓜���ܺNm��냶D�RmUTӸ=�M��6�d�No���TdT�a������Ru�6�i�73]�6��J1�#�Kws{�8�nA-�TQ�C�I����?�:� ~o��I$�O�4u�SB�r4�''z������@7۲������q#] Zh*SH�;��� ���i��樂�`�L�0��S%^������st�u��R�kyD��qR�$:�ˣKtr���;��E�3A��E��q&jc��`ܒP�DqF�P�t߿o��9��o:ƾ�<�sb"dq�MpT"F�rw�����à~^�v����}�Pn���:j8�NK~��}uW~�ﳗgʫ��Ȭ(���bvm������߾�`w�P�	9�r���vt[���;�6!DDK��X\(���w����vP�B���I#�7w7��*�k�X�������^6�
��
��υ�G�-ˣk;��m>�g׉.2��Px�j�:L)Ȩt���7I�ހ{se���f���������u 5!1uwxm=�O7Xm=��e��H�[LF�*5R����5{u�	��@N��{�A�	ܗW3u16T��`	��@N���i~M 2+�J�
`��+ �Ӱ^���~��U����KR�
�HӎN�[�����@R۬6�����50�$���ȕ�]m���9�V�r��-�2Qu�n���	�)��H�%:j8�R;7r��6��1�w�
>�5��@��N�;�f�u�t�]�k�,��waB��۰ۿ����zt��e
�EB�r�$��i�4��	����u�oG��D��i�NN�=ĵ��7r���u�&���L9������<�9�1��,>n�l��{v��;W�Ă���hB��St+Ҁ|�{��R�%Dk� j��� .b������v%�lȻ((C3���3�:ن��^��)"R�}������(=��ӵ���Rjv� �!�2�d"�)���_WrM0PL	M�8V��jT �8B�ܦMAS"l�ON�%HS���dfA�d��}dҴDk�tt����B�2#N�� `(`7�i'3*�:2

h;�Y�9���4�AD@G��ך ��H�&����r��;�5��4�f�4����C�f�KQ4��wC�Oa&u޻��0�-k��X�u���l�ۭn�&a�v�w8z���);#ר���6�x��lW	�0�[sV�-���+p��u��� ��LI�K �iCnV�g�\��K�]$8��UR���sT�ʵ(��J���[�[��'e�4����ݍ9G� W*�-쐠���W�
�vW;.�7O�rWbr��h�gtlluX�4��X� f�9v�S��ru�̻��gl
��@{p��t��W��ѽ��m�ub�f��%�8*�Ai�p=�e֭vvC5��INu�Pg@��*/.m�[�ъ5?�?}�ѥy���䖝.�>KCl�Nl�A�9]�զv5ӧBIb��P�3������76g/���u��#���NYB~gC�e�� �xM;���"7�:�����
�Q	+����R��9��7*�i���:���LcJ��i�Ӌx�J���:wIj�n�����M��K�V�b�#4�A�����m<�g�8�s��ې��q�h:�iݰe�n�5�/>m��!�nI0Y70C�d�z��	�O-���2�*B��>�n��N�2���m���Z�r�T1�;n��.x8���T8��n��P�Ұ���g[cR��6�5#
���j�@Z�bq\��l�4�H�"��B@jU\�>���(yTJn%��F4�����*��yTmC;I��D)�d�K�W)"�9v���&�Qr�͓j�.�(��  %c+̊��W9�uư����	�۵ �eU���� L�ԅUJ�C�]��m�.�X�ȶ��������]s�v�v������q��r��8��g<�5����v�s`�R�0R9ꕪ�]Z�9�jU���G��i	��A ��v�z�ں�N�=�i�7'(����=�0��/A�T���g��U�a��k�p^�����Pk�����cm-��x�:h��Kn�
��[��K4�'K!�֦��\�������m���W��R��Vf�����C����� �|����{Q�=DК�8������"u�ì�����ѻX?���A��ֲGgW�U��/;	ю�l>�kئ���5�i:�j�����S��m��{O^Aπ�u�{pv]Μ���)��i��+���F�n�U�k�8;O\�Q�5�9��L�Ԩ���K�jܣ2��@�0��8s���!.�[v�x��;j�Um��P9�[�N$���L��В$萻&��z��Wcp:�V��7;�����}�{���vL���{n�%Y�׹9e:.��3�z+;2�uN���[JhE)CH���T���΁�?~vn�� �w�&�3@�H9S����"쩻��i�4��	���$偼��IJ�HӎN��͖mc4�;�i����@ꊻ���n�6����	��@<��|�q3N	���ª2���@<��6���w�&�3@R�eĹ�Eq1� ����vwZ�ŏ��A��պ2�v͐�k\�1nж��v'7jZ�m������w�6�3@<���pʟ�͙�۽f�f������~�?��D��0�dI�HD��&��
 H~@z:��}��U]���������${U�P���4�Q�`~����@<������w�ty)MQ#�*W$�_K��"&|��n�۰�:���,)��l�9rIauWxm=�$� m�f�}�����ī6�7Q6:��$
P�7l�e1Dv�ˌ��빓^�'E��M'�w^�"R�`���@<�����䝟r��r�n�oz�j7F�I)�B�2;���ƀy'xm=�$�?L�ڧT�j'��w�*�UMuX��t�n����(K�s�7��������W@�T8�(��,����|�ݖg���{%��3=�¢M�r�@7x����[0w+�5&�@+�.,t�)��8��T�I��h\Po]�s�;b�l��(�\��6Ŗ���ۢ6늚&�� K�� ����{����1"�m1(��Js�ts6X�{���.�`
AI�J&��*�*n� ^M�>n��ـ����f���IJ�HԎN�}�,��:��s��	,"#�.�����t�j'F�I)�B�6�g�� ����{����8�QQVXk�'+�v�4��������Ѳ�u�/MQ��H�ة4'(Nv\����à���ԛ� |��	u� �t��"���+�W�Us����Jd77y��i���X�a�F�(u�7M�ހo7x.�`�W�o&�@�%� \i)�'$�=��X{�,�7{���B�%�;�.�.*� i;�7�{����[0��}��A�d#
F&��ٜ�l*q�:�맮v�Ⱥ�9k+��3��)�Y���fV����3��,��{
	f{
[��9�e��1�9�8�ч�8Ʒv�%U==�=q�v*�i@��!�����v��9����D��'[������ۜX&��v��p��Cm��rzÇ���i��;4:n��b�fUͱb��V6d�b�fv�j���mk�uk[oi�;tj��Z���{�w}p��7���\���L�G��pvI4����weY���˷"��]��g%���挵��~����%l�ܯ _&4�Jt"F�nw���čݟ� y�����z���^�F��&�I<�UU��	��`
{�`�~� |���iV!�����ӸtY���1�>n�Jـt{�\ME�qUpM�]`�=����[0>�X�U
�Bt�F�#h�B�҇���<l�מ���4�n�j����e�%ڮI��]�֦j���t�w�rV�O�V��ށ�] ;irSLNI`{2iy\�DB�&~�W@��w`���<��STH��ʕ�\���c��y���Q2no�`n��X��5��$�rn;y/۠����`�����4i��D�5�@3ٲ��d���?b�;���@�b�$�ƓFҍ6͎�T��:Ke��cs��$�<�ngЫ�Ƨr�:$b�:hQ�ܒ��d���?b�/َ�=��؅�d��NJ�r���:UE���~��p���� 䭖��˔q���)�E(�;�n������qt�ي!����������]��U����MjD���$�ԝ�{7��8΁y^��lB����߬h9�tQV�JI��,�M,��+���z�͖�75ʄ�)R�'$�i�z:�۱ڮ.<]0Y\i��h8SCw]����I��RQQ���l�k�V}���=�,�M,�MSX% �N@O��/�n�T(����y�>o�t��+0���-pT"F�Nw���`jV�z�N���۹���WWs(�W&���CT��t�}������P)�		P) ���J h
V��u�{����蛽��ª.�0��u�os{��e��ɥ���:Bȁ��r����ݎ�|���Lv6L%���e)��A7VH�j����7(Q8��۽��6X̚X��;ո�z�J��I�Iހ>N�Jـ)�*�7���<�L������M19%��ɥ���c�;�k� |���L8��w]L\U��c��~�w`����IB�����a��kD�)�I8��߷��qBS�����N������Q	//T�����"��:lt��j���V��ٻW�u���tE��U�h�E��c�S����j�G\i붩@k*qV{ݶq�Mq�/Xu�Zx�H�Xi+�q�6���n�F��tkv#�ے�je^KZXN�ن���ё�d��z��we���3��)��ö�鞆��� ܚ8���\s�kuU��-�&�S���v��q[(:��{����<|��B�9��몶�6w��c��m6Xy�2	�^�s�qFy:�:;Z[=�H�> ��^g�2~�W��!��۰߿4�'��"j��M�,�M,_r�{�� |���B��]��Y�USW��������>N�jـz�̹G�)�B#��ｻހo�e��ɥ������`g�S��J���������[0>�X�=�@�{&Zq�	(�AIM�J�]�ьp�1g.�+]�G�Z�'Svy.�2�`'۴�.Ji��:۲�]�����˰�+�5 �u3�������@s��TB�%T_���ُ��8��DD)���ST։H$S��q�f~�ހo�e��ɥ���c�3���4Q�P�s5{���R�`
}ʰ?D�_�{@?~����r&��DԒ������T�Bu�u`?7�`���|�:��U�m�omC��n�P��t:���q�0uM;��p������$�p��\�]�g��gَ��6�����@���(�Т��
'��f~�j�7ٲ��ɥ���c�=�f'��P�TD4��v ����q�?N=�@�@�R�9�kV~�5�S�g��B��� !�ZL�	����tc���I1�D�AHhbmG*�.*Q�B���L"�Sp�p�I  �zp�:�.�tdda���8o�7�&6�a�� ��)�!4d�b�4;�Ȳ��L�42�b8��G@WAT�D� j3�&�HR���6&#���٠]T���(�'p4����%4�Zv���"�?k�-��1te7f
�K`�d� 4k{5t�Đ\�+,�I��$h��
��0	l�4�I��G��Ãڤ���M	��>w����_UOS����;�n�z�bF�Zt�)�'$�73��?{+�gَ�?�!)�Ǽ��� [H\U+��},>�]3���7ٲ��ɥ�}�'��Q�%(�����V��S�I4s����uhؙ�+<���;��q�MSPI�H�������oz��΀�q���?V9��$�<��.�nn�t�w�6���r�.Oz�wX�8�MQ�X�4����	r{�����uw{yfMTe�^a�>�� ^I�>N�2"��҅ ����*�%���,�-�Bt�m�P����� �;�o# ^�S�4�o7bN���T��:���@n��F�u�C,Ņ:T7�X�#�[\$v��U�>N������~����U��� Z��)�'$�3wn�_{��7� �;��������*�4<�`�{���6�0�F&��')6�8$����*�n���@?'��������92n��$����@'xmd`��pY�ށ��r�Y���n��S���A��M�	lS����:(�5Źn�8'�)�6ax�4�-�-�
�"�����,AZ�#riZ���1���5۶�����ʘ�/;תIxSp7mvk *�;m"�d4�\,z]m�[6R���i���s�z��wfЎ]6�yM]�@zw�nkv��v���:vzl�B��"Bv:�A��	�\�H��.�kI��5w��{�<X��d�m�v�	y�/=�+"��I�5���g	�#�8{39TG$�~۫>~�`{3���\�W�ٿ����W�N�N˅�cMˮ�����ot�w�5���DDɞն�m(6�(q8����ހo��6�0>�X�B�w%D���ܕUSw� �;�k# S�U�rM�fbh�R�brKs�K'ܫ K�� |�����w1eU@�-�\�����[�z�=��#���$6%��v��NJt�PTtT��S���j�k���@7x}l�T�JVUĶ�8$�3=����s��T�^l�7}4�1}�vs444Q�P��� |��������ɽ��P=jHڢ9NK۹u`g��X�n���t���f�ii\������������8$���� M����.߳�Q��JӦv��������Ď�պ�yn�듪�]��
�vP�t��W:o����� �Y�r���)R5Jr2�Cm�;��l�3w20��8$�ꏾ���	J@� \�U)�'$�7w.��������\��J�)P�]Q �!��n�3�6�#�!�qS5{f����y7��͖��K�bj��H&�'j� �M�>N�]l���������y�t.{�;x�G.����������q���I�78�o6��&�c%�7w� �;�9u� ^�S�o&�@3u��Zܑ�Dr&����K>~S�o&�@'xG8%C*�o,ɘʹ��4Ԝ�ɽ���˭���˔S�dmJL�+����|���=�\� �}��I�%\YU6m$S}��s�w�Ƕ}j%(�#I�9;���?r��W+7/��7j�;����a��ީM$TnS����.=H\���v���ع��X�C���+��c)���R�@E)T������zi`g��z���@���@�X�f��mI+�����@j��Rot�w�%���i,C$��N�qX���@7���(���t��zǴ0<��*x���.�R�����@~|Ӡg��6s߷��5��k[�2��9,�l�W)�5s{������;��;���w~�s�Ƿ�rh�g�\���eў^�p�m�s�:�m�Ѷ� vp�;s*a�SGnW^BRY�;H>����D����bԨ a��gnȢ���n|6ۡ���c:�ݍ֛V��5��g)IHan�8�;n��$xwSmmLqńq0;��u�1lPVڰ���\�U<=z n]�t��j���ݛnۮ�
�Nݩ �F�<�nJ������֍x (���F�4uUf�������qW�-�vњN6�c��;=���6���4��s�I�$�.�+��΁��Vs۽��� ���G%�U܅QtU�E���M�>n��`�����R�R�T�c�� �n��d� ]\� �&�@"a�����MUw�w�� ]\� �&�@7xi�Ԙ>	j*QRI�tǚ������vX�M,��%
kUG��%�v��<9p��0�i�d�{F�Ś��l��P4D0��!�I�N.��o����� ���ur�c�"MՓZ͛��}uU��}�G�&�Y ".9�D%AO9�@n�O@�f��<�[b��R9NK�饁�|� �M�>n����ww��d�NYS�hRs�o&�@7xy[0W�.P�@�)�)1��������t}�g@�W�z�P�#�ДmQ>�����v��x���W;[s�v�ص�m6d��;'!����u����8W5�m�?׀r�f �\� �M�.�h@E)T������zi`b����7{��l�3O��pZҩEH�a��tș�8�ي!(�)%	@y�=�qX��ưRD"��8����@'x*jp>�X��"M�*T�N�}�,c�V|����ٻށ���~ʉW�$�P��ҍ(Ӆ���v�cn ٷ��Z���e���*��ܧ*�t�q�#qG$����>~�`{�� �;�:9į���e�$��Ve΀���ܛ� |�����:W(����6�n+�f�z�ݖ��+<�����h����iB���˰؅3��΁���@�W�z�BT�	/�"b�Im[^�Ϻ���Z���J*SLM�`{�3�잁�������9��(_c{<U�vNu��^�<r�`�t�y���Me�'F洜����q]n3��ć]�����v߿W�Ӏ{�{����58�R)(k$B��V����}�,c�Vy���x�e���T9RI;��� Ӵ`����{�	:��k\�6�9!���م��~�`g�������%|��3,�&���4):�)ro� iՁ�Ӏ/�?�3�B *��U������
��{�s���*��U���Q �@��棻���@UZ�]�������������������������������c���?��( *��������( *��@UZ?�������o���?�����U��������_�/�<t?�ο�����������UL�Q�AVIPFHDE%D� �Q!Q$%D�� aD�D�Q$H@eD�D!D�  THP@�Q%eD�"THaD�I%D��THQ Y!%D�AeD� Q!aD�T�IQ RTH!PaD�!D�FTI �!D�%D�Q"H�D�Q"E!D�Q! ��R@RI!D��Q!TJDH$B%D�(Q%�TIQ!@eD�@!D�PYQ TQ!T!PeD��"TJ�IQ �D�Q)Q"PTh	` U			 	B	
A�V$ ��(�)��BBT��BPFBEB�H����!!��@�B	��			R �d B@a B�(
B@�! d%R �	d	 &Bae"Bd��HB ��`P��B�B�A�(���	BP�B@ $$
Q��T0�"� ��%$$D%dHF�%F�%!!P@� �QaD�Q�IUD&TIVTH$D��RPT%D�eD�E�S?�����_����
�������㳇���������w�g��������������W���n������@U_�U�A��W�U��:3J *�Dk����&��p��gg������/�����Ј
����?�"��g��2>;Ͽ�����ΌU���AU��̢�����ᗝ����#��"���{3����6s>��? ����ݟsh *�_��w���������d�Mf��6X��f�A@��̟\��|�噏�P  t
�@@�@  t�     k� o�RH�T�P
�R�H�I
DTTE��-i� �QB��
A�mM� ������UR�� 
P��    z�  ���`\������u�G��
�`=� {e�,�@��{{���>��>��y�.m\  Z^�uU�ڪ�\��dFZ�V�{z��Nީ��`z�վx��ګ����{n��w� ݀F���.�^�h>PM9� �ws����Jt9�oJ)�馔��P � ӣ�� ��S�7Ew�)�ܠ�M�sJ  � ;��5�n���Jnw: w
	���:)�n uӳ�)���g���A���Ϧ���J  � i�@T��=*r┥71Ӡ�_X�}ث���`�"�(Z�Y�Cv�=<�� �;���!�4���w�;o ����;����`;��4$��Cs�����{���x  Ax  P /���J �x�w@�>���� �����<�@;`�[p3�w{��s�9ga�!��g�d{�{����0y�ry�T�`t�m  ���� �  (7��_ ���� �����
��Ά*͏M]�'��ҽǽ����6��l��c������G�7٥�B���>���M�p�{��s�f}v�97`8    D�M�)J� hǪ�J�   =��T����h�S�*&)R� �5?F�C)J� h ���ʔ�� )�'O�������?�5'{�t{��{��**�.���"���TAT�pQW��"���*
��DO���я�!�+0#b@�V �WBE�1	��6I�G�Æ�ԃ��!O���R�J���(K$�`��s6q�������η�<;y��w����N�	��m���=>N�������N�K'I�f�FE�L�d�&�P�p���) p��,��,�����BӅ9dHR�^�b��^D'5`�h��DH�r��L	��i��Kv��qu鄫P����B�](v+��^�yt#��B���e�RP�<��,,:��{74����u�H��!�D�r5��
$*@��L1�	p�İ�!XR���D7
®;c^�Z$�1�n�a�RJ��;�~�;Y�oh>� q�{
&��r������(r��%�)!þv<�mX��hG�w�y�M����m,43)O�S21��?}�KVٚ1��Ґ�,
N�yd�wn��$�e�6LIIp���[i�a�-0-�`m8h�������(B!a��/��@!�$"|@!����dF@�d��$$B!HR!��ce$6q�V0�`ԑ�A �s�+�%1�@i¦���`FB¤B��D�R�@��±&��1��[̙���������1��4����X�~���N0��d"SP��V$S#L��1ˌ�h����p��e~
�?$�O�
����M�����XY>�ϘK���f�:�H4#RM�>������7�����V�P�� 0!B�
C��Sp��P*`cF) ��ā HBMd�9~�X�� �d��bA"Dh�B@�$��O�d���!̉,�]/������K���/\V4ccI"�K
R!#K��J݄�;���#XT�������1��O�,��3�ٛ�@��Ē���B��B��XHZ�d�)r���ix[%'Zf뙁cRB��.�4Lu.�M�/�j������߭����~3LB�T��atA+�&�S	q��8�q��F�М3Y�\	B����e�������|�m;��^�o߳Z��~�g��CP�H�`C"VD�	J´��9?S�L4~�͛ѡ�F����捉�$��BV�Ǝ��� ��bI +���Ltd�4홑b@!,!��	�{�s���콺N�tu�%���a�ZF�f�S}p��(�$��JcnSr�k�~��HT��!ca�¤.������?^Mo���r4�A j5��
i䒙���,��qQAK�>q����(3V2!�?�������u�����¯����\�V1��d���^!n��������1Ќ�$䅘�hK��#.�o���7p�Exk	͒L�w�n��i�%b������l�7�	�jP����_ۿ����NE�
�
@�� �*1
��&�|;�1��p�� B�:>&���a���\޹l-�5������"DHȔ"�rȑ"�1bP�XՍ"@�H�`1�dLH��D�bō��4�\P���q��HRHH���*��w/q�~�w��<�=��n͝r0�f;
c�2@�	���aĢ$H$$HF�B%X��Ѓ\�0�D��1`J)!bU��G �IXŐ�H"�H�C!Lb��al�D��F�P�J�ȍpH�H!����1��:
$�H�Z�J0R$
$@���C$X@��1Ӆ(iaT�J�j@���n.��`�4����$�`�$T�1$V"�����B��ɩ�kg�od�,��~�o�{�~:��2D�^g�HF1aQ)��$$,
i1�Ω����'���
H���]v�o��4�#a_�����(@`D*��
C�C_�B~�U�n� H B$"�f�g별�k.�~���ܤ�~��G��1b�60��t����p+�*�t&�	 � P	 �)�.����?h�B�8a�`�H��
!�B�7̈́.HBj1�a����*A�­H�B��J$ߛ�4&�Y��$!H� �IT��$B�Q�"ń��Ʋ	�H�
����$������ Ո���"FA�����	�� F�ZuaR)��Ԍ��@�@����)��� `�b�1�(@��*X�p�2qxQ��%aBR�?���Re�ԕ�4]l��HSJ�$�(`A�5w@�H R@���e֍¶l�:���~��a,HB����Y^��$c�����B�9�	s[�ǡ�0�iH�+"����*�B'�F�h�A*w��T��X�{޲��Ed����d&��XI.�&�U�
B�dD����s�M�!
"|�dB!!C56����,�"�(@�BA�
$ HHF��٣�)�����x��q��S\J��͵L	IR0�˲��3�%ٽ�_��tȄ(@ ae�a5��I
:6���ӗ��륋��˶����a ��%8@!>�??�`�����	�!�4��L�c�L��͟�+��7�}�'�4Ja��ȕ����B5�Jf�s&��%%>��A�qaA�ė#\0�F�L����Xҁ�"P	��eI@��r�$��d6;�XT�`��T܄B�cHi�
�!B���XP�E�0!XE�3P��$�!B5`��;�M�(*#�/�����HԐs��6o�B��#�Jc$�M&k
C�ͻ���`HO��Ѹ�4a�h��%�oz��Q�	u~����2�2�,)HZ0�HB$d�C�n�S���f~B%HP��3P����#Ja�@�Z��S	s�t�C�@ B�h��P�11��Bɠ�do�O�7�@�	aD�#��H%�#� ���G�1�$�"0ĉBB��)��ke����ᔛ�i�B����H4~00#@�p1 �]pԄ��3�,���	$!�X��\���1! P7wߎsXe�ń80����$�V4�,���D��0c�:kp����Q�C���K�22�R�H��
�!e�%��Vq�bXH0b0 �0�$A ��`13X��K1#@t@� "D(�l�0 �B��alM�����!��I�*E@�	 B����E�&m�%�˶&�F�H$!B	a�H� �>C���E
1���
#�
&��A�`���`@�?Lđ�	�V]˒�J������J��0dI�+a.�&B�@�$#�V$!H��.��4�!YR�lJ$���,Y1$���&�	eHM��KX��ae	YaXRVBCD��HAla
�ic���7��xX�y,�������lQ���R�^��"�H��@�ҝ��ui/i#���n�BVp�who�xs�g�X������[ٳa�3[8�a�Gl��D�D��A���5�5�k7��B�D�$�!$�G.�~��kFkM3���1`T� ���:6���K*B$�J����(Kx�(����!�%�9)L!H��!HR!++2-"F$`@���A��Y30$�Ei�Ĕ�a]��¬
Rn\�����f�q��p!HP��@�H�j�ee!I�H��\I�twZ���a0�40a�����R5� mbU�BO�T���4����J4��dM8c���rI$!��!@a �
�[�B.�,���A�~4��Mg����m�)��p�$0I��� B4%>7�f�gX�0�A�t��SR@���\�}%5���|�>�,'ѝ�V_�����v�UU�+m  � v�n�  ,�4���B��!G�[-jN�[��mؓn��
i����`��6}[
��5T�US�eX�I ?Q!�B@h�݃�ԩ0 zzFknn� �VU��*�T��U���UUnt�D���4P9!�[:cU`Hm���l����v�$ Xi�۴��r�<��F@
Z�i�IF��$�`�m	vض�  �Ch��-� �Su�73�[��J�YV��[�Բ��꯶�b�V�M�e��79"N$�#m��)-UUF��v��UA��Q��޸�6���p��[%�]6*��yv ��lU+�b��o0%��R�/Z  [m�m�U]JJ��һ5(�e��Kh۴��ٲ� ��J�JE�.쪪��n�@[���[m�ia,U�΂� 7m&m� [Kk���M��=Jm�Ͷ �=�h�$d�ފ6ٶ�8 �� ����M-� �ko�l� �i� -�u�\�6�-���ۜnҵUT����&�LMٖ�9"@����oS��U��� %�/[yu�;om&�i-� -�[KhH$p6���AmlO����kh�J���Z�9IJ�6PT�ץ�_��%����u�m� lm��6��$m�m��m���6��J� mUTr�PlJ��ٹ{rjU�c�j��nP�Pk,�UU*�� H  -/I�˵c�6����Χ*�*����U���QJ�B5�\H�Iۀ {�=JȬ2ͮU�e�rؐ����,UP4�%�٫p�ob�+�,�n����9�p��eZj��[��*��\�T��\B��R�e�v�,���^�� mS']\m�%�Vy�%ڪ�U;`�8�-r��j��!UU mݵ�l�	2{m& �-�m� 86�m� ���*�R�(�+]*�������`�P   �Z����[a�l,� � k՛lm���6�k��ln�Fq���ѻ�2����^`8V�m���m���` $�`)L��UJ��Z�J���Uz�L�1��h 6���`[@ I��:e��`�a��@6�6��-�m�Ć�k|�M�l ��J�[r�ob�dA�E���7����ڬ�v� �Snڔm��kX�Im�;m��Å� �Y0���iz�R����kiV�8�]��j���@j�ڸ	K�{R�յ͵�,�`�[T��u�vm��H��,m+]�Hmm�k��һd��5�ݢ��\e�-A�[@ ֛i�D�WM���� �;n-�Bsi��[Q��䪡͹J���W���\���Ԫr�J�5�+V��I�`m�-��-��R�R����E�S�]�� p  m%�H�ݶ�-��'&�m��o[kUi888��:!�ҷ����n���R�;���u�ݞj����-��u�ŗ��.OMw��n�cE:J�,4��v�b��c��ݹ�(q6Z�n�KV�ڶ� T�� �6��x��A ����;^� m���m�4�t�AHvĮ�@A�d8�P]�V��cZ�ٔ��*�]n�rA �ځmګ�����AneZmؽd�    ��n�&�CV�Mmp�i6�ӆ�l�گ�7E[`�l@h�kRՎ��檇u�3�6�eH-��[���ZX��j�^hr�%ٳm����ĺga%*��t���Ƿ �*�E�J�ɠ�h�U�Wv��N«oZ�]R^��ێ$8 m��BF� v�$�c���[d�   ݤUإ��J�T�)� ���l �h�[V�%�-�l 	� p    k�����g�u�h�� �VU�< n�%Z�����eZ�`-�@@���H	p��I6�ݶ�v)���@!�c��%��j鳮H$89n�^��M�0OKz���g 8q�l��LqԵR�J�q�7^��^��}��e�༫e��=��m���R�\vn�t'%%۷[�C���5Tq5l�/ T���[CF���T��t�&� p�*ʵ����%h
���p��  pm���֑ �� m� ��݁ ��ɢ�%��u� �Z߃���	��mհ�8��n�m�@mm�	i5��``m�� ݚ�9��h�a�Uv]S�+�uA2��%��<�H�ڤ�iT���rb�xϞ�p��[̵�`stP:G	�^UZyh
���Uێ���;L�5R�+[6ݹ.�p��tv�#A&8 Ѳ��e]:�[UN�Ѕ� ���b.��p��Mc���Bm���}��[pHm�8 hձ#m�l8�Xm�6��H��m�n�ְ�5�m�M�mm�m��[D�i���jmku�m�  	  �`@]e���j��+mU*� ���&�kͶy!Ĳ��6��-�$p8���6퀑�lm&t� H�v�!snA��#]u�Oi4�*�li�5˅n��\U��	R��.!���ݒ{c�[�ܑ��bd3O5m�r��b���`|C��[�I�1iKCm��
T����8��W�|lR��Hx�2F{EF�ь�#!uZ5�WC/ ���&�lm�T��` �4\,]ZL��M� HH �`   � lq۲R�� [@ @d H�6�;m^M��H*�UVT
RZ�e�{V� ��:ۢ��l�� 	�fؐ�f8�y9����/@]U*�m\�J� �[V˱�l��W���<B#: EյΩN���9RZB�5bf��B[8i�#�^x �ì�Шэ�Pl0-�ߝ��O����u�ik��� m���o�� n�L@-���m�#�V�Id���	 H�ċn� H-�����:9��m���q/�\���һ<dm��X�����]sر"v�L,�ٚWYB��d��u����[D�ET@U*�յ.]���4k%�x�ZM��]�"�9��	��v1NEj ��.�UX��R�ՠ�A E�ciLl���$�(ڴ�e��m�`n�kX@i7V�6�� �l�uU*������)�s\����:6�n��p�[f�a֤Y� Z"�N�ݖMlj�S;uI� ��r�]�8P�2N·z��U[җl�s֧�U�(ʽcRԫJ��l5-���
��U\� �Z��˳A�UU�%�N݂T
کYUYV� �m��2M�en��'UU*�۝j�з:�րm��Ԑ٭��8 Bv�J�[���t��6�AK�c*�P@���t���X�ڶ�6�m���I���ޗ�"�Ѩ$l��` XI�  3k��` j@��-�UBF�mm��ݶ	�^��5��ö��!&Ͷ  l�h�[w v��  	�O6^������p�*UUmE�T&U[TK�� $�zP�n��C���&c3UUc��+ڸ���mX�d>��~@ey��(�ym���H�@��IgY�,HȖN�[-�	8��N� �l�@-�I�v���k��0�m��m�� B�$�e�U��U��d�6�5ۀ�,�d��m�6ض� �HM�;6��m��Ut���}�z������;2I��=�ԑ�V���;mt�f�u����pmHMT�,<]���j�d�D$�h6�v��nIl.q [[ �i�u�:��u�5���`� �FEUz��H˵R�lU۴��g�7E �
����[�5�m��  m-6�5�p='��m�uC�	�y`6ݎ	���t� �� m#m��nIk��5[:BV�m��nP8i��g  -��5�[d֕��ޫf�%%[j�T8t�[L�mm��apgK�����;�sJ�u=�A�܉����&�[��$`-���9&��l �#e1!,UUR�i��[z�  9�M�ls��֙��:� -��Al��m&[��m"� �&�� �UT�W6�� &T�mUJN�5J�0�0   ��� m�����VÞv����nA�yj��V��v7B�ݷSh [���Z)V����ۀ��md�m���[��:   � I -�     �ͮ-�kX���k��۶���o  ��j�[�6�ٛl7Uc�9�f˫�4��m�+G-���M���b@���m����n@m� s�xkrm[cl� ��d/l��� .�9n�����v� ��6lm�/Z  �Ŗ�ȫUL��U���@^@6탤�  [x�հ�m��Pm�6� Xn�`�Hݭ�� ��v�� R�W�[}@Uu�.� [@l�h�I��6�,� ~�e�@s�+J�@�i����$h�`/�kX�m�n� -��hB�d�$�l��c��˒��j��n^�H��,�T��(, ��\�2l��@m[%�i3�knZ���� �@m�[�-�� m�v��m�;���{�ʘm(�6����G�� F��� ����:�8(;�ŬDh��!��P��J#G��^�������P��(AP�������t���h����|	t�X,?)� �$`3�H(M���»��/Ο��EF1"���6��F� tT�D� ���`��#�Q#�ʩ�ڈ#�� $8�@?":Uٴ? 
~D�)�F��/�"g���Ǣ�|��Zc���������U֏�@8S��"��Pb��	�hA	��b	�� �"�Gh��H���@��~M �#�%L4���*?t*�(���]v>?�
 � j� t%6��@�tN"��Q��(���nHńbA1HBF`�`�F(B �/K�#���P�~~���� ��t���P] ��Ux ��pX�X��$d�� ��RI!!��� ��D0�� q�� a�z�@���E��ht(U4�8|?�l@��]��.�"�"	�b
4U��i_ʠL�N�TU��}I@��E fn��a��vɳ(!\)m�ݸ��pD5<r�� k�����L�H�y�s�ڦZ���[!�aS�h�ܤ��$N5���mA��̽�f�W�	�����MF�[ɱ��R2�t�j�RM�:�r0Ab��*�p�ݦ:���6�S;-7Wj�8��<ښ^m�d�eѲ�S�F����3�]&eT�m�h���l8j�[r-��ej]�YYZ��H7J�uIC,�^w�H6�j�6�8�����pyiͅX���nS6���[b�vݛZM&��ê�f݈�e�W �����%��L��뜕5I�
�.N���YG,�Km�S!Ʋy�&:�c�8.��h���,��d������8[N�z
@�DE�9��Rmv�6�ujT6"<�>V;�b�������k�mZ1[��`0[��Sm*.�-צ�M�a�9��ש)W�Bm/;F98ZLvv\۵��UW��=�9�L�\\���u�{fA��H�m�HqJ�s���*�C��.��G	�l�C�jHr�Y���q#.v���D�����y{��aZ˗n�PB�u��q�@��k5v��f���+��q<�	�����v6U�m�x���Qӱ�Ĩb�QM,��"�9�0�]���G^��57u����	#ح�jݔVh��-�p=�y9qZ�K4�Շ"��i�&���w�v�\
�mXuy
vvd)�]��]��l�[O:0J�����]4M�ϐD�N��Y����u F9��-����"ȥ�۷M��ma��W�5f��#�nA�m$H�[+�.�a˞^�,�r�A������/�.n�t��k�pl�hCX%1�7
��ۮp����K�<d4i�-c��j�.N�9ږ�; ��5Y���즚uݎc�p5&4d"8O9��$���dN6I�hM�U�cd�� Z��rcr��д�|j����(F$��*Ԫ����{�� TWb�."<��fʚ>z��E��<�?M�'?y4)�zY���W��k�m=pN�b�cA��\j���+.�W�u�ۦ�d��3�f�W�s���BTX۱�NCӪ�q�&���n�%�9��Ic`�<vX�9<���EF��Y��ݬ�-F�`R�VQM�eƠt�t\�[�u�#��N���9Yl̸�n�����6��͠�$�C1(`���hqc���f�Ui,�֩������I�fS�R�Iƭ� l[a +ab	IxFĠJ��vud�`[��ξ��_ 7������E:`��jݬuȳ�H�d��uwc�;[���ݪ��J�v���o ;$�����X���-�n�];��� ����x�`E�s�;�n�5m�ݫj�]��]���"�>��X�%�9�?yW6�	��j8���]e��h����ˎg�6]��_�Ct�(�nٸ�B�i;x�`Iq, ��]���WD��Jݮ*��`Iq,�!���nL߽��;wٹ'�gb�7h{D�tU�]�ݻ���K�5wc�7\� �K�`qWb"m���v������ʪ�D��X}��X�q-��x4��AN�;�ݷo �r,�.%��^�����oJ������̷�e��r�m1kE� �`�`ƃdvR�ڝ�i�3x�%fm`Iq, ��]���"�7���n*m���b�K ;$�Wv<uȰ���z�7O{)SV�ڷb�Wwx[<��"ü�U_��+z�\T) \U{����ܒ~���rO���5N�իI��7\� �K�`d��jݏ ��tJ�ڠ��ӵ�w�\0�K�5wc�7\��m�x�Z�̎�m)3M/%ɶ�u�m�z.��4�˖Vc���R�`��PaJ�v�� ��[���E�lŀ}�]��N��ձ�ww�E6<�*�"G�,xs� ;$� ���r��P��vݼuȰ�ذ�)#}�^���wH[�IZ�t5v;v��ذ�K�"�s���9�r�rR�NrI/�w�^����-�f� ��-� ���ǀn��{�9_,,�EB�k3e�5��3�ySӺ�մ]�z�n�-juU�7<��62\����#�7\� ������� �y���]+��jդ���E�H�7��^v<����T�Zv�	���K��\�^[<�	����-�[��+cwv�=Io���<�y��E�l{-�qWb���+n������E�l{-�I?w��䘦H����Nv��]k��i�����ls�8��ts��JפtCӈٱ�#��+:���
�*�=������3(GMD%�@�
˃nx�v�Ȃiة���0)g���Y�cqXl�����iv�������m�vȖXƭ�S��zgk����ۢ�`Z's:���pkb���3��	� ���V�;���i��٢'*K�Kr�&@���a0�}����Ni�NI t��w�2W �d��9�<�M�=mn�l,��0]9�a�QZ��f`M0e�7;�=�`v\k ;$�V�xkb�R�����Z��Xݗ��[���E�w���n�4���һk &�x���	�E�}�q��$�T���j����~�qG'����}�q� �%���	bwWl�Jզ��\� ���X6K�5n�����O����1�l�R�ѳX�����aq`�On|�]�i��,�gv�����T�Zv��=��	�^ջ5Ȱ�h��N���Z��ٹ$���[���B�4�4
V"�\x�b�>��f�v$���էwxV�x�"�>��f M���8���;�ݧo�UUK�{� ���� ��[����q݊�Z�.ݼ���`�/ �Uk���=��	6�+T��n�#���o7Z�\�66✭̭���W����̵�*Hn�k����i�f vIxV�x�`wf3 �b�:vR��n��ջ��:�c�&��vc0l��|���B�ݫN�+�;x�"�>��f͟R�T�UWj��>���uM� ��q4R�j�ҫN��vc0RG�unǀlr,�C�"vӥahV�+�`��  ��X�َ�m���|��Ԯ�)U����y�um2#4qЇ9Y8�=^U���>��Yr��ӷv�����E�}ݘ�T��GJZ���`��v��c�g����f��unǀHB�Ӎ[v[�i�;v����j�<�v<c�`�B/�7I��i[v�T��I���srO���ܑ_�h�4�i,�9��~��:��猳%*�a���unǀz�U=~����3 �$ym��=������$�jY��!F�ȶ{i;q�,��Ί�	�rGj�l"�WA �-p�i��v�RG�}ݘ�V���ذ	�\
T�cN�*��`wf3 ղ<�v<�Ȱ�`�v�+B�i]� ղ<�v<�Ȱ���}�]��N�������:�c�;� ��1����GJZ�L��+��n���X��s��������ٹ'����{ _�vBe�P΅��:��-u�IRdH:+�a���'Gr����V�u��K�cpϵi�Ԅ�����]6���q�6{[��c�����B���B	h�4�n�mi����P-h:��ȵ��,c[id"�0�f�"C��zlCH�}<H:������[6@�#�����r���C�&�R�K3\�Q�b�ͧB����� u�jTU�՗4[�̳Y��%Ay����j��nDӬ����x��ߍ��Fٱ���I�±�i���]�ҷ39�@�����V���ذ�"�;��H��*�"�m�0["x�K�{�$��pX�K����|�B�EN�'v�V���<I%ݽ��KT�<I%�v|ϾH<=�נ�t���4]0���Ė�px�K����|�Z���I.��_|������]Is��ߞ�ݿ|�Z���I.��_|�Z���I)���n�n�Ŕ�SH�]5�[o=C���a39.���8	4+N�eۦ�k�m6>�$�K�Ē]�ؾ�$�K��U|�K�ﻷ��<���XՖ��^��k��s����H�DX, ��)�@v�3w�����m����$��px�K��Ki�1&
�6[���%�\	%���}���OIww����\��r�2��� �d�>�$�9Ē]�ؾ�$�K�Ē]�B3�E�E�I+����.B�/bϒKT�<I%���}�I{�ǲ�wf�.v��#�Z�eZ�6��Ѷ�H�/=]\�:�[{-\z��sᵺWc�$�˞_|�[.b1$��'���%���z ;�O}6���Y[�w���#I}�||�Z���K�ofO/��s�qSﱾ�����]Hm����{�s����3v�S�@~�'�(��'�h9��^��@��jC7���F`�$"��BE�1BA� ?���6��B.�UbD��b1���8~�
���p��xֻ>"H@Lb��90 �D���(W���T�T�����HA�H!���޷!�l�!񠙌!a��0��$D��V��HH�a"�H�2��o�G�!@9Wt�:� �D���d�R� &�$8���:W��^@d	0J�A� !QP�����?�#���u� ����Q�*�m����"��o�s׾�<~��� ~�]徹R����^�Ur�~�Il����%�Lf$s����y�����P����U��� ��zw�ܓ�������� ~�ޫϒKT�<I%���A��whAC�eجJU�3BT�s�4H��^y-�6.nٟHß��䓓kՁ�Rm������_��$��d�>�$�K����\��ݤ��ߗ�$��3��m�驥\ހ߼��wߪ�����x�Ke�/�I-ND�\窯`�{i���ͮj�WN� ��}\I%ݽ��q?y<I%�<���I!v��Gd.V��/����}�{s޹�m��}���[p@� �  ��H�U� U�*�g�s零�����?����5�3&Mf�9e���ֽ��[m���"������^��X�K�ޙ�%�@V�6�����;y�s'9;N�kv�c�0���nb�as�����V���q.����$�l����$�ˍbI.��^�+�i(߼� {.�Q�f�[���t�n5��*���[.y}�IF���$�{��_w����⧜c�}ʲܣ����=���Ԓ����_��s�\m��?��J?o���X{�s�������ֽ���m���8s���w]˻o�L|��~;���h��sjV4��m����|�_��U���=�溒Jz��~�ZI/��n�g����/f�h�Ȣmcq�Nպ���Ӊ��\��[CX�n��\Ӂ�Ԃ�;�ն�3&^@^mb����l'���z?>�,8�L�r�Vrȃ#���-��z.���샛�vavgR�KBiڎKD�W�$�Ss��-�s[�-s�3��F�vr�ł�3����c����.�&!�ڶ��j�>�6Eh��yS��Ѓ0����'|z�B�uӳ���`��>r���2�=����=^Nnli�=�^�k��~x;�8�u,1vh��g� ?���t ~�y��`/���v�y����� y~~�pCM�c5�z ?y��ￕ�~۠�7�g��=|ާ_H�~�ޣW�v�ѕÞ� ��n�߷����9��I��~�������}�{�om�i�q.�Www�/s�ow'��������ĒZ���`rr+��m���e�l5�L�=����: ?�9�I���_}��� }��@���s�`Np�%/�:e�oaȽ1ؓ:t�Me��OFܚ�������!��A�rN<Ӯ���U���N�<��$��.�$�{{-��ܮr�m%���3��Ӂ��,ev{� =�ݷ�O� �k@�P�֥�u���p���z ?>y�����$��6���ƌ��u�4i��w@�￳�`�okպP
��k��}����{5�m��/R{�6�q��{��䓏����I-ry��I
lw�/Us�M�����I ���I�%����W��瞽��� ���� �����O7�� ���om���l�ն,E�6�a��h�9H���@�f��h�ց_�Z�~��ؾw?S[Te�p�� )��� ?~�{�� ��{_ �3-�g{��-��P��w�m0���ĺ��;��7�g��������$�����$)��z�\�m-�\�?X���]�� ��}^�Ϟz��������b��A|����>�n�?}��=����2��(�z�I"�����)��;�����>䜏Ͻ}^���а�+��q�`���x�K�Uٓ��ԏ9~0�"��ӞO&�e�`�iH++���14��U��I�0B�K6��򔶥?~�K��
wm�X��ݮ��~�o ٷ�Ƚ�|���o@���YFM=L�f�Wt�p�����??ߖ��ߞ������rZ{g�oK�e"5§@�����6=�r���s��	�~0��)�.�ջN�4;v�=UJz����7]�����V�`
|
#�s{�.��~t{���ӵE��v��췀{���>��� �6< ��KS)�nKnx8�0�	P�tgӸ��+�uvĖ�B"�<��}�rpe�\,5�L�=�OK�E6<T����W�7�޷�o=R��C�����f���*���~��W<�{��'����f�3�s����E�)��[��N�<��䷇��s�������+Z��%&]�]Yv��`z��o�޷�OK�E6<��'�&����^�����Q��ؙ�V��n�?O?���� �r[�Ns�����ֺ�]ˊ����C�s-\�ys�yX%FC��).�L���0]x?？6��6$m];=f5���;��+m;.�j��$�A6��) 겖ձ]n6�ً^�By��O�&T�;�;8y�)&� f8�8 &�m�t�Z�6zR�J[GJ���n��q�<w�a�s�B��4*N˨�62���`�]�SL�J
����99�����s���+��E���Tk3m�H�� ��tky/dH�eo9۝k��؈h�:웎�����um��/o�;���o �{��e9i]�nӷM;Wo �{�䷀N�� �lx��q:V�v�����䷀N�� �lx�ذ҇�;�l�wo)N�ŀ|�ǀN�� �r[�;�[h#��T�m;XSc�'^ŀv9-��b�>�F���C�]�I��Bk��G���y7!��x{qu����R�Rw糭B̤1:������,��o �{��/O<�����.�V]�֦䟻��}� >����V%�Q`'�d�s���z����;��vo�I�i���y4�]5ʻ�{�y��M�W*�UI{\��7�޷��h��RSV;7��$����{绠{�O,��o��+��9���w�_�^Ms3�����w�/@����������k�XSc�7�r;E�ګ����-��R���D]���!,�r�ih�f�746��y��99��y���6	G-��9$�����s� �l��\�*�A�s� ���+��t�.���ݼu�Y����W?/�������;���č�Z<�	5Am�m��<�<�	ݸ`�>����s���\���vݿ߭���� ���R���ƭ;x����o��o ���e�{绠}���6��
��vV��Kx�ذ�ǀN�� ޲�m��b2�%Dj�7%�;0`�S���5iF1�Iu�#���7e0v.��ӻ��s� �lx�ؽ������7���Lwe!��n����s�g��~x��~��N�y#����wui�;m;Wo �� �r[��+����� ��{��>�8�%m'j�����-����k����Usk�*���v��R�����rN���OR,� �����痠{9�I�?���@���� �r[�B���݁mU�t�v��=�[�����$4����E\�]�Ϥ�8�O��էm;_���E����W>A�~��5j৩5J�.�jӷ�E�w�\��UUj�?߭����`M�?s��ש�U�;uwL�n����[�'\�r�����<���<�y(ɏ(�#�2��rs�O�&��?~X��ߞ�xc��b�WLn+��ٽ���7@��I?�����_�N�g���rN����H%���0E:_�l�{p�p�M�R0HA#��>MtA�E��.���>@���!�v� ,c�V�C4"L��voi�.�	3��t����a��(0?
#�`b���504��� ��B�Z�v�#���	e�eŢ�!Q��H���J��9�6�6�m�V���(I��t�F,8� ض"�Lc)t:����tN��m��KK���;n�
����~�� �h~���}j����nь\����h:�L�FZ|g$��
�Г��v�Y�Z�������Q��Bh��\����5���W��̩ڃ8;͋�؈�Y ��(&L2Ҡ[+Yk-@��>�nzy��,�Gh1���m����6�O t=;`4���뜦ֈ^Zn!44[u��Dv�+�f�x.x|��լI��'�Y�r�9؛��/X��{	&.B�f��x����P�� �m�K�F�l� ����Kk�qb*@��Z��lS����i���Ij�֙@Ss��8�8P�!��敉�G�G��V�$|tt��)6�j�>zwO�š
�`�ݩ�&�Ԥs��PS�� �0&D8ZCf��&����ף��m���p�vv�L�Vƻu�Q B�4i�jy0Q�Yg�J����_?/�i��fjm[���d�Ꝼiͳ	:���Pc���3���*��H���������k��R.��Lj�\"�6:Ș�`�8���j��[�ݞ���`KXx��n�u�L�	�&Ga��Ie^��4;x�!��E�*Xu�,=!�4.�)�EF��5jc,�,ditgK�%Wa��O	b�+ƭ +�u���5�WJN�$���%��G0�Fmw;�u�M��v��'3@�(��[WR�/9��[`;2�֒��v��$S���=�����6��- ��K��֛!i4,�h���:. ��3� +�UJ\�.�֫���|���5�9Ui�*�Xӧn�^��=g��lU
��x�aͰ�0�<gd
z�PKF̵���\����!�bd���mr��=[�0
fW�]��56MaM�Ɗ�
�TBe�ݎ^�c�ٖtn�f�W.m]�Vs�9�ӝ��s��4���*AT;� �~8 =D��(��wK�1��E��n))�q���æ2����R��)SVyrtb��MuZ�]ˌ\R�]lu��]�,k��tkE
9����k9wZV�M�-v���1��$�,�Tt����
�m�hLɩ��b=!�� BMt�R1��c�k#[*�n�Hܷ(�1�&0e�i�N��0-���Z8�i6r{����2N�=�:��{A�ʾBc��>7i�=�:[>���u��yӭ�svː���)E�u�cx��=�U�2��l�*�S�Ms� �r[�'\���<�<����-v��Jl��}�y��I�%���� ����"ݏ?RF��X��ah���v�k�����r��� �?z���m�R�!�-[v۵��r�y�y�Ry��Kx�UR�߼�Z���!�����N��x�����������E6<t�(N�X��8��'X�a�h��X���E�4�ΣMt�8���NsL�� Q��0�]�>p�>���fӑ,K�����ӑ,K��{�͇���L�bX��׿�Ӈ%9)�NO?�����i]2�k�wxr%�bX��^��r>&��C�Ap����E��Ȗ'3��m9ı,Ow]��r%�bX�{^��iȍ�bX���=�2�.�K2��f�ӑ,K��{�ͧ"X�%��뾻ND���u�fm9ı,O}�z�9ı,O���3ٙ��U\l����/!g���=rwxX�%����k6��bX�'�׽v��bX6'���m9ı,O���`�]�C���|9)�NJr~���w��,K�����ӑ,K��{�ͧ"X�%��｛ND�,K�����{M��]�&�;fB�6�	�P����gk���Һ���;����	P�]���r%�bX����Kı=��iȖ%�b{;�f��~��,K�����m9ı,O?�ۥ̿Ƭ�&��5���ND�,K���6��bX�'���m9ı,O��{Y��Kı=�{�iȖ%�b}�V����I5�L����r%�bX����Kı>���fӑ,j@5CD�Mw^��r%�bX��wٴ�Kı?����ոd֭�m9ĳ�9�����m9ı,O�k���9ı,Og���r%�`D"X�､�B��{�=l+r�k2���	�����n	 ������Kı=�{�ND�,K�׽���Kı;���=�ô	MMI��(�E2���-�a�J�ڻ&�g����r�i�ugY�f�9��ND�,K���6��bX�'��siȖ%�b{���6�"X�%��w�rwy�^B�~�ޛ*��M�sWZͧ"X�%�����rX�%������r%�bX����Kı=��i�)bX�'~��z�M[�˨L��Z�r%�bX���ͧ"X�%���޻ND�[�����ӑ,K��}�m9ı,O�]��d��&�e�fk3iȖ%��'��z�9ı,O��z�9ı,Ow��ӑ,K�_��*��R�AdZ��1�� �s��G�L�����r%��%9>������E����ٽ��rS��b}�{�iȖ%�a������O�,K��u��ͧ"X�%���޻gw����/'�����ރ�J�7X���y-�r瀊[Y���jQ�񴖕~���f��զX�����f�ӑ,K��u�]�"X�%�ߵ�fm9ı,Ow^�� �%�bX�{^��r%�bS���{PFјZ�����NJrX��]�fӑAlK��u�]�"X�%����]�"X�%���޻NEF���'��%;=l%s��̫����bX�'��z�9ı,Og}��r%���b{���ӑ,K���w�ͳ��NJrS��_OY���;7�Ȗ%�'���m9ı,Ow^��r%�bX����Y��K�lOw_|u���/!y���zl�?[����3Y��Kı=�{�iȖ%�a� �>�߿��O�,K������ӑ,K��w�ͧ"X�%���REFC�Q��~ﭗ�f�50l�H/]Gk��dݛT@,�=]��$��t�7m-e�S$��X�Iwjۣe�����F;K«H�O(lZ�ӣ�[�,��� ��@cf���J<m�m�k�M��m-��<�
Rd˹��y�P�	�ӝ���b:#M��f�9]��;�j�麴;�G�-��Ͱ�Ȗ�[V�f���z�����K��6n�"��$�u;
"܎1	��^'i.��p��sa#����d��Ǝ4�naqBl�elÏy=���/!y?{���m9ı,Ow^��r%�bX���ٰ��L�bX����Kı>���q�P�]�w���NJrS���z�9ı,Og}��r%�bX����Kı?{]��iȖ%�g'���?laeöE�\��B����｛ND�,K��{6��`ؖ'�k��m9ı,Og}��r%�bS���G�cn
C"j����rS���'���m9ı,O}��3iȖ%�b{;�fӑ,K��w�ͧ"X�%9>��(�6����|9)�NK�k���r%�bX��{��6��X�%�����ͧ"X�%���޻NF�������s��l�9�i&?���*�>���1�9!���'761m=�^�jԉ�c<��V�k�v����%9)��������ı,Og}��r%�bX����Kı=���ͧ"X�%�����\%����W;��JrS����=�w�!�FDڔBPӸ���}�M�"X�%�����6��bX�'���m9�Y�2%����IsY4f����]]k6��bX�'����6��bX�'��}���Kı=���iȖ%�b{;�fӑ,K���������.j3!���ND�,��@�O��~3iȖ%�bg���iȖ%�b{=�fӑ,K��w�ͧ"X�%���k���rRM˫�ћND�,K��{6��bX�'��z�9ı,Og}��r%�bX��{�m9ı,Ow^���؆5��v4I�Č�Q�WSSecN7/��e�[�n8^�����~���Ql�r%�bX��{ٴ�Kı=���iȖ%�b{=��9ı,Ow^��r%�bX�~��L�K&�˭f�iȖ%�b{;�fӐ� `"X�����fӑ,K������ӑ,K��{�ͧ ��bX����ƥ�0�ˣ&���fӑ,K��{�3iȖ%�b{���ӑ,qD�D�"1U@�&ՊlW�2'���m9ı,O���m9ı,��y�y�Z�h��Y����%'8�'��z�9ı,Og���r%�bX����K��=����r%���/'����3�f�rwy,K��{�ͧ"X�%�{;�fӑ,K��w�3iȖ%�b{���ӑ,K���^���u��m�`�iۥ���]c�llC��]�s�$��B��N�0liG:������/!y�����ͧ"X�%���fӑ,K��u�]��Ȗ%�b{;�fӑ,K�����+3S&f�2Y��r%�bX����m9ı,Ow^��r%�bX���ٴ�Kı=���iȟ°Tș������?����h�][���Kı?�����Kı=���iȖ"ؖ'���m9ı,Og}�6��bX�'_{v�fx�0�Y�f\�fӑ,K�=���iȖ%�b{;�fӑ,K��w�3iȖ%��pP��@U"bAqD�w�]�"X�%�׳^�u���j�ֳY��Kı=���iȖ%�b{;���Kı=���iȖ%�b{;�fӑ,K��jz��C�V�f��;9x
�|씛���jm��x��ݠ#kj3�ZT|�'L�$�a�f����rS��bg����r%�bX����Kı=���`�%�bX���ٴ�JrS������4���:�Vn�|9,K��w�ͧ ��bX���ٴ�Kı=���iȖ%�b{;����Nr���'���Yp�JF���ND�,K�׽v��bX�'���m9�P�,Og}�6��bX�'�~�듻�^B����:Q΃� �kZ�ND�,AK��{6��bX�'���ND�,K��{6��bX�'��z�9ı,N�����E�5���fӑ,K��w�3iȖ%�b�{;�fӑ,K��u�]�"X�%��｛ND�,K���)��-`!�|Y}'2e�֍�]�Ʌ�1��p0�[�6�j,Ղ�X{e���̛��%���ڦ��01mn����"�D��VS�����n��H�N� pb�T[GB�W�vCNl=Ծ���mn��S�ڐ.� *���:�n2n1hr�.B�#��Ú<���.ɬwR&,٢��Z��:.צ+����:tt�l���{wE�/��:5n�F��]`
}��g'iؘ�����+�6aD٧6j6��h:^��Ǟ+�d��dT�x���982�7���MY��Z3iȖ%�b}�]�"X�%���޻ND�,K��{6�%�bX����m9ı,K��˙�|K�I�շY���Kı=�{�i� X�%�����O�P_�2%�bg����r%�bX������ND�L�����������f�a�\��B���������r%�bX��w�m9�K����]�"X�%���}�ND�)�NO����mrl1����rS��lOg��6��bX�'��z�9ı,Og���r%�`0ȟ����m9NJrS��{�S�ZQU\�7y>D�,K�׽v��bX�)��}�ND�,K��{6��bX�'���gw����/'�l��,�l�5KVsӌX7�cX���x����W�:�s���5�HI!�� �)��W;��JrS����|�w�"X�%��｛ND�,K���ͯ"X�%��｛ND�,K��}���MU��U]�O�%9)�NO��{v���:�mC"n%����fӑ,K���wٴ�Kı=��iȶ%�bw�v���K�f�2d�h�r%�bX��t����bX�'s��m9����2'�����r%�bX�o�m8rS������a}��T:��{Ñ,K��u�]�"X�%��=�fӑ,K�����ӑ,K�/��듻�^B����g����6��bX�'���m9ı,_����9ı,K�wƶ��bX�'~׽{���%9)���g�S�իKj;��R�`B��^<'a��ZXM�+XRY�QWY�sb��.D��	�=rwy�^B�y����Kı/���r%�bX�Ͻ���%�bX��wٴ�Kı>��ĺ��a����JrS�����m9ı,O����9ı,Og���r%�bX���z�9ı,Og������r����|9)�NJp���ӑ,K��{�ͧ"X�< t���,գ�X���QBP��SF���/�) ��6A�����z�]� }A��X ���D�M6H���Q�D�F�H�k_�
��/(.������I/�S��XA?+lx���`�+���ڄ��H?��^�T�PiF#��B�
����CI��U?QM�@0?(��TH���b~������Kı/���m9ı,N�ݾљ$ՙ�L������r%�`'���m9ı,O���6��bX�%���"X�%����ӑ,KĿ��f��]jM\�L��ZֳiȖ%�b~�w��KıK��[ND�,K�{�M�"X�%���}�ND�,K�����]MSg�q&�q�u�3v��v4����vF��t�nm��8�B5�h��֎:��K��?���kiȖ%�b}�o�m9ı,Og{��DȖ%�����v��bX�'|MKsZ��I�5�fkW[ND�,K�뾻ND�,K���6��bX�'��޻ND�,K�����r�%�b}��ܹ��5fa&�,ֵ6��bX�'���6��bX�'��z�9���"^���5��Kı?�����Kı<��;����&�˫�ͧ"X�(����޻ND�,K���5��Kı=�o�iȖ%���"  �lOk��m9ı,OOoƦ[�W&M���j�9ı,K�魧"X�%�~���iȖ%�b{;�fӑ,K��{�M�"X�%�ߵd$��}O�^\N�-5Ӹ#��`�z꒮ �(������ٽ���#;ҝ��(�kF���bX�'���m9ı,Og{��r%�bX��}�h r%�bX��{ƶ��bX�'s��h̆�3F����sSiȖ%�b{;�fӑ,K��u�]�"X�%�}���ӑ,K���ߦӑ,KĿ���Z��f�U]�O�%9)�NO|}�����bX�%���[ND��,Ow���r%�bX��wٴ�Kı?{^�.C-�d��ɒ�WiȖ%���}���ӑ,K��}�M�"X�%���}�ND�,K�׽v��bX�'�&���`�@��6G��JrS������6��bX� }��iȖ%�b{��ӑ,Kľ��5��Kı0A�C�H�{��gٚ�d�asYk�Q�p1�4�ngb�����W�78�*SVN�d�;��/4�������u�n2DÝAt3OYCPL�y٘u����ݡK� �(���gBY��GL�Sev���6�S�s���I������.�
�l��ô��v���vmTa$m�	Ŝ_E63�����D1ka�j2[d繮Y4���iYl#JZLԹ���	�e� ?
��ɻ��I�f�ImЗaź.2�򌌢Gn-�vs'�&��r,�'K����m�4��T�'�%9)�b}����r%�bX����Kı/���r%�bX�����r%�b��y���Q)k6z������Ow���r%�bX���m9ı,O}��m9ı,Og���r%�bX�>�ߍeɪ�f�5��ND�,K���"X�%���{�ӑ,�!�2'�{�6��bX�'{�]�"X�rS���=��(�-Wd{���X�'��ND�,K���6��bX�'��}�ND�,K����ӑ)�NJr_}�{X�&�L5֬�'Òı,Og{��r%�bX�g��m9ı,K����ӑ,K�����i�������o���h�j�Q�9�E��K ��43I��㒜�tGfOaUmLWZf������rS�������oxr%�bX��w٭�"X�%���~�ND�,K���6��bX�'~���Zk�֎:�������<�ߝ��(@> ��@v��wı=�o��Kı=��iȖ%�b{��ӑ,K���׽&Yf���[�fkiȖ%�b{�o�iȖ%�b{;�fӑ,~R"{Z�ӑ,K����ͧ"X�%��!ӹs3�j��Mj�j�9Ĳ��{�&��	���]� �'w��pI�?w]��r%�bX�>���5i��j���fӑ,K���w�iȖ%�b{���ӑ,K���w�iȖ%�b{;�fӑ,K��P����	O�WZP��a���:��f�GL~�l|X�Z�l��C��4��{H���4]����O�%9)���?���ͧ"X�%�ߵ�]�"X�%���}�ND�,K���]�"X�%�㤝=�j���4]d�u��Kı;����Kı=��iȖ%�b~����Kı>�}��rbY�NO7���R��5aV����NJ%���}�ND�,K���]�"X�q�8I$HQE��"�0	�ィAx?�dK���[ND�,K��~�ND�,K��}�Y��ukh�
��|9)�NJr}����O�X�%�}�}5��Kı;����K�,Og{��r%�bX��S�d���3%˙���Kı/�禮��bX�)�w�6��bX�'���m9ı,O{]��r%�bX�� 9��@��>z	ѭ��e�bQ�Ѝ��	��@����\��,�J�1&���nͣ�Z:�����NJrS���{�w�"X�%���}�ND�,K��}v�Ȗ%�b_���[ND�,K�:z����-���rwy�^B�z��iȀ%�b{��ӑ,KĿ{��l?�'�ı?����iȖ%����xF{��P�n���'Ò��K��}v��bX��s����m?D�,K����ӑ,K��w�ͧ'%9)�NO����p\&F&���O�X� %�}�z�iȖ%�bw���iȖ%�b{=�fӑ,K��0A�D��w�iȖ%�b|}!�r[5Mj��u�]j�iȖ%�bw�w�iȖ%�`��=�fӑ,K���w�iȖ%�b_w޺�r%�bX�����IQc,�,lf�v���������Ś�=]]��l��;&˥�y�s�6��b��g����r%�bX��wٴ�Kı?{]��r%�bX��﮶��L�b[�����N�!y�^O?��{�p;\�ff�.��ND�,K���]�!�*EAșĽ����m9ı,Ow���ND�,K���6���L��,O{��iXd�rwy�^B�����m9ı,N���m9ı,Og���r%�bX�����9ı,O�A��\r����y>�����P5�����Kı=���ͧ"X�%����ӑ,K� V	�3����ӑ,K������������55��ND�,K��}�ND�,K����]��%�b_{��[ND�,K�k��ND�,K���@
��O�Iy$��ΞZ�	�,�f�F�:`Nz�?#,�n6�+w�Ɋg�4� 8�ָ;Dj�f�qt8k���9]����q3�;��!]؍�ٲ��È�;>��� ��:�vU��g����]F����-�k��j��̉���#��m��3y��=�֧�z�]�:�^�r�x]7�ɛ�YWe�RXa���E�콬�Ԡ-�[>����� T!�o%�w�3Yd��f`�p�f|v'90e�Z��f�|v���[�Wd��pTßy;���/!y>��rwı,K�wƶ��bX�'~�}v��bX�'s��m9ı,O�C]�-&T��oy>��%9/���{ÑKı;����Kı=��iȖ%�b~����Kı<vC^�iW-*�G��JrS���~|��9ı,Og���r%�bX�����9ı,K�{�[ND�,K��������aV����NJrS���ͧ"X�%����ӑ,Kľ�u��K��	�=�s�m9ı,O?����M2eڛ=rwy�^B���w�iȖ%�b_��f���bX�'~��6��bX�'���m9ı,�>�Ko>��ղ���ͰE��Ýɠ8қ'<,r] �Y.a�[��c�i���f�5s5v��bX�%���kiȖ%�bw���iȖ%�bw=�f��AI�&D�,O�����Kı;�k�fYHk4K%�k5u��Kı;����8:�<l�Ȗ's��m9ı,N�]��r%�bX��﮶��bX�'�wr��Ĺ���55��ND�,K��}�ND�,K���M�"X�%�{�z�iȖ%�bw�w�iȅ�/!y<��O�1ڷa�\��B%�Ȩ�ȟo��iȖ%�b_{���iȖ%�bw�w�iȖ%���Ȟ����iȖ%�b}�k�Ʋ[�ja�.���ND�,K����ӑ,K�������~�bX�'�{�6��bX�'�k��ND�,K�A��̧2��<;w�.<]m��y�;x!.*�[���������m���x�����W����bX�'~�}v��bX�'���m9ı,O��}v��bX�%��魧'%9)�NO<|X��e­�'Ȗ%�b{=�fӑ,K���w�iȖ%�b^����r%�bX��]��wy�^B�y��=�7`]˵6z�Ȗ%�b~����Kı/{��m9��8 D B Hv�T�bn'��]�"X�%����iȖ����y���1����rwy��@ș�zkiȖ%�b{����r%�bX����m9ı,O��}v��bX�'��w��	K��,�I���ӑ,K����ӑ,K����iȖ%�b~����Kı,���+㔎R9H�Ip�um;C�$k:]���4JW[���37 <=�c���ڳ�x�{-���{u�Էh
Ds{���%9,O���6��bX�'�k��ND�,K���ka����L�bX���v��/!y��ךC-[�0�N�%�bX�����9,KĿw���r%�bX��]��r%�bX����m8rMy1�NO���3^R�j����Kı/}����"X�%�ߵ�]�"X�(�0"dO���ٴ�Kı>�׿�ӑ,K�����dֳ&���̺�ӑ,K�;����Kı?g���r%�bX�����9İ?#:T-�����t�E��D��ﵴ�Kı>��HED�XU���rS�������iȖ%�a�(D>�߿���Kı/}����"X�%�ߵ�]�"X����=��k~h\ꅙ��Ͱ#
��X�rn+lF��뉶9���>-�Ss<+t:e�W.�5�u��r%�bX����m9ı,K��{[ND�,K�k��^D�,K�{�ͧ"X�%��ڞ<a5�Y��ə�sSiȖ%�b^����rbX�'~��6��bX�'��}�ND�,K���]�"#�2%���뼗�B�����rS������{�u9ı,O���6��`ؖ'�k��ND�,K���kiȖ%�b~:ww\z�]�)��O�%9)�$��������ND�,K��{��9ı,K�{}��"X�-���ߦӑ,K��c�޺�d�3V̺���r%�bX�����9ı,K��{[ND�,K�{�M�"X�%��=�fӑ,K���<���4)�pj���'ƗWĈF���*DglC���l�+� A8������&�o�M�jT*�,dD��		�$IH��"%7��C����7�$p_�U$M���$`�$����F���?ly���2�I"BUrM�߈����$"��>y�K�iT�������"�*?��p��τ�8Ȑ*&~G���l�Y��k�B�a' ��S�Ӯ5Bu�;[����5 *��V�J)qS�Ys�[J�T��`�*t��%+`��ʀ�Fx�&�� +�hI��1�[]*�v�Ȫzȅ&�Z�.ծ�iY�7�Lt=�am��v�uf���D�,�j$�6�x+3b�j�C��S#��WC۔�e�Sح���Ge��+d�A;eX7Wl����RT\ �VX-v-��$9eeZ8�F���j]����J��.��m���M1�F�g�\�N7Y&Z�;u��]f�ɃI!�0��q"I�iwN�i�1�c���C�Q�aEZ�a�fČ{60�=��.T���v��mV�=u@\�d{0�Էu�\�S��Z��UT��,-�a�]m�㱏í����m�{-�:�m���(��u��2�Jq�����r�Bfΰ��re-�Gb+nΙn�[�R.M�"cV�kY��DW.�5�sBM���t�hC�`�r�,je��C�i�����C�Ljx���T�.sX������q�'=��T��]C��8qӢ �U���л�ٌ�Z��H��T�C�c���ע�g�J��+D����e����ָ��K��5�`,P��qt���K�3ۣb�lT誛Y S̷�jZel6���X��ո���yYƮn�)�ȱ<���6�F�5G5�%b�`�wa����F��M%��t�D�����^��n&Uu�X'���-<N��z�q�q�B¢�;<�l���!�a�݉Γ���xWh���Ƶ�ۙ�n��<(D��ji�j�M,#�H��8Fs��-N�kMA40��:�Sj���;rŭu�[)��%%e�g���'d�V(f�^JͣXV��B!�Gin�Su��ͣA� ���+j�]֛PvޢS3f��=I-��	�,�B1&ex�d�0��E�հ��d��{N�i��͔���s<��PLeW-�]S~䓩�,�|�������8�Q�~�0Ta�� U?
� >Dq?a�}{,��nf���2��n�!RC#]iM:�{Ob\�@����Jشs;u�w�f�׵Pmk��ak�u�l���.���8�m�֘1@�9[l��ғbVm�l�΢4@Y��9(��UC��x��v捓�`��\��EƓ�TD�b��+i�lV������x�z�W���.t��]Y�,�q�J�8��򂎙Ҡ`�s �_�rI엓��u{:-���`����F�ɦMg)��p,l&cƎ��j�ʻ�t��I�kZirۭf���Kı/������bX�'��~�ND�,K�w�ͧ"X�%���ߦӑ,K�����Y�:U�E�'Ò���'���y>	bX�'��}�ND�,K���M�"X�%�}��m9�ʙ��������rS��������m9ı,O��m9ı,K���kiȖ%�bw���iȖ%�b}�������2��|9)�NJr}�w��Kı/�v�[ND�,K�k��ND�,K�w�ͧ"X�%���}��¼v�����'Ò���%���kiȖ%�a������O�,K��=���r%�bX����6��b[�^O}�ڤ��fn�iŚLm��\A��X�zQG�5�2]�U�T��{A�NӃ��)%�Y�Z�r%�bX�w���r%�bX����m9ı,O���6��"X�%�}���Kı><{w.[ZmH
���rS���������O�͙���MD�?}��m9ı,K�뭧"X�%����ӑ,K^O|��߲D��
�s�'w����?}��m9ı,K���[ND�,K﻿M�"X�%���}�ND�,K�����u��ir۫�M�"X�%�}�}5��Kı>����r%�bX���ٴ�Kı?}�p�r%�`_g�﮺��*�5��x�t.�xݗ ��^:1T�*;c�e�6�j8�pT��Y�)%��؃�':�N�-��j��dR.��jۓ�y~�t��X7b�� ݗ� 吏S�e7v6ҷl���}�"�URA��+�7e��"��kiʺ��E�;n�����ܓ��f懪r��i��V�xdVȚ���t. v�^��)��G"��*��������i���hn�젻� �lx�ȰM�x��0��#U"1+��.Җ����	Gk;��kl�a	s��V�mTq��*Whm$�L���-��M�x۷)��ڂ�Vpn�WI&�� I!y��)#�_���� �n��<���8�Z&�U�^����àE6<=��Uq.�<���W�w�t8)�r5m��������>�<�t���[��;@dG�~��ڻ9��Oӄ���|�繋���m�Wwo �I I�� �ۆ��/�yy�C�6t�k�;K ��^���gD��u�/WdJx�������B��涜6���	6^��)��{����y��+g�Ĩ�t. i���p�W+�^�x}Uʪ����< ��� �v��Pv�M�]�v`M� �I I��ݸ`��Kb�v�-;x�]~�� z{׀n�� �dx���U����]$�v�l��n�� �����9{���8*��$�;a�F� D#���;�Ѳ�`m���$j	qVy}��9�,�yg`���Eh��f��8,�K��|G�g�B�7k�I�rm�s��iDH�����nM�` �$��.�̥���B�Cf��˱-��.R���n�ۙ���6Պnu���6Dq��]yx�]m�)=�"Ѳ^m�t��D�a�[����&�v��x�ZP���=��P���Jp��t���/g����l�<�]�VTta��	�\�ml�[��h�U^����àE6<�$x&��>ݺ�*��e����Sc�>RG�l�w_���Ihy��k%34uU�����	6^s�n�XM� ޱm1'��4������{��|���� ����ȭ�6�E��qWw�n�� �H�����^ W�mi<�[����J�H�v�[s������d�ԦM�J͛%��̥��qS�yd� �I M��ݸ`i�Kb)��n�e�o �I_+��*�r^��� �dy�׏_��n�+6����^��)#�>RG�Jؕ]9m�[Wwn� �ۆ��)#�	$��ۡ��Wb�t��N�)#�;�r�䷀l�w_��'�Ͼ��Km�.�,�J�j�9B�[;��:�6'Fݫ\ ݺ5�'���}�.��.ˤ�j���W��Ix��0�� �f��j��[��� M��ݸ`l�� ����O��:T[�;��wn]���>s�u oP	��,U�"�+���=��� �v��Lq�n�젻��/=����y�ݗ�n�� �N��C`�v������������.��	��:N�X��ЊJ�k�pu����}���ŹPi��B��V�e�F�YHT�X!�o�l��I��C���Ӳߏ��������?65&M���	$�ʮdxRG�v^{�R!��)[�T��n� ��y�I M�x�e`�"��umWt2ڻ�x�)y��x�=x�e`�� ,b�~Q/u�o7$��>�ܚ���[��� N��\�\������@���<)#�>��-ZN�4镄�
0�Ce���X�W�̢3��gU�ě���&]&���и����7v�Eݏ �I�_ =���[R�I� m�]�v`nǀ|�� 'd�wn��&�N��j���4��^�� N�wn]���R�Y�M�
��x�^�z�	%��69�����9�	�{ﻠy?ylq=�Z�:����p�=�����u{�x�K�7�Tv-�H�@b4��<�M���ck�e��.��iL�t<��.�ͥ�,���:���-�e��a۞��+��p��an���6%i�t����h�z¢�;FZ�����j"��Uj؋v�ٞK`��2:�.�C`2�g��gi�7ٞ�͹��-�j'n��d9�� c�b�uwN�u�ge����{e�>\&�heB4��]�{ǮJ�tR�6�sܜ���$'|׺�@Sif9�u�2� uu��6�,�z秫�m=�;a����;.�M�m*J�'g�v9�< �%��p�;�U۫j�]Ћv5v����엀n�� �r,u�NSV�t��bv����/ �ۆ��X�H��U�Ri*-��wx�e`�E�E$x��xk�����bn�줕�`G�`K� ov^$�X��T�Rn�cl�L�+˞l��[9�.�KU��g���DKx�MvIWk6`�sz�o<� ��/ �L���X�K�g6�+$��ݗ����u\�R�+ �r,Ip�RD��U�<�v1�j��������}� �Ȱwe�۬p���n�bWi;0��`G"�ݗ�n�� �!�v�˰wBV�j�`G"�=U�)���K�}Ł~���I�o�u��J���6��1��F��{.�eɣ����K��熛�\�h׊��컳�	�׀n�� �=� ��X{�[#h+wB�n� �n��X�b����6�R�P����(.��>�b�"��_��r�������6eC_JVs�5�"L�#���Ǖp �"@���Fl��.�(���(� ����..���B�@�����#}��U&�mS;��T���À)��1N��;���uP:�"@��?�	E��
uQy3���䟻��N���6`�[��E6< ��x�p�>�b�>�K�g6�+�v�{��	6�}ŀE6<{P*�7n۶�
�g�v�	VQ����Y�A��\�Ŵ�n�ڬ�Aי�tڻ�w�K�}ŀE6< ��x�p���mؕ�N���Y��^�x$��m� �!���v�v[��k �lx���	6�}� �fӁV��ݫbt���ݗ�I���X�:s���*��PȰ  8��G/o{�7$��]d�b�Qn�\@���l��>��E6< ��܌�!y/+�n�$�aVq�L3��6���㒻c���ڳ�q�!��0���I7AvP[���_�)���e�l��>�*����+j��"� ov^&̬��,�Uq#�+��)2�v	4���׀I�+ �9��_ �"Ut��n�6��]��Oe`G"�${���o�������oሸk�U�g@�����${ n�M�Xj��J��Vr�U	8�y��危a�%4fj uf�ͪbݝ�m��Z882���޸0NkL�+-+=�k�w=��ɴ#{r]�q�V:�Ԇ�j���Zt��=Sڧ�k��]b�@���2L	m�[��a�f
V:F�
�o)8ʜ���WMդ�Dgv�٭�V��Hz^��]�f��K�e,.�WhY����]��S��.I9>���8s�G����p"*�4)HҤg2;��@R]a�-��IR9\��]��:-�%nƝ������/ �fW��|��{Y)�����ձ:N�����$ٕ�}%� �ly�W���+g��
�wB�n� ��߲���a���9T�����l��]�i��V�n�젷u���U�{��~0ߟ�, ��x�2��J�ci�`��v`=� ��W*��r��~��_@��߲���`�o/��� �kmFh�lD��GsۮE �`���7]`�Y�����M��/4����ݗ�I�+ �K������*ylfeڣ.��z�~󳽒rY�& J^�?������'���:��������#c�ڶ��Ip�"���H�z�z{+ �!���i'`Z�e�f��we�l���.��� ��S�h�[�llN�����?W�=�|}��E6<���¾�U�`4��
-��hC��%�^��ْ��V����z�(��nǍ�]�&̬�ˆ#ذ��x�jZj�]�7AvP[��>�`�����7d��>�*�1����jnI�����'��w[��� R��  �F��ݛ�~��t�>�9*�bLX+v�`��x�X�ۆ��[���*D����n�t�]�wx�X��<|��� ;�绫o�C�[=M�-�K��i�������[�U��2ܒ�����G7m21��N�Wi]��v�v9 }ݗ�nɕ�wdYN݅��MYmـvK� w�/ ݓ+ ���N�i�,Vʷj��ـwe��e`wnd�`ݶҜt��t. .���2����Ȱ7���t�r�ݬ�W"$�⦕����7�nI��ڹ|][I������v�v9 }ݗ�nɕ�z�<�� i��I�M��8�����%)0�����XRX�e^S��p�t��Jڻ>|��we��e]Ub��+ �trU��5E+nݬ ��/ ݓ+ ��2��"��=��Sd�$�y����M�{�X�۫��� >��Kj+����c�+��� ��2��p�����2��)�˱զ�����\0��x�w�7$���f䟸�
n����)�]p�Ul�+g8ٽZ�9���&��É���Q!T�u+*cd-���R{$�P�n���J���d�v��r�l��b3`��y�c�3+��Tp�0u�P4��j�[�W�Q�
�!*��Ix�rK;�#Ě:
�����:�֙+6yɛ��Z���t�y��i�{7h�bÞg�A8�a5�˒etj�fbEy���9;ޑ:e�]��v��'k�<Zݹy�Y��.�ɪ�s',sۏ*,e鵵�#��0ym�~�݀nɕ�}�2��"�>ݶ�e:T[�H����&V�ve`�E�>����$�����Y��偆�s:v{+ �r, ��/ ݓ+ ���dclh�]���U-��� l��vL��ꃒ��$��Jۻ0����2��\0�p�=ʒry��Զ|b� 
ŦnuX�}��Q�X�۱�&ۢ�����1�ج\��c����j��	=���\0we�I1�Ӡ���յwX�\0�)��r�uUB;%� ;ݗ�nɕ�wt�E[�ݎ݉�[v`�E��/r����V�z�`�ږ4���l�Ӥ�� ��x�X�\07�9�������;_14�s-%W�nɕ�}��v9 n��R�^[fʉ�15�qmQc2L2µRY���M*b]�jLh��,q�I���]������.d�`���W�$����{�ci�l�]�d�`���7d��>�p�>�85I5E+�wwrI�ﻭ�>��ٹA8���/�"�iP�D&&���m�����@�LMX�����&V�ˆ��X��x��Km��[j�wX�\0o��_ I=x�X�Ø]Ҥ�ZN��y�9{66�M�b7��8�ڣ���l��(�����L�\%rt�o<� ����vL��.�6��+���-��ݘ���ܪ�x�6{������;%�=UIe���$�)ww�I�e`l�`���/ �i�]Yi�S���ˆ��X��x��pݓ+ ���H�6`��v`�E�ݗ�nɕ�}��y�{�'Y�hX�F��Q�aݵ�����n8���Bѐ[���yr�RXJ�[���%��7d��>�p�;��?x {3ƱMkշ�rNO}���`w޿c�`�p�7e�t�U�&��VӺ�>��v9�W8���`{�Xf�(�v��v�ݖ+v`�E�n�� ݓ+�UK��x�=����j����	��7v�nɕ�����ܓ�s���VF�nd��0#�B0�!�B@���B��>�$�# ��H���$$ HB����$�,i�$�22����!m�		�� @ ��B�/%�H���Y�A$$'�(m0lΨ��I��5��:����C���R$bB!�d�6t����6�#������D�v!�� Ab!����G�`�$�"D94����٨$F!		��`BB@cژ0>4�H�0�)!�H��!�T�Pb $` F|o���r�#!$?�e�8��O� U"3?.���	��ف��c��D��"�hMa��a FX�G`=���ښ� �ZT��0#�	�"���BE� @�dc �bD���$�;��E��[#"�`DI�$RT�@���aD�B0$Ed!�a#F$!BD���$�ddA��$����!�䤐��[d���)iB �	a!!HaK)
B�$a1��HB	ā�a���D"B	0!2�HB��$ @�Q�H1	 �0#M��+X"�}Ns��s��@���o�Am�%%Vmx_4�
f�ӷF g����c[p��lA(Z ����[gR��U�V�4��b�g�vtm��SV8�tl\:�6�v�vT�kR"����t�P���#�R��2�Y���nvѢ�}h�Z�W�ں/�QNQd�$��qU�-y�ͷn���SN�u;�<N.���)�ᣞ���k��:����R9�U�"j�]����*��k�4���Zve�t۶S�S�M���n�cQ��	�2��M�Ma��b|��pGHq[I�ƛ�2�n�q����@^�eM���ZH�>�ɻ��d�f�Rv���Ʈjum��"]�����g������D+A�ηh������F���@p���q6��ƒt�t�] {@�M��]�c"q����0�cJ&����k���Ü�DiLm͆:P�մ��t���"|�j�����M�*ꢐiR[�nc1��sϮZR���A.�f�Vn2�:���C�6��ԧe
����*r��\-�*��H����V�[
�vD���Y��[�5�V9]�{X)^��n��:����v0�U�c����4Ҳ�Óve"X�l<���[��/Rq�:�B�x2v�b�ax��N&jܱ���"�z�^vG=)
���7*�8�A�)�p�t[�J�,֤�)��ۖ������P��+��իQ�&6ErGp���Ӯ��ݠ4�6�%�MR�ʙz�)�ՐS]O���E��NĮ�t�nR&�ґ�c��g!�p�H\�s�;���\v%�AńA�hZ�V�.Z�����Y�n��V�ZD)��@�]QŻe��,gZLUԙ�l����z�$k&�[���xL
�T�d��Z�R�.@��V�EEf�47<#�6���%X����4�A���i�Z�(�j���G�p�m ��R�m�"&T�ڡL�tY�-Q�;Y��{f٩6�5(( ��J����� oH���9�Tz� �I{��A�	�)�_��N*��>u�����X�N��3�-�j"�l���;{T;�X��	V�)��"�]1��bs���N�k���k�x���J!����ӌ�[׀�n;�ϐ�:ӭp񶗝�!{�ѱ)��0�s�0N68*�K���u�T7a�$ڲ��GID�5�4Z����;&���+	�����]3������1�M>Ƒ��^���v�t���/g����z�}��z ��G��M;iS$:C h�k<k�;7f���bM�M�v퍡Qn�"�t[� ����>�p�;� ��� 셎:�*Ӱ����.c�`�p�7d��>�*�Sm��V+� �r,wnz�������;�_���P��)ح[��n�� ݓ+ �K�W)v\� �H����,�m]'v`�e`～>|��n�� �mmB�}t�l�F��p�`%-9h4�A|�]����@uų�.���6�3C ��2:wm��_��\0ݸz�Uʪ���V�����mÚթ\��>�s�u��2I�2��\0	�m8m7E�m�I;X��0�2���`�E�}�l��H-�.�n�vL��.c�`�p�7b,je�aL,wX�\0�z����.��/��&VݩT�⤝E��sI˥I��
�C��-]]F{2T:��6|�c�M���J�v`�E�wv�nɕ�}��}�9*�	��V���;�p�7d��>�p�;� ��U���ݕtڴ;� ݓ+ �K���VVF+G}��n�Ip��@���cl-�m;�Ur��=�0����ۆ�&V٤�)]�����,���;� ��� ݓ+ �K��.�UA[��`�m�˛`KU���F��t��[�e�	t�-m���6]��E�m�I;X��0�2���`�E�}ݶJM%E���[� ݓ+=\�9Uʤ���� �?y`�p�7b,j��j�-�`Ip�;�r��_�O{+ ���"i�$�%b�0�"�7v�nɕ�ڮ��۠T/{�M�?=�ޚ!���V���7v�nɕ�}��v9������n��k�����A܎Ҹ5�ZF�P��B�k��{	`��%.D�2�t���{�X�.c�`ݸ`H6�:M���7u�}�៪�����,d��XfŔ�]�VJ�[� �r,wn�X�\0	�l.��E�ln��`�p�7d��>��vK��v�)��[�RT[� ݓ+ �e� �wn\�Ҕ�V�7VX�R��A���
o���}��ف�a�`:�S;8kt�v1�S��BZ�#!Zr���3�^+B8�*8t�J�'��d�pD��^Ğ���d�wg�#�#�[UYQ8�L��鎤N�ҩ��ۭ���Ye��k>� 4g��z�-���-��A=�]������t	�=�vI�6�"��͵�����W����Ō*�!�J�\�e'Pn���n��QK�V;YH^ZҴ��j�-�|g���.wn�XܥRF�`�@��v`��wv�nˆ�ˆ~�H�?z�b�N�i]��~0�p�>��vK��n�lQ	ڤ:m]'v`��}%� �r,wnR0�M��M ��;� �K���X��0�p�=[� ��b�4�f��{Y$�&cy�ȳ�H�V���3v-ź�)K�L-]+��+�>|��n�� ݗU|�����=��-�m6�e���ܓ��f�]�� t՝�ٹ'ݗ�Ȱ�m�q�-ة��f�.�.{�ķ޿�~0�J�M�M]�����.�p�7v�l��R�#i��%b�0��n�� �.�\0	H��yo���J�IFh��W�]s`8�	�J��,xҰa\�e*�-��^��6 ��o\� �.f�0�E�w��[��T��2�7k �.�`� ��,)R�Km����wz��s����>�w�r��!�pEdTSc�Qbl 5>�>�ܓ�fV�E��2�vNҷj�`ױ`^ŀ}�e`�E�ld���Uhln��`^ŀ}�e`�E�w^ŀlu�!ā�j�S|j���dIp��V��ٮْ��Vd��e�5��[�RE���}�e`�E�wv�M{�)Z)7wt�I+��'\�%$vK�kذ�n��J���L�%Cv���Xױ`n̬uȰ�rR�BM �V���&�� �d��'\���Uw�ױ`�V1r]��L�M��>�2�	�"�;�b�&�� ���g�B��St�tq9�怠܌��q�,����=�ֳs��.ԩ�m��J۫wu�N��{5�^�r�A��e`���T��][��Z�Xu�Xױ`l�X�`)ƒ�M�e����M{�ɕ�N��{ݖ�I�Z-ݬW9�R���k����� ��,vR��cN�j�Wu�N�����=��>ݙX�*�UG9�I=�=,�ʎ)�lŅrL��hBml�lQA�q��ϛ�Mk��$j6���mv�\�0#q^8omq�C����hS&��tl�[DU���ӷI�Lh:v�3�.�=�C���Zx��A�vݶnй�t{ZWrݳ��t����
��Ӷx狮x4�&�\+;�~�q�Pl\P�)�pJ�&Y_=J�k�Đ�iSm-�&����p����w�ճ�9]���vu�8�& �Aac���hm/6��e^RBU�ˠl����y`�b�>ݙ_�ϐw��X�s���M��V���7^ŀ}�2���`kس��q#Ҽ���z�)��t���vOe`�E���q.�<�G<��t
�lI[�Wu�N��{5�X�&V�E��1]ӷb�j�`ױ`^ŀ}�e`�K�?~�<�E���lJ�+f��'��M��nn�ɦ�̎��s���k�v.T�ln��`^ŀ}�2�	�"�>ױ`�lR��[�qX����}�2���A�:���w�rN}�v�I5�X�h�.Ʈ�j�Wu�}� �^ŀn�� �ve`�U61��6�v���Xױ`n̬uȰ	K�V���Z�k ��,�ٕ�N���� �9��Ʌ'A=�
m��p��9�ͦR19wX9��+J�1�9�)aѺ )j�n��;'��	�"�>ױ`^ŀE#�T�cb��wX�`kذ	�b�>ݙX�<�I���v�jի��}�b�&��]�uVr�*�Ю
���\���4
T����]�^��P4+����I����d�����!�-(HS;��r�wP��$9�X���R�H�XX1 �+@h�!���y��d�w"}��&w@���l���8��ȥ �M��X!�x�1�M����Ǩ�ELUM�π�@@?
u8���`��8��h� ��P����\E�}��L��`k�g�'�(~�]6ղ��	��=��>ݙX�`kذ�Jc�E��[�X۳+ �r,�{$�`l�P�t�jp�T'����y�m�/>۱ʜ���p:W x��Ͳ�Tj��e�g@��痠|ױ`K��� ���;T���i��[t]��>ױg�#����=��V#�`�6�,��V���$�vL�G"�&�� ݨ��m�n�*�˫wf���U/o��`���5�[�[x�4��P�
�t�*����M�9{�S'Ma�r۬���#�`^ŀI.�X��	:�K��B�V#����K�����D���+(+JWtrK�(��M78�b��v�	�b�$�vL�G"�;��9E��v�ct���$��RG��V�?y`vG��6z��m
�v*E��v`��X�E����%�������>~�V���3�ٝG"�"� �.ݙX�J�D6$��ۢ��dx��Mٕ�lr, |�͕VU�N��Se9}2�B��4xA��.�e�ٻ*�O�P�|��lq�]�b�h�^:���է�Oh��T�.��,������G8K��n,	r�]
�m�g����uBWA�-�C��A��k�x���,;�F4FUF���t����(�0u���a���]u���d��Z2��wkk���"v����$!�3��;��b�1Q��䜒u'M��;M����5M���'ʛ����՚.�`�20��f�A٬�9� L�v+�v��_�n̬c�`vG�M���t۷wUueջ� ��+ ��X]��%� �\��ȭ&�I[*Ӻ�69v<d�`�2�	�<�I���v�j����K�g�=��N���69�j��Z���'v�	%� �l��69����h���b�IP�86����Т�Y0Za��Vj�Fԅ��K�ě��5:7!E�"ҥn��+ ��X��x�p�>�J�⺻�2����s����H�E`(��~M`��x�\0�&V�R�"hhCam�ݬ���\0�&V�Ȱ�ʺ8���]�s�ʥ=��w}�G"�:����WӶ��Yun��>�2�	� �ݏ �\=ϐJ�
��J�.�T�j�1_.7�^;v���̜f�����űve{-� M/�m&�E��wX���j�ǀl�s���V$^�)17h�V5j���5wc�W9�$Oz�`��V�ȳ�RN����bW@ssV�V�~�}z�s�wf���JI����`�,"�jN��F "����<�-��E�"ҥn�.�{��'���]��	6e`mJV��v�tZ�ۺ�${��&̬�ɕ�}*�XSv]"��1��jظ�I\�3hm1�����H�9P�;L���[��@�Am�wk ��ǀI�+ ��e`=� �q��I��Wj��l��UUW�x���ݏ_N@��>|h»1���[o�>��	Ň������x�{+ >�@��4��hV����,�����ܟt�\v��~�9��9���E&&˲��j�`]���L� ��^��,�Z� �[�-S��j����ڕx�x�!�0�YO@�:�|Z�,Q�]�m�t��[����ɕ�vK�;�b�:�����)�*-ؑV�j���xcذ��x�L��J�M��t�M;��&�� ��Ǉ���)/o����z��U$mR���ۢ���ݏ �fV }�/ܪ��\��'�9�+T7��]�M�X��w޿�����:���\��*���$T(4 ��B
B1(JE��Th+��gd�.��f5�c@7\u�S+:����1���M��r:��i���]t1�rr������첷7lV�½h�Ɨ�7b��.�hDڡ(뎙
tE�[9ݵ�Kb�VU�c��Ge��8��m�� �-���X��! ]�קh��ؼ]2���k�t�l����Ti��ܷ��L���f�(������L-q�i5��b�:�a�b�#����Q�[�kY���I�b����Vg	9�Z���#����c��m
dV;%-У�]��cs> y���=���=s��5l��+�\���V�=@鴼4�at��w�l{{�Uč[<�	�� ��^J�U$.�E&&˲�SV�]���&̬ ��^#ذ�Im6��;���'v��2���xǱ`]���F0T[�"�*N���xǱ`]���2��ҩiM�ڻ��(Ui6��8�L86���SQ�n`X�m0f)�@�J��9���V��b�:���6e`vL��J�F4�T�[t]��:��7�C�
�`a�_ 
� !�?KﹳrN��lܓ��ݻ�d��=�j�j�V+�v�	���ɕ�l{�ݏ �P�T�lt��ɕ�l{�ݏܮv�����"�S6���0�V+��6=� ��ǀlٕ�}�2�UUUWwʰR|(��,U.l�6lғq�k�i-��W)�]u��qn�J��⫒���j��lٕ�}�2�_ ��~�q#g�1���v�ciݼIu`g۹X��,���-����T��3Z7$���f��}۹�� � �P ��������7$�~�́�ԥj*n�wAa`��`^ŀv����'�=�}ÒpUo���|����Bl.�`]��W+�S��W�w}�cذ	H��T�ڷ`�h�(���.Z�#o!3���M��F�0mUW:D�]�k�;ڻx͙Xݓ+ ��,��6�
邩Wlt5ui�`vL�cذ��x͙Y��D[�b����C�b��y�,���lxd�`��QI���wwM]�v�%(�ǀE6<�\0=\|��uB��lJ�I#�Z�\<�<�	���z�v4��ӻx]����M{�dx��S��2�@�ۆG1	�ʸ�.`�+c��03�tS:�v^qf;���G?lvK�#ذ[#�+���<�<���V��i�%j��7�/}�䖞)�<y�,�\0�*�6�Bl.�`�G�l{�.Ǳ`�P�q����]�cذ�p�${�dx�JJ��۱��ի� �cذ[#�6m�	>q=@(� 4: �I�"I�II#!�HB2BBI$d$dY$$!	� �M�C`"�+�	=�oA@c+�π�

f������$�����ām�\��e����k�kD&�&ߒ	�$����AP�.F	��:%9^@Y��9��G`}��� N
`��	S@ ��^"h�D��_�C��+�1�F��9���'ȿSQ J�E?~��%@H�$Ua	$��!��Y*�D H�	�B�h���U�Lߗ�������غ��ːM��8l�uq����! Q��v;.� ����+)[mVp�<;`�+UJ�M\��fV��,<�^`*�`�rc�2�h�ã��Dd�����ڢ��F�ՋE;�D{�A#R��y��-��0\uUK���u�nΛ^ ��EûLK\�Ӫ���k�;���bł�Dz]�f;��Xl��˻*�qԷ0lRHE�kf�@�i��2`Z-x�;EA"����{;�ɮ+��E�VEU�t�3���˴pEh�B�n��6�&�9C�Չ�v�,r���Z�K.3�
��F7�?|����.ݵ�/h�E��I��<�V
��ڜ�������v3ǦUV�����nW���X�RqsS'(n�V�r��yݶi]� 5�`؃_VL��N�4�h�k�'lpU�v�c��:X*W.��v�@7Q��ˣg$�S�V!�X+]�U�+eV�j���O[I��L9�yZ9���X`s�y-b�̥�Y�ݕ��Ƒ	�y�gv<n� ���e�o$Um�]9h�X�\��KK�U�v��6���sl5�ip誗v9��vyطW4ZU!�M��`:퍲�� Uم[���n�!;.}8#gNq�Ŷb��]�����<��GNè��QG�񎅴4,�kr;3���i�3���SJ�4��d�$�9M����玞�uY#6���v�	��3	�nէtn���˧���<��r7U�fZvH�����6S	M�FW�� �{s�ۤ8�ӛ����9�Wt�u��9�ݕ-�1�ى�K��S�,��fx��b.�m����� � ���F�>)���S���
�kv����t��'�(ͻd������ս���]1q�I��D�r/;'Y���su��k�yv�Ӟ 떤d�f3=utظ˵���3zX�ǥ��Z�q�n{~(���6'�f�r���ą&+J�F�&^��n9�!&͸�쪮٭vN����u�O��>O ��ʿ"�� �����;H/�?�|��w���9�ɭ�h�34J���rq{!YV��w* ��5�V����.-��饥g�*\��9}��4�kۧ9^���ٲQ��v�X�*sO���sd�G+��X#���.6��1�c6��^r�^mI���*3K3�1(
�s�~���M�en8��Z�{.��)]qgsu�!DR�-�M3�j���][�� ����99<�����j^Ħܼ�	�N٭U.ڵ����=O\��Ue&5�f�Cj�p-n΁:��dx�p�;%� ��E&7t��]Z�j�`�G�Nˆ�.ױ`�c���t��ӻx͸`���Us�O9�E=�vKbR�R��H��7f�.�b�5l� �n�R��v�,,V��G�`�G�I��\0p���D�v&�6��A�f�ǘr®�9����u;�ȳڵv�nhF$��EݬV��	6�vK�#ذ	])�
N��b�Wo �o�p>E~(%@�)T�Dq"�D��3,׷�M�=�;�'���7}�Z{��Z�mh�,5cT��_�cذ[#�6m� �s�o�
�?6�L- ݟ��W8��y`Oy�6��s�K}��{b�P���wv��]�v��"�6m� �|߼� �����2f�l�jJ�*c��!pc�VN��W%��U�-6�mT\`�FƝ���wo ���\0ǱyUp��S�x�[�B�݉iSn��\3�H�s� �{� ���Gez��������Ӱ�=��5l����9����%�� � ڥ["Iam�ݬV���Xd�uȰ	Ӄ�T���Wj���2��ʮs�K��X�����O�V�ōZh��eM��<��t��*�g�G��v9���Ym۲&�u�vI��w\� �r,�&V obSLah��.�`�2��00��P����mէnݘ����e`�``��oe�%�WcWm[N���e`�``�E���UR�Q�W[n��̏ ���J݊�iYwu�vI��o\� ղ<�L���@����yP�oH#m1��v��Lom�8ck��t����L�6Yu5Y]-L܇@��y��5l� �ɕ�vI��}T�v$� l-����j�{��9č���/�`�"�;Ӄ�T���Wj��ݸ`mİ��~��<��<��˶[vX�����$ۉ`k�`I�{ oe*6�cE]ݥ�}6�E$x��X�q,�.���
� ��7��L�G&͐�U�Ӝv�ѷ��fbl�¥L	�à���.ܳ����Bۋ��R���q7��Qc\Q��v���T���lt�g&3f$^�6���u�L��ND>�\xB�NE5v�>-��J�7�s�v�Cc�2H������V˯m"�a�9.	pg����T�Vڬf�4�B�ڷH��u�<�	#�7�+L)2[4�\���	��tH�ʵ���;iMf�����-��EF0^��/N�I}���˙i�5�79��?���۠~��,M���ۆ;�1ƕ;��ڶ6���7�b���${������z{�_s��~��}U�������ޗ��\0�� �\� �jR�4��X��'i`M�`I�{���^��%�J�^�N����C�0�� ޽� �n%�}6�}�<'�JCt�N����(� ��/�n�;�-��-��da,xҐv\Ld�s�c^+j���<�	6�X�nRG�}���7��],5�r�矟-�NUu�� �H�]����T*cPm�C�����0���\J-�x�/�`b�Bcn�ʵv�ـE$x��x�q,�wS��cWW\��~�y������<��w��`I��hڨ]�Wt �r�N�9y��mֽ��S��\C"Ɲu7e<��t�e�ږUe�m�.�����@�m� �$x��y�Us�Ď��+@��h*Ĭ�ݵ�w��`�� 7�/ �ˍ`T��6!���wf��{��O�}�n`�"�a	��W7��	��`kJ��SmpWi�Wo ޽� �ˍ`M�`~�s�����?O=�5=�rh5eV��||נ}6�j�<z�,kkJ��ۢ���K��gEp+Ih%�7�8��k7g���<��[M�S���[��d��߾oLT��ױ`�q�lS(CI���U��n�T�窪�\����y`}~k �m� ��L�RwVݺV�ӻx��X�\k �m� �$xdWSE+��H��wk�\S}�k	?{��ܓ���7'���j��"��=��f�|���}��Z�[WaV%e��ۆ�H���X�\k ��Q�,T�ؗ�i���vB'%��+jD6\��.ts�e�T:N�09��e�m	���wf�H�]�����ۆ7NZs���]�շo �ݏ �.%�}6�E�~�U���ڗܻ%��5w@��_m�M�`vG�j�ǀE#��J	1��wv��ۆdx��x�rI����z�{}�%Ļ�Ʈrt�#�=ʥ6z������0�Py�j�H("f����ɭ��r������� B��m�z��E4s��n���[*�dZ��+S�f�s�]k�N$"�Y�ݝy�H�\R8�4��-X%)�6s;=JI�,V׭e;�a;@͎���	%r�r=�rob\�*�Bb�ע�E� ΜM�����{nD�a6������!b�]2�F�
۫(lԅ�T��\@�īU��kue��5T�9��I'�9};>k���5��
���U�*���c0$-�/�u�@�:�|[��Ʌ&V�`�gf� �����'v�X۷�r���A�����!��]ڤZCww�N�İ�nױ`�e�������¬J�����0	�b�5wc�'v�X�Cbi�$�[jۻ�kذ]����K >�/ ���AI��j������M�� }6^�v<T��w|
����<��\wҳ���B�V�A�tT��t����>Й��s�+��@�~J�3{��j�VW�׀j���PJ�Z�wi`�e��t|���s�C"���	�z�	ݸ�9�W)"W���)L��Ʊ��|�{z����;���e�v��ݻ���ݻ��ݗ�Mۉ`)��z�k�� �ﵖ�YU���e���ϖ�j�ʮ�O?��'��{ mj�TT��6�yD�\�'��X�(�&Ձc�iU�1�^k)���b�KQ.m�����x��^�v_��'���bI���n��]���ذ���>Sc�7t妥2�(wi�n�ϳ���9��v��bEٙ�I$�Y�ğ�`,"@ (D����� :;6��A��jn~B3�T��i^~�0�!	L�?BqBBspM�c�#T��**�{�1�9�
KF���
۲b~r(�"3��b0*�18P7r�,S�R
�7�(�H;iE������Dt*ӵ6�F�x?uO��E�'Uj�uJ��D.���lr�u�g��'�����~��]�(��5]U�~���-�����=�W9T�.y`R:)!�xi�-5wi`-������ذ�f# ���E:*6۶�hi�N��3Jݡ�[��D�v4�:�۷�&m��Εui;�U��ݼ ��x��x�f#��|���� �,cO�v�wE���� ov^���`)��{%��]%()R��H���� ��1�lx�� ��wEl����U�Yb�F��ݏ� &�^R�ڦ��O�SFA %��'	�^��������y��X��&]� ��ǀM��}ݘ� �v^����C�}n�4�*�f�U�p`�6�ラ-	E�E`��k1,ڨ�lD��`K�e��;��;'� �vb0��~��<���k�*\�hj�����y�w�PvO^�O< ���ꢒ,j�6�X��h����͗�ݗ�w���g@�~���8��RƲ��=��8���xힼwT��	ݗ�ov��-4��lv����/ ��p����>]��8��9)�Z���M��թ�Γ�r���v�ۢ�<tDc�<��V�M�������J��c�M8�4��p��#[a;\��5��VT#dc�m.b�v�ht�k����T?������B9vLs��.7n4�h��#�8v�H̰Mķ[����j�����I-�I���y��ZK]&�����pCڭt��ŋnwn�$o���'�^|ݟ	���5��l΍�O]�/[y�u��Oc��X,[�]���&��%�[(�l��<���ހ|��ǠuvG��s�d��A[��vt%eZv� }�/ �� >ݗ�w�q}9'$�	��> [�ö������7�b�7�q, �l��)�d�R|�l�k �n۷�	6^�ݏ �!n���X���]��ۉ`�/ ��ǀI�n؝
{L2�Kbƨf�1
�����v;PGgP$�=8Fp��Qfge-1��e�*��l���&�0���>���a4�f�X�9^�������Ns����Dwp�>��K $�x����;���Ӵ��.�����	�/ ��ǀvEtF"�+�T�J���wn%�l� ��.��r��,Ty]һ��+,N���z�{��	6e`Iq,�p=G�y��hM4r��Xs�twB�w@p��cE�k3q�H��t]NK�!7E�ݷw vO^�fV�ˉ`�/ �N:[R�I�wi�Ww�I�+ �ˉ`�/ >�/;\��$(B�Kj�;�i�	�`G#x;�u����C��� l?�8�L��{������N�H���Aum]ݷ�ڪ���x��.���������a4��Y��@�~�t�I����5�v^��
Q[V]�E���:�Ě�a6�&J�E�ڍ]7�d��
�f�f��:
fSG�������>��f M�xWv<�+�H)]ڤZT'o �vc0M��uwc�"��Z�S�]�t�[��ـl������f3 �l*%&������ ��ǀE6<zl�rmG@U  K���έ��kpiĽ^�1��n۷�E6<�*���e�7��=xWv<��s��� �O�m[�˛�v+� SZ�e���ʣE�����v9��Fr==��q����s���/ ��ǀE���H�`FR�j�� �����x]��k���$wa좒i���"�ջ��"��E6<=Iv?y� ��� ��2+n�m[�];I�����y`��o &�x��xdWQ �T�Zv���� M��]��	�w�rN��~:�� �ٖ���+��m4v��w@��s��-�a3m��5
��Z��-բ��*�����k�L�*v�n����-���l;���jNނʻ����*�Ie�'�E�M�[ZL����q]�"�\`��hFh�hŀ�hX���{�2�@A�#�b�E-[n��G�C`R��5�=�Kv�-:vq�%rAgL)���5_j��u0�4����'$�}�NI��u��Ϥt�G�K�6֦��U�ls�s0��(isA�6�->����4;Evx�a���}��]��	�E�}�cx�qw���y0CTZM�ww�j��Mr,�{�	�^ w�ڜM�n۷�Mr,�{�	�^�ݏ �H���0�Wt�]�ݬ�{��/ ��,uȰ�]4�&��ӻj����/ ��,uȰ	�c}�'�'���-6�hL�*F�Sp��Xv��
�x����$vd��	j��.���Z��w��5Ȱ	�cx6K�'v�8�t��t+c��`�;ۼ� s�@`z������xױ`�\
|V�p�U�k ��7�d�kذ	�E�w�9aj�����M�x6K�&�� ��Xױ��*�Pmj�I�N��	�b�&�5�o &�x�s����������'e�(-ӕqt�9�3�{j��������
6Y��;�����:�C
t��Mݝ���� ��7�d�kذԊ���wJ�����&����/ ��,k�`��iA&0�wm[��l��H�]���E&{Y�]�=���7$��׻%$����E��ww�H�,k�`^��l��u�8�.�wt+n���&�:�7�d����������<��rfji\�4Q z;`LE#X�s]r��$�3X�X6���Zv���7�d���5Ȱ��h�W`�n�v� M����x�"�>ױ��Aة(4���nӻ���5Ȱ�%��7�d� �N%�)5E:wi�n�����rO���3rI߻�nM�x�(� �A?�D@f��ܓ�{u�����ZWe۵�}�cx�%�[���E�~�9R�^8��uj���S�V�����S��.�NS�
z¤f������6Fe)�Hl�i1ӻj����޼��,k�`u�o �u]JJۦ�E��ww�uwc�&�����d��u�9NӶ;��I��7\� �^���K�:���خ	P>+v�X�ӵ���s���޼����X�B��հ�)[�ݷ��^�ߵ�o$�^��I������?�QW��QW��TU��TU�"��� ����**��**�Ҋ��� D
�D�� ��*
���H�
���@��* *������ �A �D*Q�� 
� �E �AQ��*P������* Ȩ *
� �@�� *��* �D`�@X*��
�QB"�@�� 
� �@*`�@`*"�E����*D �@D��AP���A��`*B
�
���"�*��*��@��*�� *��*��A��*���EB
�E*P`**QH�`* �E
� *H*��"�����
���
�`* �E��D��V"�
� **��
(���� �@ *b*��
���B�* � "E ����������*����EEZ**�TUȨ**� ���@"��� ����**�Ҡ����EE_�EE_��PVI��_	v�AY 6` �����[��    �     �       @ 4    ���@
RE*��%B���*�JU)EJ��AJH��P��)I��PJ��J��R��$  �   @ (  CO{�'�����w�:��l�5� v�ms�vۋ=i��o'�� �}}Kw��o}�_  7�3��0 ��zUbz+�l]i�S�#n���� 휅1iA�2d �:( �
  
 �����9o�&���Юp ���2Wy��5ťv��R`�����>��y{������p ��W���Թ5����:�{9�� z<���{�<��֯�Mɩ\ \  �    @��#6Uq�� �    @    � � @�     @   b     � �� 0 	�s K{pP   `      C Q lt 8�7��ۥ��6�Ӏ>�:S/}�U�˭\Y^۝�i��g���6��s� .OK��g��� �+6�һ���>�m�[�:���M�|�<�^�yzyyW���ju� ��(  
�
�� ='Ҭی}<��n-/[�OM� ��Zri�㺺n3����+��O�������\�� [�ɧ{w�s�� ����Ӵ��֜��y�=r�� ��{M��g����\�w��g����*oi*�  �*��ު�JhA�'�UJ�   "{J�55T�F�"��J7�JT @D�6T���������?ֱ����������{���;��Uz�������PU?�QTU������
���Sޞ�n��u���41cR6@�`����#�?B�����c�a�d��!H��q�����$)�,��	���c 0aFH�la"Q�4	B\��2@�!*Ħ�$H�`X�D�De�Iq��5]������L��R	�BQ��\HЈ-	$�!�����1��HUrD)��YxCSD���$?CA]�LS� �j�Y$���3?8I�֌�i���4�G[�Im24#S$ԁ`��_���i�H0b-H�"@t$I�D���F�O���@�ki	>��BQ$�d�I�"ȶA������b5�X��Q�X�E��~�"R�X6@��,XD2�!@ґ�I�F0�d$��hI��4ʐlj�ƌ��j~ݳ�Jh���L�0�����3���`�
�T�g�>��\HT�BH\aB�+��`T����aqaG$v*a)���\YBPԸ2��
J!XHV0�pb�$$	��*��2�$hġcXBP�R$�%!F��)���p�!f1�:
R�)��"D�0 F��� l���H�ab��X�P�@�$X�`47��5�o[l��![�]!w����|r�7z]sl��9.k�q�lớ09}��=��x}�=��C�}�'��L7	5��o{!�k���ol\?+F�串�+�,l�2�.$*`@�#��S,�@���j�&K�nZg�ƾ����q��#d%%�o��[Ʊ�� FB1��~�1�??���D��U D��]$0�K�ޏߦd7�ֺc"I	a2X#[-3L�����BD�$H�c
°,�,��A�@�$����ә�V!$̈́,�$�H1�U���a�M�	S%��i+�E�m�`D�$75�w"�78����X̐��fw�&�a���!bu�$t)�"D�1Z���L4i��(\0P��`�c\]��3D���7���7-by�߹H�	I	#�D0�LH`�	cH��1���H�4qe_�B�E6�v��A� S�Ԗ H��T`Ƒ����c"HԔ+[$�j�e>�-�ˍ�}������X��D��Hp#L�FB%H��H�-�B	HP �b�VR���C�R!0qrp`�5�`ȶH�A#%7
�`O����RI9)��jH�@�`A @��!Oƌ��~��R.$���D#C	�RJf�)ܒ5�i5�����bM��dH����f�nF\�
a�X�%c!f&���C&��3u8T�Y`X�4�h�d���I�pHȱ�7v~�sz�_�
�@"E��55�8R�f�˴���\�֩��65	P¸Fi�u��b��i�މ�,�I�$"Ǌh`5�S��J����ni6g�$�5�}��~�������S{#��۵�G!5�޴�!�S�+�,n&9L���$��~H|��W�a$21��L���~ѫ)zkXs��0CA�+��B
�)��Q�	$b�d�� �4�!s[�VH�%&��~̒��7�wCFIhO�ԃ � 4$"@"B�J~�*�Ĕ#����%LJk!qѫ.��ap@�Z�5R~BIBIa0�!f�`Ĉ��$J�`���cA��P��Y�@�9�~����w�HBHF��"I!���g#SW�&}1�1$5�z�䤔� P�#�CI,e�g߷��i��U�	�B����$)�	��40	`P15#b�
�pQ!���50�W�!VHVfIap���kd�ۃ*���@�	2@�@�(�jF��E2u�v����D�VA`a�D+�
d���\���˾YNs��'?oYWs�XXS4���}��Yy���h S �@�@#R4)c ��@LP�vH��+9(d��i����]��&�%��I�f��?B��,���X�Jbd�)"�(8�u��6H�G��sw��$$?@�0!,)��d	��,?c7����	8��(H��H@c�
aE�RʘM�a��㴊ąЄaC"�h˚%%�7�xZ�>��3L�H�f�4~kR_̹��FMo_���[$� ��1i�
,JJ�H�md�`}��,#!p � D!�7�����F���h�7�0澟��M�����M�B�`�)�2��+$h��A�
�X@0aC?�,���D�h�1�>e4K�{+������-4L5�Ɛ�E�⿈!"C`RA�1`G, �[��K$�}.LV#���,��(���	2B<-��!&���2A��lM���!�\	��H|�q0>	)���� �l� ���$"���-S��@�DHP"U!l?��|eѣa�F��F�����կ������?&#�HI@(��h@�m27�R��1�YI!N?sI�����~4��)���l.-�e��V�Z֦�t��X�#HR�.1���4��5LÐ֒]F�XQ�HQ�k��w;>�݅΄.��+��*B�(Jf�����,�5��ݏ%�Ku��{�Iw��0�E}U�cFt���(Jf`DD�A��s�~cp \`\���*]~��������v�`B'Y4T�%;�]�gw�VС��f�h$\0�� ���� @�~#de#�.kaa�޳�e?0�Z"dXi��3\�Z����>a\*��@�E�#������1�w"�!>#X�0#B1#%H7,�EH!$�"���(I��BI
��2����jV$��j@·%#Id��"@�eeE��!BR5�F0!H@�BP��p%bL��#ԃ�q��tI)WF���āG �A��M�
��\`n���c���}{ݾ�����\�֫5� ~����P��%���cbXC�շ�g���
�J$`0!�\�Q�ٰ$� lrQ��%HЂ@q17C�����81���"��BY�ԜdH8�B P	�1$�F����R������_!�_n)��˫��1
Ʀ�� �R9~���ޡ�[�9��$eB���HQ���r�֍F@��$��$��,
��� �IlѶ^i�k���ϡs�d�R�k3N�.�D�(���,���#���?~�K���L/�yù�3�l���� I!$�$+�kP�����7��;4rq� ~$��XR��3�z8B����z	�u)��4ha��A�	��u"I$�)��HJHk�f��/�6|���V�F?$cǟ;yf��ܪdt�f̤�}�ޜ7��kw3F�'�>��Կ�]��5�X̕�V��!��R�>cX@�HE��L�B���"e�y��İ����e���4ϩ9���F!$*& p�E�!B$h��! ~D��������BF(A�c��	H0��B%XXV5.�����62���̤�L�f��&�VT��E)��cq��RdىKM�5p4��SA��S��nC\)1c$C@@�����,�([3���?�#1,	 I�؛'&�ܔ�o��f��&�F�aCa$P,��I��4�5�4\��%�B���T��D�Q�!a/	�M�8MRNd2�%�W"�-B])��05.�S Y ]%�R�v�2�HF2��o�k|����<u
�H��)$��&$JJ0c���`ۭÁ��~bY#O�	�5YC5*c��nD�X�!H!�!� 09�#E�
�7���   m�  �m� �m����   -�1U
�� 
�jz7#�n�v�Ueh&�%�����A'��
�NHf(���{-V1U����tqtU]b��	��Ԫs�^VV��T
yQ;$���r� :��cE[\��Ӛ3z۶�	�j�h5���D�( ,2@#n�$ Y������i�$�bj���zg�$���QU[+�� �W��`*�$`��a���b@��rɵ�6� I$���V�Gs�m�����cm؃ �klX��m��$�c}�9f��I� ��Rʥ��[I�mW�M��&�3V�	 ��q�����5�5�G  ���M���3fk��UVCik �n��/m���,H�,1�h�H m�D@T�*Ҫ�֩U�@Zf�n m��� M�V� �\�)3�ઝY,�*А5���UJ�!6�J��km�i"��M����@����]2YG�4n(,:Km��l��
�z�`!�Z�VBSbd�*X�����az.ـ��p�k[xHX6k�  �ͶZlImm�]6��Im:�$  �k�kn�)� [m`/CB��+�8*T|0q�@��ޔZ]�ݤe��@�� ������V� �l[v�m�m�����L�+]M]{m�(	"hu묑rN�L��l�@@)-UU.̻<�U*���Єʴ���Z]�H ��[��m�  m����	;n�<*ޮ�x6V_,+��j�$H $  � ��Vڶ6}�JU�VV��*��s�$��  $�kn�R�\�Uj�	午�J���&S��z��8k��d&�ks��l8��z#\=eT �^y�l�@t�H   HT�.�g��Oeڨ
���%�U�	�T�gf��^�&�U�\b����@UJ�����
YV�� ����f���ԒyVVڶȥ��R�h8[x &�3m�-��   m[g-2+m���j����[]s)�UZ�sZA(t�v�`m���`�\m{�n��mX` �zI5�i6s "�$M6�UG��lJ���[A �g-��(ҭUJ���U[�mmP-�$�[ d}o�}&�mfӦ��M�ۂN 6�/Z�t)b�j��VUP�wR �۷6m�l5�l浀 ��[[kn@��J�M�lְ] [��W���
�S�se�,���m��$� [Nv�f��   h�Y4���U�"ڐ�'H �[\���IJ�Y �e��n,�)
 u�m�!�Ԗ��,*�]azA�[R��1�m�ڳv�)6��E<�r�&��J�n�]0��<�� 붋��ݺY��r�㴡�۾�N��]�6�������U�q��<Ŗv[m���ۚ���ު�s��� ��z���	����vZU��Z�UPr�yA��/[w��� �ݲ���%�[&��l�J�t�*�TU 9@�H�G�ꪭ��)#�eZ�m������SPh �` [Km��n�uA��UF���i<���L��i�M#��ukn�����m�;�R�U�Z�Z��V�5�i���� F��D��` �T��Cv�� �M� h�6��Bb浒�זt:V���9�*�[UPY�  H֖�ҵ�m�o�R�,6�$�o��}�u��ݍJ���!5�J���8��`�۫�6��`����fհ��m 5�ۭ`6�rqmUu�lU++J�@��p ��l���j���6*^q�.��@��@�v;U*ҼֱH��8 ���k7@U�UR u<��$ I �d�ɭ��;l-�V���Ie�Nsr��A�T��M�N4k�Z�]�,p�$ d�I�oP��v������&eTL-F�kh@�l���m[@�$��l�K[]�̆�$-�}�m�m�iT��\R��A�,���t�Ut���Urgjl�f��X[xݰH��z�m��  l��Н�vm��H���
�K��  ���;uP
�>V8A��V�WgD9�	88m� ��c�p 6�$�J��� Q�-��V��V����]&��م8� t�k�v�i6-Fڥz�\� �ETK]9���N&�%%@`  �h�����6���l�����-륌 $� �0n�:�RUUA�Ͷ   'ޝ8�����IӪL��4��� �l8���-ۆ1'��C�vT�XF��ږ6�` hӷ:If���m��`��� -�@9m����%�3�	8 �p�H� �f�T���c -��%�k��K(��8� Ҷ  �ٲ$���ׅ	����b��54jF�  l����[B��m�  �J� [�� 䄀$��m����p �j��wf�@U���L [�F��m�Ѷ���כ l-�.h�]� @��UͥX)k��t+͍�MQ-�z�Z�i� m� 6�m���c���-��<5��7,��)�-�F��]�]q(r�oQ;3:A���w�!���PYmH&�6�L��Xhݽn���C����$8��p6�I&�������Z�}�jy�U^Z��^M�/B͠� ����oo�ݷ�Ʒv�6�6  ׍�����lp��fL8;:]5��M#���=�[�VҒ�+Jn��P�V�f��`6�l Hp���l  %X��X�J����j��dm�5� ֳmm�hkE���`Λl-�qH
�5V�*�l������Bk)�`�i����6� 8e�m�D��m������ M&$$ڧUͻd�˳m*��c	UR���mJ���9��c�]KMf�mn�0�A��ā��l[@ 8�`d�� $ �ߍ�I�l5�l6��Ͷ�m[@$m�m� � nI8[%mdd�K(l�U����H�cN��T$ �6�P�l6� m��'�m�`���rN�m��H�! U[P��
�;Ӈn�����&��Z�h�Tb��`.U�O J�m� [@�=D�r�k�D�  -'���*���f5T�` I~�E���(��{ ��J�*�L�V�]um��b�� �Ć���؃�Y9�-  � m�v�-�6�hjۀ7mK��d*G�U`Uj���*�e���A��u�R����fȓZG.�[I��7l;UXM��CH&P����`�EZY9��De��	*���m�-��	;a� ��]�h��U�]*��^�kp�,�m�� [nMn"Z���m���Ԫ9laV�ڠݎ�:9��7�-�Գa[EU>b�mm��m�Hm�@�`�a���N�:D���pq�,��Zejc��P!�m�vԳ�6�� � �m�pp   0l��V�V�R[G'v6�m�� �H H@]U++\���+�M�4�j�H  H[e�W`�nU���m#���E�1mu��ΛT�����7ka���l�<�[l�
���ҭWm�/
��i&�$I�l#&�� H �6ě���PL�����'5WUr��5UP�R��0M�ä�e��6ۭg 骥V��)�󸍍����R�յR�J��WT�e��P88���cj���e��;"�N�����^�4�szM�'YV�p�rYƊ�M+& �D�-^T�yx��UÎ�6�n� �����l�@k1:t�M,��r��J�T��S��Ҡ*�e6�@U������[:�I��Ɗ9��l �� H���M&���$��mm�   ����ev_\�.�j꫕��z(8̺���X{�
R�  �\�����h  � ���"}����[Ik�I.��	ep9"�Ө�e)�ݲ���5��V��mm-��8� m�&�d� �T��m�-�$�m[��2G5�h/iG��Ts�uJы��Q�s�0�' hW��u�޵�zCN�Դ��l��t3����YN�gtG^l��Ͷ 6ڠ;iUV�j���5*�����ۍ��iee��&ٶ�U�k��lv��  ���[n��m*���Q�T U�/$��pڶ�9#u�ݚ�p   �l�k�	 $�۰�Lݬ��!&��9;k���J�sf�`mu�J	|�_�h�Uj��� �e�izS��m�Y@mf�%���-�{[d� 5� [Am�m���Sm&ć4^-�n�$m�	$m�� �Z�Б�v�`��Z�$ ���m��ӚDж� q��ia�[G ���H ��Zm��
�iB�`m� ��m��m�����amX�7o` �N�m�m� L�m��md̍�	6����� � �ΐ-�m�����l8l��kn[ɯ:�$�l�a���I�J�m���������GQ�A�?��?Ҋb�銿���U��A��Ӏ(F.�)���H� z���x�B�
�N���(���@�`S��D���+� >J�~�EM�
7�����PʧH�Ua��U�G�"��$���	? ����M?'�����S�P A E���X�?/� � ���6��� P��E�"��0�#���@C���A`�pz��aA0OÃ�61����`DvT��lb�V*)T6�@0�� �����������C���)�^
�m ⨑`������戰�]!��(	��M��@���1vO��.߈�GX�*�'�hD�� !�UO����Q��@t�+��=0P� ����L �&!�����B/�0M
?�j�b�"���~P'��D���&ǈ"�Ȍ�6�,�D( �A��c�$��?|������(�dA*"
m�8�;?����iQ4�AТ� �B";X	��DSi��C�M"Q�&��(�*�G�Ȅ� �	!���1��~�kZֳ35��om+K!q.�گ)uksg�;8䓣�vk�,�6�+��i���)�e@.�S�S/���ójȰ!@�kv����#�5M�D�ďa�g��uS��Õ%n�;��R�'g�6����Dqu�-�V�q�TH�����1p<]m�۷�3nRy��eN�VCbX�Ԅ�R�Er�QkV,�s�0cd8]U\�@[FҦPܠ/�[7/<mΫ{L�	�5��68�W���Id�n�T�dm`V�hܘ3%��O`�h)V	*"7�9�-3!3�,]7����փl�h=:� Cs˞�5���6ђ�Y�8X��G���D��H%]l:�.�f�8ɣ�j�=�N�0�˽��2r�%d8g:��<��@F@���r�M�ѬZ�Ju�鳠iv��Ўӣ	XD�'�餲�c�vrm�S��� Z�{��n�^ev
d�V^%�����H�d�u�&�a���\�z�UF�Y 6��7��u�z��y�;l���� �ڕ�%�54�`�V�9�T�ʶ�v�i\�e�.�[2iē\�X$�YP��H�<0�l�m�	�m�vt��)�ڎ3���hl[��	�`ԅ -UQej� ��m5�؞�Wh�y��^y^���<[��%��R�nWD�QE�NEO�N���&���N�y�)H� 2�=�ѐ����.�a�3rn�b���'!.$k�]�k{E�sj��^���m��JVYY��0�e����i����K.�F@��{p�.Xk��
���Q�S�,`�,ή�q�6�G%��X+qA��9�gkv%���M�1�)�Z�s���#C�hjU�Y����m=�{(��ݸ�ݞ4����)N����ڞ9��N�]�	��v���J��j�p�v�XȁfwE���X"V�Y'%�	��Tp4�\��m�p����Q,��{8W2WSy2:�r���.m#n7���I�-�-v�uU��﻽{��WFˈ�A	�h'���_���E �W�'��������2�d���u��mpQ�����[p�����)E����;Vѝn{F�L�r�OR��[Yʥۮ�J+�/�`�hf%6�Q�$��y��M�b��@Ǜ�x�q��aAoT���]=T@�\��݀4��lS<��̚���V�<�8Z�m���mרӃ�m� M�*7-n.uf�++:J�Ӊ-�%�3NjK�f�ɚ���N{��������ªv�簧�<�c�v2�(�q�&��IX�<I�_ǐ9yf��9� ߾�_������S4�w2Ay{���]�=̨�� |� �,8\Cʞ4��P�M�s@9k����W`���e�eѵZm�� �v >]�u���d���#l��<X�rh�٠q٠U�W����^]ĺ��B"�Z�����z�ũ64��;v8�J��{��M[P����5���k������7�� �v >]�r:&�n�suujBn� s��;�*H��Q.R�n|������6� 5i5`�M�&E$z�l���@�-�@���@��j��x��Lx����w��B���xK}X�P��{4��&�T��$�8�� o���� |� <u_�/���t�A��(ڞ��/`kE�v�xrE��1��l����]�񞇑���_m����˰�]�u������ˣj������ |� ��\�{�>�:��M���&<Q�4	��nI���u����H��� KR��(P���� ?��\6M*�Ɏ<&(��m�\�z�l���@�q��.D�rdł���9 9]��`V�@9+�=�{�',nm�۶��y pcY:�;s� >�Ԫ�l%��T���=tT��� |� �r �2��5`��8�%$���@�-�@����[f�}��q'�UH���^�6� {���������Ň�ySƜ<�ɠ^r�h-�rI���'Qt"�t�Aws]�*s���5�̀�� �h�v�+��� ��y�~�����o,��8;�����<�Q��� ��6X"��&d#XF�Q%Lx�rz�w�@���ʀ��9���fBr�����X���T �v ?[4g����Ey1�h���[w��)������ ��t'�L1��#���<J����w�@�-�@����-ajȜ1	8�)&�˰�W`s* ws�߿~���e��Ө�dQ�<1h\�i��˨���OY�-a�l\�]���g�_-ֺ��5,T�Y�yH���[�l������k|q�%��i̹:�!��;t�Fs%��e��.�зVw�V��/<ɳ���\��D�ְqPl]����5����x`���jZ�s�J���]��p�ļ=����@�<���ހhD�&��t���]���u���ww6��`-�<�g빭�k�r�wS��s<QӶa�ƻ]yI�d�u�Wej���n�� ������`���s@�.!�Op�G�ɠ^r�k��*�m��>��ɷx��9�YyYto��ͨ���y��+�^]�����bmD�$C��C���׀.�^�X���?k�D�̅�mf�w�� :��<ʀ��^��:!D&�p��?�\�ڥe���N�m���� ����g��s�&�4˚�]p��m��R,x�9=��s@8ۼ ׮�B_������]d���*V���X�n�������5
���?������ ׯtDD���gS�!'�4)�w��@9J�y� �W �<�]eݘ�dSWw��%
e����,e�Xo,�8��q*xӇ�<�M�2�j� ^v u+�wS*�נ���v����ۓtU#=y�6�Q�f�Z���vcO>��y;]��w�o��\����v �ʀ}}|U�x�IBD<����Y��l�-���8��@�����d�d�AG&�>;��rO��vnr��q:#�:&�n��@=��@����MX&�X�br@9�T�� 9�`R� =�[Y`�I�<�$s4[w4��h-�j^]�������^8G& �u��9��y�V��v��9�8� ����4�g7klŊ8�	8�1�$��� �h�*�ʀ(xˬ��ݻ?y�� 9]�s̨+*���8j̦��O۹�� �PVT�;V�r�4}��f6�'���ko��s�ۼIb�DB�
�q
"��k���>�/a������w%+��X�M�Д���k�ŀr۹�}r����䘙�q,̉'�J�]�kK{Z˵�+h煍���1��w���+�חU��F܋���hr������;V��3�M���MH��NM�VT�� �b� �v }��2�н/�Cwsj�ʀu����-��s�s�iı�)&hUr r� �e@9YP�u�Uw2"檮�[w�yB���w���ذ��`���;d����T<Yge���)��n9��ԥخ�ۮ����@4s��;?�G�e8�݇rmgDrVW�GY�77:v�[j;JR)7c�i�H�{6�&��6z�9�u�g�	�����1��� �(m�A!&�mt��&�v�W�6$����E��^�t�۝	�4�9�ל��$gF��5uZh�W�g�ۭ����`�kY��72�BO)� Ѐ������������[^����WAO+�;-\�sTs�rrnzFަk���J�r��j� �v�cA����F�h^m@9YP�r u�h��h���q%	�%&@:������ �e@>R�'�&$Lja�= �h��h��hVנs����`ڑcĞ��� �e@:����֛w�S���p���Q]u�׬�E�m�d�����69�f��:KzT�ذ�͵wV�m��6[u�ۿ%�A�v,��X���4�XƔ�4+k��`@��J�ҬaO©A��!G������Xۯ h9ٙM˳wK(�����.�;�T�������Y���NHܓ@�YP<ʀz���]�}��;�Y�YtmV�y� �̨�k�y� �o�6�NQ"�S3Sb ��B�e�\k���.������X嶹��zuΝJ���q%����I���������9n��˹�{xeb{&$LjxD���o���5�� ��Ł�.����(������m`�ԋnL�/{��$���ٹ��/E�.����B�B@	�>ѡ�$�uŇ�3bUi6����qш�ތ�M�D�`�QHh4�EH��$��Цo�5�BB	 @��� �0C��EH	�$!D���LX�
�C�Ձ�a�q�'�����	��:U�pO�\�? �p>����|�M*n���P�)�b2qbE�HA`ĂD�+b��-^~��Cd6w�)��� ���+����%�B$H�(`m0�?lj���8��0��B		"�@�~޵�"�H1a��0e$BE>	�D���/�> ���Ɵ���EHtT5�|*��W��"$N�*Q%�IB�������ŀ&:�N�l�VwV�9BP���� sϫ ߛŁ�")|���6P73=r����TT�ݬe��"B��w��ϱ`s�s@��5�±�8�F
x? �ۮ͵�Y���pp�Z��E��z)|̽�=���{g��iD�"nG�׽�/.��5��Q	~�sϫ jG3�*�iLՑd�Z�5�Ŝ��5�ŀ9�Հ��ƒ�KЕ�ޯ�=7*��J-+	�X��,��8tD)��v,��,�����Icj#"Rf�s�<�{/V���nI���7&��@�Adj�(�K P�T8��=B!�"?u��,���L�"JU7�U\�I|��/�5�P�K��{���ذ�ٰ�~��� �w�.��ͳ��F��9�5pn0pG�Z��,2r��4V7��ފ9�N��u7r�n�����`=x��脽@^w�@9�]Fv	D�c�"�4��Y�"��]Ӏ>}� m�Y�^Q
"��@���ڢ��iQS7v�z�����ÒI(Q3�݋ �}� ? ��J�d��d���t(�ID��׀wwb�5�Ł��Ou�N Ԏg�T��UVE�U���� ���?w�_�W�>��>��X�H�
�UUfy'bָ�gb�j�-�m�Q�s�l:�]s�m�[W"��������kb�Z1�%����3)�@���E��i䭐ҀP��x5S����#����F0�FJmbwp��۹h���4\�v��Fn�ubJ�U�6�۫0�8.맗e��v�6��\U뛣�ӴWd7#8x�+v��^X.x�T�vf�ul�mP;.K�j�3!�:��/Q�����pw�uL7nT�p��s]�%tc:ԛU'XCu�Y/6��w���7�w�r<���e�w�� n���oDG���X#�C�6�KQ�4]�{�bG�݋ ��ŀn�Ŝ�L�ˎ����%*��p�� �x��$��%U��ۚ����}�Y�M�'BG�'&`rP������(���b�;��p=	%=�{�hFQu؅a�93@��ŀz(^��������ŀ6�,���2u�x��p���&�ε/i펕6ų�8qJ���]�z�}�7~w{ݸ��l}]en���n�~��� o^,��yDy(�����b�OO��&f��DY5w9$�~����$z��@�.��>����,��,�nsм�(JQ��'�TziVAu5V�{�ŀ7��B脒�U�]Ӏw>ŀkz�ܦ\2�I���Ȣ7��nI���׋��Q���`"ޓ�j�Icj#"Rf�k�h�33�������Xz�`ӗT���(��EZћ�۷u��R`�J��6��*��M#�T��ڇ��w��5�����O	qz{{��[n,�x�B���!�]ӀyBP�w+����]Mܪ&���;��g�%	)���,��� o^,�$�Ca��.�*$��	��w����գ�����*?�5 ��C�t��S<�w߷4������ ۍE���(Q=��8s�Xm���	Ov�������q$��A9�[�4�y�����v�rjI+e��P��N�ݏ��o��ud�h�ճ����A�K��E���V�ngn�{��;�������s�_�~��{�I+˰ԒV�Ws3�H]�sRIs�;�TX�ư����$�.�f~�$�~�?~^��G���jI+m��_��r��y��)I�U� ??'z��$�y\Ի�����=�$�ov�K�_+o�CƧ�����%�ƻ/Tԕ���Ü��߻�M�b|������B���7�~�ל��_R{&a37ԋ%"��J�}�}I.�����Ԓ]��W����+��K�U&���.��s�nM��	\�D�g^u�L��)U��w31o�(�ىD��#�>�$�ov�J�j�Ԓ�s�ffz�J���=�$��.�@���'$5$�,�{���<@�UCZ՗��٭�m����s��{�w��w���������Q��ݬ4~�@I<��&fg^������D(Qw>�e�3$�����$�T�1��nG$���
fw��㜶���f�m�����r��#���O��&���n??(���a3 ��}Jdz�^L�ϔz{�zwfff}޻ə�ׯ��Ԓ~fy��ԅ��j�� ��r�ĸ�6��
.�DRL4���������<mgh�n
�p 0@�x��q6^'�N�5:��۶�Dx%�ui�B�����V��cy��E!�s<�v�*��M��=m�f*J�74���qcpc҉�]v7:�d�G;�-ļfc����ݭ��a�6�{Cr�:U�˷.�ȗMM����f�l�����J����=Q��7z�|�f\2a���sv��s�mq�l��p;9�{��b{lXy`�:z��o�9��)8
�� ?������RI+�&�����;�|�Gow&����N���<jxHۋ�RI+�&������$�odԒ\��{�|m��cx7���<�jI+��s�RI+�&��w��{�I%��5$���
�,ĢOprI���^y������MI%�ӿ����W�MIw<n����Ԓ1yj]x�H'&$䚒K�r�}I.��od�$����$��RIz�s IS�d	 ��Ӻmα�ӵ��N�H�]yы�)4��o�v�o����$�H�	Ⱦ�$��욒K����ԒJ����=m%{/W���Yԣ1��5�k5�kv�~����~P�w��7�Wb��D����I{�ɩ$����ԒJ�ɽ�3��V�_��coĦd�����z椒圫�Ws�31�.޹�!^����Iq��mA,c�,m�椻�y����ޯ}I!v�5�m�w���-�2��������o�CƧ����ԒJ�ɩ!w33�̽��>�$���5$�,�^��UXT����0��q�ogZ�]^-��������۞�A��]m���ww�S��</}�Q�
G=I%�<�3;���ϾI!v��I%�9o� ���m���kv�o̝�g��R�1�r9���B��o���fI�����RH_���I%���{�s��H2Ժ�X���-�f�m���}y�m��w5�jG����[��{���B���jI%�8q	90�r��B��jI/�/��$+�椒��i�%q(�`����I#��K�r����B��jI/yv���B��jI+��#�f)16&⍘`�"��6����.�6��)s���Z���8�Q��G���q73�RHW��I%�.��RHW��I%�9}�}I.!���%�r%��Ԓ^��=��x�B�뚒K����Ԓ�;SԒ^�X�~�5<&F��$.r��$��/��%�v��$���{�ITpc�ބjE�#��K�r����_'j��m���g9m�����U�:x0G������m��	?x��[�p�dr9���_'jz�K��f}{�O�I.�ާ�$��/��%S��~/cq�rt�=��r;���f9R�k�5�l<]yx�A�km�(�X������$���O}I*���I/���{�IT�ORI/�9��@JH#	��Ԓ�ڞ��y��3#r�����]O�ORI{˴�Ԓ�*Q��Q7	�8������羮�co����I/�w������椒��UcOĦd�ng����y����z�����z{�I��jI/���{�Iq�ZPK�K��ORJ��ﳜ��"�;�f�m����9�m�s���m�?(8@N��H<Pt���B(�b�Q")��`H� H�eW����߈|���֝+CZ����F$I�j0�~j9�(�����>��T̓���� |J���J0� l�$v?5�^�Zֳ1ڇl�S�3���n�`�N��gl5��k�7Q����
�ҽ��U���v��-��AwgvY6��T�Yvd˱�e�g�)�� eW;)�dc��0ld��;Utl��(ձgd��Cg�a{B������Sv4�N�H�U=Qc@i�jv�\�[$�^i;+p[*�-����/,�o�?|F춥7!���"k;��:I8ݹ`�l��P4m/�uV�3O;A +<@nX�������=�6��'0)���t�
���D��g4ǍUJ*Ma+�\��v8,TZ1Ru�C.T��| 'n������ų�:��mP 6n��@�A:�U�jR#+��r�;-�N�%��7�[�Wdd�k�ۑ��ٴ� ˭�:re��˳��+:�VN&w(���U��K�Nﾬ`3 H�řIGe��F���3��Z���WE����&P��9P���bZ=xQ��)�c��3[z�!�aj�/:^C�'O\]r�*Q��c],dڔ����� ��'�q��Y��U�ɡ���\�Q�fΡ��ض�6j�8zI�L9eJ����ʊs�m��6H�M����l�r�ڐMؤ�uN�'d�Z��	��-u����������۷�<h(���Ύ��G#,#�"�;)��'3v�4�4+�Mv@R&�E�@g����(��=u
�Uf�)`'vm.9H�&����N�lչ�9έ=�@��]fTQ�Y[s����:� �eS���M�^ܛ#�vq�Y���@�n�d�kgB�΀xkpXr�^6� �5�\��f�!zKc[W"mI��$�(�]�mю�]�hV"`n]]��� On�0 6�@��s�Ci���Wf�XsN^��7�,�D�|�&(Z�d�/*�Y
Z�@���K).��q�,��jm��
qeݘmر�֠W�km���N�yʶ�΋[��e%^ 	�xꧭڶ������fh>C��zP�D^�??
�#��ت� �<��|���=�`�908��f{h�
\�c�#mvCN�u9���4��Z�*�1�bW8�6�n�e�z�e���&a�����C�]W�St�3�<v׌�9ݤ�l�����Q���6m�^���{lh��],
l�t�⋣�<#͕�v�:t �C��Y(M k3�U&f�tt��v]y8����]�E����t�]��5<ey5@�^U��%/`�q��{�����o��yr�m�n�{�7mho��t����]ێc�}�|Pb�hܸV��%�t��$����I%�9}�}I/��?�z�K����%�Qu��7���<�jI/�_����!$���\׽5�33�������;���6��0/qx�I�#���Ԓ�}�z�K�]������[�5$�-��$�p��b�n���.���ޯ}BB��jI.^_s�R]�3��;��$�ᅠ��5$�br/@�s����<I����OwV��� ӥ�%T�$�	���ݻl�c�7Yq��`�r�B��2��G5n��;��ݝ�|�x>��M?��b�?Kn�u�|�<�B����Հz}xU4�TͥvMU����+S�@H�-$*	ȩK�T�B���ו3�{���I��������39֩��J	c�x���S��6w]aТe��X��x��V&ނ&5<$mš�Ĺ�٠^��h��z�{/V�{V.�����ԋ��@����;��w��/]������a��<xD�1�	�Uo8�X0Jn��Z����y���R����|�Q6��= ����9_*��埼��(����ŀ�g����IrU^�9�n �s�y� .��߿]�-�FԐFE�ȴ���/.��
?DdP�!^� ���>nf�R�\�U�]MU��%���|�_�x��8.�U������2�j�,��X��ƻ�?�;_^�^f�s(���,q��#�bx��f����v����ֆ7�]A��R[�7n���}񏐰s��bi����h�r���s@=�٠{�b��z%��6����ܙ>ŀou��\�L����*&�jE�RI�^��h�[4�%z�V�n��� �ꉺ�B�uwV�=�U����;�ޜ ��w�Q
�DBBP� �S�*�*�<������s@:��u��HI1�q���`�!)�}�|� ~���6~uUI���9i'N���]�lV�w�j���j'�erk&e���w�{���7G½�R�n�5w?�7_^�^, ��w�(��;ՠs�E�Zi��4ܚ/.��Q䒅A�޼�]����y�"L���%L�$3Uk >���5ֹÔB��u���b�?lm�ˢnfUw2����:!)}o� 7_^�^,����f��鋸�z����}�����'Ͽ/�ou��\�
",��$ 2B ��,��*��DO����f~�fj�P�&�ʤ8̬n	��{un��i�Tu�5�aaq��N��&�Y6`�ݝ��Sur[�E�ݜiG��v-�rD*v��`�g����aF+��qk���p۬���:����7QۀM��dǦ7Q�DT[Y82��F�Ե�<��{�vԖ�<rl�m=s�ل��ZG�\<.:c�N����O��Q����t���;�����^�=avg;Ul����7�	���h}����L��e�����ڱ�\>˓#R,b�O���������������/��(�y1��h�W`Τ��9 ��O]�����3M.���s� ���@<���ܳ@>3���Q�$�`�4?�篫 ��ŀ��x-�q�oM�%OT�Ր\�U��o��I/*�޿�����?O�� ��)d�X��LX������4��2n&�&���9	X�x]]���ߗ��=0XbC���73��{4r�h�r���w���>�X����9ɩ��u�2e	!�%��t)��}x�݋ ?|��$���7�)򚪀��O$�C@-��}m�ӹ���;٠[��@�����o7#R,�7$��؈A�����~���فЦw_f��<��6�G#���l�;�H�s�+*����h̫���L��r���v���3�-���@��:�ĽL��.��dԵ��Lm�	���t���xͼ]���^ h9s3GWWe��� >�]�""<��~��`�z��l΄�M㉵D��U5dW3Zܓ�{�7$����s`��)�,P��(D �z� y���� >}׀A�"P�Ji��Z��	L��׀7�� }����DN���4��$�Ҁ�ԍbiɠs�S �I(������X��� ֫Z����tk�.j2ݏv��{œx�2۱��rS�<�G���ŵ�wNU�7<��k}����� ��� ?|��B�_��� |�u���nF�Y"nI�}m����y�A�;� o�� ��w���(P����Q�n��U�wv�_�x�a�(�7of������g8�x�17$7&�%
[�� 7_^�o
"$D �V � 5�.��w�l���I�cjH#	�@>��h6�`u�0$�u�*H����1;������g��:rs=�������V��ٛ��c��N������� ��w�n�g(�����6D6"P�s$�� ��f�<ċ{:h9{4����<ď�X�.�@cjF�4���� >�]�СL�wb����ܦV6ނ1�S��qhw���/f�y��h�[4��Z/V'�y��*�j�� ߛŀrP������}8��� ���Y�a(���@��uS4�g���Xc�Z�t&:���l��ؒ9^k��5 ��ݷn���:�X�<W@4����ɢ�HSl���һ�6�l���$�\l�����Nc��mY�"�
QҐ�W+�mYv��h	�/�㜈-��[b�l��h�EM.��3�7����e�nہ�YV�췳�IE�\H������i��6�뭏;6���w罗o��>{�x!�&������_R�p;=h�k�\��Q���(��2qQ�����*ʻ�Z�~��Z� >�]�B��{�`����RS3W4L�Wxε�tDL����DB��C��� >���Q	L� 9s5K�h��D\������7��a�Jd�{� �]��>��"��p��7&�s�W�ߖ }�׀|�\�z#Ъ��^�#��(S%y ���0���Ж�������9���/�+�<M��Q���!��G����Fɺ×�y���Zz_Yp؊:t-��m@CjF�4��uޭ ��Y�o������x���UU`H�U�.��� >�]�@�c����$���e��L |�xε�r�9\�iY��d��&�y��@=�٧�Ĺ�z������˓�<���� �ֹ���xJ^�q��nW^ �$�bCrhWʴ�r�z�gM ��f�{��)�^H���2`m46�<�V�=��Z�fȶ��u�F+nRi-�ߞ��թ&kN)a�z�^��YM ��g|�:�V�Νb:�<#Y��� >���sp��g����(ޡ�)�h��d�ـ���>u���-�!��T�@EO�b�+H2~�l�]�' "DH �������QN�GUd�0a�h ~s���� �aJ�bB O�$D����f ��v���os��`"� D4s�|ኤt$CvF�e�Z[BЭh[y���2S@@�� @�!�>� ����z�@:���T:�U�@N�qؠi�D� x�)��6�P<���=��$��Κ�gJ��1�#X�rhus��@��`�R }���Hᙙ�9��7�}�,�;y�����f��|�@���mb�����M�$��;%݃�=i1�j�v{7�r�z5� z��w}���nF�Y"nI�~����;٠}k\��� �z�$wQG�����U���@�� �� ���yԟ߮�>�Ժ�Y&�BCrh�Z�ܷ����ЕW?_� ��^�n�4ML��'"��g�s��@������ruB�3믻w$�gm�T9�R� ����~v��B�?ou��w�@>��h\�����f&Ĳ��l�F=s��ڹ�M�F�����m=��Y<��ߞ�w�a<��o���9@>�{4�� ��w�!%�A�_����5VVn��y� �� ���yԀzٽ�3>�|�i���x�24�Z�>�~v�:!D���^�]Ӏ7�h�S4�M�ܪ����DzU���0_�M��Z�ܳ@�s�eɉD�wV`�o_t� �}x�`�B�(��zT�Q�TE�]MQ�.0�F�e�"j@n[�{������ۜ�]m���ݐ>\��\�]ɐ��4�A�!���厹ֳ�Q���񸶬I�����m��V��;�'A�٦���"7i�tDn�3/��b��N�SCP�v�Lv�V3qWnp����3Z�K)��z\Y0���lZ}����� f�R�켮��Y�a��x�s����	ET��I7���&�֭���1��!�ʰ�
�Մn�<]yx�A�����K^ �Ƅ������}�,�9�)��l�>@qq&�Tґ����}��do�� �{� ��s���·Q1�^6c��i�4{:h�[x&w��pu��"j�U)��/7H��`�[��; �u s�xVۀ��J'&��v���/g�r�t�~�h\�)K����z�J<�M��ZŸ�\�9������������z#i���d��zU�z唀�`:�z鬼��^���h����;�uټ0 4�#�
?��۽�{gM�r��g�b,Bܼ�4��� >]�<�@��� [)�|�^2&Ƅ����,M�� ��@;��6�J˽ܲ��� �9 ��@˰�e4�y�s�2�M�:��q�ͶϭJnLWd�e�c��s��T��Je���jܽ�F��<l�	#��/gM �[4�e?z��޽�ùqto���9 |� �:����{�I�����Xu��܊<i94^Κ\�zi� FlaD!*4E�
ʫ�b(��3�צ�-��>�UP���<s1�!�U�:�>nـ������ ���!<�QH��MǠ}�)�w3�y��@��� s�� ����"�&��~�vӴ�B�,][���68�Ɏ���v�k�Bg.���R�Yq��Yxl�Y��� �]� s���/(���������_�2&4�BCrhr�o|J"d�o� �����������O:4�hB�p�*�+�;��s�ޞ��$�O?z����>`�Ht��VAwuwX�D�vq��׀n�fB�Tou�w7$���{3u����f ?���"���-�`7l���B�ǂMe�#����]��r�j��JӣWs�Pqt�[�7o~w����;|��G�''�[��@�|�@��O�g��3�WSKA��d���yZ�9B��%T>���?z���3��	*���}D�*�)���V��� }�� .�=Τ���Y^,kjf�ieU՘�!y!!(�$�ߟ�x�_���(���IS�~��ދ��D���ܚ9e4
�����`���6d$+"��*�w߳��v�pe� �=v��N;�=�*PM��gևs�gd,̗tY=;e�mc��ܭ͡�a��qƋ��팍�[v`����v��jBv.�X
qX�n�6:���lf[d��hF��۞c�Z������*�V�n,�t�*�۟������s���;h�tz;ra�8�[n��z�L�"4��L�kM؁{KO�q�S��z�+u���{��{���{ﾕy���K�&n���3��Z�|r�Gn^5�2�9�$������{����#��),�à~\��}�)��f��,��򪤞<��NG#�>��˰s� o����~�s+/v��3t��`�R �s�s� ��((��s�$�������:���>���%�w�@9�;֛P���kw7H}�@=Τ |� �u4V\9�����@��)	�G�m�Η�<]��6���ĕ)��T�mu��.��w*�MU��v� 7x�rJ!/�0�����8��X���<�w�{��Z�Rz"ݨf�wz�>�T˩ )�:���o.�+�*���l��Ň���_��x�`q��Lb�!��y�y�.�ߖ��� ?��Q�g�L�Ԕ��5dsUk �]� ����k�� {��)G��'I%1=:�x�ih��伺�l��g�RoPL!��\�S�y1dop��r~�hr�@�T��@�4��(��2��j� �]�<����,__���w�H;�;֘���d���y��hO�w]���"H��T:�A�v��נ^�S@�2����n(�X�TݬI$�z)��x���X��>�s@=��E��I���p�>W��Ik���{�`�ـ}/]R�.�ӺQ�p�8��H��{g�����Pt��g�/��~w�k|>�W�\�?��|`�x��l�J"~���Հv�+cO������[�����6wz�`}ެ���Jd>�UU4��MQVAw5V����>����JQ�T���s��`�8�)�*��.d�����}X�_��,I%�!�V��X�@CC�'	��%y5���P�nJEU��T�\�7l�<�IG�(��|���� �^W�[��ӉyȢ)S!s{��x���]ĉ��ێ+��ɤy�==�8�t��<s1�!�s�w4�e4��}�<�/gM��:��o7R,s�4��3�Dɳϫ ����7�<�L�y����I��G���@��SD)��ذ}|`6e�]��R*mUM�`k�`�x��l��Q;]�zk������ٍ'�[��n�f��u�|ݳ �QP�-@���0���$E�	!�/
�F! _ĝ-`Fl� B0!H$ ~$O�}���!!�R1#	��7��"#/1$���>V.�7~O�g�1Tń�_�!r\Y @���D��k �r�ǅ h�d�ê	0LP�*��)��*`�~��Q(�#�??�� \ޖ��Pڵ��˰DM ��A�<ʪ����*���Y���g:갷���+G)�VSk�MYP����\��@;	OC.vQ4-r9�gn���d�ù�mF���s��(��\�j�M��JYdL�)hл��8[T�9�݌ɂ�U�[[���T�=��m�.=��B���M�`��H�d��)8U�Wf��Pнn�;�6(�lv���/v�[=�4r�k���.�=�+gE4�Q�`PV�W�%��kX�6y��l��W7�IeK�HH��b�[�5J�t2�.�ڰB��8]՞,7����j�s<q�#f�yL\�Ƙ�h��>��طm�k�)�
�nT쁫j�t�헔9�8�� �S�QM="�8����٩gC�W�r	�i0�:%��ݻ�6�2�٢;5ݖm<��S���+�.Kv�nU�����i�K������*�s0��b��Ɔ�s�^\n6j
a�hh{,85�{��l!N���I5����e�fqC�F��lc],���a���)����" 6*�E*�L�t,x�,��bmP�t��֙o�����t��>]����Χ��Q��x��Ym��MB���U�ؐ�Uy�*��6�ۮ9Bz�vl�<��<Q��۲d�͂����<��+R����;m+�+�kaX9�q����7T:�����5؝WlAX� 򠝙���g�:0�9���l�v��=��@R��7�s�)bgu�M�U2�����&ڵȁ��J�l��h؛T��!�џW¹�^y	����qe�ی�B�5��Erѝ�uӍ/jx�q�N���r��(�X�2,T�!����nYh���#�8X�	�sy_`��ϴT�H�y��\�Qq�lTA�����n1�����:��Z����
l�r��Ֆ	�SV���n\�ef{e�\q ��mΈ6�K�r�W[,ج�c6�y�`��k
[o=.ո�)=fL�]L-�>�|��)�U�!��b@���G�t�j(�� �@����O���7){S����B�kC⽠��Px�݇\��X.JV�"=��X3^���9��G���[=m%��%�a������ �s�<�^.Z����ۗ�5t�НD��x�*���	�l)��Ƶ��5�2K6S�k#�����Z�:�{/��W:��uˀ�9�ʇ\�O�.QT9`z��v��$\v��*&ًvX[�55��0�5�nd3Y?(�(��s{m�~�sPO5��wH��O �Q�Ee��,>�zY:�[U�;~w����<𹷵V�]�}/]`ͻ�H=�ŀ��0Y��"C��>W��[)�o���7]�=
#�U�\�I7%"���q�����h����������ˑ��Lq�hw<W���7����u���vq�7��&�T�M�ܪ�Sv��l�=	B������0��X�h:��Q��"�N{'nzƔ��;=mͭg��=�"5J��ٙ�i ���I��G@����>nـo���$�H7�� .��ꋺ��
-UM�`7l�K��K(�G����3@�;:h+����m2�#fT�Y�o���7]�����Հou��q�Oʛ<�#s4r�h-�X��09%?>�������B$�3&j:�f�6��bX�'����ND�,K��ߦӑ,K�����ӑ,K��}�M�"X�%�߽�I.��ݳd7�k#��:��7@��-�����ŗ�����ŭш�e�'1O����X�%����M�"X�%�����"X�%���~�C�,K���{ٴ�T���$'�����%*�E���2�,K�����ӑ,K��}�M�"X�%��>��iȖ%�b}�o�iȥ�bX��z{%�frK��S5�Y�iȖ%�bw�ߦӑ,K���{ٴ�K	���!��9^��6��bX�'��p�r%�bX����Y�In��f��k56��bX���>��iȖ%�b}�o�iȖ%�b}�}�iȖ%��#2'����6��bX�%<���a&���Y�2�Zͧ"X�%��{~�ND�,K��ND�,K���6��bX�'���ͧ"X�%�{�M�n�C�=�֙�l9�x�ӴF�㋡�1w��:!��M ��ٍ�<>�&�m9ı,O��m9ı,N����r%�bX���{6��bX�'}��m9ı,O�N�م��ff��j捧"X�%��{~�NC�@c�2%��w��6��bX�'����6��bX�'�w�6��bX�'�By��̙��fkSiȖ%�b~Ͻ��r%�bX�����K�dL�����ӑ,K������ӑ,K��ݛ����	��e3WZͧ"X�����M�"X�%�����ӑ,K��u�]�"X�h� ��} ���Abj'���iȖ%�b~���Y��,�4dњ�jm9ı,O��m9ı,O��z�9ı,O����ND�,K��~�ND�,K��v�8���=�Gb������՛t��)0�h����p���U =n�N^��G3�6��bX�'���iȖ%�b~Ͻ��r%�bX����m9İ?�D�}���r%�bX�u�'���V�3P�[�ͧ"X�%��>��i� �ș�����iȖ?�P�Dȝ￸m9ı,N�W�ٴ�Kı)����$�d�2挺ֳiȖ%�b~����Kı>����Kı?w���ND�,K�}�fӑ,K��|I��\��e֭�[��ND�,�`dN��ߍ�"X�%�����v��bX�'���ͧ"X�%���ߦӑ,K��'m�L-��sCT��ND�,K�w��Kİ����f��Kı>���6��bX�'�w�6��bX�$�w�יn˭]j�P�c�)b9�$1��!yc<n)*^��r�T�f�ScmI���4��^z[�W�c����^m�;'Y�I�q�K����֧�ݎbƏcz�ӎ�.�2#��@c��P��A\K���( AL�;qṗp��0t'4��Y�;�۰�p�
F�p�t�Վ{м�t����Ê3���nλ���@U����)�'Wk����g��ލ�t������ë��ex�{e�Y<�A�nǓhr6���Z�ND�,K���6��bX�'��~�ND�,K��ND�,K��8�_�RB�����M�H��U2fkiȖ%�bw���iȖ%�b}�}�iȖ%�b}���6��bX�'��m9���,N���Y��,�4dњ�jm9ı,N���6��bX�'�v��iȖ4X�'��&��!��צԐI�=附�L̹ff�pI�>��~�ND�,K���6��?�dK������r%�bX�￸m9ı,O���d���Yp��e��M�"X�%���{�ND�,K�{�M�"X�%�����"X�%��ݻ��r%�bX���I���P�r�ՙU��`2�G�'��1Ԗz�%׎�I6sp]�!=��.\�s3[ND�,K�w~�ND�,K�}�M�"X�%������r%�bX�w��ӑ,K���I=�K�}2]j�M\��r%�bX����m9�������9����iȖ%�b}��iȖ%�bw���iȟ��2%�ܞ�ff���0�5usZ�ND�,K����ͧ"X�%��w�ͧ"X�%���ߦӑ,K���o�iȖ%�b|}�N�I�̹�嚹��r%�g�"w^��m9ı,N����ND�,K�}�M�"X�%��ھ�m9ı,Ow�p��Va34L�j�Y��Kı>����r%�bXQ����Kı>�W�ͧ"X�%��w�ͧ"X�%����OI��j�5��2��nD��١�g]u�wl��X#���7�}���+��R)lg��u5��w�{��7�������r%�bX�}��fӑ,K��;�fӑ,K�����iȖ%�b~��d�%����T�����Kı>�W�ͧ"X�%��w�ͧ"X�%���ߦ��~��,K�o�m9ı,O���2j[u�	��[u��r%�bX�g{��r%�bX�}��m9Ǧ�H�D�@�Ø������D����r%�bX�wW�ٴ�Kı)羷�[u�K�tj�Zͧ"X�%���ߦӑ,K���o�iȖ%�bw����r%�bX�g{��r%�bX���'�	s/�K�[	���ND�,K�}�M�"X�%��{���r%�bX�g{��r%�bX����m9ı,N���l�)=�2�˚��K��$��웬�����'b�+�mq��J9h��U-�YsMK��jm9ı,O���ӑ,K��;�fӑ,K�����iȖ%�b~���Kı>�j�R�e��r��j�9ı,O���m9,r&D�>�w��Kı?w���r%�bX�w��]�"X�%��x�����	����]k6��bX�'�w~�ND�,K�}�M�"X�%����z�9ı,O���m9ı,K��w�s5��ѓF����r%�bX����m9ı,O����iȖ%�b}��iȖ%��C�H���#���k���Kı>���L����T�����Kı>���]�"X�%��Ǻ���i�%�bX�{���ND�,K�}�M�"X�%���%�N�C]�F{Y!8��P
��1����}\j&oa�L ��wN5���VG�nEc�w�{��%��w�ͧ"X�%���ߦӑ,K���o�iȖ%�b}�w��ND�,K�{���[��fdѫ�k6��bX�'��~�ND�,K�}�M�"X�%��{���r%�bX�g{��r%�bX�Ğ�ܾ�]j�CW56��bX�'��~�ND�,K��y��Kı>��ٴ�Kı?{���r%�bX�d�nfR��0�5usZ�ND�,�D����ND�,K��fӑ,K�����iȖ%���P D��{����r%�bX���<�-�˙��ˬ��r%�bX�g{��r%�bX����m9ı,O���6��bX�'����iȖ%�bm�<�����$�)����L2�fe�3 ���)��携�g��:���ӝ��2c�6:ȨͱG5:�%l�˶y�K��EӦz�V��u�=��%;OMs t��n��Igî^�V;V���jm�NI ,rk��gv�a�d����9�1p�	�IT/��5Y�3ͥ#��)��78��Vzi1ٺ:h-�+�\�:{&*�x��u���ww���w���=�q���]X뒒�#��sK$���)�*΅w9�����q=2��Z�t��S5u��;ı,Ow���r%�bX����m9ı,O�ۿM�"X�%��w�ͧ"X�%�OY}u%�f�Ն����r%�bX����m9��DȖ'}���Kı=���m9ı,O���6��bX�'��L�\�WZ�jk5���Kı>��~�ND�,K��{6��bX�'��~�ND�,K�׽v��bX�'�ϼd�Kn�asP˗56��bX�'���m9ı,O���6��bX�'��z�9ı,O��ߦӑ,KĿ�z�0��0˙5&]kY��Kı?w���r%�bX�����Kı>��~�ND�,K��{6��bX�'�v�1����K��l���&�l�;&4���X��G�b2�R���;v��n&�����w�%�bX�����Kı>��~�ND�,K��{6��bX�'��~�ND�,K���L��'�L�P��3WiȖ%�b}���m9|�_�$�~���'�,O���ͧ"X�%�﻿M�"X�%��k޻ND�,K�Y�)o��j9r�jm9ı,Og���r%�bX����m9ı,O{^��r%�bX�w�~�ND�,K�z��-�L&f���]k6��bX�'�w~�ND�,K�׽v��bX�'��ߦӑ,K��{�ͧ"X�%�OY}u%�f�Ն����r%�bX�����Kİ�D#�z��m?D�,K�?���iȖ%�b~�w��Kĳ���߿�����F�m	��ݸ.qWi0x,�-�4L\�\]�y�8�v7���#Z�jk5����ș��w�6��bX�'�fӑ,K�����a��L�bX������ND�,K��ږ�L�桙�56��bX�'���m9ı,O���6��bX�'��z�?��&D�,N���iȖ%�bg[����0�̺&MkY��Kı?{���r%�bX�����K.�� H0I���J�|o���p�R#$!B�V1a �@�H�0#^�II%��I�XF���G�ĐHX�h��7�^��c��p&�I/8E��1�$X$���0�F}6�����@���Sq�~�V
H��X�&� A�$��H!�$��%!�cA���, �0�!b��!R0�"�R$#q](�ӂ��$F�	���4�D� ��h��b�z�ʈ�"xȜ������Kı>��ٴ�Kı/�=�,����԰�\��r%�g�@ȟs�m9ı,N���iȖ%�bw;�fӑ,K�����iȖ%�b_���[3f��Mk.�6��bX�'��ߦӑ,K��w�ͧ"X�%���ߦӑ,K���o�iȖ%��{��?}�� �ͣѠ��L)az3���S�=$�딛���LV[�:�zc���\棗-֦ӑ,K��w�ͧ"X�%���ߦӑ,K����]�"X�%��{w��Kı=���=%՘L�)���m9ı,O���6���1ș�����iȖ%�bw޻��ND�,K���6��bX�%�}=e���a�5!����r%�bX����m9ı,O�ۿM�"X�%���}�ND�,K���M�"X�%�ߡ�0����֩�&�SiȖ%�b}���m9ı,N�{��r%�bX����m9İ8 �� $�V�]F��"��/ʿ&���w�w�iȖ%�bx>׌�Զ�.5̹���Kı;��iȖ%�b~�w��Kı?{���r%�bX�w�~�ND�,K�{�m̾%Ѭ��a�hЌg�q������u��:��,sƍ�U�=�����n��ˢdֵ�ND�,K���M�"X�%���ߦӑ,K������r%�bX���ٴ�Kı/�>�.{N�5,!�56��bX�'�{~�ND�,K����iȖ%�bw;�fӑ,K�����iȟ�9S"X����[��WXj��֦ӑ,K��w�6��bX�'s��m9ı,O���6��bX�'�{~�?���ı;��r����ur�jm9ı,K��kiȖ%�b~�w��Kı>����r%�`2'}����Kı=��M��Kta34L��f���Kı?{���r%�bX�}��m9ı,O��ߦӑ,KĿ}�kiȖ%�bk�~�͓�e,��O8t�i�\�mq7u��wH��A��w%E�#�-���,����2k�g��l=u���!n��;b\�gp�f��ۓ���r�h�-v�	�H��PL�H1���^u�ۮz���[#S��>�
�e��ӂ4l��̷&N����zV�z�g�����j��j�����N\Y���}��3H��-�Y	pє�|
�L���&�����8�4b��2r�S`�et��j䋠]�Wj�==�v��2�m�������ou�b}�o�iȖ%�b}�n�6��bX�%��{[ND�,K�{�M�"X�%��þ�0�����T�Y���Kı>��~�ND�,K�����"X�%���ߦӑ,K���o�iȖ%�b_����Ƭ�˄�L�sSiȖ%�b_�����Kı?w���r%��2&L���s�m?D�,K�����r%�bX��7���u��r]�f���K�ၑ=����ӑ,K����6��bX�'�w��Kı/�{��r%�bX��{	�=�S3R��h�r%�bX�}��m9ı,?�T#��y�6��X�%�{���m9ı,O���m9ı,O�w��=���.8mř2�$m��kE��E\�����%���+r]���3��z���r%�bX��ۿM�"X�%�~���ӑ,K���{�����dK����6��bX�'��6����ur�jm9ı,K�������t ���N���K����ӑ,K��}�M�"X�%������r%�bX���ܞ%�0��&SS3Z�r%�bX���p�r%�bX�}��m9ı,O��ߦӑ,KĿ}�kiȖ%�b~���{5�d�ѩ˚6��bY��2'{����Kı>����ӑ,KĿ}�kiȖ%�b~���iȖ%�bx���2����T�Y���Kı?vk޻ND�,K�w����~�bX�'���iȖ%�b}����Kı?|{�$�9.f[�Kr���<7;t D�'�t�s�T88ƌ��T��*V��ďfˊ>�~����{��}�kiȖ%�bw���"X�%���ߦӑ,K��f���Kı;�o����32互k3Z�r%�bX���iȖ%�b}����Kı=ٯz�9ı,K������bX�%�{������԰�kZ6��bX�'�k޻ND�,Kݚ�ӑ,v�""D��b�����&����ﵴ�Kı?w���Kı/{o����ڹ����3WiȖ%�b{�]��r%�bX��ﵴ�Kı;���iȖ%�b~����Kı=���}3sQ�ɬ��r%�bX��ﵴ�Kİ�H���ߍ��%�b}��]�"X�%���w�iȖ%�b}���[�̤�e�>v�>�qN3�7p�-�n�"m08aZ.^ɥ�`J9��q��lk��vN�����oq���b{���6��bX�'�k��ND�,Kݚ�ӑ,KĽ���ӑ,K��d=�/��L��jBff��"X�%����ӑ,K��f���Kı/~ﵴ�Kı;���iȖ%�b}羳0˜���T�Mfj�9ı,Ovk��ND�,K���[ND�,K�{�6��bX�'�k��ND�,K����<jˬ�L�3%�]�"X�%�{�}��"X�%�߽�ND�,K���]�"X���G����J����܉�7���9ı,O��,���[��˒膳5��"X�%�߽�m9ı,O��}v��bX�'�5�]�"X�%�{�}��"X�%��g��?ٙ�[sY�n�F�a�K����x�Ŭ�*������I2sv�n��S3R�I�k��%�bX�����ӑ,K��f���Kı/�ﵴ�Kı;��ͧ"X�%�{�왅ˆz�55).jm9ı,Ovw~�ND�,K���[ND�,K�{��r%�bX�����9��f	"|��f���j�`��s�^(@�-���n	"D��w�iȖ%�b{����r%�bX���잲�L�)���m9ı,N��siȖ%�bw�o�iȖ%�b{����r%�bX��w��r%�bX��><{.�MMf�!33[ND�,K�{~�ND�,Kݝߦӑ,KĿ{��ӑ,K����6��bX�&�H&��#�F(0�@'ݳ��}u3VY�Zk52��\�0�����c9�Ia�u�ǰ�U��v�<�v:�i⻮P�%X&ǷuG�h���"�!Ԏ���:�H�H./6���Ƅ���d��v:���mk��\�]�V3�m����*�UnG�@O!fx)W�l]m�q�]'r��)�u����"ۑ�g��v��1��Ҳ4Wm8mL� �:zِk����{���v_�]�G�S��qk�ի�k*sՋ��y�v���U�ׄ���]]j���֧�ؖ%�b~�׽v��bX�%������bX�'~��m9ı,N���m9ı,Oϧ�,�.��3P̗5v��bX�%������bX�'~��m9ı,N���m9ı,Ovk��ND� ʙ��v����.�33%ԓY��ӑ,K����m9ı,N���m9ı,O���3iȖ%�b_��kiȖ%�b}���fe��55��3ZѴ�K��RD���6��bX�'���ͧ"X�%�~�}��"X�%���{�ӑ,KĽ��.dɅ��jjR\��r%�bX�{]�fӑ,KĿ{��ӑ,K�����iȖ%�bw�o�iȖ%�b(�=���L�?��$�Z�W=��`�n���s�pmZ62W#����햡d����]�Me˚��5���~�bX�%������Kı?}�p�r%�bX�����r%�bX�}��ݧ"X�%�ߧwd��h�fh�ML�kiȖ%�b~����4�n1�H�~QM<�Ȗ&���6��bX�'��}.ӑ,K��y��/�)!I
H[Drk��ɲ����ND�,K�{~�ND�,K��ޙ��K�Dȗ����ӑ,K�����6��bX�'����.rK��S5�Z��r%�bX�g��ͧ"X�%�~�}��"X�%���{�ӑ,Kȃ2'���m9ı,K���,�.��5�,��ͧ"X�%�~�}��"X�%���{�ӑ,K���ߦӑ,K����6��bX�'��5b���`�ۘ�Ƥ�P���#`$gp6y��\jۗ��qp0o6쐨��k3Z�~�bX�'�����Kı;����Kı>���͇��"X�%������Kı/�?�2����jXYu�m9ı,N���m9ı,O���3iȖ%�b_��kiȖ%�b_�{��r%�bX�����2�}r���njm9ı,O���3iȖ%�b_��kiȖ>xA ����A"i�
6~��%�����"X�%������ND�,K�j���[陚��5���r%�g���������bX�%�����r%�bX�����r%�bX���fӄ)!I
HOG�$��V��eU�B�Kı/��m9ı,?������O�,K�������r%�bX��wא���$)!sMP]U"I��n��;���[:��Đ��!�";�m����q<V���.��Uk!~!I
HRB{��ӑ,K��u�k6��bX�%������bX�'��ND�,K݇}�p�����T�eֵ6��bX�'���Y�� ��W"dK�����r%�bX�w���ӑ,K���ߦӑ?��
�RB�^'�OXd�.�UUwY�
ı,K��kiȖ%�b~����Kı;����Kı=�w�ͧ"X�%�����2�332]�f���Kı?}�p�r%�bX�����r%�bX���fӑ,Kf��D���w�kiȖ%�b^��ٙsWZ�K�Ѵ�Kı;����Kı=�w�ͧ"X�%�~�}��"X�%���{�ӑ,K��-��I�0��x;=m�������pu.]���@[g��e��f�m���a:���~����%����m9ı,K���m9ı,O�{�6��bX�'~��6��bX�'��{a��a�5\�kY��Kİ?�Vg�����%�b}���ND�,K�{~�ND�,K��}��r%�bX���rz�f�&f����ֶ��bX�'��ND�,K�{~�ND��"{^��m9ı,T�w�!~!I
HRB�#�u]�6]]����iȖ%�bw�o�iȖ%�b{�ﵛND�,K���[ND�,����~6��bX�'����[�frK�Z�k.����Kİ?�'����f��Kı/����"X�%���{�ӑ,K���ߦӑ,K�?
� D�~�l�*~	�0b�#���"Èh��0��$'B��u�� �BC��
��@�	��<�H`�R!b�� T�"Q$B���T�]F6E� ��!	�I�9�@���9�?�� ,X�-Ia&�B��ݳF����@0f`����`&���#��,�BF$HE�6����!$## �%�BA�F=5���p+$�R"�X2H1�0!�	�"�	����@!E�U��p�_�����}�d��,X1������ "��f�6�1a @�,��$(�Wq��[;�ֵ��ڎ-%Uu\�u�9�d6%�oe�y�� \��\���N�:d6cF����-�xBY��m�61ŭ��n��܎ܪ�V�P�`&��� �h���0��S!i$B7S�s/q�6�y�{E��h^����vju0d��`��C4��iP����d��e�&y`x���J��.V��-�h�'W\��v;��kW9اLhm��qu9��SH��Ⓧ�V)9�5m�m�q�F�Q�m��3�1���9��s[(`y��X&yZ�;%6ц�n��y�\�k��<=t2�at���#C�c�Wt���	����a|�h�c�YX��"�,�$m����x}��\��J�!*���#�*��b����x۬E��ږE{�7<
�Ð��V��(0d�fz�Lr�����e���xꋬY�m탔�goc�NM��v���5�jL�Nl𜱱�J��J�H���4��v�n�ظrLAPj�j8��gWg�Gc��۵�4XՌV�� �K���vR���ۜ��R��(�r�F7�r��*֡������0��R9wR���mS��1�ᮔ���u�x�yL��@Y&�9nV�MU+l�$�d�ˆ��6ju�CE�g�`/G�����㚐B�Pو��-��v#��rYTΰ���C�}/l��E�Y�H�n�oN]	\���J�!E!�j�aѱHQW�[Xz�y��i-q��rK��c��7(a6R�y��m`N�fl��v�e�gYڙ�E�/D��ډӻNd�BzuK˗hNq=
K�-u�&\����Z�&�.F���Mg�����}��d������]�!l���o��1J\�H�^����L>`��t��1��$�F�\`������j
vi�tl�@5�1%�6�3I,�CÔ7��@��k[���s��2;:R�/cL;�GF��],�w��M� ���8�t�c����F��2�VjI4f��~h��;"���!����z�ĩ�Q�+�V8�h/_��?
? �D�$���v�ֲX,��+mԮd5v9��]X5J�vw�Tۈ�cp�{DmQP*.��fm�b������v.z�óP�[��]�A�[k�z�ϋ=x{z�8c��f��T��ZNv�m��xPm�'�63^w%�
���6�r(��{n�ӭr�����6[�H/cZ\3�˸����ք�ձ�ݧ�3Ā�J��e�y����
in��	�WZ��!�ф%�˸h�5�&l\����<��yX�{g��b���L�n�u��uذ��ʴ�{���oq�X��{��r%�bX����m9ı,N���m9ı,Ow]��iȖ%�bw>,;�L��\���f���Kı?}�p�r%�bX�����r%�bX���fӑ,KĿ{��ӑ,KĿx�ٙi����lfkFӑ,K���ߦӑ,K��u�k6��c�*�"dK��kiȖ%�b}���ND�,K���&2�j�j����r%�bX���fӑ,KĿ{��ӑ,K�����iȖ%��3"w���iȖ%�b{�W�}3sQ��f��ND�,K���[ND�,K����"X�%�ߵ�]�"X�%����m9ı,K��i{L%���Y&�nL��p1ˬ�Hx����^���W����nOBY�j���\�2����ӑ,K�����iȖ%�bw�{�iȖ%�b{�ﵛ�@��dKĽ������bY
HN�����nn��D]լ���$)�����Ӑ��"/���<�Ȗ&{\���r%�bX��w��r%�bX����m9ı,O�v{%�39%˭S5�5���Kı=�w�ͧ"X�%�~�}��"X�%���{�ӑ,K�����ӑ,KĿ�K��%ԸMh����m9ı,K���m9ı,O�{�6��bX�'~׽v��bX�'���Y��Kı;�}	�.��34CY��ӑ,K�����iȖ%�a��b���?����%�bk��Y��Kı/�ﵴ�Kı>�~�|�jey`�gάkVv��:�՝c���G�YP����h㓍*��(7�Fӑ,K�����ӑ,K��u�k6��bX�%������L�bX�w���ӑ,Kħ�o�L&d��V�h��]�"X�%����m9ı,K���m9ı,O�{�6��bX�'~׽v��bX�'��{a��0�5\�kY��Kı/�ﵴ�Kı?}�p�r%��B�B� ��D�L�z�9ı,O��}��r%���vh�"�T��EJ���ВS������:��@>��@�^�D��8�7sj�Ÿ��� ���>�ʀz�8,EP�dc��Jƌ �Gq&��y4\n��v.�<�M[mo�e���r�v�g;��; ��*��Z_b�\�Q6I�m����7�"!B�>��X���k��6~Ka�Dx7��27&����h�ڴ���}yf�}q��yLq�L�7�np��� >z�TA
!$$�""�x�:�w�7$���fa�d��ڽ͸��� ���>�ʀw�n g�B�.�1�ȰnH�9lgs�݂7�:��E$���0u�n��nK/i�o77r y�`ye@;ط {:Ǡ}�
"��ǃs�ܚ�[���
*�u�8:}u�=w�}�	�RH�QFL$s4|�Z��@>��@��w4Åb`ނ#P#NE {;�y�����[�>��q"i�`�r= ���߭��9�h��=����fGB!�QS�mt���܋���9յ��8���Wc�N;c,�WY��C�.�fu��(�71s��v���ru���Gd�K�p<�F� ��X�tm�$ۆ����	GD<i���ֶ�IL<�KЊIZX�0T/n�����4�����`%��$��I%'s�2V���Na�z��Tv�O�˴�����[�������������ӹb�^ۈ؟c�s�����ֺ�hڅXoa����th�o�F��y��h�ڴ���}yf���ց�)�H��NL�9�-��w �v��T�������<l}dK�1G���c��,�=����;V�~k�b�bND��<��,�{�gc��ڋ�S��7&����h�ڴ��^�}yf��8���1�3Ț[�
n��s�«[&��{Y�m��.�P��(��x!��A28Ʉ�g�^>�h��� |��D~���ŀo&uAU�%�Ԛ˚�ܓ�g���)T�1��"?�W���Y�I��>�e@;ط }��q"i�`�n= �����Ӿf%x�ՠv���/��eȅ�na[�� ��T��p���着{q��c�cR�'&h�ڴ��r y�`�ʀz�@,�,.��Q�ٷNn�[�,m.Q�N����fv'�7���a�(6���QŠ^>:��; ��T��p��]Ve�e]柶�s7 �v�,�{�gez>9pJc���Y��>���	���n�!�Ċ�('� ���<��Ͻ^����^���Yr�A2=�h�ͨ{�gc��; ��s@������F�!8���^�y�`�ʀw�n ��*̫���\�����B�K��8��v�qs��c�gv��qPm��eƺ����,������=� �b���r���֡A��L27&����oؑ�:@/z��p�3��7�1G�	ɚ��n �v9 =˰ye@z�̰x��C@�Z��@�rנ{�x�>��?EN�s�~��m
��Jf�������� �ʀ{�n �v9 �ZV������X�i?<���ܛk
.�Wo�V��	��(嶣�&�b�ݓ����7{�`m78��u�_�6_uhQ���)$#��H�hqڴ����� �ʀ|�8^d7/Cr�v�gc�ܻ ��T��Z�ƕb,�L�Mǡ�<��ξ��7{�`m78��u�l�r!A��@$�h}n��K���@�u��ܶh�fg����q`�P���s�cK���p�7m�a�c�RC�8!'P���[��JE��)<�v�R\9v�&D��1��v�y��C���uaP�ktAsR�f��ީ˴u[ą�U��"���uq�`]�s-��i�WI��?����}'%�++͎D����ڶ�B�9��Sv��%��q��v8:��J��� �V�^�l�m�Bvd՗Y��MY�� �3{�CY����ӡ�<J�v�I#�$�7.-��v�cqqu���L�ݘ�<�u��<a�������O�{[N�^��%��v,��GQC��1Ŏbn-��נr٠}����v��Fp�ƺ&$��N7�k��Ň%	L���9Ӯ���X�1������h}n���@�|u�9l�=�̹qG"L�3h�ͨ�[�=��@�����s.5��Tm��(�mx%�7�uE�1+�u�ɹ������5Pb��r��m�%���ۀ=��@�����qn~�X�(�$��q�9lۙ�	z"P�%
�wذ�]Ӏ=��X�p(D(4�9$�>�����Z��@9�f��ex�L�(�XV�� �p���ܻ ��f�W8���d2A7�x�c��� ��x��78�$��dUU�g�����}lu�շ8w�V헛'6��8�e�Y<�A�s��a����?���??/���*��g;��^�e��e���@��)�}]�@�|��9l�9�f\���&G0�C@��۹'~ϻ��џ�1 ������6���5 _�� ���4B���@�B�πB�H0F�� )�v=�B$La~	�$����e΢�؄d䜹�~~I�Z"u �H��$"G$Hi�!��>B ��V H���L�q �	�L�К^ |�F7I������Y���S��?	$d�0
i���ӱ(@��"�'�&Nl�G4�M|D��Q3�!�y��?���������&�Tx�w�>����@��4qC�:����D�
i
��)��x����]����پ�}zgX�7���ӑh��= �]�}� m� �eݵc�w�xn�e��@�`ye@y�}�&�Pq**��0��$!����N���̓�<�c4]U �S���9��1�kh�4�9$�=�����Z\哹�{٠s����gLQę�nL�>t��B�:[� o���7� �4�Ƣ��&��*�,��[4~���ڴ
��\�&$��R9&BQ3�������s��$�e&@�9����ܓ���v�mф��5��M߭��;��;��m��-��s01�D"mF,q���rmS�ރ8�ے�mlr$������X�o��:�k#��H�z+�V�Q�Y�r٠_���=��'��"54�ZG8�=
&C_u��ذ����3-I`
	�c���l�/��i�3<�.Wޭ���@�����
a�wv �e@=ط j������g<N�cr$�6ㆁ��@�8� >�� ���p�A�M�˩�5.6�E��Z�!#d��1)����!ՍT�ܧ���v@P0��:M�(�綫��ε��n��W&�wlhWT��!����r[����KP2�<j�����bb����2��H+�	qk�+BY=.z� v�eUd�s>T
��.i�4u�2�#:�vz�[�^�7 �i�r<���/j���X��mt�s��v��G�LP]߾������9���h�{���68�Wd�g����W����z�f^�^e��
L�.Mu\,~�߮?o�@r���n�Ÿ�W���h����d�= ����>U�}�j�=��W�s�GRHS	��I&��7 �b� ��̀��v�j�$I��L�8�?g�f.Yޭ�[٠r٠{�Jh��F����r\�;�����ڐv-�:�� ��0B�<Py�LbQ��W�GQ�LE+��DӦA�cy�Vذ����ܻ ��R�ſ꯬=b�l �)N�c`�$�@���ٞx+� �����P�g��]��r� ����3�'S1�k�� �[�}gs�ܻ ��R��elX���b���C��x�e������rS@ⶽ�g��Q�K4����� �v�v��\�}gr�癞z��q%��i��K2")	䐶�c�M�O��17�i�	�t����'��x'0k!$��Κ�����@9m����e��28ɒ)�۬興�>��� }�x��fr���>�t��xނ#P ��@��z��� ���*, 7قD�9, ~ �o���nnI�｛�s�+���1��zį{٠}l�q[^��.r� �)J�hQ�Ц����9�Z� ��������I��t Ф�S cF211�Vv,m�:��n:���9����$�6�s��������֮@>��r r� ��R��eO��$X�mǠ{���{�DD)�}�x���n��&O��K��*��Y*�u��m�r�Q(�{٠}�޽�X�I��d%��rS�y� ww^�M�x�lB�33��ݗl�-g�.F�J�L�H@]�}}|� U��j@;ݼq��ݮy��2m�nn-�67Kɢ7�i�e1m������Ҽi�<�ƒڽ�݀}}|� U��j@]�{��%qQ&I�iɠ�4o%4�f�����p�X4(�iM�]���� n��B�����������oR �J,m� U��{��
����� 5�f	�uH�#crh��Y�w{��@�]��xP�BI!!B"$��!(E|(UB�@� �h@�*{V�$d��0�gk��ǱfUd��j������ѻn���g�ۏ\s�ݺ�
ú���';5�
Bh���K��'h&3�;3��O&쎿ۈ6�|��*Yn�E�jj�g�N�C���6pح���C�s�M����2���SpV��c7p���t�� �!tg#:pk�K�B���x{I����Al9\X�"�l�W�:�=2e�0�e�b�y\�D,�ܗ���n�=p�v�h�W�#��ön3ӝ]F�I�.`��:�>K/oE���m������Q����wu�J"?H}&���[�I��d$�@��Jos<������׀�x�BJds�5���q�$R����Y���߹)�_�V,xމdj����� �v��R֮@>��*���2�,�����j@:����W���"���d#H�Ab����㺃�u�lu�#�z�C���Q�{�s��hQ���0�$������ֹ^�r�4�8�"�aXێ$�����&�HE�����|
�H�5����ٹ$���/ܔ�ٙ�g�;[M�0]R<��^n@=���d �v �� j��_,\�6���(�z�l�/ܔ�8��C��>N���;��Ԓ#	�2�M���Ԁu����r r��r��Z;�ASj�Aj�U�W7h�㷐�rYC������	�6X"��g��\K!�̘ڐ�
�޽��@9m��-t�Ď���,xނ#P ��@�^�{����� �W z��v��i1�i���٠[�M+3�<�""�"�@��@���T߯=�ܓ��{4�e�
	��L2I&����۬�	}N__��
"e�u�#o���5kq�@ⶽ�g���z{����M�}@K��,df��0�����i���y&n�{0�b;]yq1����M&ǂ�G�iǠz��f�r��>{R֮@>�<_aV���i�ov�v r� ��HZ� �����3;Ω�$)��d$�@��t�:������W`�bQM^�j&<QHh{���נz��f�r�6M(��A� JA�TR��~Jj:�y�>�J�K����w __; 9]�|���\�{������&�PM�1�E2!��e�a��汱�v7����.* z��oέ�a)I3wx���?=�`-��P���W�@>��Ġ�OI&���ftDD�绫 �\�� ���Mׂ�?#�$�6ㆁ�mz���h-�@��S@>�Q�x�%T�24�܀}}|� �v�ڐ�r�Y��X�M8y�ɠ����Me�X���x��bR�p��$Dt*�5�K��d� �o�W� � �@�6>�C(9\�0%��!�T��"C� ��!����s����5����x|
 �8�L����s��O�e�'\���0$�bDO�6������@@vj��#X�߻��~ �Wl���|��pN<@"`8�O߶!��Ek�kZ֤Ռ�j��c�Gk ��v۵*u�n���&�@٭����#�.4nIΫ�����bN�n��@�3���[V�g�I����X8[[n��q"����4��,e� s�c��Q�u��L��`�L��$���q:����m��n�uZk�΋nz�6�t��%��5�me��@kX���G�Vf:�Y�Վ����Q�U��ඪ��x��-9��<�a]�!֙�[$�- F�iw^���X�l��m���E�Y�vZ2�N65z��C�,�mJ�)1�gD��Ev�s��܋�v=n[���P�gu.�D�rt�l��:�M���m;<�=���[eF���r	�OX��Ku�L����ΖT'�tr��E!ɳ���y��%�A�F��
� =>3�A�T�޹���X�]tS�9��
��{mW^��K��<��ϯR�͔���WA������c&�	��e�PV�R��tL��fy�2���`���Y�CAm!l��В�0v �lZ7�p6ڥK&�ũUYn�T��+��7(�o�?? 2�.P�sQ��eej�c�)l책�}���-��ZY+E���GFݶ��mۜ��Q�Ɛ�7�n�h
�͵�i�7;l���9I�j*,V^)6qXu��YI r,����F�.�:'�*��B7W���3����64;`�ukv*�[�s6�S"���=�[S�k R��v���z� �f��)!F���-�n�m� ��B��d+���b��W��ɬ�WW6��M&� �j�i-r�T��71��؃��}m�hQ���(�_N�&�ubtk)pY.K�9�7<<9�bM�ڳ���S���G�}m*���["]j��A�Tѧ[r���pt��&�^���V{S�ܲ���m^�V�֒x�z���@��fz��%�m{����0�xv����r�B�� q\l5M���mԮM/*�*���p��̯@ P[үh@��6ն��3Y�LQҟ��������
�U ��	�P:)�qBPWk�?&�����M�/�'�~���us8�vb���
ո�nc�]nm2b�Em��j�N�^��ֶ�ܲZ�R2 �li�7kv��ɮ��%�.wY�N���X6�
lG;d�PCzWuf�S�ڷ=s��Bf:ɲ\th�vŸ����J�K�ݭ`��˦�[N_l�M���
c9�k�2t뵐5���/W!����l��Զ�v^��8/�Z�h+ڧ���f��d��"ƦF`s7���!��G����Ԡ-�b�g�`�3ctE����Q9��p�%�j8��	)��d$��[��@ⶽ���4�٠|�a�n!�c�/t�u��������>{R��V��F�AI�����l�=���8��@��b�X�8mYw�����j@:�������J^%�x�I4o%4�r������'��V�^e���l�s��򝶸���yB;7aJ���qu���L�s0MG�P"M6ㆁ�mz����W`=� <�_e�v��2:���f䜿_����p��"�B����q� ��ґ�Q����&�ߵ�'߻�M���y���#��ŝli�ȤNM ���������W,�;�wY�$�<�5�rOC���<��n��8���ӳ��9D(���, ݓ�.St�&<QHh+k�=\\�@�-��=���9rԶ<��m3���F�9��-�4�kk�����s���"��\e�<��$z���h廚���~y��.��@���.�; R'	�JI �YP�Ԁz�������FX�Ŏq��=���>Vק�HQ�Y{.s� wb�6X6�Z�ƦA1�4����.Y�s��h�Jh*�ǂ
�di�����~���W*�ڐZ� ��g���nbg�l������qvK�V��W��jNuA����.Fފ�݀w,��j@=j����`�e�$�<�5�nf��䦁����`�* {�%^�m�n�U��Z� ����rʀ|��ۜ+<oA�RG�z��f��w�7$�~�f���,i�5�;�=�g�\e�)��%$�9�w4�Ԁz����� %�u��ʼO��&��7Ńp\�ס�S g�7/KPs�q�2D(7�9&h�Jh�r }�; �YP�����jdq�@�[^��<�ă�^���s@��S@9V.<�+"̍4���k�u�Xt(����oWt��υ�b��Ӈ�894r����M��Z���h�2�S��<ڀ<��-�>��vܲ��<�	��Q"�� k�� ?S��sa�����c��p���@�ӹͮӧ�������.��7���ڧº����t*X�=q۷s[�Cgq�)7�.%�+Gar��l�7���ݰD*6��ˤ�yNL�,���	��Kq���N�e�=�j���-��3��7.�g.69������z���X��[��&���rkg���@�癥pV�l���*�v�:ZWs_��㝏��|p��ŷ3����{T�7R�׫Ya�q"CŜr�{~�i��psvx��\Kֹ���{�OӀ~ڝu�n�� ?=w�~kGD�����Z>g+��f$[��hݽ��ڷ�y�G�f!w���{Eٻ���� >y��[�w����]fX��c�G$� ����M��Q��9D%-�~X��	�^F�7$�/�@��r���� ���������Lx�������6 5vx�\`��C����z�f^�_S����s��247���z9n�{yf��v��g��1eli�ȤNM��,i(�Q�P}z� �Z� ��:� �Y�`���n`׉������Zw���z�{��ܭpyq6�j�����܀yŸ{rܲ�זh��X��ق#P!�@����$�o����>��M��W�Cv�o�벌�	5�r:��6�X��tP��e�˴�ڱ������ � �* |�8� �������Ux���}fv!F���3@>���>qn���� �Ap/6�ne��&��v����4XfL3�3�|�)!D�L/�K���ŀ{� >s�/f	Ydhn-���4[w4��4?y��w�@��\b�ؓ��Iy� �e@�v�:�����wn7�����h��Rl1ե�<�9�94�[p\icթݖ�\��v�]���K��nf�{yf��v����;�{����Ty�m��Bc��@��V�3<J���}x}ذ��x�tJ��`��G"�=\\�@�-��o,�>�ՠ{�:������b�h����]�:np9DDBbpRH \ �By.DSC?�B}��/�4��Ѭ}�F�,p䙠�v��__; �YPݩy��w7mg*V���\�7;��^y���k=<��&	��h8��m�ÞZ����[�}}|��e@�� ��̣�VE��@�U�4r����^��v���$|�໌Y�Ɯ<�D����T�s�8� ���`��bH��&�3�����^��v���]�t%�K}ߖ�u"���ɏ�M��Zs���^�@���������	BJ>��L��Wjh&�'���]H�uI�c������[�c0h
��d�ݤ\YX������X��^�Rmτ����q�0g�k���Q�v�j����U��.ۊ.��.B�Ge �(�]u��z&��\�k�����L�miS&�Axg������`�IΗ:ygS�W:Ӳ���(+��]JP8T'��^�`�m���kF�\S�/9�,9]I�VRj�欹1�۶�l.-I��T
�۱�8�\�Ŷz��-�S�9<�bDƠB9����s��h�]�"I~�ޮ��>Z�URu�]�Y�e���;�T ��`qn���4|�\t�I&h��hqn }�; �e@:�\Ϳ�{[w�����s��q��9�T }�h�*0U��#Cqh��+* >�`��j�z��݅p��Q�\��w[7��������ڀH���ܗ6�;u��q"6�2W�m��.�8�����(��rh�̳Dǉ;��fhܒw�{��|/�|��M�9���[x�Т"&O���+������E$�/_z��U�-��o,�=�J��dĉ�@�n- ��w�k׋ �x	K�}8���*����Yq3sw�k׋ �P�B������h��4�pU�<y��")42cs�d�]��,d���ۨ9�Kك�B�7`g�!X�
	�8�L�yf��<��}O� >��>ŀl�wQR��D�x��@�|�@=�Y�r��h��@>�Q�0U��#C�h���$��wf�'��uF)���ӧF�"��-C��X��CJ��;޿DHG�RȌJ��X��N'�1�h��~N+Cd �����ѱX 0#6S Fp�6����3�F��f���a�@淵���p��z/���,0��@�~��S�!_ڄCfဆ��1�0T�Na�$_�	A���*�؂8)_���	�(+�������b~H	�Cz �(@��@�?�t����krN�=�=�pW��4��5&��˹��]k�BID���׀s��fK���j�ۙ� ��s�� �m�/.�}�.e�Q�L2cK#�c#r����|�y�w8ጱ��a�(��Ȫ"��E$�9_*�=V�4^]������hw:u��ق&5���n�9�T ^v�sp�����a�D�<J)4^]� ��h��h��4��%�࠘cɄ�v��w�k�sߤ����J?D(" @�@H�� �����./����������<j(�O�h�7 >[v�2�����v�1�gn.踴�n�^�����Z`�sي��u���/N�u�8S�4��f�������^, o]����p����ŝli�9#rh���ԃ����Z����D	$LG��Py�9��>��`�*�YʪƛQ�Ǌ)&�|����W��h.��h���o,�=�J������4�͸�۰y� ��s�v�I�C���MK�;u0��̊%Y�Q5�Z�vB��`�4��G�]L*��r�֝;]�@.];kp�e�K��7&gZq��i��Y.�I=uC�D�NY8�]O�g�|#��WFڨ���+�%�!Z��gn[�� ��r�&��ڭ�E��)�y�Q����>�� ,aK�m����1��$5����z.^�L�Wi�qN�d�˴�©H�������q�>�N�������C'9��b�
sX�rݤ�rn��.* z���94Hb�8O�N����������Q���� ��6J�S73@�Z7wv��s��-� �S�<���H��w����QF�x��@���@�݀>�T ^v z�h]��ۛ�Um�nn@�݀>�T ^vWܯ@���,U��cr5&�~�* /; o�� �m�w�?^��m����S�g�`��gn�(�3v�#mE�vm��"�k������^7Kw�m�?�7�r��; }̨�g6�e�M�eܔ��������b!BMD]����<ʀ��>i3�E�Yz{{� ���>�T ^v ?r���"�&�H���QI�_�w0�w��w���x���R��Q&�a$�= �of�_�f�{j�@�r�h�^����x�(G�Γ]��r�k�6�g��Փ�t�� �gÉ��rݶ����Ģ�4�I'��{4�U��.�� ��q��*�dL�M��`s*�W ��U����\GU��V�y�Hܚ�.�����]x��,c�Ԫ�?Σ�=�女���M�Yb0X�<h�##r�}UVZ� .�Wv �2�b�xQ��D$C�G�_����ξ��zm��궽�&Rdf9�q�c�n�w�q��Z[�h�7[6�d3��v�������I��NM�l��� ��� �v �v�ayV��n�՗�� {�P�\��`[d�9�Ն;�D�cɄ�L�
��˰�]��ʀ}h.an(8&�)$���@�[d�/9tܛp���R��!Z��� �����'�>�����U$Sww�~����B������������D-�A<RO5U5r�k�7[gu���k����2��exvZ��s��mb1�Oy�B9=��s@9�Y��f��-�@�t2�<h�"f� ��`���+���?�RGع^mDBD<QI4��f���a�L�}� ����?4�j���Ij�����9$�D*wu`�b�*�� �[4�����`��Ņ���e@W ��V�@>0H�O�B+
Y�Kӱ�pa��p�[��b]X�m�{r��=\m��R*��8�{�gl�#�cd��^�-)8+�p��v�K� ۅ�d�-�]�{���M��|Ok��˲\��"K�a�G�R��=k�w3�I�h�6��O�ٝ�]��w]l�2���ݣ�8Lu��[)~>���G�\<.:c�TTV�^G`x����4MY��o�(R(�{�����kY_$>��Z7���1���j��T��6�r�SA�.#�=����U߽�N�Հ�� j[u���`Jz��bp�A�4�H���f�Qm��.�U���W�T�D���b� {�P�� �v ��GB�:UUd\�uw��DD�� ڹ .��8�6i���F�h^m@W ��b� {����:�1�X�q�� �1�"��3���'C������ۛ��}���v�q�<t��!"
8� �~�E�h���Vנ{r���f���(��S��B ���0*4 ��*(q��~ŀ}>�� �� kh҆�r%#p��I4�.�U����h٠s>u����a$�����; lW`�� m[��	�
G��Y�T[f��׋ r۬�
B��3B�:�]����!A�un�e�U�qc��i��f^�_4�����������h�� m\���g5�P�ff����݀>�T �v >�`e�h��i�XL�	��[f�?��B�Ny$�D�I}׀v�ŀ{�5��M��Bc��@/ܳ@���e@W`)N��h�k7(����X��s* r� u��3��<�	eh:L���I���5�ǫs�j��`Ÿ#�D�QxYe��h6�l��9M ���
I����r�4��4"�4g�<Y`(7�<�I$� �v~ }��:�v ��R�~�B���⃂i�RM �r����=�*�w4�٠^i
�<%M���6� {� kn�'b"`1 � `$X |A�B��33�}�}�h )�Cïp�(G&��^, ������6F��P�A�������=���n�.�hd/;�mNGN��Ft6�jwe�.`���ݴG#���5k�����w�l����7ش���:F�x�6����z�Q��h����l�=�������r���݀u���e@W`��@�q��,Q�L@���.� �v >]�u����ʺt.�&I3@9m�W�g�q�$���nI�
*����*����������U�QTU��EQW��EQW��U@_��EBBBEAX*��U�TU���EQW�QTU�EQW�(�*�¢���B����
*���*�Ң���⊢��EQW���e5�5�P24m� �s2}p=�@      

� k(  A@�   T����RT(�E�
J�$Q  QJ��(R�*(J�(��R�	)AJU@
 ���      �     ��{�_sw�S�{���wR���zU��Δ�|�\Y֝�������4�гk�ru� ����{��� >���.[�5�n���wo-y�����Ҿ�w�u���O'�ٹ{��  P@*� � ﾕq��c����F���.�]Wp ��:����8����F��g�/x k��ڍ���^���� 3w���k�x������y��כ}j��u��&��yޜ����)������������y�ɧ���@  P   #B��|�s���<�}zye\���/}� <��O].,������si^��>@���ݻ�W�}��� �ɧ-Ž��� n�j��U�Ӗ��t����|�z �\v���|�sɪ���  }�@�   V�ޟJ����޷W�J^�r���2�,@ni�)e�LM(P{��JP9�� �B��)F&�i��Ҁ )K1M�����v\��Ѧ��Δ(7Y�(�R�0 tΊR��蠣J)K�Δ���M)� ����%AB�(�� �R����M(��,}������AA]��NN�o[��w������+� �=��W�޶���� �����|��/t���K�)��e{�s�ɯ6�/�{�Ox �)�g�g������W��yҼ ODRy�J�L��S�*U  D��R��`h�D�*��j*��db41�BT�ԩJ� h ����$D 4x�?�����������ĝ��{����* *����PU�"*��PU�e@W�
 *�NOi	��H^��&�EJЭ��2(ZS2�YHkQ��m�Y�c�g��,)�� �$YaP�	
ID �,a�2�Z��ͿK��Ɗo�K	bsx�	L�?}�s<y�r��O�,a�8��.B�"�%XQ�l&tX2R�d�1�]d�s���0��Ӥ�#�a!O���(`�R����2�XL9!)�*�2��22ᒸsY�s�u��,~Ӌ��F5$	�aB4
H�)`��
�dj* @����f�!��Jk
B%�1�!�d#s�-�\�(B�n2B@�!�R1�H4$��h�,XGԖ���$9��q0g����g�7w�k4%#Ijb�2`1�����g��c�PH��X8�;W�uv��T��2p%3��zޝ����F�����q�!�!�R�(@��Ƅ�v��WG�P!X�R ��!,��6��jӃ�BSX0���)��F�$�H,��� �ԃ	�#��0�L�j`Ȅ
�rl��P��Єi�3��*10��0�@��#~�u��	 0�+0���D�H$`�@2�b(@������J0���X��@h���d��Ib�4A�A�F��#\!+��%p#T2��\�$�8b�XE  ��D���!L	`q"B	AF����h���@�a��fB0(�8R�	&:��f�R����F0J�b��$S)@ѳLr\ÇC�>�����d ���\3�t�0�q������f%��"50�$X\d�1��(&e�Ļ�ۂB3(��@[�*��.	I��Vc,�8�jC
LP�ZB�;�ɨE��W[�ш�q2H,#B0����Dp�?�r&	!aTJ���4�V5CE%"Q$D4E$G@H�A��	Fx��$��XF,�dD�$�"ŊA!4cR5�!P�#H�H�!@�RGv��0����.�AC,��,�D�&!
U��1���)��$Z`�AÃ[�nXev� I�ԁpK��I0a���:l���I8B�	��`�2������&�R9���#�~����ce%�.�0J`�ź38ozɴ�1�\H6)Zp%0%�.ZW40��)��c�֋4r�7�oE7r�2cD�!��q�,�24�ɔ��FK�%�a3�\���s�h�&$H�p�@�$�`�Q"Q(�Bq~�R�x���Mԉ&X`�ir����c�,)�&�\gL���&�p���e� ��	����!!XY T� 6o{�a��}�a��2Ja��e��BSk���B��X�
c	.5����FL2�|��1�3�"E�"FA�\e��g�q`��M�Y����"H��H% PJ�%��y��F#!pFE� D��c>0�t�ۂ<,g3�Z&u��D��N�����n1�Sa�Ѣ��>�qed����|�b�V,��X�\C��YL�I�ư�F�c07O��_~|���n	9����3D��HB,+����&!�����c�.��6HGp��L�JK5
@,�lh��&w�C,�O�64`GH�B�E� �c��U����
B�F
@�[�ovE��S�"H�q%2mH>X�:gk2��Y`��a4H'�
$
0��u�ǖ��@�B4�R�$d @ FD��~>��Nh��m�sc���-�$ɭ�!B��Dj����r�r�{e0L�.�k0���#��CR-(JV!J�
@�t"���R(�HV�%�ϭ~�T ą�BH��Ja�
��&~ZֱR ��3.6��=�w�ДÞ2�N��Q%��00 ��i)�$��Bw��V<AXXk		3�2&)HbR2ST��*�B˱�A��Z�bň�xL��%�R-���f�������X8�Ɛ
|�bC�q��Bs>�l����b8`2 ��G
Ĉ��� ��M�3�T��!�К���+BM%���*Yx�w�?��cL3�2�������$�ږ���
��$��bF%%�X��5aH!	�!���H���VH�dbA���I ��)�5���24#H��2j��
`��I1F�`:t��� �萴/%1#��ga!K�zB⹸�$әXH�P���D��M�
��s��C�5��"p ܌�q���o4�e8SP�H�!o�1���2e�)��	Ą��! F���!���
a�A�������2��f�11J�$ 
�*�p�S�qD�i1�����"ar�'���#$�D �H,�̲��S3�|ى�z%(�CB� ��
2��w8��6K&"�X40�l��hd#LB���1������qa��p�+��C �#�~ѓ���0]>�20x`�5���;)�4c\>	!M�����F5�YHX���L�����S(�?��v���T�..�Q1�5 X�H � �!��Ap��.�5��Ire��3ht���V��_�JX�NLP�$�h@l+�u�R-L<z�F�ɣg��v��ddnM�+�xa�$�&$(����	*��~V������YlI���42I)��L��c����)��p�ˀ�F)"0 e�BL~//k�3���D
a1�1N�LI��0*S8�1��pXm0S1����J/��8du���	�>�;�I�. ������]�!7bXr�dK��l���Y�2����,d,�y�w9��c��:.���'>���l�0�9���7�hC
Q�l$"@�`�B�2p]
`�8���$�H[#rZ�,L+��g\3I�m� R��X�JG.�����.4K�6q��G;"}���
�˨� ^f]>s�J�U�O�R���	�P0���ɔ����##!bE0�
��5�!P�#�$3�W��f���|��iX5jGxv�j��+	�$1���U�p�c�, "�,"�E�"�h�"`q�� �b1A�q`X0aL�� �~�Y>0?q1��+�R�0a F���6%$�"T"�!�b�:B@�g�+�e�i�.��L}эV4�
�5���ϱ��t�n�XR,ay��@k�c���޹mq�o�%ƦϷ�3�ĺ��h�A��GI�c����(�P�і�D�a�%
�ys��~���M组���B��R�\�@��4ČJ��)��VC.R)$HQ�� FtLk��g|����hB�"SXe��e��q��"�plɒ`���Hd�d�Ʌ��3�=�	B��l�˧0e!H��£�n�\:,ѳp���pƸX��F�)�:�Yݦ�BS��*JƑ�jb�o��p��2dы1m�
�u-v��
s�R>!��֑����}�\0�@#
���ƙpB�D˫x�/�jG;9��.s�^R)	!��i ��T	��#�f2R;�d⟶l�H�萡�b2@�N���FnJ����&�����iņN�F��- 00 � � B*t:H1j���cC
bH$r�hE"������BI[X�l�������H�X� R��+��`c2����0ˍϱ2t�d"A ��]4��"э`ф-B�1�$`�CH�I"_���js!�~�>Y�c��p��\��j@ W�Ra$R1i�dH��� �BF0�%`F���)�xm�đ(`�L���z9���r        �À  -��|  � m�   @�`��nju��&�4^ I��   �    �� $mmR��HUҒʆ�8}>��e�m n�Ւ΀� Um[G�&�`�M͸�KӈM%�n�0֤.�m%Ε4+U!5u���� m����XÖVV�	���,�� ���r�5������G �� %Y~>��U�jG�m�`+<�F����M��b�	
 ۶�u���!fٕg�j�z��hc6�  66� l H�Ce�j��q�n�ηm��e��h��$HƎ ���f8h BV���5�r����h��Dr� m��I��l8'�Z�5IN�kM��;mۥ�K-)j�� ���nٵ��ȕ�����`)���\  �e����a��n��޺M˒�m�    u���ͬ�����C�)���s��K [@  p���` e�h[E�*�j�$(�Mr���U��"��K9j��hz�vȠ[Ki:8�m  H r�ݖ��m�44�wT�˶�[@[;M���́�j��  �� [vݜzK�l  �a���e��m  ?�m� �$�]%a79����QEPMU���`[I,���` 8�-�@  pݰ�� .ĵtV�ڗ�3@,M�:ImF�-�� �m�:�[@p-�m��      l �֊h   tQ%�6ܵ��­<�WV���5���T�����lV�]��9��:H�5� ]�۲�am86�	өqNv�M��F�۱�-�k�pI�l��AKUPU+ʀ��E�d8/M��-kx� p6���ܓ�f�:�izYv��\�m��^� p -�����6��*�m+]m��i��h�F�LR��a�ܐ 6���i�j�	 �%��m-�d��	e㭼m[ H�`�t����mp�Rq;U���ة�$��c�lI�N��;V�Q�n�v�"�KHMU\^m�t�`rԄ�R��gs�mq��L
�u��;n�j�j���Km����v˴Y�O�D��9_n��	If��H9-�U��8Jvez�$���6�&}@�$��i��b��2F�]���"An���̪�P'�qU^�P����`ym�I�*gY�6�v�[��@���  ��x-�9v�jٶܷ�Gc�~�K��	o���V˵J�HSu
���i�EKX�,[>�į��0��p�WU�t�M�d[x:NH�$[m�Zm�)^kl�8m�>[L�@�+�TF��hm��S` %��  m� $��v�H� �y5m���[@ �okp6�  -���lI;`�޻O����ᵴ 6�i$�]5�j ��z�p�uY��6�j�U���n���8�H�^��
�K%�-ɷ� $ m����ϧ�4��b�j�TV�<*��� %kR�*�l�$[�Bjڨ�[�m�VU��^����l�	  ��97F��k��eZ�u��m�[szܺ����l�lT�-t�rVt1�n�M�m���[M� � ���д� ��`m��kM��OG  o6� ��H ��lj@ֶ�v�m[u^� [@-2�X�{Z�J�  H�6	�8���v�:l[B@��5�浲�l�@ ,-�[zN���d �Y��m��      m�����Hm�h�z���e/Z(^�[h�ƭ! e�$<��˧^��d�'bƺ� ���h�u��xh^-��'nJ�i�G�i1ѭ�/a�������g��!mc��hL�ܽyj�Nu�� H-��U*�[2B���w��t��� �l  �hhr@IU@X�*ÙXw]�n�:�m[m -�$[@����B�j�M� \  m� 	-��6�H��l���oQ��F��v�f`$8��KָK%�+n�G;*��J�8�v���!
� -�M�.��m�زL��g3����N��:l��l�M�]�8  �{[l�n 
�6��$� �`�R�&���$��y�P�iV�U�
����5U[*�ekOA;�K;9�B0���iJ�v��u�s�&V�vxع"۶�l  �Epz� l��֚��`�c����C��H 8[Z
���i�٤�m����^�iyjU�@5�m ݲ�m�����[M��ڏ�l�:HI�ɶ�ݰ-���pkZ@�	-��-�im�8e皫�l�p�IeBK�H�l5�$��&5[l��C�ۢ�]*�K*dΛc7�m�-����-�   8 � t��p���mz.�t��  ��l k����`�j�-��  �I�	l 	-���� 
�c<Vv��;�^h/�R��U\��#[;`mfsm���6�ŵ<�f�R+�����UMk�,��I�p[�s��e(q,�   ���];mkk��&y.P,�Q�W��G[��`8m&�$ H�B���� l -�m �` $ h  l�i��۶� 6�8lkXֻJ���2u\	ְ�J�� ����-�   � �T͵�m��6� � �5�m,��l�٤���s��R盵�V��X�%�mS�˦�t� t� "��[-]��f ����j�U^y�Jm��,�'m�Z8�!Լ�ev�E{eZBh0����Y@j�Z�%K)� -�*�'U�+p���\aڪ�� @m m��2I���!�8���f����S��;�5����3H5�Yv[�[ߣ]6��8v��u�[@�`ۮ�ڒm\첧5*��@\׮������Z�k[��  �����l�	�\8ۥ��hm�I�\ ���vq��m��t��n�h�^�\�`n�v�Z�����Ѣ8
/��%�e��NIBA .�iu���L �CvA檝6p�� �lm�Ԃ�(�ڛnll�#j���n�nb@� �� �հu�T*��WP����L����K�:� �z��mv� iUUT�)T��.7�uR���kj[+�	:Y%-n�9�����Yx$-�8�  ��.�aF���
��<�6�[u�  l�t��	l	�:P�۶��I3�T�h�ۤ�,����5�Yv ��$� ��皪]�
�� ���J�LU�:����[�J	�]nh��^Iյ�qm[@��[j�P��` h��xe��1ș��UU�S�c�#UkST��m�� 6�	   Nڶ�m�[Cm�[@d]'N�p�Y�u�l	 �55n�ʲ��jk��`��      l�m�[v�iV���m��k�]uΝ&ZI5 H������}�����t�p$m�8�ޤ�-�[�km�m�G-����l �fݰ� A�e��\���x`UW���m�v� ���,I�m� �,�Mk f%S�UUJъ����L[@��ޫOXj� s�6I%�u���T�ĵ *�5Ɍ���a�s{Z�"BG�i ���u+���	�
�i\r@�}z��o��m-�m���Ãkn��m� �i�	n�	�ʖ�e�kq 
Hmi��6�  mr�m�~>�� ,�hm��^� ����m�m6�V�WY�g2�@T,3ԩ�jZlհ �@�lۤ��� 	l�@  m�;tP�fΒ_FT�S@�o�� m���(!ri.�K�Ā>_��-�������kR`�2�h�   � ��F�.9I�ms�:l�l�RԪuU*�F 
W� ���mۜ����j�$!oP 8�6��`�7I.�f�Nͻk"m�D�"ŋ���0  �p U�K:�am���`m��	$HڥYgf� �$$-� qŴl�mH�ic$�ܬm�v�8�Z�"BM�-���e��`p-��  m�m��gYN����+���Um]�C$$nm�ݰ���� �Y�a#�&�y�Ā
Z��J�K�Uv�V�R�9+3m��f��۹*@Cm��K3a&ݰu���:��ܒ�e*��n�=Tl(�F�P^��t�t� m�]*ҭt UJ�Q�)�tJ�mmu],m[D���M�  9���n���
kp  �(P�����ks�[���l۰8�md�5��u,��L�l��	�6��d�'2/i����^&�n�`b��E�0H-̻p�I��� 8/G����m8H��u ��v��K�m�m��p:C $��K>���� -�\�V�9^YZC�m�UV��6�lm��pm�n?����)�b&�@؉��A���iP)� B h�2 M����t"�T�:3��� 1�WJ&	��"
�Z*�@�Р8�4��튧8 :O�AT��~N�� hW q@�ED���D �9�	 RP"9)�P�!���  ��KUBA i ��S������P;�t>�1�Qz���mT6*�8�Q��ñTx�@��W�@��ڢ9Qȣ)��"�`;E���']�A� ch������p<Ut�Ep��^g�:�	����UMV�=D��a�.jS��D���*�x�!����L��P��$ T�J�8~�`@Ȏ�j@���hT��;�XU�a�����t&x/ 2 G#�"�(N��\5b�Uj+N��~: ��h�dP�R�T�|��A*�Tخ�=v���: �(F!He`E��H���� �$D
p
O�# ���	פ���� ��X���*�P8�.�X�`� 詥�����ʄ�B�х$����(Ֆ!"Ђ��� ��  ˥v��XX�H)$"��U+��vs=AL���D # @4*め4UTp��T*"e@6�AM(��Qj)�遴�u@W��,("��EH�Ȱ㻿��UTjnU�j���1�9�Z�U�p�ye'7�[ .1v�@i�^J��q�x�����.�zm���ʨ
���Z��+i���&�ܴ<��6v�� 
��8��U����q�q/]Z�W�Ȧ��$�a6ڝ'1�;b�@6gi�(���#*Ba�Y(.6��;�JCfFFZ�e��3�8qW:!�ݍ!�몵.��6Q�M��÷0�tm�d	c(�AAӛ'�g�va6.gGnŹ�X�xX�hM-ڈ�k^��L(@:�ַLX/^�IT�a�	[$�r�N��s� �1u���m�6�q�I�˖�$�^��z���P"r8����.{V<-�R�!��ݫ��m�fx��rq�{/M!f�mm��ftYPZ���1�)6œ4�`�;-UT��:y[^��%�
��)�[W\���E����-�;w;.�Y&��:Cnj 1��pL�:Y�q��ɕ���BCn���T
��:q�!ۆ��L��9�f$��@9���Fp���n��p�M�d6X�n���궞�i�U�P���Vs[��\ۮ@!u�c���5m�
݆��f�U�UT�T��y�Nâ�k=��)�7th�U[�:������څŰĩ�R���Kh�sZ�	�[{e�x�Y����� �۲���狀nr.i(�[iٱ0F��4�ڶ{t�v��p:5��ݹWLg��4���6�S�r�Is�$d��|���DN����cn��HԤ��t���mW�E@�ZV8�YEP
� ��εZ��-���청����ڸ᱑�S��l=rg�<=���ݲ	%,kl��l�]�N��,���Qr�Y���3ͦ����h���U��P�{8��U��
uY�
3q�VXyRP��
#�l�p$���YvZ<��:�5plK�I�ں��pGjk��s�btUv���A�Y.�BOjV�s����m�Vkp�t^aI��A��"�m-U�+�Sbb�8�q�eS��!�?*y�Αt�*�z�� �G;�
mV
w�B� 
����S*1R�P�yfi�\Yq��1
��:%�9��t�����^h��	�-]�Wkc`���:��m�u�����d�m�4��7��ݴȉ[,����C\q��j[dz�W��飣��R���np��u8����dt&�ޮ;	����]/mǭ.��n8��p\��Smճ�+;5�a�93;\�^�t�7I�.�gg�7b X�w������2�*;ě��c�&%������/��ɔEL;�8�wnP�v�ll��/�U�ϷZ�mi`�����������ym�7�
L�9]�$�٠w�S@�s@-��A85�ª�P�v��v�6� 1�r����15r#x��rh��9m��9]�C��h��D�5 ;���P��M� �n��؀��sD�|�Sn)nˊ�ՀS�P�y�e\H�e�MկV�n ��k���[k�\��䚸����ݠ7]����,�\�jH(�ԋ@;�f�����E��"_���*=DNro������9]�@��
(<Qc��E]]�7]���u�P��@s���F���m���������wJ��:#�:�}ޙ��&�&ۉ&���~�h�;۹�r�M��`�H؟�c�|I>�0��M�N�ڭ�κ�81p�uY�ƻ1��0q6��,���n-��s@�{w4[)�~�h:|��	���x�&h�Z�6� >�nP��]27ܽq7".B�wk ����>��^����DC�P��{��ԓ��{5$��.�\dx�L�!Hh��h�ye4[w4�,�\�jH(�����j�؀�ڄ:�(
�$�ۄPh�"X��lJ�,�ƼQ=vd*:�KQvd���	d��$J���n*f�>�_m�@c�r��mB��b� ����l$����M�ϳ舙7����(@n;b�s6�.j-F�I4�$4Wڴ���=�gؕ留��ƀ[]p�,���n-q��l@c�b�ވ��DLF �P0�0*.﷯]I6^�7�	���x�&h��9_j�9_j�9��ŀn�L���5i�r�ڛV=�P4��VΞ�ŭcK��qT(X�	Y���\L�� 9#��;�|�Wڴ���f~A{��@�*a�dx�L�)$hu�Pcj�؀��t�����Ȇ���8�ܷs@�,����K���@���
v�(�ǒ575p������}Hu�Pcj��m%$i��;^��Z��6����6
�"=誓����������z����9{��f�ilwPu q��NΎ����'a�sΟj�g��4�ܚ�K���izD�B�G��>��I��V��j��γ�[���Zwg�n���+��s�NID���B�w�}��^2i�{f�����5�L��[,n۱k�����=Pk�2k���u[OT�v�7G�I��&(�=ttu� %�j���K�����������{�����o��ّ��լ�'"�x���-�ݛH۩��;��ϫB���q$ҎH���~廚ye4.v� ��'�%�$k�ۋ@��T/�2=��������ĶzjnH����C�4��h\�z+�Z�[��w�������8h{�z"'k_Rz�J�mBq��ο���	�E$�@�}�@��w4��h\�z��;����L�)�]#�]�dRV�+l��:aæX�N��ٻN��m6ǈY>��Q�q~���4��9��#���>�8�"n���3����&������/"U�Sh=L@O�-�}�I7�s�RM���ԇ;jŤAIG1�C@�j�9_j�?r������T�Yȣn	UM����z"'z�J7�Bq���Zm�O�1,r,�n-�-�@w���������"M��3��XN��n��Ϸ\��2Q�rtX�����r��ڍҞ�4�e�5�m�����Hu�Pcj��\M�o��4.v��G|�zx�;�)��T��#ǂfI#�>�9۩&���jo�G� F�Q�=���4�?+k����q��r
,nI@|ݱ��tܠ1�r�!���(Т��!8h��;]�@�v���h�v�6���ŉ8pp�����֩]�X�;^4��֤L	�o4n]qB �����	!�v�V�̮ՠv�M����IJ�'�F�I5]�!�r��������_tܠz���%�`�1���e4[)�v�V���hz|��"#k�9!�r۹�v�V���h,��}��`�: �Ш����ԓ��ߦ)�<Q�n8h�ՠ{ﾹg��}��@�s@���GqE�(�Ld<s����'N�f.-3XmYXz�u�+]�ۍ;F��3	�Px&a$Zs�ՠv�M��h�ՠ��"�q��r
/��h�S@岚k�hλV�e9��(Т��!8h�S@�v���j�;l�����ZD��sy��v�V���h�S@�s@��(R'�F�I5�hζ�ވ��r��7�� 5�r�u�,��� X 89��1.s�q�8�Yΐ� �k���[s�Խ;D�6.Y�Y�2�!��Օj�7�8ln��Y�3zi���HL�q\K�Z�w�/�>�5�nn1i�AĢ��L&��9�*޼�NY�ٮ��b�6�.cm�����r3�ia:�ŋb�qų����Gd.�3�L�\�b�.x�+�y��Z�������Z��=��h�-�j�^�9�d�/��T��r��K��ٜa�n��ܚn;�c�ѡE�=���F��NnA��\i�>'�|�X/�nE�=�Jh�S@�v���j�.u�|�k$Dmcx���7l@k����ܠ5�b���1LQ⍐q�@�v���j�;l���e4�������D�hλV��e4[)�v�V�~�!_�5#�Q|ۋ@���\|��C�r�#sbi�UT�Ep/5q��޻*��4�e��7Vh�C	s�����0��
4(��#M��w�S@�M�!�sޏ{�����%ZH�����	!�v�V���>Ϯ|�������%�(Dq�����{e4��h�%*ȞEq$�nE�s+�h�S@�l����Z��X�O��Ȱ_܋@�+�Zk�h�;V�qw��ƲDF�7���ڴ�j�;�v���hϾ�Ξ��Bck���e�6�3�.:���K���:�ѭݪ�Ǆ z��<Q�mH�|��w:�Zm��9]�@-�0���	�DI���nP�b7(:{��W��z"&C��/}�) ܂���Z������N �%N��j��h��
A�,B!e�f�I�(�b&�J���$$�td�� 3�pP���D`�.XU�HY �dI�! `�1�e"FE�e1���H9BP��#�0H2P���ۍglx�oD��U�e!*Q��S&��$Jp&0G}&1���	�;�cZg(5��&C)(���!\�a�D8t� @��őH�!&�	�abu�^�
�̋ɜ-M��+����#!�1s��8Z}�bB(�NP�؃�49��õ��Wh�S��Ð�B�8,�h�k���A��6ANU* ()�U@���=˩'Ǳ�]I!ӽ4(�m!8h{�ϕ����x��޼RK�T��{�7�i�l.F��R@�� �gz����.-�������������B<ġt��n6C�+��������.$t�:.ýv*�8߽�w��}��C�+ �����w�wJ[� 7]�������P��t�Ev��R]�����J�;ݽ0��-�]�}���]��Ѭ����QUwb���GL�uwJ�_W-y1LQ�Ń�8h{�}=�8{�ԓ��{5&PO�V�\��Qu-T��*UU�������Pm[.���gz��U*^�K����7}?���P7�L���D%���汉��θ�<WY��q�:n'v�gE��>�t�q�߽��q���I�_7"��?��w�S@�v�g��s��hx�
4(�MՈ�l]��G��(��Ҁ�����UJC��4�#n��@�f�}~��-��RUJ�}��X�ޘx��n+w$��v���ڥUT�շ����,����ԕU$����onh���+��`��x;���=^T�{����7��xWgz������ŗp�x)9wW`�inV��ơz��hF �+����>�d�``\�n%�y�M�a�箅�u��iNv)8��=mAtm)�l��2tғs�K�������dX����Y�6����0n�)��l=q��4�f���7L[my��#sss��r��a�Yvz�]�ip/N�u��=Ztԙu�M����O*ͩ�-I8f��j#`�z���{��������b���r:�z�t떼r�u�'�N��TqmY�of;xٻ/�?�?oIֺS��n�������nP2���} ��B�r���Q��HMH�v�V�#���-�{�@��o�ă��ƌ=�����D��[7^���a�������7��x��Y`��r4��9��~���������`kշ��i�գ�'mK�q�������=IUWv�_�jپZU���@�P#�|"1D�X��.;v���ڝRM&�nPoX3�@�ûZ���m%��H�|��\�h}�g��%��o���n�ո�ܒ��.n3��'O���El~���Pi�j�K?��� ���x;;מ�^J�%!���tU���+�o ��z`��^J�*��;�u��7^��n5e��E��`m*UT���xvn����^�$�>�ݘwoEi�r�HMH�v�V���>�z_/�U�y�vs� �$��]{�dq��wq\�%�ln���"ȸ��G�sn���Ӌ�ۈ?��R�yb1B�m����پx{ـs�o��J�aݛ� �*���m���9-�ӎ�忀��ٞUUI�����;�u�_�:�j�M��}Ѓ�;X㑤ӏ@���;]�K�/��}sb�@0*H��� V$S�WUmR��Zɼx�wf��:�ȭ�m%�p���f+��-��|��k��}�+�o���)�<�6�M�5w(�Z���C�\|޾ݳ �RK��M#ww �\j9c.�I�r���*�V�d�<�3q�vs���������K��j��.'�K��z�`���s����K�\�� ��:�ۍYj�Eݘ�ݾ��U�T�C}��uw�� �{)�����H�<d��6F�BrG�_�n��D���� w��1P��[n]���>ssm�'}��jI�s=���v�U���gJ4�J�@H��@x� imR�ǟ���;�6A�n�h����l@t{͵��>����ܠ=[�M����H&'���1�di�08�s�]�2j��4�uf��z����o�������,���#HN������e4r��3��/�<h��,בm%c�4w��?�RJ��*JC��������;��o}�}�fcg��)�<���M��� �6�������*�J���~0����r�l�tT���$�x�I>�����s����U�T�S��޷�yn�#����"��v�s�� ��%[�}�����vw� UU]��52	��<�Z�vu	��Z�R��ˮ,2��!l�Ok³�n.2��+9uڭ�gCY�E��^����(v���u�3x�8�pR[�m�'��7k���sQ:S���keF6,gj^W�X��<f�ۙV����+@����e��t���<;�$�6���ݮwS��۩���B)�]����A���]�Ywc7ks�o���U�(��,��q���#�8� G�7n7}�������j8۬�릻�x��]�g{Ok��ґ9z�wtϻ��h�$'$p�s��x�9�,Zk�{3? ���y�F�F	�RE�s��o?����<wo����f��ڣg�����$�h��Z{�M<�������ZXUܸ��1G#��v�=��������r�oR}��z���m%m8h�S@��]s���P�l@7Cv��WsI�^�d�8�s�kT��E9�f�6�]������Տ�t�}���*@�4~m������nP�l��A�wJ�}rzm �ƇA%��9�޼�W?U4��uD�E3\�2 CeA4��d���CJ!皛���ԓ�ǽt9e�}���L���Bdi�x��h�����w�wz�� �����)186HȒrGg�b����;�M��s��xJ��>��� n�Q�ڻ`��%$Z9e�@�g���}=��l�v�M�ƺ�ȜS�bJd�狍���uÊ�2����t�e�\LwG�v��y	?}�w�8�fBb$n��E���-����9��x;��䪒K��om�ѯ�T.Kwv�B�����^y/U$�7޿���s��y��f��4�#n�Kr���� ���}UI�>ʬ@�LQi��T?���~�u$�_���/jJU�&ۉ6��ϕѮ��Pmk�/�p��w��(c�`��h�ՠ{9e������;)�~�uw.57���7[��K���A�],��vƜ�,�7��k���ş�w��}65�%����NE�W|��)�w�e=�~A|��v�g����FFܑݼ����y%!�6�`��<�Nu��&�wb�F���[n]�xv��9�޼<����I͛�o�~0��"��J515�$4=����>�;�';��ԟ����O�iЇ�)Z��I!*�_��oLy�^P�,n]�!wo ���x�IW�U���/�z��Ɓ��Z:�kClmbqb��v�pu�+Z�r$ �j���뮡�0�[��8�}�`���H�6��F8�_����4�m�t��{��}!��J�L͝m�rH����~9}3UU*����x����9��mUUSf�w���ƛY�wf��>��^��&�����g� �ޟ;�o4�ZI*U�UJss|���� ����W�RS}���;���ӖH]��rGv�w�ŀyU*^���߼~}=�}�νI2�9mE�шg�aDē����q��#0ov����}	)�c��uR���d �I�&���$�$'F�Bm� h����)Є0d�XЗBSa���9}2�%�0ͤJ)Z�M)y��d�oȹ_�a1��qP3�k?m� [C��`�l���:�U]��x���kp�ՠ�]jXP6e��qq�2��.�Nvq�FkV��췳/4��h���6٠-mS�H�q��Wkl�tɽuJ����{K��ܽk�6c��D�ڝ��%����}'���� �DvS���jд�:���(�8CB5��Yj�jU��N�Ν�p���rܺ$ws�����`��y�g�Ǌ�p�g��������PS�v�ւ�Ŵl�4h�}��ɭ��-��T6{WR��֬��v�{$��^ԹG��\��tg�]p���ֺV�����;�X%_LvN_R��;1
x%���c�喹�\[�7د�s�GI�襹�*�l�X �Z��9gQ��U)b@j�,���+� �ia[6�[m�	u�e��vظ�]&��;��`�
�﯍�۾~M´�F��Wj\��p�5m5�Kn�Vfg6�F+��%Xw<�Gn��#kZ���:ɚ��#� �8�9��!��)�^)�<�Hꭎe
ϵ��
�dz�-U���AW�j�����S�.�6@
c���^=�Z���Y1��t��PPj�T�s���9�'d��9��K��m�֮���B��xr�l� d`�����;4�чnŵ�N�&�Q��qnj�؁�렞, �'+�@ (�q�sCZɊ�iQ��Ʀk��O.P��a�ggk�����SO+��\��n�[W�$�"7NH�\u�j�q�ط�b�R�pݪ������<�\���6��URIymX�
����U��MX��:x�p�MUv���\�M��烔�� �ꚪ�vӹ�nب�MA�J�NE3.�j�ʛF�[)�)5+Yy`*P���P펇��r�Ϊ����":,������c�����!j��#D��s��đ�ˮ��C1��]�b2l����kn7H�%b��� ����溃���)pަ��֜��J�dL"ҵW�H܉�%w���wws��Pz	�M@>4"q�� \E0
���C�\TW���	��U�L��?Mf���v��zu�ָR�p�0Gb2�gn��}i	�����U�U#$;\��ME�՝dt]�������O7k��Q�p��V�ǂ�-���k�ɍY�ۛj��<6�!;����+mms�n7<�,9:5��`Es�;�85��8tg������i&GnE�`�2í��M��>�'Nc�J�gN�� R��U
,�WY��7���~w�����~n�:���Onc=��k���i�V�Y��u�m�ی;F�����;}�v�v��u��@}��z">�}ܡ�Ƒ�?mF��$4�j��3>��!͛�o��X?���I��:�B7��"H�W|��w4�ى^�<h��Z��ZD��j1�N��T���,�;z`��^�*�w�@��J�<���M�����%ޒu�m���R]���6�;/G������������j���7\B���� ��g�(��� �t��5���ӆ�y߽�{���v��̬H��~I%}=���Is�QjI.�/R��RK����w�����*z�Wl�c0b�9�ݶ��g��)��G
"�B`�$Q��@j��Ԏ���3���ｳ{��v)�$�l�_�{>ϛi_L�1H�2!���������$�zIRԽ��۾�����s�ԒJ�֒��#̉&�}�oUN�����v���o�%�x��/U��}��ͷأg�<Gq� �����|��>m����k6���~_|�|���| ������s�Ù��#۱;.�݆�Xku"]��꡽d�{G�y-��}̍�'!#��I.�<��������$�8K�������o}{��ͷ��4�J51��ĵ$�oo����fcmZ�����v���o�.��z��+�o۾��B���j$�$���I{ß�Ԓ]��~���T>�HQW�>ϳ�[�m�����ͷ���B���bK6��IW�*�w���>���n��6������;����zo���������N�J9�k~��\o�D�W��>�[y��I{�ORIw�i��I\t�\�5�1����:�=��o,\u"�D-,lq[���ַ�	��{�����n���S�*P~ ������� ���?���|�s��*_�F���[��oz�6�=�&D�s7�I\o���fgʹ�����$�\�$�-����g�|�]x�+y��Q�GԒV�|~��W�T�/f}�������$��;��$�lw.27��rGv}�oj�M�f������/�c}X�;�j���X�A"5����!P K<dS��"~����OߒK���� ���S�pZ�K���}�m�W�RU噾��m��g��m��]���\I�E%���X%㳎8�$'�vzz�]AĎ�3�+�e}v��x߾�����L{�$m��j(�s�K؝�z�K��٭�oy��_(��b��{�7�m�鬁`)q4؅$�1��9���ު^T�R�����m����}�m�I�ɚ�RII �~����'Q�9y�ߟ������7������T��j��&6��w4���}��1H�2!������}�}�������Iݓm�Ο|�ڤ���G��������0L�&�~��WekRIbI*��x�o�/����������R�n)(`R�׼��/%�qm.�ť��S���Wn��!s�I�Z[��ę9��C�pg�� ��n)�\�k���8l�]"T�-��`�8�����p�s]�ca圝sD����b���E�*�}[�	�U��^�ͷJ[h.'dӃl��ˮ_>��[��@vy�*���+���Zs��9V��;�G��������C�ܴ�@n�a�,��`�q��c$2p�	��]�_�s�3��`~ގru�s���s�[�ۀ3]7�uF��v�۩��������9�������@������䒽r�RIr��?�9Ȓ�;<֤�����dn	9�R�$��Z�K�����I\}��I%�ݧ����U���iLKr�l| ?;�������RIw�i��I^�E�$�ږ��<���M�9��$����ԒV�|~��W�QjI.[g��%�����cPX��7.<m��w:}�m�R��>��6�����4���ZԒ_��L֮)#cdkq)�Z;�\��Okn��N�8\'Tu[َ�ݗ������X�9$?~I.�7I%m�����;+Z�J۴��$��~���,�1s�um���vo{�ⵤ�z�c8✾Ǎ���3��6�;��g�$�)#g���@���Nã+w������> i�}?���Z�L��ww���3.���j�$n�B��Ǎ�$��ߴ������1��{�������^�Y�6���3|E�n	7#mH~��]�n�J�g��%�vV�$��i��Iq�,R�M��.�<v�s��vY����ᒩ4���#y���zS�Q�q��ķ+�� ������ߒK��ũ$��OߒK���RIs�Xt�ܑ�r&K������m窩*�ݷ�{<}�m�x�m����/�m�ܝ&@17�A9����?~I.�7&��h� �E�J��V !�`�y�{�����y���7V�o;�_;�Lx���%��}��������}�m�����ҥ&����6�ݽ2b������RI[o���$��fv�ͷ�m���>�����#m���Wh߿s��lga��ru۷�s̎m��,���gGn4ru�F�u�rH��vY~��|�����}�s��6�9��yRK�~����w��������P�3��G�m��Ο}��R�>�o���w~_|�����^��Uwm�l�#���$����ͷ�����}�{��窕$��fޓRI{���$�U�đB��m�XcoR�U&����ͷ�m�x�o��t��n�C@`	"OEr
�$�����cm�wt
��H�*\���IqRjI+n����n�jH����>���~R)�PDNr|�qt�<^��e�+NC3q�l��k�ֶ]��{���G�,䱦�X���=�_����X{���U_0�7�xޮ��q��\�H���P��]�;{� ���kz�ʩ/*IH��+N�!l�����ذ3��᪒������w Z�41_�`�ۙ��ϾU�����Zon�yn�WN�6�	�#�B�������5$�w��/��n�ԓ���Ƥ�Edb���v��CV�]�y�b�v9�]����.�q�*�ڎY�N%j^�^t� <Z6B�\���*�N��+[r�Թg�k �4��]�p���HK�N��q�\1k!��R<��q��T:�1OJv����ݛ�n�h����|����䳍��~�x^6�\��{q���qI�2�,ؔ�r8�7)Qq�e�L��[�N��ⅺԩby��H'�zC����ّ�[�k�F�̉�3W,%��m@�ԕ$�&^��c�]څ�z��P�xڄ���D{�Hs�Ҁ�nax�#hQ���I�廛��Ďw����/�{f���wjT�l�{��y�j$��I�;��Z��Z}����X�w�q��E���4�W-�m$���x9�ŀw�{��^��:��x����Ʈ�r5"�Kx���DGow���]Ҁ{Z���s�.���c�Nvn=��箚0�/b�q���^�[n����\��Xw�6��E7(��z=����h��8�"s4��j۟�b�B��"�JX�? s�����R�����,�J�5���&�F�;d �[�7���߹�Xz�^��I��ش���@��v�}�&ܓZf���@dN7H;��z'���Ϫ�� ��F�rL�/-��=��g�������3P�n�i���L	�
N�9:N:E�Z�&t�\��$�]�2N�3��Nn�>�~����[|t=J�p�j�������(�j:#�菤;{�h��"���,A�h��h����;��ŀq��n�ޥT��7V���d���on-��ۚ廚,ߌù��Rw�f8����9��~��#�@Ћ�C�d�`3�� ePbD�$HA�1��Ʃ����)枭Y��;�.D2~�bk0�V�x�6�Ej��ā1�t&���@"n�pJ���H�\2�ä~O���LXҫ��L����� l~>�KWXf> �/Z�����a#�8�0��Q����j|u@����i~6Tr�}�TЁt)�p)ׄ��=¸z �*lP\"&j�j� �9C�t�Z�U)�}�.�rw^ }���v���p�Z��T�=��� ����޻V��v�h����<Ȇ��g�@w��~����@���������·X��w]R�L�6ؓ\�N��4�U��z?�wr�����Gq� �����=�s�;� �;�^���/�5�޻�:׍�\�'$�������@l�wh�ܮ��2Uڱx�#hQȓrI�����ur��%IR^J�Ol����b�;ޱ�^D�(ۉ!�$�}�gʾ��h��Z�s�wF��qDV
Uw����UsVE���,X�7$�/]�@�J������7���?�������V��ٓ=�Z8|Gog��ݤ�\LSZ�`.^Չ{y䊰V�v���ww���y�N�Jr��owذ�ŀq��n�U%U���Z�e'�#d�1�3@��s@����i�@nkP�����wOVԸ���$��u�v� �'z�ڥI$�o�4[<ht�Bn��Q��d�wx^�T��s�x�}� �9}0>[&��e;F�Q�nI��-����5R����>���xN���yR�ww{���[����p��B�V"M���%�3��
t�V�p:�ݹ�:�68�	tg��ڝ��[7�iIu�hn۵�@��v��õ�B<nm�մ�i.�$C�\[��rcE;g��9 05̈́�ŉ�f퍪J��m!�1qͶ�˭��:�>�3�̇v��m�b÷�@�[��Þ�]�ƨ��n%2���:�$������AҒ�Z�Y2+�����Ew7u�ٌbc1.3K��gްs�V�J�q9`5r#���]�"�5�<ҿ?{޿i�AB�D��L����4�[&��;V��v�h�%*ȞEq$7UV 6'�ވ�������B�3i$��LNKi��wxy7^���,?����;����x�gW�ƲD(�or-����9{)�ur�4=���z��?`أSEU\ 1��q[�_ ����Z� ��cw!�`��'�Li|N�|�q%\6����ì[m��a�ݟ;Z����\��؀؜n��ܠ1�Q��Cyߍʕ�7�J5̑�4�ڶ��"":D\�  �ELbq���;l����d�?,��5�PȜ�������B�8��r�Z����AB�D��L����R��ݠ3+K>�P��ٙ��57MĐ�nW-�@��@�;w4w�� �[������-K�2�2�5������r��n,��v��{uӆ�y�=7loG� ��?z��w���/e4�[&�^gW�ƲD(�m�"�;�� 1���ݠ7)�_�d3�	�b�Q��Ĝ���Ɓ��d�~>tE�`TEa`S�DLCj��Ј����q�]I9�{F����1ߜx	�4�4�[&��;V��v�h{}wƁ�JЛ���fK��@nSr���=}�|�8�ށ)�����Ɔ!	�I�F6��v.yp`hh�vFj��S�ru�+qn#^��ggVO�4�E�����9{)�ur�=��~Az��������r$ܒf��m����G:�� �����B���H�Eq$6ۆ����4����T�o����9��0��p��b�Eq	�˻�T�$�y{� �;��&��{5&< ¹���9Ԓs�v5�!Fcxۑh�n���ϳ9�o��U��4q���^��F�nE�����;��\�^�\�"�X&�0b�%۬O�T�^oRT�)��'&'v;��r��~�ވ��v�̭s�=���� ��j\@�mGv`�ۼڪ�^IU$�;پx{�ŀ}���=^T�$�<�؄����fI$����@�;w4ܲ�W;d��ۍ|�8cnI1��m$�'�w~X�m�q��n�<���*�����5���\��rո�]��v��k�@fV�@fkP��=�{�(�
��t�������7��E�:� K��V�ꎰf񝽻[h��:V݀Ca�B��˷6����ټ͸wtKb�a��8���)�#`�^(3�J#EKc�7hf�.yVӭ����J�� V%Ř5���k[R���Rg�:�5���}������`��*��`N�H�if��l���zIv���wRX:��ێӠ癋���W��T������ww����Ո�,�;�vq�ŵy.�O-ur�ђ����2y#WX���%E�o-�n��!$�@��}v�̭r��֡�;b5�\]@D�+�L.]���Nu��UT�{�ŀs���v�6���5�ۍ]�ڄ������B�v��k�@fSr�>�j''S��i��kU>ssL��ۼ��޼UR����wߖ {�H���q�&E�Hh\�@��@�;w4r�h���J��"!�%�2&bz��fE9�Ԟ�j��,	T���[^���w��Ys�B�1�$�p_���9���������^��5�}w�:o�t�Kr�8�8�ԓ��ƒ1�~U~�o��@}-��e7+�&C���-�NdN7&h留�vɠs�ՠs����IJ�'�F�I��8hRT��)������y��s��<��N��x�;���V�'�!0�ww�~�;�@~�{5����| 滴ޏz!��{�ݪ\�NV8��Gt����]�P�9n8{Tz�l�ua�����?I�b�/+W?��B1�9���M� w�6�)��I��9�)�Ċ�}w�s�u��s��RM���&Ը�㶣�0�wn�ߧz��Щ�S��4�T�U���B��<�}�@[�M��hM�M�(�d�I��UU�U;�����`�v�`y�s�w���?���rG��-����?�#w� �_]�3)�@l�.\�6T`���;�^;m\3Q��fr������[�8�њx�߽��O��%�&��m�޾9���Z��G������IO,�䍵cp�:��&������{� �wذ߻}3����L�X	�+�L.]����x���,6��*�);�_��7�`�:�v�Wlv�"���A�;��B7��mk�A>��#��"�U�9�:tz�o�c{�Ԓw�1�t�̹��a\��}��� 򤒯*���O�w�|�r���ߟ]hk��r<� ����jyv�K�GX#���D��Gn��[�ۧٳ�o3�&��n:�[�9�ڴr��g�留ʕ�7�M��"Hށ���^z�W�;�{���`�9�3�*h)Ob/c�4�$Z{�nh�e4�Ļ]�zz~����6�j쩩����9��@k��H��(?G˽��f���<D�Fڂi�8h�k�@fV�@f6��;b��г�G��1��T�UМ��e�V6 ���A�`�\�h����Q���^�6��:I�G%!h~G��7��i,'�H�a� 8F�"0('�I��0��"A ��!(C+�Z�dR{��>�쨟:z$b@�3�29�4�sa_�" 1�HF� %4^�IP��/694pg/ƪ�).^�
B �dc��}$j9T9��v�}{s���/{�����j�����m���,�#�]��8)v���e�]ll[u@Y���C�ɴ헲��ŔҨ��bs�vԨ1rw �1ky�6�;(X9��bjU�f`��3*��;�n���]R��Z�]��V�\	��{d�6*H10h\jhxD�I&�6�ځ�b-��h*s5J��UJaUa�6��tL�xX��n��c���
�duXс��]Y�h�Kx����4� �.)\�Ժ�r��=�g��m�չ�l�J�I��[��r0��K�V����Τ T�t�c�=+Ӑ����|aR'(��lX��y�j� @s�s����׵,����0+�)�U&��Vȼ���q�&J�.GV���n��4b��]m=t��5!���R[e+]���P 
��J� W�-����ܙ��;ip釖ǲ+WR��۲�H�������c���A��u�I 6�sY@�<@h�� Ÿ�Bڡ�;
�g���Xx���ɰ6-����ȏ\pq��uXꇈ��1�Aݮt'nK3�aj��h۪�-�i6�N�bĻV���8%�r�va�ܙjCru *�jiV� �QP�!�PY��l�l�Q���N�B��Aڢ5�8u��L���"s�,��kvӧB�8����JEխ੶�F�F���䞎e��Ė��<&($�2q\-��i��UƟ�Ͷ���Xknë��6�qn풭�������v�<TOQ���ܢ�8�U�������%ɇ��\�U �n���n����p���-�����=��v�8��ŗ��d�G88xݱ�E^8�e���WMOC&�iV��:���6�&"�T�K]���K��e�����P@�O9FA�F����UmY�F�PuF�t�����6��We��)�Z�q�;*-�C���Nf6�U�mlڕ�j���B2a���#m!1͝���kN��K��+, �zz
y�s�3��12[s�3�ʸEN(�X���QN�@�u@6m9���'ΰ
�( �S��uPv3%@�3Nt��:��ƹU��X�ݪخ�Z�*ʘX�9�c��T ����*�`�sⶭ��җ��K�������d�;<F��\q�=<�m=�����hN���۳���F\�d��9͞����t��q��s�;�X�n�t�z�t�Y��Di�t�[\�z�NQ����2mV炌Im��J�䍧m�n�v����O;<��jԓ�`+��f�����w��}���(M�����s���ؽCIWNg.��Zq�l�n4ku���~���6��m�s��ܕu\mwJ1���?G興��ߛ���_?��H�1��QǠs��h���~��d�?>w�=IR^IT�����y;��v���������� ��k�9�w4�G�w�	5#p��z']��@l��@f6�G�_.T�	�lP�b$��Vנ}��G�7��6�� >dT�k�Ի����������I�õ�6En���-��7�\�vid�����uz�'k��o����`�o��������|ïwf sʿ�6�jA���4�)�Y�/�ވQ����>�@d�u 3P�{�*�䍵��s���������P�}��7X�&���$����A��뻩�ܡ����U��U󱬑
c�ۋ@�-��9��h��o@ⶽ���UTȞ<��,�䷷Y�[�zX�ɼY�Z|MС�v.���s>xۘ�jb1'3@�l��ξ��+k��g�ｹ�{����	�d%�0ܜ왪��gwf�n��9�)�Uӭ	��B1��7�r�Ƥ�}��Ԩ� ��	�c�Φ�ξ���r��"�Id����@f�b6�� �z"v�u �_��6�jA���4v�h��o@��@�-��/]ƓĄ�"%$�s���Q��R*j�ڻslڇ�����'1�sϫ&�JE�<����cN:�[�8��@f6�����\\�D�R\�%M�� 2u�]�L�����@s��� �ү��d��cx�q���؎���κ}T��}Ԁ?V6�)��I���|�}�4�|ޒ}y��Rs���HDpb�b�`-L�s����{��}5$�Ώ�~��4@c�:�[�8�k�?[w4v�h;ҽYj&c��s�g�m����m���\2��\�X�M�c�(6����(F1F�.��������k�� �ŅʌS�\�K��}��mUU6w�za�$�vnɠu{�z���$�NcN)&h�؀�M� 2[t���� �ff�D�Fڂi�8h{>��}=���{�@�m��;�)�v��y��LDb�U]� 2[t��z#;�����@k��I0�z�@I�i�����pd�(��"6ro\I���mVPɉ+8�fr�* �[�NN���n�T*#a�R�X6������s��ˎ:��5��q9��/�����u�Z�LL���>ۣ�k�y��p���A�Z{	 �t�K]@d%î7���Z낶ڰ� L*C������{/m�����k�ڭg-Z���a渎H]�Uٺ�yK�m����e���ߝǻ�o����̑v9���n�W�8\�Wós<���$̭oWk�'�VH���JG�r۹�w�S@�v��q[^�^_�6�)�I��z�t�R%�H�jD{�'m2�^�G��8h��o@ⶽ9��rِ��h]���р�P��e��P��v��n��3��1��$i���۹�s�S@�v��s�ՠ/h���8�Q�`�0g5������ӎ�a�Am��\��ȶF�b�NG&h��9_kz:�Z�[��[Ԕ)���&ƚp�'���cZT����js�֮���;��s�S|��{؞l�`�!E�hu�(���� 2q���5�tk$B�on-.w���o���qr���h�~x���j|�NB5�8�H�nPcjkܿ޷tٹ�Z9˷\�;Nn�f#J����6��`c�M��[��m����l&�s6@d�e 3i�@}��@f�bgMhM�IE�#��9�j�bG;�nh��4.Z=�Ď������G%���~��,�;}0�%K�$R���aQJ��J���0 ŀ��Xb!Q�]9:���|�V�~���mFӌM�U�?G�_.:��m7(?z'w��ީ(x���YcM8h\���#��~w��k� d[/���3�n���n�lO����Oe���� �gmM��]�w<�y��]��DU�����nP�؀�v�����|R {>�ᬑ
1�q��r�h��8��=�v��}�A����
AF��JA���Nk)�M��v��c�_�yd8�qr���h���Ԏ�A��mP,A}��SRJ�Zw�QF1H��uڴ��3yq���@d�e mӸ�*jbq�+n��'�ػ.��ZQ݁���jy��;�b8�����4�'��Ƥ�7�@�,������R��b f�&I����q���4�즁������M�����"�򇈜���&���l��f��؀�6؀�n**��`�!E�z�s�|h留�ܾ�T�$�';���vU�#Wh�QPU݈���ָ��}����f��, �"���0D�n���㿟��o����4tE�d�MxW"�:�A���s��A��l��㌅n��g��騽$�����a��ظ��Z�c�%�k�^��Z��Zջp�n�d.�6���h��ؚM���
l�E�vRHI�nLO[��]��s�^z���-bM��=),k��Ͷ�P	��Q��6ƺq��[IĠ۲�����i9擭�aV�cj�!��	I�ʿ���������;�?+�&��;�Q�dpg�vF�M��eQ%�Ɲݪpפ ������%!�9})�qr�z:�Z9e4�G�H�&�q�@�����]wJw��k� 5�I5Wi(���z:�Z9e4v�h\���İ�~&69$�8�[�H������N7��6؀��BQ5N19������8�ۏ@���h�e4tO*rcJAcc\�9Up�����us�th�HK�r�$j�4�u"�"r6�D������z�vQ���m��eER�"�
��n��1�&��{58W�d �¦�."�_ׂ�v�N6R�z&A�uz�d�F1�䆁��x�?s��-��������a ��BRٶ�Nk)�M�1�)�^W���p�8��=�v�y~��� ���Lj���X=�[�XИ?��'���f�Nz��M���mv�8X�����Y9#����66��E������h庰����$�`s���>l��իd�������cj�؀35��Hk~���Q5�&�4v�jI>�����M�x�3Zm�$~�4�I��A�	 |B�B�F
�(@+�4�HȄX��!X�!��A�"C|�� �C�H�0�3��21�I C$(Df&�1%V|�gaʤ���B��CRB���C&�E`�g$fe!F	@�3D*D8�w�cd�&yN��݂\�b����0o8�8��q2�|+�A��M!! �#&�@E�Fp��j�)R�y2��O�ʠtG���V��uQC?��p�%�x"�ұD�s�kWRN��ѩ'xU
D�m��<m��C�f|�{|M]wJ1��l@f�
�`E�36we�3i�@fkP��v���&�{r4\$����i�ǐ�2u�����Q/#X�퀺��z؍�́��O���D�9Z9n���M �;I�s�ՠ��Ⰲ�Q�$���s�Qw�!��Z5���tȯK�X�Lc��v��?s������;)�Z�ZsТ�q�2h��{5$���Τ����ԝD��H��(������|gP*�[�2dC���4�-��v؀35Š>Ͷ :=�йAwQS'g��ۂq�q۶�:��ԋ��H��m�Z���u�.h��6�,���=U~m����� fk�@}�l@cv�m͹���m������qs������ܶ`~���T�$���Y`+���v[���k��ݠ>Ͷ 2s\R �-HƲB&��rC@?r٠~�e9�)z'5�oz���&웫�n���f���]|k����RN8(Ӯ,0+E��j��w����߉`iۮK�%����86����݊�TlI�]	.s�+&@�U۝ח�'�8nq:ym��Rh����X;3�=A��/�q����l���Y�su��)Vnm���rU�NL��{Dg\Ŷ�+7/���cb3Yɮ��m���&��-Ǒ�����-�Ә��G�k�ʣ��8ۛnK([�bL1��K6B��\��ޚ	[sǻ��������=��o|�N�۶��3�{�]���ܜ�u̬m��g��ݺ}�s��s�*�π�k]���b �n�"=�;g����CS"ih�)$z�m� f7h�m���t�����{�T7�Hy+V�w#��f s���~����UUM���n|;7^ t�z�;#�.7���j^����}� ������@?r٠~�B�9k"x�Ny9ۘ��*�UK������׀~��*�]QGF��$`��c � �<]CN)��])�\�痥6ƍ��a������JȒ��#�9�j�r٠s�S�2���8��& w���R�n6E.�I&��s�9A�Zd�@H Eg�;����>]��)�m� <�6�28�rh��M�����%���@;�zh���W��������R��b �n�w�9�p��~<��ȚB&)$�����?����w�'5����Q3:�����3��i8�y�̯Mn�ٲK4(0���n�i�Ș�d̙�m1���4�m���W�����@>�$�)D��I�M�;)�qs�z�vS@9�f�>H����D�m���lI8i'/;�I7�3٩�,SaD,��h�DR �EA����u$����9��y��	�Ic�A�{1s�p�7{��m��Z��u�g�&��rC@9�f��}������|ށ����?\>eC�m��n��n���n]��&�7X���� �Nk\M:ޙ�{ҽ���D�8�M��v�����~�e4�-�k�?��,q?�1��\���b ��ٶ�Νh����(�nE4�즁W;^�����{T�ܣ�2dC��ʺ� �5���b o\���Da�>Z��!��U@���T�$����wA����ˍ�]� >ݶ �͠7i�@9�t���{��c���x˗v�ݞru� th�]�CJs��*N���p����Հ�t4����V|��m�M��k�7l@;�<Op2D'�%�9�;�j�*�k�9�)������fgͅ�_,��6��yv���� ;�uM�v� ��6�28ő��v�h��h�h/>�=�~1���c��"��� 7�m�M��k�k�) �����, �,l�{j{]t5T�N#��by��l�F�;��vm� =���h˰ho&D� �P��;P�I�)��'�@3a�-����{���	)��͒wS�9���`ѷ5U<�;���Rvg����O<�l �Lx����ݞ�z&��ֻ<�����ɺ3���Fۂ�g\�������A����Yԓ��-n/a�g��w���v���n9���+Y�۝ũ����S�J�1tvZQse�m��ހO��I���̵���t��@f�b o\��܀��L�r4�qH�
���v�h{λ�>���UT�^�<o��;##IƓC����ƀ^����gؗ;g���=ڥY���'��$ᡵI*�I��;�9ݿ_9ـ}��� ����f1<�D�E4�즁_9ـ}��� ;�u��J�l:�j.����lu���m�lx2�q�\�j��z�6���]�O�7ix�V��~�� >Ͷ ���f���v2Ւ���r���_L���RJ���Q� ��m������dW���?�1� ��S@���i��|���z;g���h�ǉ�"F(܊hyzs����w� ��/��J����� �{�_�D4�#C�k�h�ݾ����� ��/�滯u'B+n�wn�p�V"���]����ԦJ��6H-��ך��&Ph�)�����4��M�;)�v�ՠ[T��q��D���p���4�즁��V����h��0���B$r)�~�s٩';�v�l�&:0���tiZ�A2���1�@���\��:�����w��s��R�r&�%݈u�Pmk������b x�۰D�8�I�"�?u���[�)�[<h��h���8f)1̟
(�����]>�F���Sd�z헬(��1D��m���'Ѳ錊E��h��M�����9]��8��&�F��
7"��m��z"&G��P������G��G=�,���(�ㆁ|�ֹ@�͠>ݶ kpI6T�II�1�����h{j���S@���yN�����{q9rHչ#�� n�6��v؀�Z��ֹ@}�Pƾ@�(D�1�#�8(�CŶzz���͔oI�6s⻶�wnq�[C�S�����۶���(��� �nm s���ı�#x��䆁��}/��9]����4�즀~�1�a�dq��qh��V�w�����3�Ɓ|��v�c�_�d��@;�T@}�l@k��DDDN;}(�uI�ƢId��M�{)�v�V����x�����$�j"��@���"M�MX0�0 �H� �0��|��G,sR�� �+�0� 'X�T���"B0IR5 � BL�"E!�ʄ22�,�7�� @b���2`�&G��@�T�j(�[FM�0�@��0�0Г��*qm��F,0ax' )^�~O�'c;�};�Bf����T���P�AHF\���ѥ
��|Ȥ9t�ORV$0"A�0`X� p�(�>�ň�)1�Ȍ@"Db\��6���H@�2���{G�ㄨHlb|XF�Ϯ��)��L�`F0bB�|3�,Gđ
A�E�a��$�&&�@�d�d�Hđ"�$8�f0�!Fb8��S�։!L?t��Y����w�{�Wߥ� 2B�⪪85�-΅@n�gq-����F�	���⭭̲�ٶ$��rf�����|�m����z.L�!*���ULn�*�isv��
D���l�vF�Ic7�g9�Ug����S�]���^z��c���R��tk��I��AvE*�Xc�M+-��ڝl�g6�!vZ)��@��,�W�����s���t��s���nݲ����$�F��u;�˶�.zw;Sr�69�t�\��fJ{�8�r���]E��h����9�'�N��Y䮎��v��s�U�5���1�A�8�n9��:�%�`�k�Z����l/7m�{{[��2���y�]l�l�O�,a��:u���$`V�"� ۓ&��S)���7Hm�@P!�UU@W!�4&zN��n��M��Dq��ڪx �y�n��M+��MSp�)e��3q�[�|�
d���e�ݐf��ؓrP�n-�h{M����k���٧=�����l���$.�w=�Ӯ'���rl`jYt���L��t֩�sZG<$ʄ$��nj!���vvٓS��FE�&����U��@9�F���:-�Zi[�۞l
����ԘD�vu5��e%�Z������]KB�%��;�u����մ>���KJ1v�^����n���^��yW�����r��j�����������n	c8һ=�d6�cv�y�v͋�6L�۵������61j��ڱՓgC�s���l�
9x����@1y�4F��ۙΞn�ؐ��J�q��G*�rm���t�l�sۜ��7.Q�I�nk�d�)GYEv�H���M�z�֐�^��2�r���S,��Ҫ�p[6Ûr��Ԥ���lꮺd�'��9.���@VQ�ٕ%�xp��*W=�<��{c�.���-�����e��W���#m��i6�B7��h���@�h�vĐ0<�5��	׷-�Y.g�g�:2(����<�#�D|�Ĩq2H$B"�:#�(���^� x ��(#�C��5�)���9WFʞ��/*�nd�I8�6�%]m���8�;=�F�����\����I�W�7m��I/l����Q����k�vv�Q��ٷ�7.��=,�a�˚t���MF�S�9ݛm��ūPqڶx�X6��u��Ӈuz�s�����	��[�mڹ�싙��|��[(sx8z��8�i�v�s��j�������N���������/�.Lフ[ps�ݻ7�6+kTn��fk7Z�k'H�'\{Y>�L2<�,�LhjH�C��ڴ�9׀�z��~����7|v4F��o�h��V�w���~�e4�ڴZ�u��m����'�n�6��v؏�����}(t�P�WTL�Li�Br)�~�e4�ڴ�}�@�;�T�s��ؖ9�oTwb��H��v�~ ��6��vS@�g2缿8�6��2(�ƙ������]6r͖օkM��a�My����չ� �5#��w���@/mS@���%�{ݘvh�f��Y*�-ݼ �;�x���ժ���c�/���v`rv���H矚<�j$�H�Q��9l� �H��� x������~�hi�F�4
��@��ڴ�-��r��;�#JF6���mk�����;��1�� �[�n�����Z6gv�ƹ�m�6�j�j��:����:u�����:�}�>~{2��U�W? s��@}�l@9���G����=�,�fEy�I4��ηH��� {��2���BX��X�rC@��@��ڴ��߳�� ��&U�D��po��I��=��)I��;�G6��X����̥�I�����N{^�t��bX�%�����7ı,O��zi7İP�=����/�L��L�ݽLڹ�V�n���bX�%�{:Mı,K��^�Mı,K��}�&�X�%��s�]R���L��]Zk��FA0l�����H�=Js'`�C-�t��Y$7^��ŵ������y��;ldh��]�R���L��_��zi7ı,Oc��4��bX�'��}t��LD�,K�����n%�bR�=�k�j29v\d�fR���L��{����? �D�K�Ͽ]&�X�%�x��:Mı,K��^�Mƒe&Re'�7A������F���[�bX�'��}t��bX�%�O{:Mı,K��^�Mı,K�ｍ=�����ow��~�'�̮t�X�7ı,K��t��bX�'��4��bX�'��{Mı,��S�@�\|��_�g{��Kı[�5��Aq�d���)|Re&Rq>�u��Kı=����n%�bX�w=��n%�bX��=��7ı�������T<�NZ;\���u��![l�h�ա��)ּ�k�;�F1O�7hm�&3��&�X�%��w�Ɠq,K���ﮓq,Kľ��gB�bX�'��4��bX�%�Lc�.L˜䘹�3�&�X�%��s�]&��B8���%�����7ı,N{��4��bX�'��{M�Kı;���r�B���_�I��I�V��/�L��L����2��&W�
P����n%�bX��}��7ı,O��bX���N�EwyK�)2�)~�sf�q,K��;�cI��%�b}���I��%��X"c��߳��K�e.o�C^�Q��d��,�_�I��Oc��4��bX�������%�bX���߳��Kı>�u��K��K+��4���MR�?���.�`���i�Aպ�CΓn��]om�۫����r��驺��=���������]���a�mokSc���$�������^Y�*l����1�Ͷ"�ck�����gl�9��4�εg$�w������.�Hpua�l�w&����#8�����c��˘{oecAk;��
��<�D�ٚwS
�WH�j���	����&6��c�J�.6ݵ9��+mH�k������o8�8��3�[�6����c����&Re&R���^�q,Kľ��gI��%�b}���@n%�bX��}�i7ı,N�x�?veS�r������7���{����gI��%�b}���I��%�b{����Kı>�{��Oኘ�b{�5�� ��卲\Ww��)2�)19�k��n%�bX��ﳤ�K�,O����7ı,K�O{:Mı,FR|���Դ[���̥�I��Jļ�}�&�X�%��s�]&�X�%�~��gI��%�X�w���n%�e&Rz���M�j�wh�n]�/�L�ı>�{��Kı/�=��7ı,O��zi7ı,K����n%�JL��IU.�%���-Kv����Ri�	p�����Z�{a�L�[���۞����j��Կ�I��I�W�yKq,K���צ�q,Kļ�}��'�1ı9����n%�bX�����1Gm�6�܊���&Re&R����I�o`�(t@�s�3��9ļ���&�X�%��g޺Mı,K���Γq,K�����|bɌg3,�q���Kı/;�gI��%�b}���I��?�����y����7ı,N{��4��bX�%��%�37��Ų�9�n%�bX�w=��n%�bX���t��bX�'��4��bX�%�;��7ı,N�z���qrHչ	#��R���L��O���/�X�%��{�M&�X�%�y��:Mı,K�羺Mı,K����b�3
Y�F�n9�"������p�]9��C�=	�5�kXN�:��#Ў'��n%�bX�w���n%�bX��ﳤ�Kı>�{��Kı/�=��_�I��I�sv(�Դ[���3I��%�b^w�Γpı>�{��Kı/�=��7ı,O���)|Re&Re-�tR9�Z���%��s��Kı>�{��Kı/�=��7��ߨ� ��L*���N�$(l��K?�ksI��%�b^����7ı,N��f��\b�wo)|Re&$�K�����bX�'��4��bX�%�{��7ı,O����7ı,Nr{E=a��mĥͦ1�&�X�%��{�M&�X�%�y��:Mı,K�羺Mı,K�����bX�'<a1{�F�c���5�$h3�F��r�vFdZap�5�];V�N��M{I��Η��bcc8��}ı,K�{�t��bX�'��}t��bX�'�=��7ı)K�{�e/�L��L������D�&.s��7ı,O����7K�9Ӿ�j	 �w���)"o��U�-)2�)wMxin]��!$r[��Kı9Ӿޓq,K���צ�q,KĿw�Γq,K���ﮩ|Re&Re.sF���]�,nGm\�Mı,�9�o��n%�bX����:Mı,K�羺Mı,����D׶{y�n%�bX��=���&n-�&3��&�X�%�~｝&�X�%��s�]&�X�%�yӾΓq,K���צ�q,K���)��v�����q��=�(�rm�����Wlж�֍�oL���'m�ޮJ:e��n%�bX�w=��n%�bX��;��7ı,O��z�? O�b%�b�7޼��I��I����g��.1Z�79�Mı,K�}�&�X�%��3�]&�X�%�~｝&�X�%��g��Mű,K���Xb��q)s�c39�n%�bX�s>��n%�bX��{��n%�bX��{��Kı/;���7ı,O����Lc9���c7I��%�� ����~Γq,K��s��I��%�b^w���n%�b؟s>��n%�bX�����鋛�p��ۜ�:Mı,K��}t��bX�%�{=�&�X�%��3�]&�X�%�~罝&�X�%��P'{�w{ۻ��߿��2]E	Xj{7?������ ո�휼���ڎy���졻 n�i�66�l��Ξٶ�J�S�@��Xh��b�lL�!��6+�r�Y�a*�v/F����-��Y����m-'p=;�7nmip�Z�=k����GF�S�HTm�%(y�f�9"<=;JԶu�^��j��v��7=Z 6���vy^���I�1�^�k5��������>��x�E8�'9:ܝ�&@�j��:Q���Z�)'gM��9;���]���is��Ac��7���{��?���t��bX�'�Ͻt��bX�%���t�Q��LD�,N�>�t��bYI���������p.Yw��)2��b}���I��%�b_��gI��%�bs�ﮓq,Kļ�g���O�R��B�)>���F6��nFD\���X�%�y�߳��Kı9���I��?�����{�O��n%�bX����)|Re&Re-�褚�v�w,%ی�I��%�bs�ﮓq,Kļ�g���Kı>�}��Kı�n�R���L��_��Q3j�.1Z�nst��bX�%�{=�&�X�%������>�bX�%�~Γq,K��3�]&�X�%�㞅���1�����&�nqjd��R�����3�$mc/��[7o@ZWn���Î)m_{�7���{�O��{Mı,K��t��bX�'9���7ı,K�v{:Mı,S)?۪!��Q��d�ܹ��)2�(�/9�gI�p�P`#
ҌQ�C�F�t؛�bc���I��%�b^���n%�bX�c��4�)2�)2�_��c�;pr�iܻ���Kı9���I��%�b^{���n%�bX�c��4��bX�%���t���oq���������is��Ac��bY�R"c����&�X�%��w߱��Kı/�����Kı>��^R���L��\掷�m[�%�p1��Γq,K��ﱤ�Kı/9�gI��%�b}���I��%�b?�շ��)2�)2���^Vy�y4K����S��g;�< �[
aB��뇒�=���i�3�ͮ����)��O����%�b^�߳��Kı>�{��Kı/����7ı,O��{Mĥ&Re'իI&���	c�yK╉bX��{��Kı/����7ı,K�{��n%�bX��ﳤ�S)2�)s����W!q��v��+ı/����7ı,K�{��n%�C��B,#�M 6�g�>���$���'Y���mt\sW AF+�"5)���FE E���X�!�}�����>5����HM-Xy�01é��a8+�s(��B2�A����`�%M���# "�@�*0!�a �T0j����A� ���
�V?TЫ���&�"��G(R�4�8���S�&�C$p���C��衕3�Q�"�Tr� ��b�>A()]��*
tP("D:��Qk̀�D�K�}��7ı,Os>��n'�T�Kf���Elpi��ڻ�_�I�����~Γq,Kļ�}�&�X�%���޺Mı,K��Γq,K������F]�'r�R���L�ļ�}�&�X�%��g��Mı,K��Γq,K������Kĥ/%���.@�Ib�*�ٕb)^Χi�b�%н����F���cM6�%�3��>�bX�'{�~�Mı,K��Γq,K��3�]�g�1ı/{���n%�bX�����f����Ac�w���oq��������v��V8���'��߮�q,KĽ�gI��%�b{�ﮓq,K��::߭�]�,c�.��R���L��[���I��%�b^s�Γq,K��3�]&�X�%�~�gI��%�b^��L�ɛq�0��8�n%�g�@����}�:Mı,K�����n%�bX��x�t��bXj&FT�`Ѐ��	������3�]&�X�)���)&���	m˼��I���'����7ı,K�:{:Mı,K��}t��bX�%���t��b]�7���s6� ��1�]��u���zUuLW�RIzK�F�G=n�c��3��^�g13s���Kı/����7ı,Os=��n%�bX��ﳤ�Kı=���I��%�bw�Ň�&�q)s��&s��Kı=���I�~H�&"X�����7ı,O�Ͽ]&�X�%�~�gI���W1ļ���Z�%ݹݼ��I��I��{���n%�bX��{��KȬ1/;��t��bX�'��߮�q,K����=#.7(v�˻�_�I��Os=��n%�bX��{��n%�bX��{��Kı/9�gI��%�ow�����ӡ�N�+{�7���x�/�����Kİ�G�׿]'�,KĽ�gI��%�b{�ﮓq,K��$dg���\YpdɌ�%�t�k����j�7��M��H�=\Ϸe�ū��-q�s볣F湧�ղsnܻL%�g�m[b��uisZ�a1��u��iq��l�VR��{n�M�RW���?㾱�kA�a##Vgt��`�W�=�5�ZB�ez��21:��!��v�)ۣ�a�j�՛�:Tdv���5[-���t�:�q��b\M)&���6�8*T�V�Z19�h���4˅�6�f��CŶzz���͔�gd-⻶�wnq�Rqw��"]��JL��L��_���%�b^s�Γq,K��3�]&�X�%�~罝&�X�%�y�{Ŕ�L[�Y�\��7ı,K�;��7ı,Os=��n%�bX��w��n%�bX��{��Kı/Oz�=�\��8̘͸�t��bX�'����7ı,K�;��7ı,Os=��n%�bX��w��n%�bX�w=�<܅�XB���_�I��HJ�;���q,K������n%�bX��w��n%�bX��{��Kı=���ŬDV������/�L��L������Kı/�ﳤ�Kı=���I��%�b_��gI��%�bS��=r�C`�V��}�7a���3�l1X�7Z�k2��n�ێ.�y���:�ɳP�}��Kı/�ﳤ�Kı=���I��%�b_��gA�'�1ı?w>���&Re&R|����e��&��9�n%�bX��{��6����l����6)�q7ļ��Γq,K��3�]&�X�%�~�}�&����ow�����ӡ�N�>�~d�,K���:Mı,K��}t��c��"b%�}�:Mı,K�s��J���L��[ө辸�w����q,K? @�O�׿]&�X�%�y�~Γq,K��3�]&�X�%�~�}�&�X�%�y�{Ŕ�L[�Y�\��7ı,K�;��7ı,Os=��n%�bX��w��n%�bX��{��Kı8x���f��9�3L�����v�R�Б�\�6XgK`���n�t�����)z����@�����7���'����7ı,K�;��7ı,Os=��n%�bX��w��n%�bYK�o���W!q��v��&Re&Q~�}�&�� #���b~�}��7ı,K���t��bX�'����7��U(Re/M61y����ӹ$��n%�bX���~�Mı,K���:Mı��"5�b�L0�"	�~Q:	��!�q>�����q,K���f�q,K���5)�&,��܍�v��&Rg�BP�9���/�,K������n%�bX�s�٤�Kı=����n%�bX��t�_LY�Za�ė9�t��bX�'��z�7ı,O��l�n%�bX��}��Kı/�ﳤ�Kı;��XǮ.Y��!�q�s�q�&�˜�CM(�]K��[3�e�]�ݓl�8(�iS�EE��ۉbX�'��i7ı,Os���n%�bX�����n%�bX��{����L��[�����E�r�I.嬣q,K��s�]&��QX�&"X�����7ı,O����I��%�b}��f�q?b�"X����a�-1�6�+�g7I��%�b^{߳��Kı=���I��?��"b'=��4��bX�'�g���Kı/Oz��;��V��_�I�T%
^���R�Kı9�~٤�Kı=���I��%��nqz0r!��S��D����&�X�%��g��|��gfLL��Mı,K�w�4��bX�'��z�7ı,K�=��7ı,Ow���n%�bX�;=K�o���38���6���ڲ�=Js' )v긍6�������I�O�vz;8�n����oq�����t��bX�%���t��bX�'��zi7ı,Ns�٤�K��K��`�ը�]ۑ�wo)|Re&%�~罝&�X�%��{^�Mı,K��i7ı,O{>��n%�e&R�PǤe�Ԧ�K���I���'��zi7ı,Ns�٤�K⊐�LD�=��4��bX�%�~Γe&Re&R�xin]���Y��ı,Ns�٤�Kı;����n%�bX��{��n%�`~���߾�)2�)2��y?�q�$��M&�X�%��w�Ɠq,K��q����'�,K�����4��bX�'9�l�n%�bX�@@��Z-��QH ���� {�[�ͺ
��V�X9�������v�@jw&�p���м�e���c��Ӄ��Mi[շ4[q�L�X���l���'kcƶ�Ӯ4��^]�ݔ�k�T��fJ��m��)�v�5�a�. v��X��&�#pۇz�mv(ݖ��n�Hj7�Ԇ��C�t�K�'7vf�gi	حU*�3u�H��v���~��r�ڠZQ�,9���&����>������w�Qwn˧a:;r/us���N����Ψy��fۨ��k���>�C/�nB�L�8�8��bX�%��糤�Kİ�1����4�D�,K���ȓ�J�I��o�2��&Re&R�<�)�93-0S�t��bX�'=�zi7�q,N�߶i7ı,Oc߿cI��%�b_��gI�����'sz)Oj�.2��K�)2�)s�ݚMı,K�ｍ&�X�%�~｝&�X�%��{^�Mı,K���[Km;�KYK�)2�)vw}�&�X�%�~｝&�X�%��{^�Mı,K��i7ı,Ot��֨�]��v]��_�I��I���t��bX�'=�zi7ı,Nw�٤�Kı>�{��Kı;�����)��=�ҩ���m\�U�C]�x���4��'�����Œs�LcΓq,K���צ�q,K��{�Mı,K�羺Mı,K����_�I��K�k�jܻ�5nBI.34��bX�';�l�n
 b�����Qt�&�X��}�&�X�%�y�{:Mı,K��^�M�^T�R��)2��y?".�2Iy�M&�X�%��{����bX�%���t��bX�'��4��bX�';�l�n%�bX��ﱇ�c&,����t��bX�%���t��bX�'=�zi7ı,Nw�٤�K�� �J[����I��I��Ox�����D�\g9�n%�bX�����Kı9��f�q,K��}��7ı,K�}��7ı,O�(�����8��s��C��݆P�C2�.YY�^p2�"�|P�����4u�zy�[9�~{���7�ı;�~٤�Kı;�{zMı,K��{:��$N{��j	 �zl�`ȇ\�Z�H ��w�KQ=ı/�����Kı9�k�I��%�bs���&�X�%��L�y�K�n����&Re&R��yK�,K�罯M&�X��:�T�jD� �*�q5�sf�q,K��=�cI����L��oPǤw"p��.�)|QbX�'=�zi7ı,O��l�n%�bX��}�i7İ?*�Ls߽yK�)2�)oO<�V�ܑ��8�x��n%�bX��}�I��%�a�A�s�߱��%�bX�����7ıK���)|Re&Re-�;5F�#v�L����Ӛ�K��uqF���i�.KH���ӹ���Ñ�֗�Zn������X�'1�{Mı,K���:Mı,K���4��bX�'��i7�e&R}�vJ"cR�m�[�s)|Re+Ŀw�Γq,K��}�M&�X�%��{�Mı,K�g��M��t�I��Ox�����D�r]�/�V%�bs����Kı>�}�I��%�b}���I��%�b_��gI����L�ͽ֮�]�2��+ı>�}�I��%�b}���I��%�b_��gI��%��`�uT���h��> �l��/�~�Ҿ)2�)2��|�=���$��n%�bX�s=��n%�bX�����n%�bX�s���n%�bX�s�٤�Kı>�&K����b�sm�(n��l��]&z���4ș��Iuvcۨ.�s����ը�]��e����)2�)2������Kı>�u��Kı9��f��"O�b%�bs����KıO���Gr'\�w.��&Re&'��4���H�&"X���l�n%�bX��}��7ı,Nc��4��b�ow��~�~�*t*��~oq�X�'9�l�n%�bX��}�i7ı,Nc��4��bX�';�zi7Ǎ�7����?xw旨
�����{��%��w�Ɠq,K��9�cI��%�bs�צ�q,K���MĲ�)2��{�Q��lj�˙K�ı;�{��n%�bX�ｳI��%�bs���&�X�%��w�Ɠq,K���>���t}Ӈȟ�@މ֨�:,(�L#ڟ�~ʧF ���*i�/�����&"����n,HH�n�Uk7p$��J���ئ߸#���m&C� P"�A�e��#ɤ�w���FE�;��&�I����5DH�tu�o���$ �������<i�$&��{��	�*&� r��B���!��R1�R��:�H	,A�'D1�Y�r���h"�l��ڿ-���`��!*���2�E¼�3�����m�m��$��
U[�����G3��Ӽ5���@�Y�he��>��꭪H�A����E%�ڤ �^5,�n����T<XӘ��0��@x��� ��d�<Ԥc8�T�P�4��\L鵗FL[�vFv�!;�S�ܐ�9UgE&m�L
iQ�E�Ks��!�#�# ��޴$���M�KS7v���؜3�oYJ�-�9���c��hL���Y�G
��e_����^�h�}p�j���A�@�z_��`� ɶ�{>ݶ�d�!��bx�:�CmRe:Rܗg�n�4���r�C�)�����g�d��	����q/<ϳ䍱�g��cUN�ƒ�Ch�@�s�ywl�u�n�j���E�C��V@�P-m�4�E�KS.	L��f����p��N�/�����L�M�y<7O�jM�����ٕv�u���!L�nڶ�,q�S]��pF\b �^�xV�=K�5U�����'����,��:ZC�1t�Π%'V�fh�)��l&�޺��ɲ�#��r���jLZhkn�g���JL�f�!��]�N��v˹��̓t�J�m�Zle*خY���ʵ�lZ�j�����V��g:G���� 5�&�&�u˳5��r8:��F��sѝȲ��nϳIt�^�ٝn�3��-����,���Jܮ7S��N�<vj�CɆ�n�q�̓�.�7fN�U�ێ9�\v�X�v:�۰����
�^�:4�I�wd�$����[uЇ��Uv���ᵩIj�lTh����P�Z�0�j�}����6��NϠ���Wp�v��m*��ۥ��mT�/@e��B,c��]�+HH/K5S�T����$��gG5�L�kC��-�=HN�c
���E�^[P�����F۴˲����t#�H��M�B�af�N�5#���w�E��@]����e~��D��X�7]`d��m!`Ik�����*j�Ü�3-�gP6��<��P0���h � t�-P8�� �T4Uڣ��
�K)U'�_��7v�e�rKL��v��tc�M�����Gٸ݉;$s(ø�)��k�on׭PVBut�yu�3��N�-�r��U�3���ˈ���I��Pm��K[7�떇Vhf�1ϖ�hD�4����8�r��K�+6@ѩ����]xߡ��E/f�gr�a\�.�荤6B���l�'�z�X��5i25�٦�gF��$�l��������o�~o�?�8a�6�N�nc�h@�v�;*�n4�ū��z���-ݮ�N�E�#Q4仟ԼRe&Re-�L��Jı,N{�٤�Kı9����n%�bX��=�i7ı,N�>�3��g�13&&s��Mı,K��i7ı,Nc��4��bX�'q�{Mı,K���4���T�K��/�O�C���$����&Re&R��ze-ı,K�罍&�X� a����~��I��%�bw��l�n%�bX��5��0�v8ݗw2��&Re&R�罍&�X�%����4��bX�'��l�n%�bX�s=��n%�bX��t��N��r\�_�I��K�;�Mı,K���~��}ı,Nw>�t��bX�'��{Mı,K�~����6Qq�z���td
֩� �^��n�V�ܛ]Mu��]	����:G��[��Mı,K��i7ı,O����7ı,Oc��4��bX�'��i7ı,O�{��ng3�q�����4��bX�'��}t��P
e�?���L���j T+UxF��\~���'�~���n%�bX���l�n%�bX��}�I����B�)?n�J�cR�m�;�o)|%�bX���~Ɠq,K��;�Mı,K��i7ı,Ns>��n%�bX�1�F���ə�`��1�i7ĳ�;�߾4��bX�'����&�X�%��g��Mı,� ����e/�L��L�Ϳy��E��I�1��fi7ı,Os�٤�Kı9���I��%�b{ﱤ�Kı>���Kı8s���3Lc8���M�۝�� �ŦX�+�g��ҥ�@�ͷ7F���Ŷ�ٱ���[��~oq��K��}t��bX�'���Mı,K�{^��	>���%�����I��)2�)o���W�dwv;nۖ��,K��9�cI�~A#���bs��l�n%�bX����4��bX�'9���_���
L���?܌�ڎ�8�n%�bX����4��bX�'��l�n%�P���m@ш���g�]&�X�%��w�Ɠq,K)2��F���.�\qFK���)2��b{���&�X�%��g޺Mı,K��}�&�X�%��{�4��b]�7������w旨GR����{��,Ns>��n%�bXq#��>Ɠq,K��=�Mı,K��i>)2�)2���{��˅� uwn<F�gbm�`�հ8)�@<�i���>c)[����"&5.6ƮIo)|Re&Re-��̣q,K��=�Mı,K��i7ı,Ns>��n%�bX�1�F���ə�`��1�i7ı,Ns�٤�Kı=��f�q,K��3�]&�X�%��s�Ɠq,K����s����$�?��nh�hs����:�ׁY��Ě�&��2����H�lA���#���DB .1H	B��/��~5�ǂ��Ɔ���D�ZW;^���S@����9�ڴ?w���$1D�^gG`���
��W���b;3r�e{	D��u�E
F��Li�z�YM����9�ڴ�v�򤩚ڑ��7RK0���UUT�g9;� ��vh�e4g-I�F�D�M2G!�fV�@9�t������� ��6cB8�B�ۋ@����,��{�M�}�@��>M\�Mcŉ�����l@fSr�s���";����
�T�S�'���d̙�9�x��hÝT#q=t���V;�L'=�$%z�n���Y�:�L�:�H��w�����*R؍&Q��-�$ôz�d�����PR�$��f�n��i|q+���Q�̎���ԫj���Xv�s;�E8��Ϭ�t4�vY.�I,�d�:nsi9Rqau�kF2��1{=6��<�.�XԔ�l��`� ]c:�p����V�˸�뻿�wx�~��&ִ�=���.�q�\�W��%��+,������^���T���m���&�[:�}������ܠ�t��mBe��P[h�%ـ~�;מ����|ݘ�n��;�_Lڤ�guD5��2;��m���{��ڄݶ 3)�@gA
�F�<#���ܷs@�즁���^�UR��sv`�m�B�8�$�������8�V�W-z9n�ކ�� ��d,Dq`��j�pu��!譖wbιҦ���6���6�p�K�I��r8�ZW-z9n�s��4���PƄ,q�����Ս�ȏG�"��HV҄=� 3)��w+����X��܏@�-��1�3�]Ҁs�Ԁ�u�\�,#DI&h���9�j�:�k�9�w4�W�Y����!�s��@t{އ[�_�ܡ�m���\�l�����m�p���1�u�)�*7Rj�u��9�:�<���c�\�*�1�8� 3P�Ƕ�e7+����C��!xj7��Oq�ｹ�r�S@��@��@��*b�H�Yj���@c�b2��L,�������?��:TRV������`����>����bo#I��qHh�h\��廚�]��K|��X�I#ur�����ڄ=� 3)�@d>��~h�T����VS�����v��.��A.�e�h'�q�]r>��I�Q�9V���@c�b2���A��R�����$�4^�o��ϳ7k�Pw����@l���
�5�m�h�h\��廚/gL �SC]�����v���U*}�ݘ9�� ��_L
�T�UU%>��$C 41z� ���ﮤ���BcQ�L�O#�9�w4ײ�8�ZW;^�yV%+HmȰQcY�5�t�3�bw.�S�f)�λ�K���svwn��I��$m��x����즁�;V���^��[��~�k��4�M7sv 3)�@l�@f6���b�z1 ��PƒŎ4��6��*������ 3+\�2l�j\]�uRQ3Wt��mB5�ݶ �G��.��=���!�#D�4V� ;��k��r���ڄB���B$P|� �y�SݥĔ��1i��t�!�K�3�(�.�@��1�����{�9��p�5�9yV��Q����n�ؘ�6�yz���h�����e�s���t:ۓ��tn��ʽKѰ�ۈ��chw@O1�e]��R���]��Z3s7i٤.������Q���n��V�nN^а�\=	-�T��� I�b���A�{d��R\�Kף,��/���;�||���Dx�<�Zm����]Zs�ey�������]�ݺ��y����a4x�0�MaNg����4�������UU%�n�, �Mmj���ɹ�������mBj�l���(5��O��?v��j�l@l�@}��1D�.�nj�����mB7m���H;ӏ���i�1lPO#I�6�s4w����H������.���oi�kx��Lt'H�M��ꇞLFm�d�c]����ņ-Ɍs c��������7T 7v���2�@lN?MK�./)��9Ƥ��{�]EO�!� ֧;��X;��~|�fmU*�����l��˩,(����r�n�:� >�w4�S�V`�&���3@�{(�������{ӽ�� �&;�����ݻ� ��{0���������{s@�{)�qpI.��G��O#X�"��ّ���fr�5��܆��K�y�̳IeL��X܄O��?v������짳�
���_xK�H�n8Ɗ��6� 3v؀�������N֖��4�Cm�3@�{)�qv�jw_*��>]?i�Q�� "�!.x�rIa32��r�1L�����p��i�A�0�Du0G$:�%�ʆ0�k��B(�їJ2��
H�b"�b�6�@���lq��Zɸ@rq+�I���FĂB<�"FL#�!� c�@�!p�#��B2�E!a�hN�e�&M�o0���2!�H� 5�0Wp� it�pT��!�HaS�)�Ӡ>�8v���\\���[�ww w�ۖ+c�������:� >�� 3[P��T�;�� ���N=VZ�R&���>�� 1�����ηHpC"�l���6.�s�=إN��1p�ف�8���8�U
*]3����O,�Ʊ&��HcmB7m��n��}�{��O3�5�m9�;�M����m��9m��q`��q�� ��Hh:� >�� 1���m� i�����$Q<�@����������f��� @���pB"Ab#^��B�)����Ҥ�U�J�����L����x˹$�.�������m��n�f�m����d2lʖ�,uk'I�B��QS��Q\��p�G���Ν�<���(Qa�&�J������w�g[�٭G}!��nh��E�Y �	$4���i*�����X�w��_L�٩�RM{!27���z;}��^۹�~�e4
�k�9{w臄h�$����z'�wЀ�w�ηH�Z�U��+0pX�XDә�~�e4
�{0�s���ŀ?Ԫ��֚*���=�?w�	�R�dv#[y�z�B�:�N��=m4n�l�F��{cLgj ��vC���}�6]�tl����/�G���bZ���.���s�8N�H��qz��=݋�
�b��A�׷Kvvpz�qQ֝��Ě�8n�q�J�EY#gs�������G\w%%���:�a��sA�9rm�G]��E�%�MI���"'�:�PeB���R���#�%Hu��|�9n�-D_��-�b�^�k�Zh�P�2�b.-��{WJ\󶃱�c�\�;��wvh���L���,��q��_~A���@<_{(59&(���kP�xڄٶ���K�#�&;�=iH�N9���4w���?s��]�z�v�h�����<�'������b��٭B�j{� �H5��I����;w4�w4�즁y�����50w[s�B�n�vyY]&��6l�Kl�sr]���bS152#x��I������/-��?u�������~�xF��9�MI;�wF� �O�(=8{��]�)@9z���P��{5�t@��&��nf����h^נ~�n�on�[���I7"�*z���P�oZ��Z��0ۂI��X䈏�����-���?u������5*T�v��Dq�li��P�N^C�R���:�.��u�"{v��,q�#B�A�93�������h^נ~�n��Z��$�&ۈmB���ֹ@9z���P�oZ�� �� �H5����U�z���5<�; b��DO�70����7�A�9��9�RO�c���..w15r#x��I������-���?u�� �-�on���l�˻�@c֡���;}? =�ۯs@�r���A�ƅC���1]�W���Mu���`��wh���޶������S�Up��k\�����P�ǭf�[���I7"��٠}�� 1�P��k\���$�T��]�G�G&���M��s@�v� �-��v����#II����sI>�;۩$���u&�
+樟j��Q��*!�U����{5!���h�D�q�G3@�v��朗��v|{���;�XҥK��Ư]^wc�	�n�g���l��őU�� �]�ৱ�����Q���Y;��͍����؀�[Q�HoWt�:'\D����,o"�=����۹�r�V���׾ϳ3/��臄x�d%Ո}��Gz=靖�������t��쉸�l���T�6�Z {�h�l@c֡�a��ISwd��Sw(q�@}�� 1�P����n��Z �=10J�1�����6��k�#�GRi�n�"ײ�������v�^8�̡�qڔ]=�7K���"\æ�y�l�-Μ�]�M��l�!��M����0�����k�(�1v֝�1����1�Y�R��6M�Ӟ1v�[sѭ���=f�m�P�+l9��tU��=�:������j�+�h�m;g\m��[�!dr\��vK8jW��*�{�����w���;���}ߟ���N�n����N޻*��N9Yb��m�v����]�#^�WGgx�����&n���ܡ����� �m��ږ��$hRB6��4[vmk��ݠ7]��9��aQr�qₓ4Wj��٠w�S@�s@-�8A,K$"�`܋@;������tܠ6'DԸ�do7�NM����[��r�V�s��@�>��3ϧ��i������JӜ�H������dS lt����moh��xCfoDL#� 9#��9�{s@�v� �;f���M����Y��#i��'��{u��j*< D��1�R��C4��@��T��%�R�������=��߻�X���I�h9�4��h��h�ՠ��tTx�9&)QSuv��v�6� 1�r�7[��ږ��#i) �	!�r۹�r���9���v�`�I%����f��6��cLvwā�K�OMdcq#���4tu�A��Ɛ$�zc/+�6�ή�@��u��P�t��ı�,ȴ��h��9m��9]�@������L����iɠs��f��w�ѩ�81!/*��̙7�������[-�E�]�X��ڄ:nP�v��u�h���Y�D�	��?u�� �n�n�m�@~��ޘ�eQR���?����n�����ko��75�<VKg��z:R�=m��c�\�*�(��o������P��ڄ�Z� }�i,��Xܙǎ94���ڑ�n����h{l�?vԵ(�6������q���ֹC��h�Z���n�@�&ۈo��~��Z��4��ѩ1��y B������P�(w�g�5$��q�ffZY���	���P�v��u�@cmB�Nu��T���_�q��n2�I%����ҍ����8,Lꃗ%T:���ۄ.W��o
�	��X�9?�}��r۹�~��^Ͽ -���{�o��l��$�jzd�O� 7�h�Z��'K1P=��$�	��9]���٠w�S@�s@�q��q�� �C��Aމ��� �_m�@c�� s��Q�p����{e4	���ܓ��fd����I�T U�� ��� U� ��@W�* *��PU�Ҡ���TA_��@ *(��"�X�,F��"Ŋ"���(��","���"��"*�"���, ���"��"� � ���AT�T U�( ���@Wʀ
�T Uv� *��PU�J�
��T UȠ��� _� ��� ����d�Mf�5�L��f�A@��̟\���      �`�� P   "�$  ��@(<*HT!@    *�  
�Q ��JH� ��A UH��*% � H 
�    �  � ��� ��)J\��R���(�iJ)e��\���JY;��x��qez�紫��������{5<��   q�w6�뗭��t=3��w�}<}}:=j���͹�Um��ܩ�r�ז^^^m�{w�J�x�}�   P S� S�J���ޯ3w�]�Ҽ������|����]������j^���kT� mSldʺ��N m�U]�� ǡ�oZW6��u�Խ��{j�����ҷ7U�n-_^�}�ק9��� ��T  �  ��K��e�9���{�ݫ��/r��B�G�����f��t�iy�ڝ^���}J����  �}��ϛ{�r��w� O*����/;W�95;9rW��>���U�T��yo������mx �@ P
 (c� ����R���շ6�mqwM�z S�����}�y���,�f�+�P�>���Z�6� ��6��ܲ��}�Rͽ����W�v����ү<z {�.O�+�n�o����[�z��x �P(   � ��J��ZW{��5���=�(p �Δ����QJY�:)��4�
^�:R�`:��Q������Ξ� ��唥
Y�� ΔҎ&��G�
R���M:�=P4�Ҕ��(LM(����F&�� ��)��R   ���6�*Pd ѡ��=U)S$�P a "{J�i5J&@ j~����)P  ��M�L��w��+�W�M_��mJ�wwu�����rr��IAE\��p(
��

*��U���
��4PN�<�!!�,c! HB#�+ �Z�#�B$ Ȑ�	?��N#R"I�B͇�+I
	#��À�\,$,HA)h�J�BE ��"�G��j�#L)��(a`�5�
	\��j�8!X�`Q2"a!3+|��2$B5`�D�jH�ɦX&@�H���,L�I$Jk��su������,������:6�%i��& H6�0$$��pa�b��_���		�K��
\�?oGC	B.30D�Z�@�`b\a�o�鲗�\SK'�H� R5 Q�@q	�)���C_K7�y��!�pd�LB4!A����3�Ipd�,�S!n���-Z��)�#�����W�:���1�$�5"P�BHIF)%YF�P���0bH�&��hb$�2 ъD�1bG#
�A�a�+�K)-~Ӊ�-�4LZ3n�J�"�JT�n�1��D�h`2A(R���4cI"a�Vb����5. �/�`�!P$$�	 "20Ŭ�ə�&�	�9K�@�`2� ��$� @!���d#�F��0�W0��)�$��gl5����H��
S�/(m��~Hs�}p\c��k�J8�)�"���jl��s$!�!
�H&d+
0"���\�/F�a:��S���D�`c`ܻ��/	N��$Ca ,b0b��.$$D X�	� �:�7��B����%0a�0��+�9�H��@X�	 ����$K#�F\!�H�	i�4�dBH@�B����$�LBc	�@���:㯳&��o&�	y
q/>'��q��\�*BƄ`@
�Z	�t�{y��`�La�q
bSƐ`��P�d7�g�4�=�<�Y`HRFH�h@a�qfLy��[��jSŀ*��b[3���x%.}c>ί��8�}������wj�V;;��:��w�\/��4+4cf�0ه.���vo;+��v�$���a,�P�5 `�����0&���s�Rı:���M}�ƨƱ���B%֙�M�Bm%̦�ܝ���P�H�~!su2X\�s>x��δ�` @��"FD�.B�܇8�1h���H1Ry�����+)�6h	����ۄ��$HE�RHI�H��@&�8ˏ����N �bA��B=��%�B�pBi8�	�b�T$_��>�I5�vf7��Ա6PԘ�oJ)�C��@��f��1��f3��a!�b�4�N0j2|X�DBKW0NuO�ɂ�j�:_&�2gt٭]ld�d�a<pfI0$�L��F�U��"0�I�\�������)���q�!
����M`40Y B!�L�Cu]�HP¡5�s���z��vt�'�$&���4�aap`�p1(bcw1B���0`��3�8"�&%�0T�iɍe0�4�6ĄB@�2,+�,0)�r1*A��T�Ha���3��daXH�@�,HpI>�ìV_��j�#\$ �bXA�i�$�X�S��Lf���e0R�ØBHā!G.R2H0$X�0ϭ�!mוO�
󢘌Jw$ƞ}��~_��W���XP!V� ��_k]�$�L�ԍX���˙�fC��}�S D�lH��1dX�X�	 �
!Xg��.22�0��� B��)(`��&儎� �dB) 0�N`����!$ �0�
�$l��@g�%;��4���;4t���B�i�%C�3M+�o�;��60�5!Y �@���"B:~S
���9�B>��`H0P*�!D�H����%�/��w3�}��S����b��g4�@ �73�Q� ����%�>-�vƄ#���P�H
E�t��FGa��)P�
B�I	 ���w��K���0m�x%�0�O�\��Fd�1��ƌk"F"M�$��L����X�HBB! @�nx����H��Y)$"BI����"l`bQ� ��+da	)8�� d"P@���!\�%"4Hb�H��#\,e\!0����7(B�!�!pdcH��\���S ��iw�E�`0���22W���D$�D";$b�~�s�A`G$�"�"�JF��@�-H�X@�0���ֈk?|jA�2p�6AԀ�Ø�Nq����%� H#����$�!D�q������|<����R	�ԇ��Ć��8���+!�Ks��`%�a��q	0����%H�"��HP�0F
Q��*	�MN ���!�5����/��������f���8��5��	~�RM�589&��a�b�[�>J�he%cR���X�cX	#R0��2B]�<SP1��r�0�չY%e U�R"��mɋ�������@cv�t0`@HT�\$.&��l�hPw���ݪ���G� 8�%h��檸����� �bňI8�S�2pe1���C:7ψ`�#2�� � � �AB0N!(Jl�1��!X�e6F�#���rXi%0�*J���R4��Ѓt�>7uu�� �k����Y8��%L@m Q"K�%8"�`����A���&3�����˧g4��);a5��l̺��Mˮa�2��$��!H���,�-�#򒐿|L�>ɒH��mC2F;0���2�hƬ��2m�0� ��B�H�D:�d�'؄7��`a#��10�X�aG��\��B����{�a�	3��l����
�5�����v8��RS.P�$�`�d���~�S�FeHP�R!����*Fg���%%��d4aXu�YS�У���q�cI��)���-.H��s�H��PH��=�&y#�f�2JYI�s��6i>�	>!@��hF>)2QB�Uʕ���7���d%!hF,�b���5O�� ��� BH�����#���0�!B����(H��),������:��-M����o:LI H����6��2�)��6@�RX���H����H`�wxc��H$H��� d���\'1�Bc:�5�ݐ� b#Qi��1Ef�:!�F� 8�q!pp�'8&��\-��*�LfFG1l��B5�Ɣ�I65b��fD!c	�InaK_��Λ���c�*K����	��F�G'	��VVc�0�"B4��[�BHBaL�8H\l�j]��XNs�\ޱ����j1(}^gY��nϋ	x	L`C+l�F�&2�3���9~�~2B�!�`A*+)�\]l�6c$H�V2bޓ�B!
�����2�HH = T�X�����'9V���$~�7��f�3#�F�:�]�>`Cf�T#^�2@����u��@$b���@��FBSQ���83�m"P�[!C0!����� �
���7�w���8l ��8    � �   e�[@im8�?�m����n�kn��e���lJ���5�S���V2-V�b�e����n���:ʶJ���һ���l��)
m���v�i[ 4\rF�Hl�րlm���I��mI5V ڶ$D���m��[Aa����m��m  �V�d�mݶD��m�6�� $�`
�X��h*N��/5HM@`�ejBj��_� -�t͛d� A�j�K�k5��ie��0RD�U�/R�I�8�G ��U+.�l�UPj�;��x���m�T�(u�N���cX52@[%6�+I�J�` �A��a�]ݘ
��@��V���6ݭ��ͬ�  ���ml���t mz݀49�m ]ێ�m¹"M��s@WU��m*�Wd]�T��_'ݮ��X�h�s-!)q��������u�R5N�Z�U�\�L�R��Ke�l�� ��t�� ���Im��6�h'�|@� 6�� �h 6�am�m�m!m  ����A�[*4���w) ��UV��4�Kn�������(96��� ��ඖ�l$�` �5��o^�n���`m�6뮮�H 6�m�ic�����g  �$ ��\�@l�ڤ�Z��u�x ֤�   ��$	29m� �	��v�[��Y5�	 w\�t�m� ����b�@�H-��H�\,=��h;n�Hm�im�6� H/[��km��s��  � �	�E��6Zm�6ۛl�koH  m�Vl@ �$pm:�L HvҲ��ˀm�m�f��"K�ŲP	��}�� -� ��h�� �,0 6ݶ� ��K:�kVe͖ip�@�J ��v  &�ۚ�$���@ �ڐp$�lq��N�h�ݫ`m 6؛\m��  m�	i�  �:�m#lk6�Jp^�� m�Zl&�h�M� u��	 �`    6���@  ���m��I�6݀  ��6Ú��R�  �`�m�P���� �ձEזXF�Սh 8m���mI[  jh�a �l�6�f� ��}d��� [@��}mm�e� jE����@�uɳU@UP P��l+OdݬT=��k-��tab,���s�L�4p: �svZ'D�  6�m�lVҭv�m*�H�P:�� m�հ v,�V�PN���
9Z��j�����R(pr�Kӓ��l����M�  ^�[@ [@�nH�Y��l �nm��5�A��ِ�e��D�m� v�ֲCm�[Al�հs�ZXmjL��	�\[Kh8$6�-�qm8  m�m��a���l �  [Ki�ְ   !��[&�� �m� �q�lm�4Q���k���I� �`6�n�` ��%p�v��]��qm  �l�����l6�m�m�m�lH[p  Ѷ�� �i ���Ͷp $��p$��&�m�  mڶ�m��V�,�մ  |߀ �z��U���%�P@�   �x���ivG��j�`��h�m�m� &՛`�l�b޲h  6� j@s�  kn�Lp m� ��5鲶�m ��� ��E�Ӕ����`*�����ibt����P M�km���6ؽ��ն��� 6��kmT�,ݪ�b�M<�5]J[+(ն܀�cl�*]�iT)T=���[]��[{[w  ��n,v�4��үju!��\vݦi[v��v�M��3l��-�n�`u*@�m���M�kC]2F�Mmm� �i����$  8[E�Մ��-��m rE�-� ڶ Bėl/@�.�UV�-����č
n�#j�]Z�Q�kY��1 ]�ŊN%]����e��z��KqS�U�b�H�k2g����m�$֋  Hv�6�[I p  �k� � p�,��`-�� -���    Hm���@   l �l ��Cm�p��m��� 	�� m�m��` lm�#��#���&��v �@�m[~-�m � �H@H���0psm�lm���  m�l h�`  �`   ���M���\b@V��Wf�m���۰l�m!�[@ �  -�e��N�6ؐ �mH �]�I��� $	$��-� �`��l�%�:)�U�����$�{nm���v i�l�6��w m&��%F�u�5n��-�U)r�ƒ��v�Ӳ�;Q!� ��p�zr�m�ۭl�!z���cm�1e�u�	-V��N ;2��T����	�(۰[IkW�-,b 
WWh8j�
�ʵU�G�:��A��А��fm���ڹ��� E�6�I]��u˪��d��`�(8��$�mP<��G���]ձ���UU��p[mP ]�6��m�۶�"hl`�F⺀U�v�ٹ��������IoP��km� ����	 ��H7e��H >]+o� ��6��ͫv �[��m�kn���� $[C�	    H��\�l��YR[��l�t�!����Hi:n�l�m��6^�&�&Y��*�J�v���U�=m����Cf�8�ԫKe�2P�N1� �[�R��� K��pɵ��8([n��Z��^�7n�ѶŴ �$����mm�-�R���[WJ���ȁ@�q6a��m�  h  6�u����m����$���z�6�o�f��   �]$���[@HK��2��MUUT9lh�������VeP�j��kj�p�;�-@=��  �N��%Z۷imHS�5Z��J�1[=��� d��q]J�v��quQ�M��
{A�ī@UU�Y.&f�]U��;��u} J��q��[`[D�Vֹ�  h���엉2�*�h qa��q�m6�]�z��q  i�Ui%� "�@ h���ٶ��Z�X�����Ό�M��	%�䑦� ݥ�:m���͔�I,�߻TP����.���n Y��-^��m� �m��9&�� [�]J��y@C�m��� H�x[MwN�� �i��Ҭ�+�xh
U�Y��'a�L�nH��pKn��g�E�gI&�rBA��Xamm�۳0��6|�B�A:���P6�z�-�p��-�خ{T�=@�2�mljhx�S�������8�^�2�Vq컙��۶`*�c^� �`l$��'=qJ�Uմ�U�����x��@e���i;q5P���[�`Z�H-�M+|��f�m���\�[��:R	Q�暀	� �T�^�'��`��ڪU�Tb�hJyi�Tq;n�m�B'���m*�Mk���� ^��-�� �2�&�m��qe�    �5(��b�A� Z�� ��;m�-�hm�.�3�0 ���ָ6ۄKN�D��A��lI��km�-�@j�I[TJdm\���m�5��U�%QY��t(�e�ӫ��� 3ӆ�  $��V��5��[oZI�bM�� ��;EH$彭Ą�6�kf� �8 [F����nz�/���\�� �-��J�,��H�m�6�a%��޶�@m��n�`��m�kd` ��H-��p $vG6�ˆ8	 �$K�P�*��V��� "��uUT���T��W��m�"�6�  h�р[BFN/,6�&�L	lv�n�:�V� -� �hZ%��M�SI� �iw9.��[lH���Hh�l �t�� I m [Ɛ���p���gN�N�O��m�}�π�^�VH��ۤ�x� �m�*e���v��Z�V�c��jR_*�F�
Iϐ�e�����A���MM�mjf��fZI!"N $ ��a�HH�6ۍUf� ��Z86�� [RK�np�sn�m�h�K##i�"��lɮ�&#&�p�Y-��is�J�6�<�`pt��d��ݓN���m-���nݺ� ���K�bU�j1��ݶl�6�j��ШqsØ�$q�kd�6^�e� 
[A�[B��Ͷݳf� t��[m�$  -�p[_��%�}m��b���ll���m�'I-�   �Xcm� hͷ� �Ӡ6�H �� $$    $ �h$q�hi�-��KJ^���[�I(q'-��`���H �`�`ٷ`��[n� i�� [V�t�i�j�(LE�VQR3Kmo:�m��� m�9�d��
�)��.�~'�UL'� �`�|�4r����81QO�]���L�P�1	�@�K@1�$(���QUPJD��
�"l:�:`�RE]�H�������
.���5A^�X��� T��@���������S=���8$U;8�ހ|����_��P�<I$�EM	/DC�Q�Q�����P�c���"�EG �+	�?* ��G��8�@:��Q:��k�ܢ�eb�#)�xw�28@b iS��8��q� �D�L
�
��P�dP�\�Qx�ARA@h�o|uT�0��G��|"� ��+�&V:A�Ǡa &
�~��p�qڈ�P�� ���~G�U�4`.�r�)���Q>
������G5#�W��D����O�N�#�.b
�(0A��00�|�E��\4��CW*��b/C	�@��$`D"�$VA4
t ��(�U{�8����,�V�$� � Y��~EN!v&Pt��!�����j.����q��2'T�&�P��� �S(n!����i�a> 6}�O����� �r$��h`B��%��IEĔ�I�ʪ��m��m���7i L㶝��mf۷^jh��py���9Ȍ�g���ʑ�u�kxm��0Jh��.T�Y�nd6���;v�Xɷ:�T�2��Y��@n92,r�e��2m��eB;e�L#�g�9��tra�3��Fu��+)Z�q�5����s��5����p���d�Km�vV�ZNnٺ^WIZ�k0� ��*�*��5��YX)weS�
MgR�@P�\�I�yU�j�v@C8jԶ�p2ֶjܳ ]{i��]=fv�ݕ�۶���Mk0��$�v�R�1umή`W�v�8xU�^�-�a���:]��UN�q�74�Y����rܦ�%�a�x[m�T�U���d�벹t;m̪t�` -Zl�ꁮ(U�$:,����nxK٬�m ��hm�n����f�v&�<�;9y�l#�Fm� ��uU�*�K�ne�'���R���ΐz�-`���X(cU)�.�b���<$A�g���LJ��HJK6q�6[0�U{6�D��	�C���@�{yI�ı/�ML���ƫ,Va�_hk�ku-TL���k�Y�G�#m��rr֭(p��v6m�a��ZBz��R��,�ը�Ҷ�#ʑ=+��n��^s�V2��U.UYV:lX��P)W��#���֣�`��/mv'PJV�ZH����a m��Tݩ�^	p*L��6) �3vV��*�t�<�m��N�ݸ�֣n�}�A�FK�61�:N9�ѭm�5���u�(JulwcTL��N�a# Ȗn�I����H^N.�9��v{v�k˛D�n�	Av��5v�<¼��d���+)pt�GT��$�#y͘	&�Mo[,6i�i��N\� I3l6p(�
C��.���M8f�C6�p�����Ƅ�]"����t��+WR�WoE���x�+(�i�ج�a��W���W4Y@=�;f��X&iZ�)ƸB�f���s���U��"9߁]�T ��G�꣥�����DS��0� *�Q�ګ�AH@^�6�䋩U�5D�,!�%��j���9ч�&X�w
�v�Rq
���T���f[�8��s8���Su\�Wg���p��\�7Pv�s.�K�T"��$쩡��NAr�[��r��m	���`;9��p�n5�1ӡ'bv�r��5�q�7=AD�D˧s�4s��IF�M���Ns�:�-��n��*��/jY��\�t�(���@�ṫf,�ø���=����^�p��8�p�8�!ƅ  zJƨ�����F�d���X�A7o9��Vz&"X�'�﷤��g8���#�$b	mlT����Kı/>�s��Kı>��q��Kı7�wzMı,K�L�e4q3��L���'�8�l�Ie���X�%��/{�&�X�%����n%�bX?rg�)��%�b^}��I���L�gv�m�F�Ukj�d��Kı7�wzMı,K�L�e5ı,KϹ��7ı,N�8���L�g�u�O���:�+e�/�X�%��f{2��bX�%���t��bX�'y�v��Kı7�wzM�3��L��M�l82q�������W��J���jn9�V z^y�ƻm=��8��h�7B�eeP#%/L�g8�~����ı,N�8��%�bo�����bX�'g�a5ı,Nv�ɔ�t�;I-�/�8���-��C(�Cɑ������&%G�D�K����Mı,Kӆ{0��bX�%���t��bX�Ӷ�1�N���[�É�L�g�ל_��,K��{0��c��"b%�;��7ı,Ow8����%�bo'!����!e�8�L�g8��0����"b%�{��:Mı,K��=jj%�`yFb'��}t��bY��'�l�#-��n���&q8�%���t��bX�'y�v��Kı7��I��%�bw�g�	��#8����ק�+�BR��9X��c��CE���L�E�z��[/L�w/�7β��juu-�),���_L�g8��y�,8��%��睺Mı,K��=�MD�,K��w:Mı,K�͝�qLSd�l��g�5ı,M�<��n%�bX����j%�bX��s��n%�bX��q�SQ=���bs���1���-c���ל_�&q3��^�_�Q,Kļ��Γq,j䂑P"���"�����q�SQ,K�/��^q~8���&qw��D�++��qf30��bX�%���t��bX�'y�v��Kı;�w��n%�b�Že�qa��&q3�~w�9]&q)�˜�I��%�bw��mMD�,K��{�&�X�%���=�MD�,K���t��bX�'y-&{1nr\�L���Z��^^�f�W�0�Ij�[sz��tQ�m��=�:����}���,N��4��bX�'yf{0��bX�%�;��7ı,N�8��#8���j;$�E�%����g�bw�g�	�y�&"X������Kı=��֦�X�%��s�Ɠs��L�g�]��H�Kcb��qdKı/y��I��%�bw��mMD��1=����n%�bX����É�L�g����Y,�),�s�&�X�%��g�5ı,N��4��bX�'g�a5İ:(>H-؉O&Gq7�k��n%8���/�Y�c�P*��0��Ň�bX��;�i7ı,N���j%�bX���s��Kı;�㶦����&q>�|aݵE�qRXu���,n4�v.�n��0q�뷷V�
�>���TZ�YK-�8�L�g8��N,ı,K�w��n%�bX���o�6��}�o|�C���J`쉁;�[^Ɍ	�J�T�NV��V�ۀo�u���0�o۪��o�p���G\A,/
�`z��痽lIK� �"`K��5騑1Z�G%x��������1�͊�s�������W7�p�nf�	&�q\=e�ٗC19Y�c���tۧ��Vk֞ nWh&��t��^zm���34���-��j��
���L�!�Ϧ/��{3Y�[( ��v��wA�}��OK�K-l���-;P�Vg�#�r׵��q�`�<�ݖ2�99Ѷt��XmLO[zMk��������qy�٫��[��:�.����Jv�ř12L�8�9��]� "�N
��)�<e�wE�[��u��R/*q��(��ul�:�������n�8ݭe$@M�`N����ݥ���F�dT�X���p�n��M��^����ؘ�fŗYu��+/,+`sb�n҃ ��L	ٺ����R:�[t)\��ޫ� �D���-�&Il�-UܬR�b��+�$�09{�d���ޫ���%ϗw�n��;mV:�%v���l���ܐ0a�ճ^^̝"b:��^و�"���Ӕj������7f��?w�������{� ����u���3��RN��׸�$�1�냢p(�*d�	�3z��T�@�٠>{��Ը�y��"b�!d$��n�� $�09{�d��:B},̲��!ح0=Ēo�������7f��?w��o��D���K�[n�ݘ��$�7iA�I"`m�ۺ�~sh�q��`�u�u���[NZLN%��׍��D�㗜F�99��0�4��&Iln҃ �D����`w�2���ZۡJ� ��K� n����v`�n���Q��b��ԣ%(��h뼚�S�Ha+�L���N2lL��EO��#1��1�J�T�n*գ���ݸ�ۦ�I�x��n�u���%��c����t�-�n�L�D��6`,Ol�p�������}#s���L���tn�V��7nT��^õ�۰���շ2E[����޶��0��HO��1X1�+��ݹ����w���>�_z���>��"�EK%�K�$�;$LlP`n�Il��0>�k66�P*��:Kn��t�;�;۩$���u&�@z$@eE�T���k�s7.l�?w^���T�mТ&$�.�f=����3g�-�v(�'L�6�9h����#�[X�H��0�s=d�Kl�d��+�+��ܡ�Ms��Uv�.�+`݉�ےc��n���Zڪ*r�j��p���6(07k$��ؘ��ں�1X��c���-�wv&绳 5uhIZ
X붘z�v������1��J�T�2�Kcb+V׀�v�K��{ޟ���Ϧ���v�I�O�*��p����;�JPĥ��tfΫ�:���mӥ��=e�2TI�M��6:�����a����u��v�L[3=]�!�����+u�t k��[c�b�5^�VW���_���c`��v�YV��I�ד-��V[M�I7"	ȇaJA��ELr�H�l�0�%2�*u���;���u�6�EH�8WNvģxs�k5������l�2��L���� ��U����!�`!�%&;C��3ĸ������М���Μ�ӚO@��g���9�K<�U��~�c�(07k6[ �ؘ�A.��և�ـ~ݺ`�׀�v������̵��
�
*�0�-�n�L\��A�7EYf�X���Q�׀k�ـn��7����M׀}�ֶ������`�Lܓse�7k$�쎘�q�L�ߞ;N�8]HIiDvT.A�M�9R,mq��Є�<%�^�2ǢI��se�7k$�쎿UW�\�7��`�j�9-,v�^ީ���>G�0V�!��Nޓ��Ln����-�/J�d���1,�)�[vGL�D���-�ީ�x�{���R�b�9*��"`M͖�ݬ�l	�09��]�'�KZt��{;� �T�~�ŀ�v��_{��'�-�V�AP֩���ڋJ�7 ���t#,�ؠ�^�g��@2I,�ڜ*j�W��7� ߷q`���{;� ���3T,VVX",�l	�?UU�����L���f�~I.%����5�*r�j�ʰ�{�ԓ��;u8d�N��	#���gvl�!b�m]���� ���`� ~@��8i08P�}U5�Pٕ1�D9�6R9Ä́T�)�d0�Z�0mt��8 �?2�[Ȼ!�ME��QW:���lVČh���@��Ak"AM�a�` BP��!#�b�� �F.%�B[�	I�nB2�b`T:��(���;�U�H�d���� |�NEځ�A�mm�ĵ��1�$(�#�x��8V���"i��@��{�|H� }�g>�)��� u;�S�A>����<�xO�h���(X(Sh+�ztB`"�d
���|�E"a��� OA�A����B��`�`�`����4 �666>���˚`�q2��1�gw���}t �666=�MzhA�lll}��f����A�A�{�΄�����������s!���9�n�������M;����*{���;����ﱩ'����I�9����<qp����]�	��^��L�2tK�m�'C����n_A��.˿��{��]�y��m�e�O.�K�{� }w�@g���9�d����;����&"aD8<J���kY�d�m�k��S����\̹�(�0�wu.�$ˏ�&b���>�S����o6���ؠ2�|�2V�N��9^�8�۫<`����|�s�2!� ��R��M
%Tb�~C�{��u$���&,����&!D�z�k�K�&d�7��u￦���@��:��#j�eMX���n�^�:���DdG��;B=�I��3l���,�����(�XIW���� �}ٌ�=U_rû<�=^���`�
� �����\�f���wԨ켚�I2J 4;��DC��Kʈx��7t�(�yJ�d��fw=��@|�����T�8����HZ`y$Uo��lԒ}��:�v���RyQP��� >��jzªY,R8ܫ ?ovh�fIt��x�'�=yJ�y?q�����Z��i�9�f�h%&,����7VP������r&�$�+۲Y�ݦ��=;�B�ݹ���Mن�Z^��nX3r���:�:"^�`y��vM�	3sN�=������1ɖ�9z3�=�L[+�U
��(ԣh�%b���|LrRѶ3f
�[jE���]"���[�tS����WsX��J�hQ�N7#p���޻��U�$�x��2f�Ŕ��q�c5O$�I�=:�;k��E��a��+��{7n�w��M���"����%�@�}��w�.��������\zy�C-d�����V07tP~����:`��`K��~�=�U������=��, ��ɣ�Ds��P�O���Tď(��`y�����w� �z]0=���,}�G�a,,�]������3.���<f�* �/&����ԅ_��}ñ���m��m�ǝ�×�f�M�A:^m�6��ڷ������eGt��swI��ה�켟�ܓz�7��0Z��<83.�RA2Pz�e4D���]�Z'�O���צ�׽ؠ.�+���rfL����:`�$�L(��T}�4��ȡ��s�.q��/���`/�Q�ȫ䶱�Im���9�q$���LwK� ��w�Iq&�����_�2V�NJ��07tP`z����ܮ w�Ɂ��v`�\]Sͳ�^kѵ�����$�i{N�z]0��Ԃ[\VEV��b촉����,X�(eVVU]���w}�� ?ov�?�#Y�e���@rLͻ&�ʔJ��Q��*���q..6|���zOy�����..q6{�TO@%��te�ϻ�}�7^�H\M4����"�X���|�A7�}��X��� :��H�]R9e��{�w^���Ҡ<���L�����o=�8�����I^���,Y�����y�6(x�Ǡ92e�hP��s��bッ�M�v[G;3�3�s�l�J�lδ�mֹ:�\m��~�u��Sk�] �ߓ�ݘ��L������z�F�j����[p����q���޸��b�>wfy��k�Jܩ�J��1,`�����鞻���`v����F�ڬ*�|dV�q����@�٠>^E�o��d��e��33$��$�%��3�W�.�_e�D��/t��T�9݉����g ;�<�����?�����YT��mq�7F�7[ske�{Mg��U[����z�M�h.K����fv���ց,ĸog����l�;���Xw}pC�S�8�]R9f��/"���&\� �ޥ@��@|�����a�{��`KkhLNS ���X��&�K�%o��@^-�(��N�&R�b���`y$����|����W8Ps&\̚/7��]Һ�:�^U����I09}ٌW�wj?�<�~��pēG�n��+��@ѻ8��4l�a���8�RZNx�φ���m[Q��h���s�6z��i ם�dg�6N�s�VR �c�rdx%�g�ơ���H�V�8vM[AU'`E�m,�����6�om:^_mLݫp��F���@�L�Y�l-�$ad]2\��8q�vH۞�qj-l�\��@�lpƃK��[Ci�ķJq�|��T� ��ʊ�AB�5X[5q���<X��ڗv̑��%��e�tCW���m��l#�z�{��]�qʹ]��o��~^��L�ؽ�r÷�����=�<����Ҋ�`����&������`�]�g�7a���Ttr�Vf*`�����f3�]�j/�����lB���-�`y�;��z{Θ��L�vc �$��x#,�j�/0;�GLwc�o�1�������������І�G0vkq���uH9S�׳�����Nui�;�3l���6̕�YiS������`r���L ��Sl*���#*�>wf��x�8���ҹ;q�Q
�������I;���jI�������[j5J��mYl�>}�L��T�����Θ{=�	���+�Uu��1,a絛�^~��L���K�O����=��p�ʝ��!j�>��*�&nI��;��[��P�2��lװvWvښ%���eT@��륹!la��ٯ���-Dܗ�u������ۯ���:9F�$��>�� �������Z̒d��^m*w	Dl�<�/��Ȯfe�&d�n�J��ޥ@~n��I���G�H�H�]R9�jI���F����ѩ���X%!Ux�����xP7���xԓ���5$��݃�	mmuʰ<����� ���09}ٌ=�_d=�`��+<�T����,/09}����=�I~t���w׬�C��DA4��*�gcu���.�]p��#�u��ϷQ�^����@rR�v��,Y�;{=�ݸ���t���ݘ�����Tԡ]D�`�|�\�z�iP{݊���W;��!�^QYY`��X��b�??�f������b�;�.�T"��*Մ��9����b��ٔ�9�W�C/U��D �T�E��k��ԓ�?L�z,,�W,�??�� �Iq/���ݮ��ߝ09}�ܓb�b�.�ߤ�}��Ҩ�3\*�8����Y����]���yo�E�"�8R1WS��7�?�`�09}�=�g��4+������ЙIV�wqg�>}�� w}�}ޛ�<�M�}�&�VUK%��T��ｌ�"g����CΘ=�X�;��mF�\��e��\�8��(���3t�T�2�&nfIE�wL����u�XJ�[n�zn,��3.d�7���nF���2h
T��C�|�O���������$Bx�������X2�"�"�,!6�,J�6�s���Bf�S:{HNT��`l"E`U �q��g84�$ީ(Nv��i���0���X11�^! C�,.�oc�0�%��;���3��[v�[j�m���:0k\���u�����Ҡ `x퍭��fӕac<,���!�!��T����:E\|�+�����$8;k��v�us��F4݊�8�r�{gZ)�j^�\%�C$l���M�F��MIE!91��u�sOK,t� v`�w�0�G�e�L��d�m�U[p˷)�˰4���[Vʽ�l�=����C���Vöƚa�H3k�B�n�l�-:��f���P�]�j��Jl,&�"�-ku ����`K�!t��jmns݋�UgYpC]W�b�Aq������+l��@*湠��\M7��@UP���3r�VX4�KU��@.L�x�P�����1\��C�X�R�wH-UpqTv�A���tv�su\���UZ�+VH��� F&퍸�ё����4���T����>V#<����V��<�u�,Jf6i�MƦ�v.���g^Hb���ࡍUR���*��$�]�����=���c�کIb����/+բ��r	Z�ge��lr���ur�ٶ��+hp݇Y nEI�l���L��k� ]C�EAQ�����c�K<��Q`UV��]�m���K��E��K���R�i��.��w&z�"���5�s3'f����n�V�0��̸e̶�d�b3֝Z��tqd'y�J�nl� eR�ҁ��/F�[�G��٭v k ��P��D�06��T�-I��#��Jv�-i���˼y��+��*��f.j�[s��l5l�V����%1UiKt(�t4�����֍����.��v��ԥ�"���j���v��gh�j�dѱ`2���q����)ږ�e�)���{/;A��1����۠�4cð*�6�[��m�s���jn�.��;�ն�;[�$Үͦ�pG@q�C��`J݇�@k�����r)e�,-���T��!ܮ��HB�@���p�^��mה��E�&(�8��f�����N��݊=A*��~N!�X7��ݲ�\\�W2�Ku��y1u���ð�4�\�t����u�3�GI������d8�bc���;�*�jWt��h�m�vK���&�9�mU�e��x�5
u��/a�V��l��
�:��`2��:��6[ݲ�k>x��Y㛚+�ݴ���bѺ��Nn���-�ԉ]:����I��m)YWnj�U����ʷQ��ɛ��0��L��L�nnk\�J���y��ɂ�3�:��O@�롗J�s���J;�S��fG"�++e�����T�/�=y���p�鴨�7]T*��*Մ�`�w^�.qqH��@^qԨ�yJ������}p&!����=�����(��h���X�{��W^��EH�]C��$�ץi@{siP�zd��/6(��{�q���ЙKL��q`�+ꩪz����;�m�e�̲�S���I������y�][�z�V��dM�Eg�g���}?�5֖y��@e�k�����a8s3.I�z�z��{�m��
A��,� ���1!�U*�db�aD�Z��"I����By�S���&���}J��Fc�3&�fM^r:"��x����w��3��@}����fN�q��>���wc�U�����U��'���L	�=l������r��'��VWGj�J��;� ����7}~t���遳,���]�,�)VY㘱�9�f�.v�Aʴ��+�n.=.xy��zt�n�VG`�� ���0�׸������s���<V��I"�b��1c��096:`ose�6��+y�@`���<8���t3�Ī�z�I9�9۩����i�< }��z�5��ذ��q6muR�b����2��7+y�|ފ���TZ�E�����*F�T)�l����]k��9\��t����`vE�V\�I,2�7n�h��\��%n��箃����@�aeU6��*�L-�V�t������LM����~��XK��`wk'��*���XR�ʰ��Şl����5�}0�׸�͝�7�Z�Z�$���������g��}~t�利0'bu�@Y�t#��q���`wǰԓ}�tjDP4~@*��+Qh@ ��{�\�AN���������ط�)$j���6If��7������p	�=l���v\w�ե��G}�}m��:9&�p&���[L0<JN����<�� H?��.Yːq���ЙIW�_oR�/�x���#Y�I|���iP��g�*���9Vߧu������2h�_7����Pe�*�d�3����HԊ� �m�W�k��`}�����8����b�7��x�ks���ʋlv�.%��|��`{}� ��u�{������;�7�Ȫ����G*�>��T$�6�w?����>�>R�%$D\� ,EQ��^L��\�4��֞��%a�ӻQx���f���l�����=�.zwer����ݞ�����6�.���m���/@W��{R�`yie�k��d��:�a�	���;ٞ�-p=��laefVmq�8h���j���q�GgpWn^ۇNs���{W4�]�{NG6z�ݵgf�fuѬ~?s+#���vݎqU���"��V�(ԵXGbrПg;�s�����n�x!7=�cx��ڷ%��ȼ�؝�iG��=��åu���6L�
�BR+U��x�O�����`w��rþ�t�����
����-��l���{.:`rlu�w��y��[����6If���LM��빹=ll�`*T61��)*�?owߧu�~����, ��\M�S��� �U~�Ǡ?��sz|g?R�>��TS�'�]��S����%rW[T�vt��H��\v�,U�s�k��v�w:���'/[Fj�Ŋ�6y09�q��c�W,7�|���71�U�����m�Os�EUʢ���}��=�GL�{�����3���8�����V++*%��Z`w�Θ��l�w.Ocw��L	g��Ga)��J�?�8�{۾x�f��c�*L��ߕ��ja��
��k�6�f0;�q��GL�w^߈�oc-Q�eE���P��>$�I�M���Nċ��u��y��i�<Vտ�}w�<.e#,���/t	?_�LI07�����k�����^$R1�G%r��̥_��2nQ�o=���@{��K<��\M���Ke�r�{7�	9y��S �T�F5��j�~����,��b�;��V6�T)�l��W�\�=��_�09$t��U}W5O[����v�du��Yf����I7�w��q����"��Q��3���w/W�����a����a�\�7T�y�ƻn�c�����T�g�5ٛ#w�m�?6�~�Ǡ-�yɒo�.����^�B��JEj����N��s�\�l�y�@]��*켥\��̙��:������� �����u�,<�K���{�m�uv-؜��V���b�S3$��}�P��Te��"P�@�A4}��}�k�cRI�{�ĊF��\� �����7[ovc��s��]�����Cܻ��fe�v����t���u�vgg
.{\d��]�ֹ��ٮ�덯�������7Z��8n���}���w�-��tcV�w�ovyS�m�����ow���mF�R��e�6޾�F5�Lc��_l�����f������{�}���{���������d��f���y������o{�fj� �;���{��_{��/���"���YH�_�6�������m��}��oo{��ۿ�{���m�'v
��nR����m��wn�m�c�ٍ�m�{f�m���sum�B` GA�4>�Nc�Nj����������\\e��6���ٞ*.z� ���XFä�rܩc�Սg�g��N
\���΋<���L�pe:9ر�#�9�gp�(�`I�0\�E�m]#�Un�K�A�6�L��k�=��˺�[��K!۳���ga'vGqA��Cײ�b��7l�ht�`M�6y6�QeYF
��Q������;�����Go��!J=x�r���fK��6^�v��������뭑�Xd��aK��8HfR�Pt#��������1�m�w�vov�{��7�+�b��g޿�6ߓZ����lr�������� ��-�s�������~�ݶ���1�%�#o�w�ĊF��IW�Ͷ������w_������^���~���~�1���~]Z��9J���w�ܾ���oo}���߹;�{��O��o��m���/�ڍP��8�,��������o��=�=����}��x�o~���������َ)��i��EYi���ĩp��]�)�7�mvxڈ|r�p �#ђep����߻��/ߛm��k��{���%�ѷ�}�cm�����JE]e#�͘ɽ�m���n��j �D��O)��{����.�m������߹;���Ĥ��S}ʣ�r�Er׍�����{��^wF5o�S�����}?l�����W����7�!�UB;k�����:�wwsvr�˻��Q[��UW�Y���_?6ޭ��nG
����Sm�{����o�����m��}��o/;���~�{��%�] �[��-F��h{:��nׇ!MŊ"rEKU�7S'�8��)V)�B�ʾ���}}^6�߮���������&Lޙw~���;����?L���(H�m��u���}}�Sm�{���Ͷ�۵����9mowؿ�j5B�H�m��n�m�������s�7����uD�"LQH�	����(d��a2�"1��Z���1�e!�*d2`M8�Q���	��@,JR���� P�J0� �$F�cFv[�1f��2a	��}���J����O���0�0�����#!�oC��D��G�&.xx�I��"�"hPٮ�AP�kc�Qȉ��.~T������)z	�8��� �¯�J&
���T����~C*�_���߫��m���ͷ��\�[U���	j���8�R{������}��x�ov�ߛo���cm����cr��*�u�ڿ~m��ݯm�qq{s�|�z�ئ6�����~m����"�lE"!n7E���#�],�B���[]N�\Dܗ�u��{�}���EF�<��������� ��tcV�{��g�C�!�f�{�?�um����O��YT��������nI9\����(���܊K�=���f\���܎'+��ʦ6���/ߛm��k�"+�9��~��ݶ����j�m��'�B�ʿ~m�.$����m�c��7�m��tcVޠ��
s{���~m�����Z)-�;k�����{����}������7�m�w=�խ����kC<�W�ք��
9P�1��nV�sЂ�[�@�bS���8Ԋ%�'n,m��+�#��e}�m�����}�w������v�.s��#o�_y���~[[���⬎�HKT��}�w������v�m��n��������{��RF������YS��*����}}^6���u���ĹĤ��ئ6���~_�6٫w�q�)Q6��ӻ�\ə����������Ԣ��������m���x�o���c���������������߹2M��j�����������{��ȚB"�_t���Y1��R['i�F)8��&'�X ���ܼ^�էĪ��ʅ���ڭ4�����?F>6]�;2��8�"8M!P�+��u�e�gn�-���\g���ܭ�n7 ���ꬹJ���彗���cJ����#��p�p���4'�����)�hP���ٵ���jݼ�a��j�1�2l��΢wS�G`�f���l�n5λ[`[<��ήq%�b�.~��ܭJg�dW����Ϗ�?`�0��Ȫ�uݜ�7���v�_��{؉~ʎ�}�� ���߹\����(�����ɜ�����X����Ϸ�"q�-)\����m���\䑿N�����׾�1�����~���$c�p~��IlP��^6���?~m���(�ә�f{w�_|������������v�T��H�~��}}�Sm�{���Ͷ�۵�o�O^�������ߦGdu:BZ�6���/ߛo�w���6���?~m���)����]6��"�8���жm�nH�������/]]8�\���{n}��z5�k:n�~�7��~k�gd�r��sc��̻�I�S��y�¬�r�En[�k�vc_s���,8��I/��Q :��ޟ���jI��b�ۻp��qX��/#��`�096:g�����������Ri$p�9]M�U��=���v�u���{���{��q�-rYi�rH�}ٌݎ��0?}�W��\ ��Z�$T����<ˌc���zl;](�tn�;tVxvy��)�ȖV����{�096:������ڽQ�WKۮY�w��X&�L�D����`J�]̅�^R�:�!-X����ۻp�Ŝ�k���TaQL��d&�
1��ɓ&�fIf����E{�J����9]U�P���X�wn��v`�w���~X��oUdr�EnT����`{�{��=�Θ$��U\I/������lh�j��h�t�i;c��yV�m�J盋�C�5��K!t#_e���g ��t����od_���\_@��L�d�ð�	��lr��c����	��`K��`vlt�8t�l��	h#�ʰ�n���ׇ�8�}�����X_�p"{mmGlXbX�}�}W"���y��GL9T&B?(�k�'{ܝŦ)�],��+�>��,�\K��{ߗ��p�w^�u�����%��
�:��艔���z���f�,��g�\o��\�V�fGdu:BZ����X~̚�/��p�ͥ@b��<Kʗ%J"ba�U _�&�3&nd�f�7cy���TٙJ�.fL�D��Х<þ#++*�1&���l�GLI0�ݸۺ<N�Z݂t$�����Ē���*��� {ٓA̗&d�7ky������'+���X��ŀ�d�qx���J��33�%����*#�I�A2�9��1��bс���]��N:#`)�n��^P���s�@I��ia�y�,��V�M۫���A�4���w�>$0�s�Z:��"bG�q������mJs�0���l�npi�-d�]v��]{p�E˶m�I7���6�[��X�iv э�v3m��!�mۭ(��Esm�`��kI�v�;���@���`:ٜfb�ˌc&n2� �Tw�����.]��>ֺ�dtuYB®^�yc�e:��v��,*�����\IY��)D�GرT ��ߓw6[����GL��p"{mmGlP��p�w^�\�L� ��@_wR�{2kY�w72Vú�P��9#vW�w��,�����ݸ{;� ��7٤���:�$v�d��ߕ ]��w�Aə$�{�*Wa���YU	]�U�}�p�l�{#�$���ܹEY�I�����{n�U�h��|�6��M+�]�B��_ø���ENIo�7f���e*�̥ɓ|�]��{��A$-�'BKk�>�wg�Rē\HI	��c2L�$�dM�J�/3&���ǮM����!
�U�*�>��� ;�?Uܙ=l�y���l���ĉt�ɉT�ə����������Kˉ����u�\�U`��(KeL	�������\��:`쉁+���͸�����|�۹�Y�T�tv't7L
���j�E=��ֳ���M۵���7|�'[1�2�b���:`N��w�&��xWѾ�$�U���#�`��,�v��`zd��;�?U�+p��X�2��c�U��p��:��s�h@����C �V��k>ލ@���,��S��H���-���d�(��3;�P��T�fM�[��Z݂t$���q`^��~ �}�ogu�w]oc-�v���~�#��bnT�ss����{eqKL�n���<V֗�xA4���	b��J��Ԩ�̚./�2o�.�iP|j� �"d�N���@�d֥�D���gu*=�J�3;���l��D��r&bf�܌נ=��Tk32nf���@��� �{V��j������q>�w�@m�Ҡ{2h!$���R���I҄�|�DS#���RN}�y��!�<�3*�3ٓ@s$ɗ&Q��>�7����)P'�wHs!�Aq�Tr�=d)���O��P �W��.{m.:�o'^�Z���YUQ����n���׀}��/.~`}�z��z<(;��(O4��*�d��Qgu* �� ��۟�.6wW�aZ�+�N��U�n�Θ$�����7}���y�iA���	bLJ��g}�٠�٠2�)Ps&Ow��c��A2M���I0�D������� ��jI�ڹ Sh�P�4IJ�	��A"�((u�N$x`�L���
�D]���4�p:C�JJB�d$�Hɬ+4�=%O��F��F1 B,H2!]%C�!�$خp�w�#����U�YA�����>>,��А�XBc8��;��W/ȚB?)����|�l� ����A�0��6l@�Bd �	��n��@*��y! �$ ���n�������[Rצ����8C�"�;Q��谻t�<�0��P9�B鲑b9�d�<<�i�.=svu��tm�ͫn��.ڱѬ�ȳ�[0��t�S��s�ܚ�wS��S�5��dt��-��ʘdt,ۇ+�e�UL�4O@4�6*��ʌ�^��̑ k�MV�T��j�d�J������hshq"vK&!s�L�\��mD�۶f�@H.i�[v�Up��r�茆�Uljdu[��slN����L�r[Z�6ޤ^�ٝ֎G[�6�P���k��W,WF�TkLp�=�`�YR�5&F��0����W���O�cS���;;m�R�H��ٮ@���.��@M��bۃ�W�1�Ҁ�t�Π�;Jk�9��P˘��](
K\v�t]��u�#d��w"�aNMڠ7
���+n�2b�TJP�Yv��[ ��Z��=^g�K����՝�t�Tc��<�T�J�E+�e�Ɔ�vD���t�e1�����RZv��D�QEM�u�T6{l܀�4�r5e�71��d�n�f;
�4�s[rv�95�����:͋�=���u�m��D��p��GřʫUgی@��*����H0+>8�40N�ݜ<Yx�;�����i��;��v*�e�v�����r�J3�n@��
�m��mŴ�}&*�*�\<ݠ�R:�. e� s�+��؍���=�9%��c��m�f^�jy�+l�6[`��q˰�)�9�$��`�����Rk��-��mtl�h�=۝�H[f�]�4�l�]�����ð�j�E���j���wp�ltT6	�����R�#s�B���hǷF{vC��*ڍR\�M@b�G'�@꧝�����`�f�'C���:������$�77dfV䋲�\k\3�ծ9�A�J�r8�L�v7/3�,�泵n���"�"p�M��X�lOZ�n�	^3�Y�5U���jW�+c�V�(&����>.s�I�8�"=z��@Qx�*@6��ڊ<z�P>��6��T~:��^�I��8&39��@f٨ho^����%�(��C�][���^��r�\�\�P�����s�H+n0Mldض���*����N8v�O:c.��R�Ì్��jmNz2��8���G=!�+�u�	hӴ;y����l��3�M6�9�Ҥ�v��̖�4�"��ӺI�������c
���Z��r0�@9iS��.q|s��_���~�Id#��8w.�2En�vư�5H(��q���ֹ�񛧪r���@�ʬ���l��}�z��fR��d�.^�3;����]�5B�`䍹V�۸�~ݸ�ٓ@e�R�I�7(��]GD�̧�S�Y�����0�D���������K��lU�X:ܲ�.&��z����{2��gn����PҞa�$�
�D�wyJ��d�ɮ�~_ }�z��n�]	e��	�Y8r�LE��/M�Ug��U[���[�&��]�7����
���:IW�;�{ o۳@�d�37�������E3� ��@fd�2��RI,I%����8�<�0;�0���2���ut�I0�D��b�=Uw��:`���>�t��X)e�%���.>��※ݥ@�d�s2w�ݚs%l;�j����Z`}�� ��}�������t�>�m����4Ln[�87ͷ��n2�Ld����F�k��Q���Yc�����V }����ݸ�d�ܓz3���WO(���/.<�#��� {ٓ\��w.�t�.�iP�̹��q6{}铕;��(������RO��tjpH���!Ȏ�1��:��ݸڻ�(�'Ubtv�\I=��ʀ.�f�=�ɠ�Ow���"65��	bLJ�{2hI���ˀn�x`w�:`	�,T�-�,z�ís�̏n��
��q�nlS�������T����5Im��ݸ�j���ת�`n�Ɂ���0<�]�)�A13@{�8W&M�gu* �� ��ۀo{V��j����Z`}�J�=�ɣ�&M�gt��<P����U�����V�w޸���ԓ﹞�IO�Ad0�'!��@d��! aX�q	ߑ[+L�:�P�t�"f���x��w�&{��GLvGL��?x��:}M��Dx�#Z�r�MlC\�S�и���/lꪏ\�6y�3`w����dt��dt�;���(�'U�t#v��n��丹�!��J�&I's3�h��(�����rB��{2� {ٓG3��Θ{�b���Z�s�%U��%X�I���vh��({2�$��w�@[ц���ӕ؂[-�>�n���+�ߗ�]�Ҡ{2hf�ɖ$�#;��[Xe魲݇;T0	׭YG^�//ix続�%\읺�ݔ�1I�W��ώ����j#��yvy�%��]i[.�p�j�Þp��!\�A�+m��N�8�Y"*U��u��F��n�C�S"��&��qXM۩8�:���F�O3�Ac��<�����ۮu���e��� r����V�v�@�[�7N84ܪ5m���X;�yŜ��8������?ɍV;�9�.�!���+r�c���lK��ݺ�ڈ|r��'[Q8Wf���{#��ȽUU\������v�zGj�%E-�U�}��, ��ɠ=�(˜+�3rd� 嫧�x��WXꥎU�����>�n�}�7�ڨ}�� ���D�5"��J�8������/�GLf��ݕ1Ю�Ux�ݦ��� �\������}���v�wgT[,U���HG��|����1K�f�.q����B+��Y�g�����n�ݣ���qX;O�}�{ w{� ���?�\_�o����{W�np����%��b{U�Ծ�ꨑ'"���ş�_��$<�0�g����v ��p	<�����dt�6lL�U2�F�Z��%��Ğ�s��}�X����t�?>��v�Ua*)h�C����U\����x`l������7m��T�X,��9�'.�U�T]���е��+�]h3r^۞��dYz#ZE��\ ��L�T5C��\���ذ��y*�IJ�vKp��� ���ٔ���k�� ���H��L����2P�<P{2�nR�3��"�j
@H��ا�1��w� �t�>К���
�V� 9� ٱ0;�Pa랏� �.��������v� ��n�ݺ`��0�۷ ��챧c�X�����P��e� e*^�7�
N[���G��+\;<ɍ�[ci��A-��}ۦ��� ?}��07��n�^���	]c��`l��Ș͉�����t�H�+��v� ?}�p�ݸ�v�w{t�5t6�RKb���专U}w=<��x`l�R}W�L�2��f_}�M��c��$yR�"&hz�
�2IrM��q�/;�Pw�p������j:4�8����wg�H����Un�.�{]>�g�';^��E��}v�.�3e�9�0����;ݾ0�OO*W\(NXY^��0�����o��]��~1zF�!*�6IV o�� ���0���۸���5�lm9]�%��e̚37�(��z�fR��d�;�� �ڽ��k,�IZ`��t&^�ߗ���@e�R�%��c$�cB�?0;�S�\Y�c96͔�M�k)$�փFyg2��](�]b8%�eZ8C���M۵�GV�][uh�q,l������V- 킭��m����ZVb0U�.��V�Ѩ�u��+vtVt�������!�v{�rFI� ��.����nݨW:� Vʛ\v�mpl��صkeN.�p%���몜�u]���M��!���)Uu��:�Ľ�Cb?~R����t�d�t�[�)���99��d�]�c�M���^��)*�FWZ)h�@��}� ;�ۀo{������7�|�]F��d�*�.+�x��l؟�='�0'�z��5���g�7�̔D���%��}���6[vGLf���!�����ff*`l͖���� ٱ0�ˏ۾���m����P�"���~�� ٱ0&�t�ٛ-���R�,Z)�n���+��zP��q4�͵ٹČG���n4KB��s����H�D%U��*��{�`M�遳6[ ��06���Mv�X�[-�7��Y���$s�/5��y�2�ڒY�d_��.�f�//n���W��X�e�I#nU�o�������]��Ɂ�t�����+.���2��I[ �ؘ͉�;���$��|�]Z���؊VY[�U�6&��l�+�Od��	݉��|����.'�/U������\�צ��P]<��=�.MҜ�M�[V�ٱt�b\�<遳6[ �ؽU���zz�"�R���Imxvw^ N�Lf���ݘ��iE�yx �!L���� ���<���I���Z��0X�,�]Er��6�b$#!�\V�(��3�	�B11'�(�F@�$'ÄM�q�
��Hĉ�)��t2��0�E�!��K(0��# 1�md�D�7�`��$`F(@��p���w�8��0�]�D�,D )f�H����D��H�a	���}m��!(}���JP�T�!C�z7:/X�U@��'�K�C
lP2�uE�Ă|�BN�P墋>QC�� ��9��ߦ��׀��������r���������;�Ɂ�6[ �v&_F��`�m���n ~��p�l���Lf���r�����*K�v�+U��{�̊�:^�e��2"&��K�N��qX�V+YeRI[����x�� ٱ0wb`sr��Y�XZřN�����y5�̝�76hכ4��WTz��lE+,�Km�;��0wb`l͖�9݉�;��tbTe+T��!�/�1��6[ �ؘt� �}TJp�� �q!
�F �D�Ni�36}�~�V�EN����;m�w6[ �ؘ5A�/�1�ݖ���bSgVw�;�{5뫷*Ln�$�GaE*��!u�&���",��*�znh�� {g�f�0vD�ٛ-�r�p��������Xw�L ����;���ﻷ?�Iq�^�D�u2[bb�H`���ٛ-�s�f�0;�j��V+YeRI[��{�=��< ���ys���Q��@^���9.���2�0���wb`l���L';�v�I�qB"����2		+�qq+�ޓ�R*�j�,
V��͊�թ���Y�c���.���0�Q{]��>�qյ���OT9n��\� 
�y�M�6ͮ�șYιr�:ƫ2Ol��0s
W>ќO2�36�u�x��,�+�&ã�g=$��n��6��*���]��l6����dֹB�ҏ+N��u�P�+7\�wWd
H.^7m� �����0v�ps];7*ݟ���{�����=���j{0	خI�p�hn�i[����ү]>�.=K7���v�_}-=Z�u�,�to�� ��v���ߘ}��,��4J7S���n� ?}y4�^=��)P�8V�K��;9t*R�$��Bb"f�ލ�>��*9�Ĺ�7��� >���oQf�\��8B�&%�5rd��{ʀ���>�����x����p#�V�� ���@rfnM���7�y��yJ�=��q
W7<dr�<�M��,�T���׎u6�x�k����z_\mՍ�+��f{i(`���ٛ-���u�������x`ov�Gb�Z�*�Jݷ ���ϱbI�3  A�&)��/�Lo���;�0ﻷ �ػ�b��Ț�ZJ�쎘5A���vy0'�z�]Fݲ[j��\�U���۞0�vhȼzL�{�*�2tD����wy��=�ɠ9�l��]�Ҡ;��`|k+�;��Q+U�HX��أOM�5c����Uy:-�#�:�׶c\�k�%v��3`l͖��dt�٪��0;���;��evB�����쎘5A�w�fl����<j�$p#�V�$� �m�}ݸ1PL#���")B ���p�n��:�&�=�T�X�0�ؘ3e�9�0�U��G�$U��V+YeRI[����x�����������ۀn�bln���O#�I]�nm�H�+q��Iļub6ݮɶ����Ee�5 � ���,�ۦ }�v���x����%��YH����P`���ٛ-������I���W�R��⮪۴��}p���쎘5A�6T�B��X�]�K1&��lvGL��ß|P��<9�����\������:�~����d(NXY^���Xw�L ����;���.q'���K%����E�suOZr�Mbʆ�q��p;�+���d����DuESd�~}�� w�fl�;#�ޕu*�T�e�H`���ٛ-�;��f�g�s��^nDԌ��	%}7� �ݪ��~�0����b}sT��"��-%l	ݎ�5A�N�Lء�j��؅�K*�>ݺ`z�h��(��*�Rf��3���<PcJ�H �1�ns��Y+�͐Ѻ-�8-Cu�n��H[���:-çU:˜:vA�F�<��ͤ��v֝��� ����pݺ�E����#n=:Uy�g0p�]�
�Y1���3�Pۋ�p�W�׊�M.��^����;qtMr�%8����Ibr���d�qd5X�*�ۘ����W����ĵ���Cہ�n+B��Gr7�e�YGO��y1<E��"B�
&��靣N�k.9[��5�<���gڭ��Ur^��	�5)N*ꭻO�wv���0��� �v�wul�6�!U���Z�݊	ݎ��A�N�O�}vn�_[kvB����`���v釸������#N����2�SUU}�^�?�<�ؠ�����>	�Oj������wk��09ݎ�����z�t��W%=��^��l���g-a��R��z�v��\�I�^p�$��nU����v/	ݎ���Lwb`N�^�E"��Ț���wq`�8���|�>�����UU6=q� �D��uA����m�Z��u֥�`�������U�vy��<�ɓ%�X�J�,��Lwb`s�:`N�t«����;���#N��B�-�?}�� �����t�'v&�ݏ�Y��/n�����>>������9jE;������6��nl�Tj�+��8Ed�����:`w�0	݉����v�l332���ay�����Lwb`rlt�߻��ϢkSڭYb�V o��u$���O�����Tb�U�P*є��Pb���hԓ|ﴰ��l��"��U$���{���ߖ�t��v:`�w*��Veaj&!:��Tz���+��/ voN���,�4]�Gm�:�
�B�-Òjr�uYUE����#pۄ[]X��{n}�I*�Uұ��b�;�� �ؘ�ƽ�����ŀw���jR:�U�\r� �^Mrd��6���J��ה�S2I�}�G��8B�d� ���X�c�~������L	��c�e��|e]�T������t�'v&�u��{�~۞��F��I"#�*��Lwc�;�09ݎ��0'���d�G��*ˏn+�@Y2ӌ�/j��WN[���#�k��d�u�P��Wx��N�Lwc���^�vy��ڼ�X�e�I)m��_w}�~�<���t�'v'�웕r�ՙXZ��N�"U��J��ה��ə;�y�}��,Wu��+��e%��V��t�'v&;��UU_�{����?1�BTE]U�*���p�wqa'~�tjI����R�Ţ��<�� ��D�F��7�;�@Z�1 º��F!�G�E��sF��� ���.L�T����
|p�N��߷ߜ��I��h��`E��1�)V�+� �L�8��B����bt�MpA�����4 h`�P�B�-����pHBMd��h7�� ��	$��^��������d0!>��M�@7!,�"J\� 4y�~D��(����$XFC
Rcj|�<+����[$���u��κL���be�2t6Q3�V۳�,n���uӊ�\`
��RX�$k9KmR��g��j��Ӯv}�kf8�:I��Y�yP�"6�	��9L�v�G���疂�C �pM��1Բ�v����x{)k(�`Pvt���og�ef̀B��wm��v*	�WQ��r�zD��O.�=򨑙v��`���^�%v�r���Yt��I��d�f2e]��wX�WfU��V�K�f�á��I��-�X�v����=�msn�j�z����69T3�eBȅ�ֳvV�q�-�H� x j���]�cZ�	-�杳����6ݢh	^.��R�O6ByT�VR�r!AWH�kU*c-:.n
K���͙u�vi�o'=BEں���+t�]�*���n�A�2�Z����Z�g�d�H�bk�	�0�u+�k��w��T� �R�ީ�Ɗ�D��&��)�`Jyj�egy�(�q�R�lp`�xP�cs�+����Ns��X$�n�ӆ�3�)7����ݗ�J�6�f�v5-�!$S�"œk�-��J�<s\q�(f������nȒs>-��w h��z�̞!����
ѥ:{iKubZ�,���:eg�j�Q����Z���np/��Zq�g2�+5]��*����F�G.�V.ݐ\%�QI�oVG�z�S��[^�'z[�"�f4+<���C�@�'�8W��Nd;k�p�ll��ۓ��t���+�Q[v�]�`w`j��@��Q
7[�&�e2/[�V2ۇ�A<�&�e�j�J˭��C��\pe��$UP
wDWV�x��d�0UU���B<!8u-h���C�E�de�.��-Ʉ��#&�n�#���rvHzM��$�[VXl!ԯ,�q=i�ٸYj�* 'CU���-i��Ի+����CR���c	���z�୶��J�����8�AgQ�'ʊe��P:**l8�=e@�Q `�|��>� Ҩݨ�~\��Ŀ~W��8ڶ*����B���i���a�q�1��
��t�5u�e�t��h��Bpj=���Jl��u�1�m=�91R�:��ts���l��Н���83�g+y�,ҩ���b�������;Fٷh"X�l;��cX{s�!����96ݭ�;4q�8��n�qۮ܍������l���K˰q�H����v
�l4u-e{u7��=��w�.$��ڈ`d�u�i�N1XCb�֑s�<J��k�e�F������ת��ݜ��%���7c���Lwc�W,l��=�k�%e�/�v�~���9ݎ�����v:`��̣- T^e�;�� �ؙ諭���:`{��X�Z��[b�ؙ[�`�b`s�0'v:`�gv{���z�����fbI���t������ŀ�v��^�X�=��t9n���鵊���N���.v�fIgkn�6k��6��@��(;�HU�w}� ��w o��������b�<���=+��U%ʵ����N}U�O���������u�o��Xwlzƥ	Quʰwb`s�0'v:`s�06J��X#J��%�����;�������w}po���K!
�M�V;������W =�Ɂ��t���u%�&/�_��t·��[,g9�-��utmr\祘�1�m���y������eWgV�aF���ߝ0	݉���u�}\���:`.�3��1KlL�ʰ~�����LM����O��fȫט�,��X�"$���=y����JS)d�d��}�r�ꯩ�s�� �"`۳b/+�y�""U2L���ߕ��Ҁ/�ہ�������<���=+��U��X�����ov&7c�&�L����퇥㗨�e:��5��0���
1��^�V#A\�)$R�qq�dx&�u1W &�&7c�&�_��d�������*�:�n���Y����{siP��T~���I�����*d��xD۵`{}� ���,?�M����>��, �wI$�B��e�n�L{�09�0߾�V��Q\��73$�����
ֹ���&&H�ov&7c�.l�7c������ڈ�|X��kl۱;��(��c��
�t��X�V�S�k���k���r��Ln�L\ٌn�^�������:���(7]`HU�~{ݙ�ə��fҠ�٠>��U�&\�4A����?�e�T�Gl�;�b��ݸq7��`?o�����BTEZ�f*`݉����˛1�����W�/w���]K��L�u!33@}w096:`sv:`݉�����it}��~�����4���7@F�9��(\�]�g��g������1���J6,�"�Wd�v��-cV�7�-�X��� ��.	�sۓ�cg�lr��՝A��ʹ�b�X;��]���4��թ5��=u���A��B'm�\9�^xY��q�WPp��vъ��wjwD�\u��t0��j�]��l�Um�K�m�Q"�ۅ�p�n	[�~z#�>N�n���>�I6ķd�3�t��*i���/]���Kk@G+D��׳�W~��J���)Pz�7���Th�$�%EC�ʰ������pn�L	ݎ��_]����<�YV%��$x�@y�@]�R�����m*�w���rZ�T�ʤ�����ŀN�t���W�W~���4۹�^VjՁ�Y���;���GLwb`w�����$����1���N4�3���^�s��g6Yճi^z�����Գy:�.��YT*��;*�}�b���p�w������M��nЕWQdɩ$���u�P!�I�or�������#��S��U�H�L�y����*9�sDgwR���n�[&Wd!B��,� ��q`�:`�&쎘(��//00�B��/0;$t�'dL�0&�ŀ�^��+l�NrGev�[�wB�s���M��'Z�v}u=덫qɨ��V�@��LvD�ݑ�n�L��X�ڵ�j�R�*�R�p�wwc�d�����:v�b/+�j�̬�T�����#�]���V�����ާ����'��jI��v��B�K����ŀ�u07dt����&m任H1Q��1S �ؘ�:`N�t�������E�M����ڪӵ��=!4�m�E������#�At��1�6�g:�:�Y�07dt�����#�;�07M.�Ia
�AeX��ş�g۵P�v�}ڨ!w���	QQy���ݎ�쉁�#�ݎ�E��mu��^2�U��%�߻�\Oy�n�L6��ﾽ�0;5T�ĩe%b�Y���07dt�����GX�n�~���enTn'�S�]��H�����!y��6�\<v��v�E�av�YY����v:`vH�N;�����,�w���,�:�Qb�d��쉁�#�ݎ�NɬjЕWQd� 7�ۀw���	�0;$t��Ɇ0Ta�U�J�ē}�}UUW'��`zO:`vH�O�n�iv�KP�"*�7��Xd��쉁�#���U[e�++�+�b9&�aգe�,6��Jm�I�m+9^e�(���<�n7ڞ��۠�6'��6Njv::E�T�[wGA�T�VY]�N��A�nv�����G.���u2�r��e`i:}X��lq� ��v�t�[0ꍎ:+[�lr)@vݞն���ym�Ս���wR�h۪`8�Br]=�i��-��Nx�bܗF�kYjӍ�¡�5��www�.��#q�Tʺ��h�0-���㪬B��DRn��˛uZ�8*�h!8��4G**�U���� ��07du����XzO:`���u��K�Q�`��p�w����>ݺg�;��KU��YT��L������Tk$��vt��٠�͝��Pv;"�U�o{���T쉁�#��ك�X�X�ի�X���#�;"`n��7c�����,��6(��V��蜸U���.X���v����
佳���vyZ�f*`�&쎘v:`vH� ���:��F��[p�w5��L) )!6�C����RM�w o۷<�8�=������xJ���Θ�:`�&쎘�-��h�Шr9V�}�~X���vGL	�046Ȭ_X��"�S ��07dt�����#��\���3Z�v�YXV�5d�L=g�i5fqup��Ɖy��]�uϴ��vy�tuRV,U��X� ��:`M��ݑ� ߷n��gf�5�X)��{����vD����+v`��W*eV;����q`��pũ%@�D$`�ut��� ߀
�dЫ�S���O���7��p�1�L0a��JT*	��c"���%���o�J�\(�A�>y-��0�&��4��a���Z��l.�MCJ��,��l&�O�FX1��UӜ�<ā0�r FBH��2BI(��"��*a>0b�b��D6#�$�����M�(��_� �^*�Up�w���Q�� �p���'Ȧ��Q�+�B�Px��"PE����C&MLɒ�����yJ�̋��92	Q��Qv�0	��#�ݎ�w�� ���:��F��[p��t������� ��0;2VU��Y��B��~�c||�lP�;+(���u�ٕ惴qS����j[*��xDU�n����� ��~�����+ҽ���G*�>�w{��w޸��b�7��Xӡ�me�-���KLvD����;�����{lr�j��U$���{�\��}�� ��jI�9����Tv����"�����}���gRO{s��2�a��̬�T�����_l��p��\�wq`�4]�Kh2��@�ֶ�F���*����ٸ�l2���]��a�-��B������q`��pl��v:`m�d�ā*2��e�C ��?W�]���Lo�遽��I6w}�&�!j�Ul����;#�z����o����&;.�X� _@�Sl��]�l����q`�iծ2"�C�J���6D����6GL�ߪ���{�v����Y.��,�V��t�kf��Zy8��5�m�A�y��\G;T,p��L�Dz�8��м�:�;]FV�_����ۭ�ˇ\���&�k��%��+*v2�b���c������q�um��@�%/�%�iI{u��*-v�OnӶ��N��C��p��qҀݣO$���=�4��{�{r%�clV�دh��pt�K=U�o{�����������\��ˣv�y�e��]�]v..Y�[y}���&�Ѩ׍Tq�����`vlt���� �쉁�{V�-V+\v�%-� �{���u� ڛ ��0&���f]`��e�u����:`]�0	��c�Wwc�X�X�#�`q7���`��`�l��}�*���K�f$�&Șf���#�����7b;�4�v'#����fvųH����U�X�v� ����N�l��h�%Yt�,I0͉�6GLjl^�X�z�o�wҲA�/�v�{��T]�EAC��C�or*�D�$ؘ͉�r�mK��E�f*`Sb`dL��Wd��`{}�Xӡ�m��+mi��-��9_Uߧ���y0&��mvD����7*uZ�,��[�ov���X�� �b`r`���˫UFz�Cm�<���k�\�a��L�m��N���r�5�Sn:[n��ŀ_n� ���%���o����J륬tn�ڰ��۞\I����������ˉ6k���jЕ[j�� �ݚ ��&����63-I/32f���� ~]���wT�[e!j�Um�0��w�<����쉀I�0?}���$�(^Gm��w ~_lLI �v&;�
we�.�/3���s���l��V�K6���K�I�cb��Y�y����Y$ BУ�J� |��\ �D�;݉�$���%�vRJ]9L�fd�&d��w�4��* ��s͛�{7*uZ�,��ۀ{�@f^R�Y3��7f�7sf���4�8@�Tێ�[��.?{}�`�=��I;�w:� �J0rSFή,���p]ݍ<��Zƫ),� 9�D�&Ș{"`M����y턞J.�!Wv�h1g
�MÖ��{XM�4�1i�vʑԓ:n4d�� �dL	�:`�"`sf�0�����m��ݸ�w s���Mؘ��]�w����VZI0'dt�9�D�W��}Wg��`����N�rF�B�G*����Mؘ{"a���ܦ���e�����-��v�}���زI7��s�'B�p�4T������"�H�A�5X��=�kZ����nX�W�����9x���&:�.�u�<OS����Y���r���������圩4���ɨ�'#��F�����[l�VC�b�.Qv�ʓ�x������X�V�4�i�g�S�`��<�>�	¶Ls������ڇ/�s�j��;��iGa1!l`���;k��T��7�����}��Kt�\ӑd;S\�K%{�����wq�H��b燍�B��i݉�MaE��l���gSդ���}q���%quel�� ����~_ z���I���l�����
�M��%����<�8�ú{ɀzO&�Ș��e��+.��Ŋ�:H�݉�w�&��� ��z�u[l%��ؘ{"`N��s���͒���U�J��I�w�&쎘:H�{ݸ��E�7juKm�������l�`[j�8'����T�M�[7�ު�nKn`���X�B��;m���b��� 7�ۀ}�p�ӫ\��+Z�Y$��w��M����
������#�ɾ�Ԓ}��:�w��~DE����z������[��z�{"`M�� �I��VKJ�RV,Y��Ę{"`M�� �I]�w� �G��J��I-�7��L�$Ln��;��_}_}+%]���Ls�ȝ���q`��fۍ���\�M $)�]>�=;A��y�q����3�$��&7b`�W,;"�/�{GQ���[�}�@?~�n�H�s���͒�!%Yt�+Ĝ�}�{�I;�{�S��PbD!��P�$ �(�J���
73�M�:�N�v����ce�(� ߷q`x̥@w�A��&w�ݚ �i�\��+Z�X��X��O۾� ���vGL���1e�Y�����a��Pp���ۊ�\�ۯf:l���^�U���фe� ��M�[��ۀ}"`M�� �I�c����+,�FbL��0&��s���M���6o�=�J��I-�=��S �I �"`쉁+��SYi*J˥b1b�Β&6D�;����1TIA�Ԉ B��q�>�}�RO��&/L�\��X$�Ę� �dL	�:`�p�׹#���LRX�D�I_,�e�\�H6 ݪ��\�!ֳt��6�ѵ�*˥IZI�w�&�0t�{�������� ����*�YxE��y��S2fwY�4��4�fM Z4��H��-v� ��p{ݬ��0'dt��ҥKXP,���e�Ln��;�vGLt�����"Z�V��$����n�~�t��I0	� ����_V��[�]Uuc/�&Ρ��.D l)b mX��d�4�F�,���Z<: �#��4����aL:>�H�O��y�J?#]8w� o
���P`�P �����&i�GB�v�Tb5����~"�4�XL��d���t�sp�������|7̙7���}�������	S3W\;Iي���hX�ô�#���{c���2r�p�P��VRU[Ѥ�&����05��V��ym۠^τ�(��m)�H[z�R�8�Lu�]�{F�vܜǁc\1H 1e�-U�NƯg��d45��ؖYk�A���H��N��6�%���2<���.N�!���2�v�Dn ��7Ѿ��dv�^��H܋*��ni��Y�eB�gE��¨��E ��f�SgY'SY��ZI��`���Y� ��K`��#8^ �7j�@j�)We��ΰa�9�n���"N�j��K.̡XL�M��
��Å�b
����U�%�b���t��`m"�hmY�aJ�&���� ����XU؇�Pګ^��A�:��X�����v�YT�!s��@�i�udq�B�%X�t4R�fw��=�ة���\\�\��b����5ݶEԳj��zU��Y3�łA��v�ɤ]S�ѩ
Y�+���U����&8!�c�k��x9U��y^us韱���r�d^Z����Lu�y0��D��l�3u����c�q�֍r��֫y #��Q:4�6�	�*��8bi0����VI0�T�g�}��6^�p�
<]�v4�J��G-�n��⼇ �DDn\�;Y���3�::�W�9�V�e�MWd�/N@9e���j�l%�9NKn�l���n! b�x��$.�7���5G.�3εj�(rL�kg\�7t��[/mL���j��Q5hj��{lj��m���6�A�3SVN�&�s']6��f�ݚM��s�n�:e��@'�c8�HJf�0J�*��z�[�r���Ij�ݒ�ī����<)�^z����GP�$�G@S�e���&ʖ��}�â��z�Δ6��Sr�fe���2�ケ���VQ�����*����yV)�@P 8�a�i�d�[�v+�ۮ�7}?|an�΁�P6(p���yEG�Z =ZA:��&�M+�U8��3�E�,����bѵ�$Bf�Z:뉹R�3�(mt��$N���zT�� ��ٞ�\��l\�V��Vx���m�l�[�t��[�g�'j�]y��:n�Ȉ���&ۉ������J82k��rg=u��c����W\��!S���gX��Om�xݬO/�����K
�X�ֈœ�X�.��++��C&�� �]��6�Z�k��xV����{���w�:����At��÷�r�W.�Ҷ�z:I��u�ey�d�2*�1[�{��,�$t�&�L	{��fe4�,���wh������݉�/vc~�ŀ~z�7���]N��9V o{ �dL�U�߷�t���6J�b�F	at�e�L��0'dt��I��{ݸَ8��Q�n;#�:H�Mؘ{"`vU��3����c��=)�4"��V%T��5ev\��7#�5m��YQ�ӳ���:H�M�0�D��#���V��Kơ	n owns��%�B���j!��i��(F; �yhy����Τ���Ѡ�u��6w��!�j��Y%$� ;=���#�����&Ș�f�J��I-��9�?o��`����ہ�s�\o�����F�WmV�V����;� �"`�n�, �N�tj����d�yH��U���z	��`�g,rYx��^�D���%R�e�X�ZLl��sdL	�:��`}�~���)0�)`�V;n sdO��}����:`�~Ll����{�〫/����}���۩��_&�{����I'��s�$�n�G!�Y]�`����v����_wf��j�[a��x�1ZLl������f�5�=s����ۀu�:��mQ�F�B5���z��=Z�\ܨsy�N[�k�n����ó��]]V,Y��Ę6D���c��P`�ۀ}���J��I-�5�w�ڃ �"`����{.���KX�n�Kfq~8���&q}�y�8�D�,K���t��bX�%���t��bX�'��{Mı,K�L�K���]c���q~8����ĸ%)��߳��Kı/=��t��bX�'��{Mı,�0F�Cg�'�>�O����&�X�%���{��c73ĦL��9�n%�bX�����n%�bX��}��Kı>�n�4��bX�%����7ı,Oc�0cLX8�.Gn����]B�vT���ܶ΍J9����.
��G�I����=7j{�'�ı,O{>��n%�bX�s�^�Mı,K���t��bX�%���t��N&q3��<yz9$B��YGk�/��bX�s�^�M�� �LD�/�߿gI��%�b^{���7ı,O{>��n%�bX��'��3����F��3I��%�b_{�Γq,KĿw�Γq,$1?~���I��%�b��y�g㉜L�g�}�4KU��Yq�fcΓq,KĿw�Γq,K����]&�X�%��;u��K�g���_�&q3��]�f��BR�.&f1��7ı,O{>��n%�bX�s�^�Mı,K���t��bX�%���t��bX�'�0@���B1J�H��,���d�\��\�܍��JJ7]�wa4�Y�Ur�4Z������vJ�mѱsJN�V��x��u/9\Eru��4n$Ƶ���Ok
��[��rnc������(��t<ueњK�/F\�2��W�|�_v�;���N�[��mɚlWY�rR8�ӳ�tn��9�7�Hfݭ�T��8����7�����f.����`Wr7�2�����o=;��v�L-�^$���J�ѹb��vE��ݫ:c������]:��T鉵`�Q���oq�����~~�͚Mı,K���t��bX�%���t��bX�'��z�7ı,O�_�uWX��i�_�&q3��W�����?�q,K�~��&�X�%���~�Mı,K�v��I���\Q�C��[����Ⱅ�U��m�/�,Kļ����n%�bX��}��Kı>�n�4��bX�%����?L�g8���~�c��/�����ı,O{>��n%�bX�s�^�Mı,K���t��bX�P����L�8��N2}G�"!
`�S�˜�&�X�%��;u��Kı/��gI��%�b_��gI��%�b{����q,K��=u���ɜd�*�\��muѺ��!�yꗵtɛ��x�o/�@���(6TP��%u�']�q~8���+���t��bX�%���t��bX�'��z�7ı,O�ۯM&�X�)�[����-V�Ye�RKs����&%�~｝&��Q�L:���'��n�7ı,O�ۯM&�X�%�~��s����&q3����+j���33��I��%�b{����q,K������n%���"b%��߳��Kı/=��t��bX�'�wئ�R�������q3��L�����q~8X�%�}��:Mı,K��{:Mı,K��}t��bX�'ܙ����GUu��\v����g8������/�X�%��X���:O�X�%���}��7ı,O�ۯM&�X�%��f���y�:�q��M*
����\�<��3S�vdz3��NƋI��Z�1f��s�&�X�%�~｝&�X�%��g��Mı,K�v��A�},K�oM2�e�e�N2�9߾�x.J����s�&�X�%���}��7ı,O�ۯM&�X�%�}��:Mı,Fq?�޹���g8���5z9$E#�3�˜�&�X�%��;u��Kı/��gI��7!��(P�qf�}��t��bX�'��z�7�&q3�Ӿa౜%u�2����Kı/��gI��%�b_��gI��%�b{�ﮓq,K�;�M�)��'8��[��!2�T˓D�:Mı,K��{:Mı,K��}t��bX�'9ٯM&�X�%�}���/�8���-SA|� �DMޱ��,5��Jh�t���Ƨ�f7f�(FGf�ѼH�	Ό�Yk�w�{��7���{=��n%�bX��f�4��bX�%����?蘉bX����:Mı,Fq-���~��KX�e,��㉜L�bs����n�c���b_߿~Γq,Kļ����n%�bX��}��Fq3��_N�F��U�:�ai�_�%�b_{�Γq,KĿw�Γq,K����]&�X�%��vk�I���&q3�����Fܮ����v���%�g�X��{���7ı,O߳���n%�bX�w�^�Mı,��?��""ЋV-R��L!��@��wȜ���:Mı��/����������8�L�,O{=��n%�bX�w�^�Mı,K���t��bX�%���t��b���/�{���@݄v��U����E9	%�:e�̼9dݫ�.�;����v��涠�nn�\3�3.s~ND�,K��]&�q,Kľ�}�&�X�%�~���&�X�%��g��Mı,K�笞�2$J� V;L��q3��L�~����,KĿ{�Γq,K����]&�X�%��{u��O⸩��'�~��QڬV��$���㉜L�g����t��bX�'����7ı,O�ۯM&�X�%�}��:Mı,K�����j���t����q3��L���}t��bX�'��צ�q,Kľ�}�&�X��b&9����7�3��_����/ֻ)kUKmy���bX�'��צ�q,K�������'�,Kļ���t��bX�'����7ı,J��C�$D9B��Ƿ��^C�n��&�v�r�b[�Zn:B[�Tػv���ҭ�g/��'��)l�sp2��6�&�`�/n�N�HJYK�Q����l�cdC����`�b�.�
ؖ�pip2L�K8YT΋�EE�d�t��}�gC�j�a�6�l�n��X���[l�c�nrѧ�#'��u�y�@����s�vŤ{=��Ƒ�u��6f�[�k*㥹J��vq�{��w>�z�����gO%�51�P�ԩ�f�㕺 0�<�Ոݺ{�q��V��ԥ���ı,K��gI��%�b}�{zMı,K��}t�'�1�q��qL�8��N2������b^S&qq��7ı,O��oI��%�b{�ﮓq,K������n%�bX��ﳤ�Kı=�=}w��Lٓ2��3��Kı=���I��%�b}��zi7ı,K�w��n%�bX�{�ޓq,KĽ!�g�3.st��bX�'��צ�q,Kľ�}�&�X�%�����7İ\@˧���|2q���eч9$$D���8��n%�bX��ﳤ�Kı>���&�X�%��{�Ɠq,K����=t��bX�$C����8�=uV{]����֙��؝��\�36ikfc�I梺��eS�jsqc6ɇ�{�D���SPI�q��	"��ܦ�z%�b_{�Γq,K��s{|W$
�c#M˜_�&q3��^���p�:` �p&�D�K[���Kı/��gI��%�b_��gI���G�&q-���~��JT�U,��n%�bX�����I��%�b_{�Γq,KĿ{�Γq,K����\��q3��L��w�h⬩���&�X�%��{�Ɠq,KĿ{�Γq,K����]&�X��b'=�G=2�d�'8�;�G�;�K��O���I��%�b_��gI��%�a�������>�bX�'=�c��n%�bX�ǽ�i7ı,N�z�^��.��[�~u����n�7/;;E���+�jy�f����m-�m�
��]b��{���,K����t��bX�'����Kı=�{��g�1ı/?~��e���N2q��r�"B�!�ď3t��bX�'��צ�q,K��=�cI��%�b_��gI��%�b{���q~8���&qzt�y����
ǜ�&�X�%�}�{:Mı,K��{:Mı�x^��a�6D5���K�$�f��:�!�]�G蘊7�@�ֱ� @pd�� C��jUI3�<��� � ���"*�ft�ʄ�qBJJ`ҏ�UڻI���*B�V0UO�8���w�Pq8�P~ .9����$��)"?�9�!O��d@�aC�n�:�w�s�L���&�B�.D��P^�D˔Hà�� �E>Q6.�C���S@#�>��S �x�N��3��&�X�%�����I��%��-���pv����)%����g8X��{��n%�bX��}��K�8�ُZS/�N2q.I$�t�tS/�&q3��[����q�J�GI-�/�,K����]&�X�%��{u��Kı/��gI��%�b_��gI��g8�ų��{=,QX��7)L���n�$n2�r7dn�q5�y�5�ۧl�|/^y�e-cET�ל_�&q3��_n��7ı,K�{��n%�bX��{��~Y�LD�,O߳���n%�bX���23�Z8��uFܦq~8���&qz{�Ɠq,KĿ{�Γq,K����]&�X�%��{u��Oȸ������~�nWI`�u�3����&q8���_��q,K����]&�X�%��{u��Kı/��gI��%��/u��$�V^WP�q~8���+�Ͻt��bX�'��צ�q,Kľ���&�X����C�&bĂF � 2�@GdR� �H���P��>��w�&�X�#8�Q����
����fq~8���+����I��%�b_{�Γq,K������Kı=�{��n%�b������Q;-N�`�2A���&�5���{�W+�kۚ['%�l�:��w\b�]�q0��y��^8��N2~��_�%�b}�{��n%�bX�ǽ�i7ı,O�ۯM&�X�%��w�.%�I���)%����g8�����3��2P2q�GwE2�d�'8��^��n%�bX����I��%�bs����ƠU+$�8�L�g8�=�cI��%�b}��zi7ı,O{�٤�Kı/�����Kı<{ނ�k�����;l�/�8���������M&�X�%����l�n%�bX��{��n%�bX�ǻ�i7ı)���'��ⲱ�r����g8�O{�٤�Kı/�����Kı=�w��n%�bX�w�^�Mı,K�T$"�`��ޘ���1�ۈKtpN�q��[��B�� 
��F�&����=]d緎���p 9�Qɮ^�m��؝���%�ʪfp.	�<g��ǵƷ}�s���Z�qVmC
������s`�{b��ӥ�Mqh���g�3[km�p.����mOg7u�֎���N��6��9���u�f�6z:��&�A��h�S���ݺ�\�N�Z1��Y'tItQ������֏��T��qNÃ��rAm�e��Y�l&����	�BC���׶m�U�WI`Ӱ���i��&q3�1�����Kı=�w��n%�bX�w�^��*�蘉bX��{��&�Q���e���D@䴼�bf)��'�bX�ǻ�i7ı,O�ۯM&�X�%��w�4��bX�'����&�s3&I��@��Z�8�"B�&	s�&�X�%��z���n%�bX����I��%�b}�{��n%�bX��}�_�&q3��^�<e�,�\\�i7ı,O{�٤�Kı>ǽ�i7ı,O{>��n%�bX�n��_�&q3��[����v���ɂ�d�n%�bX�c��4��bX�'��z�7ı,O�ۯM&�X�%��{�4��bX�'�z���q�n'����c]u�1�pXcd��5�'�u���sۢb�����v��d�g�w�{��7��=���I��%�b}��zi7ı,O{�٤�Kı>ǽ�i7ı,����D��e-c
�m�8�L�g��{u��<�o�}�D�K��{4��bX�'1��Mı,K���3����&q3�ݫdG���ec�6��Kı=�{f�q,K������Kı=�{��n%�bX�w�<g㉜L�g�[��m��*��M&�X�%��=�cI��%�b{ﱤ�Kı>�n�4��bX�'�7�L�8��N2�|���x	rZ^T�3�m>�bX�'�~��i7ı,O�ۯM&�X�%��w�4��bX�'����&�X�%��}�ۿ�ns��xxs�;:'���M�:�Ń���+��K��^ˬ�{t���)�{���7���u�i7ı,O{�٤�Kı>ǽ�i7ı,Oc��4��g8������X�R����8�V%�b{���&�X�%��=�cI��%�b{�ﮓq,K������n+��8���ɨ�V*[,R'%Y�q,K������Kı=���I��?���O����Q�Q^!��T�Q9_�]zi7ı,N���i7ı,Nw6wٌ�
�c#VK3����&q3�޻牸�%�b}��zi7ı,O{�٤�Kı>ǽ�i7ı,O���J�kn���^q~8���&q}���I��%�a�Pc�?��O�X�%��~��Mı,K��}t��bX��{����Դ�Ҝ�am����
:��g��Mt��:���
佷1�����g9�.s4��bX�'���Mı,K�{�Ɠq,K����]&�X�%��{u��Kı;�{��Ÿ���LRg��4��bX�'����&�X�%��g��Mı,K����I��%�b{ﱤ�Kı>�=u�\I�2���s�&�X�%��g��Mı,K����I��%�b{ﱤ�Kı>ǽ�i7ı,N�秱�b�,+v���q3��L��u���q1,K��}�&�X�%��=�cI��%�P�Q`�o@� @���,F��Рp}����{y���g8������X�R���9�Mı,K��}�&�X�%��Pc����O�X�%���}��7ı,O�ۯM&�X�%��A�Y�B���c%�1ہ��$<ct�Wg���7���v�v���Hxvy��rWOZ�嚯׻��bX�'1���i7ı,O����7ı,O�ۯM�},K������q3��L��VY@�V25d��n%�bX�{=��n%�bX�w�^�Mı,K���t��bX�'���)��.I�;(8��w@��%�wy�g9��n%�bX����M&�X�%�{��:Mı��D�Nc����n%�bX���~�Mı,K���`�32`�3fq1m�f�q,K?*�1�gI��%�bs�~Ɠq,K���ﮓq,K������n%�bX��=��7+��4ZInq~8���&q}=�LMı,K�g��Mı,K����I��%�b^�Γq,K��(;�D� 	�&幘)}��f�8�Xn��Wv9���<llE�) ��l��30���OlS���K���;(��!�ȉs=��Lr�٫nmv� �x�=��\�GH�/Xu�sh�H�� ���}/�l,��*va#g���gs �����s�mغ���mںك>��#Z�������*�\$h�<c�gXj�"v�:0��Ff�n��#��\g2c��:���1dş6�S��Ӏ���4���RrtQ�F�9chۧ���x$y΋�k�X䮁�=��{��Y�������n%�bX�w�^�Mı,K���t��bX�'����&�X�q3��n�$�B�!a[��㉜LK��צ�q,KĽ�}�&�X�%��=�cI��%�b}���I��%8������X�R��)L��q3��b^�Γq,K������Kı>�{��Kı;��zi7�&q3�}�����Ke�K-�8�N%�b}�{��n%�bX�{=��n%�bX��f�4��bX�%�;��7�L�gv�޲F�Ukl�Y,�/�ı>�{��Kı;��zi7ı,K�w��n%�bX�c��4��L�g8���SВ��U�Я�j�K�r�&�`9�s�!��c�^�V3Ӯ@:�]-m��VZ����&q3�{�x��bX�%�;��7ı,O��{Mı,K�g��Mı,Kܓ�,�QYY`FJg㉜L�g��&��2�(�B ���z�B�_���E�,~��KX��x�n%�bX��{��7ı,N�^�Mı,K�����[���g�9��s��Kı>ǽ�i7ı,O����7ı,N�^�Mı,K���t��bX�'�$��.)�6d̹&s��I��%�b}���I��%�bw����n%�bX��ﳤ�Kı>ǽ�i7ı,O�g�1��V,+v���q3��L���3���bX�%�;��7ı,O��{Mı,K�g��Mı,K�s���*q��I"f�Mͭ��]
9L�/b�嗡���,����Ʈ�vy���I��cn�����%�bX�����7ı,O��{Mı,K�g��Mı,K��3����&q3�}���n�⥲�%�s��7ı,O��{Mı,K�g��Mı,K��צ�q,K�{���/�8���.�f���U��S8�q��Kı>�{��Kı;��zi7ǈp80��%P2��&�\�^Γq,K��9�cI���g8���5?R�Z�+(���ㅉbX��f�4��bX�%�;��7ı,O��{Mı,K�g��M�&q3��^�n'<�b�������%�bX��ﳤ�Kı>ǽ�i7ı,O����7ı,N�^�Mı,K�#�ڷ�,Ű���ͥ�N;��A��:���DdG�[)v����K�E���"v��+��i�Io�/�&q3��]��~Ɠq,K���ﮓq,K��;5��Kı/y�gI��%�b{��OGZ�X^�3����&q3��g��Mı,K��צ�q,KĽ�}�&�X�%��=�cI��%�byM�Đ�V,+v���q3��L��vk�I��%�b^�Γq,K������Kı>�{��Kı=:x�Б����R����g?�1���t��bX�'1���i7ı,O����7İ(TtF
��E� 1G�E�AT��r(�@18���8�L�g8������R*[,RY��:Mı,K�{�Ɠq,K�������bX�'yٯM&�X�%�{��:Mı,K� ~3�}��2g6r��gz��K)�$�D�T�;U)ݦ�^#Gf���$�"s��N�^��{��,O���zMı,K��צ�q,Kľ｝�g�1ı9�߿cI��q3��[���R~����R�.q~8�K��;5��Kı/��gI��%�b}�{��n%�bX�ｽ&�.%8�����_ҸX���d�&�X�%�{���7ı,O��{Mı,K�����Kı;��zk����&q3����r�K����n%�g�"s?�~Ɠq,K���߷��Kı;��zi7ı,K���8�L�g8������^ۍ&�X�%�����n%�bX@? �����$D��߲��H&�{�hI�?�������

*�U��((�AAE_�

*��PQW��AE_���E* �"�0A��A"PTX � B"�2"�0 �R"�1E��X� ��U��((��AAE_���U�

*��PQW�����U�(�����((��((����e5�c�!-� �s2}pC�     J}     :    r  �  /Ң�)@  
 $�)IR
�
@

 � (�DB%�@P@RT@��\    �P  Q@
 w ��K=�֕��{�����yoU*p>�D��E��T��:���P�Ӟ�*��� 9�Y�P��jP �Y` � � � P�@@    �0   T�ҽ5q����4�,�J���'U*f�R���*����-J� �
 "���C� Q:U)��LMQUe�TSR o�[n-�t�ͺ�r�=��v��@>���{��k���s�wt[����P:|�������8���bOy���}��|���7��n��Sӏ`�� ;�T@  � 8� ��}Q޳��ycѹ�t�w�{l8 _o9��vS��|��,����Ǽ� ��>�qw�yyn� ��n�����k� G�E}�|޻x�{�{g��כ�^��
<���]v�ɯ��������� � ����P  bȠ�{�Zrj�qj����쫋�V�� ﾔ徽��g^�w��{_wy��>� R�{m<�{^�,� �y�]�y=�-� nT�w�ݷ�sۧ�z޷�g}�� z6�eqg/v�i{��MK�� �    �n����=������N���u{{� ��W6���}��o���^mͩ]��{��w��Vl� ��wm������@�}���Z]��嫛)͸�}��� zS����g�>�t���-�� 4��T�)JT � O�G����!����O��*�C&�d =��I�JPa2 S�	)*��db40�!IH� ��'@���?�������J{.���m�g�����EQ^�j��AEv����� ����AE�*�Ȫ(*~�����4�It�0`c�C!K���d��,����������لg��&��0ׅ�,c�#Z��`�X،Jc��cm����s8�����,����<5��lK16da�����!�X#0B0�4���Ph�UYM4��V�B�I�!y��EEx�ҍx7���MR��,,d0(����J��5�pI �`i�0Z��()��4��9�{ �0#&�`�\d0��y������cg�f��l3Dc`�!��ry��:6�d0ԆK��N�d�,��f�LAYh�kc�:�&���>Ԕ�@C�������8�8$�I!),��?Y��M�ha�J`�	�m,�:��.g�:�{o��c`AHKE�Jњg��n(�׮� �ĉ8��B1���{��D�|	�Dlla�l�V�� ��u.A��D�Nd5�/)#	�Ҟ����i������_:�?A!��H��M!�<,�7��o{�}��[�3�	"L�#��eF%f���3[��3�k6^��S����ю� �,S1=���ɓ5�,�}����35�e�Lj|X��"XI�-s�v��(��%])�j�0��V��s���oy�f�'���t�9Ae��L�Hh�����5���IACAL�������}���;���Fi_ �C,3���j]ӆ�$͎��� �I�HF���[�ޠĵ��c8eC�� �P�)P���I]��s���R��!K�0#(|�}� ��h2��D����o�y6�n069�mv�7� �Xa��`� j�$�*T�!WN�T$�Pd&"RD�!N�0tSSFI�6��g;HH(� �*��q5I��>�$p�ou��z��
פy��
�,����8c�p�Gi��`h(!&�3|ߛ=���C$l�u��!�*���B�cς#�͆���
��s�#Ӂ�����H=	eѣ�MckF�$f�搌��5��;�7��,�l	��`Y��Le��p�^~�����j��V��Ă��7���C�J��O����T&xxW���Y��X�b���vW��k�R	#0�	��m�r����hH�H��B�������Gi�io[�0�#,����j���o8E�����&��$4�R;��c�������s��(��r�qT=�>�ޖ�c5��%�NKZ���o9����c6�ky�%�D[�!Á	8b�a��#��K!A�2��7�f��G��7���\ׇ�e�ś�TAY�de7�02N�Ѽ����*M1X	#,��J�#3�`��!����a��7a��Fo��a���ȍ��LƑ�R3F�>��l��5ݼ�&{�5�f��g��_{�h�����<�x���wG~C�O��x|F�[;�i�v�n$h��ᡳF����fw����zִi��p�dX�x���Uy�ߵ����39����|}z�oI�@�Y��H��8���������w��
+���' �JJ��Y�՚�Ȭ4Y�3M�H��I�1h#���>!�a���ֱ������3Aa��Б����;('�-�j)0�3a�N��IKLB 4c���4&��s�e��3��y����4c��c	1$�3{�xg6��=�I='Ai�
�Uf�Lg6Q{���y�ԲF��Z�x�᳈xl=cs^�[�͙������z��#�'0J������~zs�Z3��q6ID@Dh��8bV�4�#E&i�	>OC ;@Q�RtÀL�,�8)$F�B�	2 � �I��c8�XSD2�IA��ɉ�,`�N�A*�`hٛ<��,����Ȭ'y��p	��L��IB0HB��8/�ᤃ4o�{��	oG��6�h	gdΜ$��<cЌ9��f�G��c�<O�RIp�勪�s_S�p]|�.Pn�+QW[UG��g�L�#<�C���@1<�c��>�L�����0�t�*PH@i�8h�����HF��i�0֚�Zcp�t��&sxy���a��8�@4B�H����o&�֚��r,B��ph"q�\p���$�&I������n������d�LXILGJ5���^i(Fhזkj�:9�ĵ�(�y�m��C�1�y��4:�~kFk9�q��p;1ɒ`*  ı#�0��y�y�c���o,	Ōv|��w��<>9s�%����69�0��rp���D�ct7:��pc4n�j��2ĸs��� ���F�%�M�g48�;��p�4;_ 04e�4l�#4l�����Z�"&\)�e"^�V�K�{�>��F461�iI�� 	��Ā��&�cQZl6k�7���"3�٭�Hխ�͒��#�c&� ��� qcf��4�݉���@`$;x�,tl�Ӭ�f��p>x�<HH<6�2l�ы)a�a��Q�:u���YK�p��5�p�9kZ.;܄A����y����XϬ��%&,��̤�0�*��,U!��4F�Ȋ�R�Jf
 ��7)��,��U����=kćv���EBb(J���Ф��ic�W6�M�{�����$!,0x�J�1c0I,=6N�`DXi43���8���D�i�Ih�>�Ƕ{�
�zu�=>s~e^&�<Z��F������O]Nj��a�߮}���
@�			%�Q���4�� ��g�LN�OBՆ��1����=4k���{�ckD�:LP��#��F��@�a$����S�2`�D`�:6�!� �t<
�t�d�7�O�<��I(��!&��2����s|x�g�f�a�{��2Z�F�,�N��;)��|�	N:p$�Bd0"�ϳ��|ᡳZ�/�a�,�ݘa�6���@Fb�+�W �Նl�)�N}�C����8��|�����<a�p�`���:�F�6s��xsE�������b{�WS61>��@��)Ă�(�!��ך��Fpc#N�խo�e�6�`�g��=�y��,�ψ�Kl��ѐ�BI��/��o}��4�5��6��a�ı�4K�&l��ۅ�}(�N��p��G
`��I$ �(G�����ǌS?]�2_������bȐ�(�դժ]��&"!�F�dh֎{{�xq��k.&�P��I�$0b$ ���ɖl�׾d��ώ'7��cS�=�<�?o?�D(�orkam�dd[��a��7����7��g Ԏ!���h��e$�p4{B|LU8�!�X�7˥��pa��3-M��Xh������Š��8���F-��u�����<5�1��0�c�O��jsLf���K�g�����i#-Pyf_w\�\��)�[8�.��#`D��k7��Z'���d�4����:7�����h�ĝ:�t����hT�,@j�ÍC�S b،�'d�h��iiv�jٚ��Q,��
!�C	��0 �2�3V���߯<�So�2�|�����1�JX����{�6>�z��F$�:��>�݉�����e�0Ŋi���X/o<<�ǃ�hPMUʃ�AP@���j���{$�m��[d  '@d��h  	.�$    � �۞�l�8y7]m��)��YՓ��5U]-�r�̭PQ��UI�8�ŽV��U�l��:�  �U*ԪE�S���N��o���m�2iZ�T
��)SԀ�u�P
��U*ܫU�E�Tr؜��ue��[dH�m�v�3VEP-���]�ꖡ�1ʵ[+˔���vV��\  ���m�����j`2�U*�v�T��|!�-�6ٷ���z�Ȁ @����ٞ25mJ���h���e� 8 $Hpp�cm�6�I�`��j�UQ�K�� �l9���t��mx��( � [B� $� ��@   �@�Բ�p6�m���p 4kp-�M� ��	%�fI��	mM� �8HA��H����(    �`  H&�ոդ�m�� �m�mض� �ڳV�m��$Zl �  �`| 	� vݰ,�qL-�6� ۶�H�v�ݛl� pӣm�P  pu�kָh ����$�I�m�rW�Iڒ:Vic$�N�����  �l��ޠm��F�l���   nδ [@  �j[Mۚl-6��lm�Ā $ ��[2�Q���V��6��-��-� -� 5��&�p�� ��CE`�@m�tE�miz���y: 'E�v�˚�	4�J�o)��BVR�;�}>m�A^�@u�Z������`  �`8�k^�n����m�u��T�H�x�B�Q�@Z�n��ͭ���Z�=n��p���se���h�	,�󍣒K� �h�m���L�� �\���-������jU��{���ʭ ��l�Y!Yv�f-�A�{j���vZ���2ùF;O*�*걖�h�.i/].�7���M�n� h��r�[�m�6�  xx ��K.��m�؁6� m&�k�[t�I��ڬ�  �uU,T�N�8�U�gEUT�p�T&�V ;˰� m�[m�@�9  �[&	6�6Z�V�ZW�Z��آe�� ���� @!�vKom��� �m�m���ֲ@��� �-���z�	 �f�H ��}�  �� ��m�n�tݶ-��m�,඀�V���!�l�kX[\4R�  m��lH	<�lm� ݶK(�q���$�R����ry�+��m�Ĵ�5@W�����M �R�R�] ;��­ͺ�Aa��8A�z����u�]1ĉ2��[����6�*U��(�7W ��WJ�Sh���PX*���p��!�l�n��U�8)yG�̠5JK����iV��<�K<p*�9��ۤ���.����T2�HQ�N�d��j�j�i����t�E [l�Y@q�\�;l�@X`2UuR��U*!L�Jʬ�Bک�6�l��jݪU�nݜ�K5R�,���YF�"�q�%y��.k[F�-�8q� rC[#$ ��$�m��nܺku�� m�j�k{e��6�  m� �[@��*B� ��fV��YP  浀 6�?B�//յR��	�*� N�$�bK-��D�-�`X֖�m&m��6�٬�p
P ����i0��z:���^�B�����^.��U�h+�s`3;��v����%��m�5O���,���U7HR�UT  ��  u�CD�mRY@��,�<��V�V{s����`� m^�m� m� my�� G p[c]��	    '�I(�hp-ɚ^^��o ݶ �kKY������ m�rM� 6�6��d��`�ki6�[���	  �ie6�֭�!� $Y�r� ��V�!��$m����UUP|��@5���h�m�h�� $HhY�R    ���l   m���9�U����i�m�@U@�۰m�  BM�8$�m��_]�l�p����"кl-�m�f�@-�� ��j�y�`()U7�5��i�u�H����  l�Ŵ�Z��&���Զ��\m�    ����A'�����:��[\ݴ��/C�βF�W�ra��#���8]��+���Z���l6�@ �����6��=�5���� @	��*���mI! ��λUIp[B*E�րky���\��%������m��l^�tۣ]�@���     6� %����BMɲ�U@T��m� �I�E�d��T�$$  �UT�MT�ݫR�T� ��X�ɵ�m��pm�M�{l[x��ku�M�cm��& �k ���6�^���v@��Q��Y؆�p�l���էN�8  �]�m��m�V�-�K��� .�H�@�m� � ��l��6�-� m�v��[V�p$���4��}$�w� ��`@�ڐ[G6�Rm\<�*��-UU9Hrѵn�+iJm�[N[�8���;pa >�����`ڶ ��8-��-g 8��6^Z��ԫ椁Jmckt��p�mEݰ�`rE�Si6 	  ����Km�i��Ԗ� �m� ��ض� -� �M-��Rl�:V��-�&�dIm m�0m[I  �[4�Ad(K<L
O5g�� ��l�媶%+T�U��#Y� v��*�Yb��0A�g��.�g n׫eP��C<�̮�F�s��[�ںI ��P �U�
�x��j�Yd��-׮9��������뭠��`H��A�I���S1�	8[�+�Q��EJ�*����m]*��Kt��P @3���?���y~�K*�`� ����j�e��تU�U��������9j���� 	 si6xmz�h $u�d�V�KhI׫@  ���m�y���[Yv+���N�X��$8R�j��ަ�l�� I��m���o0mm�m�H �r�:I�jF�m�� 6�Ҭ�U[R�2�� 6��\�[UV�]�m<�W+��!Yz�ʰU�
��H�`�d�A�:� %�m�V�0 ��M���H!W.Ĭ�X�� A�n��pO@m�.� ��   �v�@$��+M�C���k6�H ��9�l#��%�S^�Ƹu]@Pp-@UJ���VWm�A $���),:E�v�uvdP�m��Ùt��^�2�z��[9���s�mI"GK(y�(����3K�vV�g6� $ �i$�{at��m���޶� �'q�1Tpm>W.q-e��W��XR����  ��u,���	6�4���߾�&۳Y��8�lνh   �40-�����6�̒� ��lŵ,���L [u�07ԭ&�|m� v�$�h����$�7l h H6��i�t�\]6  m�  ���e�(m�` m{6�Ti�`U�\i\��ݝ� /.�]��a����V��g����>_*��P:(ڪ��ˈ7d݃c��Be@�^Y`kj]�u K9wma� @���m��U]u�y�=&Ҙ@j@ ���CD����)핶�޲$�����L�`�����M!�L�k��  n˲[(���n��$�Ѣ��wm���+@T��J�UGU��hI:6ڕ&N m�;!��.��8 ���䍪� k�O��n
Im���
ڐ���% �T��IX�ˮ�u�� ��R�e@�UV�+*8 𶂺��ao^�mm� �$ڷ�M�sm��v�  ��l � ��-�����^� �6� A��o�|�`	8���'E�v�۶ݎ_Z ����&���� ��7j�  $ ����n:�y���/�����hHm&�I,�j��nt��8��.I�Ƌ���@�M�o����I�R�l��I��im m� � -������ 
�]/<��J�ژ�U� ���fӦ��-��aض��@[D�ioP�n�z][s&��55�헩[[Y8[dm�m$���l`�  gD�� M� [BG �:�8m��8��x�.�bn�5�ga��m���#��y�s���7c�%��������a��f�pa�J�,ړn୕V�P��b{��T�W]C��������q�W���&��3kh�^��J�P�V���U������M,��7R��P6^� %��ۿT�]�����z�k�TU8��]�$Q�`�(��?�g�}]�qL]����x"m@1�"p�b$�tC��Q8��*���0
=Lh.��L@�����4�? z�I�fHe �N
�(T>x*qp�+��*� ��{��"��l=@�x���S�`�P��)�i�N"��
�z|����z*��đ:�� ������<^����t��`�\�QaX���">��Sz� |����>:�;� z��࠿t���!��(}:P@(�� N�tq�=Пʠ�W�i�]�����V�>��Џҩ�x�� m�x#�@��<BP��L�zP�� G���� =� �� 4	z���W��T�m�=�Vͼ:x��u2�$"#@��)�P08�=��P��x�����A4��3�s��RL(I*�P���0QH�4+��(oh�*�����8@$�*�)!,�"�J��&�Q�S�>��P)C�N�}����0J�� }X �����>�p8mq4�I ��y���� =�)����0PpPҨ+�*&/  �8���!ꏒ/R�� ���+���(03�a���y����w�{{��*��Z�8�m��sk�$��L�D�mhP 
݀ҙ�4�ut�Ĵ�8����x�h;@l;�@��&��KO;;��`� )b-����G��[AY�k��cj��S�24AJ���[�p٢̹��j
��8�Wd�sbIv	���\�X�u�X
��m 
�U��,��pζZvm���<i��-�Ҋ��M'h�EӣZ��#l&�1ۥXcs
����*�Y�%����v��e-K�2�A=�`�s��َ�l,�Um�)�,Šu;�I*�I�N��h	.jӬ�&�;D����Z����4e�镪��sU����z�My�R��(�uH�`��!v�ta�cR��0�H�x�{Ojٮ������4k�	�>e�ǔK�����J�[� ���0��@��j�F���M�y:���eE+'K)�2k�j��U�5l9B�Hԅ!�h����L9��n�UVѪkY��l���k0(2*������f魭�����^��aV�s��vV�SW[W\1ӎv:�dܽ�I��E�u5�Q,�}��C�;K�ٽ�]��d!���\�4���T�㴐s�5�v帶޵*�$��#����$<N�������-�7=�1����@܁���h�#��Wg��pܗ���Ucx݊&��/=n���JЎż��V�s�󳩅n�#�Q�ָ�6�+�6�Z�x�AC�5�&ͭ�3�CP�`�Nl�!gqvvC�G4�!�+sv*s��Pn�*�ػf��gZ۶���к`i�R7�q�զ�:��y����"N�&ZS;Omj�ۙ�5؇s���Z��Z�PqR���˻u*�Q.�Sʀj�i���`�`6U��)Y�iKWS���q�RїV	lX����gz)�s0�]r�U%Ŏ&�7=���ls�/-�DOS N2�˱;�dV�Ԕ�����uIS���T�ڮ��ߠt�v�
����ʇ�'���SJ x��pU>�[t?�Ms��t<a蜣�Bm��2cGF�L���\,j��z�l]q�p���Y%J��;���rdM�>f:�"v]ul�1����.{x���`�yj�E�d5�m��b8�ø�{�NƮ�Ț��rANX��6��6z�&9#�
Uq�jX��r���ka��`|�d�Ӻ�	U�[tb�
�6'i������~*�����f�լ�јk+5#�/g��{r���@��d�)ɱ��g���y;|u�m����λ��Ur�_�� zz���R������W,���vq����K07lT���&�v^9hq�@q͂�s�"54���Jq�`b��`s6i`b��`wj�;�+[8��F0#����Ɉ�r��� �3v����#��[S�nқ�fS�-�2j�v6lZ�.e�6h��s:^�[̶��@w�1׎Z��� 'e�1')�NH���W+����T��L ���S�E��{�5�32i`b��7kM�A�R�JNGKsmێb�l��o���=h���J%9N	�*���l�����`wj��}�����=�^i��D�p�v�[��׎Z���X����T6JQA�)7)4�nq��dny�R���7M�{�֓!��l����ȟH�q�׾VV���Kw]����"i�1��������`q͂�d�^9h���.�l��,�%��?{�L�������R)��!LH`����U�u�s���=��G$�RHX����r���8��;(����.�k7+7wx�;1�@q͂�dŶ��ܟ���i.��w�'2l6����'^�FG	�:%�C�g8u��{.-�gY�����U�m�;q�@q͂�d�^=VR�h����	�`s6i~�H՞�3^�X[��3kRmF9Q'�+�pY�;��U�������v��oN0W�a��8F��K��u㖀��1�6#�W�}���T��((.��?��y�U����Țmp��8�:�5�͚X�����V����2H�i'"ISn�E����;-����f�1U��Ύ:�w�g�/��ة�&�1�|��]X���(������B�R��?w���)K��CW�6���R\�©R���yT�JO~ϻ��JS�����)<���VH*����;q�n�j䗕H�����<��=���qJ
@d�7�UaT��k���R
[�M�B娮��ƫ
�J�K���ʤE'���k�JS�����)=�>�
�K���G�pw��^U �D�}��y)@~g����qJR���`�R��;�u�)JL@�!/`���=ۻ������ ��j�{g�vv��1�iA��c��.yfKn�v\��Se�H��9��Ӷ�'�9�m�m��A�f��ȕ�ۢ#��`�v2�ɚ܏*C�6��_�cD�g,6⻅sϠ+��X�j�u�z�3���&�'Vmnd�7&�|sX�mZX;��]Hc�W\&���ld�z�15JWJ�f)�\�fѼ�f���{���dGȩ q����w�ςnv�q%��l�+���]����]���{X�aݘ�ҡv��-�"����oW����JS�?~���)=�>�%)O~�{�R�����k�JS�ca��� ��K��H*�R���Y��d������)JO{��ג��Vn�������sA�&��B�8�JR����8�)I���ג����{�)JR{�}�JR�}��Z5�����-��WR�e/7�UaT�O���k�R����w����k��)JR�ޖ��޵�e��7�my)J{�w�┥'�g���)���s�SH)~�vUaT��r���c���Gj[���;��C̭Kٞ�h�H�n[!�֓\@��uiM�{V�#��S���o{��}���JR����8�)I��������AT�{�yT��.��K!r�W[�췭��R���w��<�>����G� Ъ~��������{�k�JS����R��}�w����+��q\Wq�;�*�U ��weVJR���)I���py)J{���*�U U���wnYq܇��eW⨯������)JRw���<��=�]�qJR����^JR��]��5���)�/*�U ���j��@��'����┥'��~��R��>�u�-�v���~�8?	(l�W#;
��A�u�^/�I�YoN����n�;�f{r�ͳhG<�7�v�z�%)O~�{�R����ג����{�)JR}�}�JR�}~�Z��1�v�yT���ۻd~$2S����┥'{����H�_��i�H*�U~�P�Ț�r�qFM�c�JS����R��}�w��DdIGB�O���F5)�o}��)C��ǒ���|]�[�[���H�IyT��/}~�U�R
��~�n)JP���c�JS����SH)n�6Y����$.5XU �^{��qJR����JR�g�w\R�/}~�U�R
���;�q@R�N {er�.z�a��9��uύ78�ki�>�8ӎݚ"XEpww.T���ۻaTR�g�w\R������<��<����R
�
��[n�]����>��ȫ�T�Os��� �P	�JN�;�����w�)JP���c�JS��wv�[���f��޷�)JR}�}�JR�{��qJR����JR�g�w\R���74"i��R�8��>��﫝�ۊR��w���R��=���&*�y��*�@�Q7�'���
©R���Bյq�5,���eR
�����^JP�g�}��┥'{����JS�~�n)JR}�ڵf�a���B����-,��F��gr�s��q���;vz*��n�^�t�:�ʙ�3��{�"�g�w\R������<��<����T���ݕXU �^��7B��n�&�k{޸�)I���py)Jy����)JO;��y)Jy���qJR��;vY����$.5XU �_��i�H���ג�������)>�>��R
��~{��q\�]ˆU �)<�{��)�{�u�)JO�ϻ��J�~�n)JP�ޝ�kY�5��k{��9�/�����k�R�����>JR������)I�{ݯ%)M!_W~+ﾮ�� �aQ�I��
@�ۖ���#�� =��حǉiSF��ӎuI��3�^#Zu۴��W���Z93ZV�r�|e8А'F2�܂�3�km�:�a9��%@+�u�hWŜe�e�*q�b�s�zzD:��v��佛�F$�kK����v��l	�yv��ݤ���y���g�#AO;�ĺ�3�5�i�۲��a^�xC.�v/'�������{��w������G6�nG��}?�l�q�1E;�8�F�
�����m��3=��=p������[�T�)?��߰y)Jy����)JO;��y)Jy���qJR���ع��ӷ!dr�U�R
���f�T�JO;��y)Jy���qJR����XU �^�}�jڸ�"���2�QI�{ݯ%)O3߻�)JR}�}�JR�{��qJR�ϺXw{2����lٽ�k�JS����R��}�w�������R����ג���|]�ܹc��\��R
^��֫
�Jy����)JO;��y)Jy���qPU ��7թ���+q�WwweJ���i�v1���n����swb�fP��<ju��V����-�x<��<���┥'��v���<�~��$�)I��`�AT�?w��"�;����AT�<�{��@�!��bTG�>qJ{�w�qJR��s���)��2�R
^�c�n+���>o3*�JR�����)JR}�}�JR�{��qJR����^JR�;��j՛��٣y�޷�)JR}�}�JR�{��qJR����^JR�g�w\R���sAȓm�B�#����>��ܚ_�JRy��k�JS����R��}��U�R
��^v�e�[��VGr��l�Xz�%[˘.���l�]��<���OZ�ÎA�j܍7"���?U �AK��XU"S����R��}�w�������TH*�{�kdL%��).UaT���=�����JN�;�����w�)JRy��k�?
Jw�/ܫyr��+�\��R
[�y�©Q�o����T&��1c��z��5�����a�H��K� �����gA�<ӱ>��1�0�EhCi���`F"2���!#%+X�!�FGq� 4���d�P>u>P�s���{�>a+E���l0r��;�h�D�HH󊞙�
hc z�����C5��� iM�g=%�O�&�����ހuE:"��x$�����.HC�=N�D%��Q`g@<�4!��\_��I�?~��R����ʤH)~ե�oe�di��2\c�J�0���~��)I����JR�g�w\R����I�����<��?��q�+Q�d�pʤH)n��XRP��u�k�R��%	BP�'����	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�w��<��(J!(J��30J��(H��(J�m�@��
�*]�j���nD�NF�X�t=&*���sHN-plwPZ6Aˤ���bUT<�-�Ȯ";�R\X��
���0J��(H��(J���(J��"��(J�}����(J��"��(J3�(J��J��(L���(J��~���(J��0J��(H��(J���(J��"��(J߻�מ	BP� BD%	BP�&��(J��J��(L���(J������(J��0J��(H��(J���(J��"��H T�W��ѻ,�$Q�._�ʑ	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~��߰��%	BP�f	HBP�$BP�%	Bf`�%	BP�	BP�%	������(J��J��(L���(J!(J��30J��(O߿~��(J��<���(J!(J��30J��(H��(J��_w���J��(H��(J���Z�(J��"��(J3�H T�R�x>����ڻ�Wd��	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'������(J��J��(L���(J!(J��30JF��(O߿~��(J��<���(J!(J��30J��(H��(J��_w���J��(H��(J���(J��"��(J3�(J���_�a�(J��<���(J!(J��30J��(H��H T�R���j܍7"���?x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'����	BP�%	�`�%	BP�	BP�%	��P�%*���N0��W��6���%	BP�%	��<���J��(J��(J3�(J��(J��30JT�RH!y��k�@I\RK��(J��<���(J��(J���(J��(J��(Ou�k��(J��(J��30J��(J��(J3�%P�O߿~؃�4>����44 ����@�@��{�=�oZ֮]�+�d�#=OJ4�E�G[ �e��%�nНjӸ���y��}��gs\��?]�Д%	BP�%	BP��%	BP�%	BP�%	��P�%	B~��߳�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP���~��J��(J��(J3�(J��(J��30J��(O߿~��(J(O3�(J��(J��30J��(J��(J�}����J��(J��(J3�(J��(J��30J��(��.#/��!n䌗*@��P�f	BP�%	BP�%	Bf`�%	BP�%	BP�'�w��<��(J��R��(L���(J��(J���(J��?~�����(J��(J��(J��(L���(J��(J��_~��<��(J��(J���(J��(J��(L���(J��~����(J��(J���ar��(JY�P�%	BP�%	BP��~��"��K�ߕ T�RHP�%	BP��%	BP�%	BP�%	��P�%	Bs�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP���ߵ�P�%	BP�%	BP��%	@�	BP�%	BP��%	BP�'����8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	������(J��(J��30J��(J��(J3�(J���~?k3yl��y��7�o�P�%	By�%	BP�%	BP�%	���Д%	BP�%	BP���ߵ�P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B~��߳�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP�}�~��J��(J��(J3�(J��(J�hL���(J��߹�(J��<���(J��(J���(J��(J��(O�?��f�Y��vkv[޷�<��(J��(J���(J��(J��(L���(J��~����(J��(J��(J��(L���(J��?�U\��(O������(J��(J��30J��(J��(J3�(J�������(J��0J��(J��(J3�(J��(J��=����<��(J��(J���(J��(J��(L���(J�����ʞ��w��\겹�5nת���;�ll�0@M���ծ4�6;WjJa�ⱊ����۱�	�����[�W]@\8Tt�ջDc�4U��Q���7/; 8��ݭ�ݎ�-#�4����g$q��d��jl���Ga�ª: �^��/��;���U+Z�y�n��;WI	�=�+*�çIlͺ�r�N]t��9ouvghY�.���%��g��K���6}��}�����w�q~�d�̷]�˺���f�^�y|��e�uȃ��q�qM��rw�ww����\��Z����(J��<���(J!(J��30J��(H��(J����?�<��(J!(J��30J��(H��(J���(J��?~����(J��0J��(H��(J���(J��"��(J�}����(J�R��J��(L���(J!(J��30J��(Oߵ����(J��(J��"��(J3�(J��J��(N��Xk7�37�lլַy��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	����8%	BP�'��R	BP�	BP�%	��P�%	BD%	BR������P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'����	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�w��<��(J!(J��s0J��(H��(J���(J��#��,?on�۵�{޵��P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	���y��%	BP�'����$?���R�w���)JRly)J}���9.X���/*�Ure.����JS߻���);��c�JS��ݼ�AT���Z[68Ԅi��2\j�)Jy����)J?��������)J}��k�R���w�<��=��sF��wT���lYy���7<��PL���Vl9ä��������ػk��4ͿJR���~���)�{�u�)JN�;�O�G��e)O����)?�g��m�EqF�X���
�K��ݼI4��p] |*��ԥ'��?`�R�����R���{��ȏ�:��_/�7vԹ �$�*�U �����R��o���0'�߿ly)}[�|��>����p6D�lN2�7���R� 		�����)JO߿~��R���}��'�@$��?~��T��z�x�#M�-�-��*�U N����R�� ߷���)JO߳��©R���2�R
_%]���\O8]��)8.�vm�^0ڭ\�%Fv��cg��w'8gu���w��?}��ױ�Z����JS�u��8�)I��{��JS�����$�)I����JR��k� �K��q\�\�*�U ��֫�,�J{���qJR���~��R����^U.�UM� ��.->���7rl��x<��=�����)I�{ݏ$<�6�'@��(jGçW��ʜ��
1�O{�~�)UH)v��
�K���DV��;�ַ��R��'~���)ߵ���)JO���%(?"�����qJ�AKu��n2+�7r�%�XU �^����R�����~���)�����)JO���y)J ������,ѽf�<��$�8�;r�NZ�d�gm����ާ�@�]��c���B(�c�G��v��I�����<��<����)JN���~���;���8�)I�ݯ��f��Z�5�7�z�%)O;��p��1ԥ'����ǒ������qJR����
RJ�L�^�7��r4ݶK�>)JR~���ǒ��}�{�R�ȡ�~���`�R���w�qJR��zcW�r�I.�*�rT�T���R����?~��)��o��z���8����$�����}ʩ*vR��ȫ
�K���中�٭�ַ�qJR���{��J������R�����ǒ�����\R�
_*�8[,',%���K�9�c"4� Z�t�k�=N�ݭƦ��8u<"�{���q�q��6;���
�K���U �D�w���R��;����%);�?~°�AT�O���Ej+���%�*�U�w���?�_�ԧ�����)JR����VH*��ߺ�u7T��������b��*�U/w^U �AK��{����U�R��k��qJR�����
�K��r7v�rX���H��A�~���`�R��u���)JN����R��S�\_�����)J����_H���m;���q�©R��}�┥��	�������JS������);��py)Jg�;�ִY��~RQ\P(Y'�n�X�����6�v픠���>O�i.^D���{�*]8nަwg��t��^D�+��6Y��:4��si�-���ehݧTv��,�g�E/E�6����wd��rY)�'�I��#$���l�<Z���e��u�F�U|��ƛ�r[`�}ç,�pg�P7<<� eq�)t�)�"f����V��F���=�`��7�x{�mI1�۱Y���lLv�ݮ�h�ձ�d�:���g�/���v����.l'�6x�)I����JR�g{�qJR������)�뿳�R����X_D6�,�K�qVH*�绷�/���jR���?��y)J~�����)JN������
�T��; .�Vȥ��r_�)?~�߰y)J}���qJ@aK��*©R��u�R
��z���\j�7rD�ƫ
�|�.��U �)?����<��<���┥'����R
��~{�����8�yT��}��c�JS��{�)JR}��py)J}���qJR��}�2����Vo[{!v�b���JmL甸�9��h��:7kg8�V��Rܶ⸣w,���
�K���ʤ
R}��py)J}�����.JRw��AT�ի�7vԹ ���H�������48D� |��=�`�!��Z- z�~�U�I�s�7ۊR��}��p�AT�=ݼ�\�R
^z�t��ݖӽѽ[��y)Jw���R���{���)�~��qJR���������m{�v5q��%���U ��I����ǒ�������)JN�;�JR�|�i�H*�U{���M� ���'����߻�)JQ���������~��\R���{ݏ%)O�}�њ�Lua��I̲�؎Ӻ9�W���C�t�ƅ쥫*l�}�o��e�MY�#?�)JO߳��JR�{��qJR���v��P���=����)JR{�������Q���K�VH*��{4ėԃ�qԥ'����ǒ������\R���s��䟅�%=3���e�F���c��H*�R��AT�=�u�)�Ә��h�� ?(,�����������\R�����m�Ȯ(���aT��RT*^_o_�);�?~��)��o��?6����*�U-�j�خ\�9Gs\R���s����	����R���~���)�w��R�?]�3��6x����W�M�����u]��oms66�Rͷn�;�f{r��0���7N��rR��߷ۊR���{��)�w��R���w�<��<�Gݭj�[�5�oU���)JRw��Ǒ�Hd������)JO߳��JR����qJP*�{�kdCNA�)%�U�R
�����)JR}��py!�#%>�w���
[��VH*�����	܊�%�vk5�qJ_� �;�?~��)�{���)>�{��'��'��=PG�T߅�T�_�;�┥'����\M\�չq�q�©R��f�TR� &?����e)O������*
[�u�©R��"��P���ι��
T֭�9r;N�|mhܥ���*۬��rw��i���Ej+��˹p�T��.��JR�g�)I��{��/%)����*�U ���u���b���R��>�u�?	9)I����%)O�����)I�{ݏ$�����dn�%� ��^U �AK��5X)J{����)��d����ǒ����וH*�R�z�����]��(���rR���L��y�qJR�����<��<ϻ�qJ�T�ԝ�hy(K޵��j�n[%���H*�R��ǒ���?o�����)I������)��o��)$:h5ւ�ON}��v�LD��a���ӎ��J_���`Ly��=��R�ߠ��`oz�[<6�C���."���0��}���M����³�&+:|�by"9Ę����@��xx�d�*��1S'��gj;fB	E�{!�4�lo���<�B5���n��hf���X���7����>����X��C"���wL�Ny�m�l5
  �������oF�o0�{�m����6�%�rF^�^�� (�l ��c�4.ۙ�k��t��M�m�X�$:�4�*���A�ۀ1�_mW+h�l�C�lk	h�k`82+(�v�=UUK�)��B�AÁ�4�Al�݌����e� �]�ʬ��gf�^���\9�.v� @H#���8(w�Z�ez��q[�G��~^'?U;�6���6[�{-�	W��m6Jh�[�Y{u�s�]`�B�	U	U�N�Ij(��S�|Z���2�I��!�q�]�F
Z��UH9+T��*�ͱ�50m'I�P+{k��s��9\��\5&�'A���ט�N-�ێ�H��b����tl�:q���2�nA�k�o8��7F�ϖѦ�ݪfr�㋠ąS�v»Jgmv ꍹ}�L�4!0�K�E��ۂj���z{`��T�U2T��J��we{V�Z���u�ү��B��@qښ��R<��lmI�w�6���MJ����o��䎮�z�iym�- [y�α3���)m�ݶm�h'f�Vm&9�\N�N��H�id� �&Nݔ���I�U�؂b�r���8�v.s]+:��cg0��J˹LV��-]��;l=�'��g���@u�����xM[��J�l�Q+`�������p�v4�y�s�%���v��jp݇H[�.8٥��c���!�۩ù�խB�`����A����N�]�nX夝�Ü��K�kg[��څ��ʌ�&F�m�NͲ��GE�e�*�A�A4[P�Z�DB�p��]�[�gk8�F�K�F�I��X��{ki!�l�Æ�g=R�R�m��;7H
�hn�_:�0v�h�çh(΀%3N�j�H���L��jv�o5�ڬ��Z��h͌N�J���,�C宎076t�l�O��hγb��d�t���l�������u��j�j�u#��B�S<�]O�t�9Ɯ3qҤ��r1���d%�\�ػ1���y�E�SO��J���qg��x���#�x����ʙ��4�_T~�u1sz�/�&�A�l9zƔs�+������Ӄ[���5�N��1@Cs#�z�p���-ƭVe�w&���q��}q���i�ր���zIP�Kʻ6�6�n6s�2 ��8��y�k�f�ۣ[��jsMk��<�|��;%X
]Em2<z���vXN�nq������GX�Ru<��ъa46i���3��[ݭj�Y��*���?�My���W5�X��XD��$&;[�KX����`��ў����w<�}]�+ٽ�Z��)Jg���)JO���%)O~��8�R\�������R�[���	܊ӑ�v[�yT��/M��G�(���jS��p┥'����^JR�g���R��߭��j�#wr⻒�aT��{�ز�%'���^H~EH�Os��k�R��N޵XU �_���DV��;���.)K�@ �;���^JR���ߵ�)JOn��%(?
K�����*��-��2+�7r��2eW�R��u�JR��F{~�����{��8�)I�~�ג�����f����7lލ\�]�z��7�:����Y���t�m�zfg�9�I\X�Gwd� �.���AT��߻�C�JS��)JR}߻��?�s�JS������):~?���k5�ֳ[�l���%)O���8x�a IlC��
�\ 	`w b0̰��}4& ~�%)<���%)N�߿k�R��]��T������*��k��E�ܶK-܋))JO�߿����<�������;~��%)N���qJR��t�;����$RK�U�RI!R�������w������}�R��d��ҫ
�KwQ�!;�Zr9wcw/�)>�}�JP�g�����);������<ϻ�qJR����7.�ĖٹUu��Φ��cuR���E�	��	OQJ�?��3���n��x>JR�w��qJR���ݯ%)O3��\�S�R������%)OS��qZ���2�H��R
^�)�~��?~��)JRw�w�%*�{ﻋ*��_U]� ����XȮ";��˜��JS���渥)I�s���BC�\<UP16#���Js��ÊR�����%)O}:w��kV������H*��%�I4���>��©��~���)JO��v�����#��wJ�^�]|�n�.��W$iUy��P~������=���8�)I�s�j��AT�u�Wh�\Wj��]�.9��a�[r�mri竣	��0o.���c��������n[%��E��R
[�ҫ%)O;��R��w>�'�Po%"�n�bʤH*��C]"w$RK�ג����y�?	9)I����<��;����)JO��v���Bʥ�����`�q�reR
�����y)J{����)��@d����\*�U/7�2�R
_�Ke�Ԅi޷������������ӊR����my)Jy���R��?�Q�䂐?�"�J;}v~ }RI|�X�W��aT��r~�İ��Zݚ�Z����R��w��y)@~�u���qJR�����y)J}����+��߿��ߏ%�+���$t:�h�8C:� �q��X��.��g��{��|�8��ܿ�&UxU �^����R
^�}�JR�}�xp?��%);������U/}\�#��]�܃%ܼ�AT����w���"������)JR~�����)�w���(b��?k��݅�q�+�5XU �[�ز�R
�}ذ�UI$ߏ�� ޽�~�׺���%�,n�X�R�O{{��<}�x�~���UI*{�ߖ /{��H�n�E$�� ��v����*���ǀwwذw�ŀe*UU?5{�?��ƌ�U�6g��Z4�<p���[,v؆��w�g��F��P�ndǢ6����r�6��rnm�tm�Ҍ�Oc,�)�W�A�0���FRŦ㓴�C٭���,�����ۄ�nMv�NWX����pVħ3���;�hz�ͤo���'Sz9. x�=����+���g���\�֊ZiX���i�f�ս��|��O/<��淭kQ�V�E.�d�X(��9��|g�����;�X��';+�����I%s0BwM�r��w/�<ޟn*@8�W�\�����}�l�^�V�iy��W��� qR�$�7&��#��}Da)�N"9%X�ʐ�&#�w=7�I�H\��ldWn���d��>~��}x��0�۫R�o�Vez�q4�9 ��@8��'�\zyR�$�����k6k��]МŮ��@:���5�#9��_E��w=Sj;����?|ag,n�3t�O*@8�.I������:��t�rU���uw�:��!�/^i�(8Wپ��U�~�nU���,�*I&�{܆�D6\VH��q`�{؀q���I�H	��H�N㉹.]����|��O{s�w{����:�__�ﾼ߾#,�+R�uy��W��� qR�$��4�9���c$NR��bpJXy�Ek!v� щ����
�a�$/&�]5����m���HT���1 �� 33n�-�kX�NTI����]p�{ןʩUU��t��;��X����M����q4�9 ����l�`ff�Y$��*�`�*X�%JWW�ٽ� ��u��٨M7Ci�T��,=���r���X绷��Wԯ����k�Q�Z�"Y.�X����:�u�u�{g�36����W�k���"�hq�Hع�f�a��us���]����t�9�:ے�JJ��$9L��rG�:��;7&��l��I~a��� �GA	�8��r7Bn;7&�ﾪ���O�o����v�ꤒ��U+�߾#,�+N(ӻ�'$0ߧ���v��I*M��z��`��ݎ��"��IwT�I=�޼��׀{��0
����*��Q��T8~QD�~��ʻ�?k?j�f�m�n]bK8�OZǰ@N͂ߛ��*��������Չ˖������5	��-/-WFA�����qkP!m����w��竉�#�J8����XݚX�ݾ�I*_�v���<�N��n�8���!�o�4�T�$�5��xm�<��i�*���U�����rԸ�c�p�9��^�ߺ��IS~��0�� ��C["��ԗr^R�}�y��| 'f� �b�&�U佫r5#����������U������|��k��*��6$*�"�����~���%�8�*@�)5�Tq]m�.�`+B\�5Iw_N8˱�ƣ\I�ĸ�l"փ�������v�}�^�uS�a��<�5��Fz��m��l��S+ s�"W���QuX:�����<yΒ[#�L����8�d1��*mh8��=����6�O<;��3�:�%��I�-��ۛv:�۝0&]m�iSP�lT͢���#�`�ER����U����JS��ŜV�9�J��Iu���G>zۭƦŀp�.���RX��Y�Z�F�ܑ9!�;��@;였��}U������B�F8����٥���k�+����l�?�%I6x�m���\Q�������u�� �}�a�J����秋2������A%V���v�{ӌ�6i���Wʕ���<���F;wh�₊�C �6i�u%��q���x��� ��=���ܖ�tKnI+��U�zt����Gny�����s�݄;"�nTS�$JSN7R218��7=<X��x����U��{ӌ ^�!��w,�Z�\��ߺ��}�z�T�I�3�V�� �"pS����U!�?O���q�{��3���u'|�wr�-7w���|٦*��UW}�O�����H�6+R�)'$��,��,�ɥ���U�R���8�<O���8�h��Iw�{����M��=7�vl����8���;�L�B�ͬ=���S���.�h��,k��n����{�����I�q�n���5�3@����x��� �6i�U*_ԕR^Xw˧�ܾ_deȜ�9ܸ�=�vlS� #�-z�諭H�mz�M�H�
�܅����`f�o�-��|= b>лb۶�M,�����D��0G�}�����h�٘���i:�b0P	�6�=P>��� !�P�����<>���.�x�Y�hIҞw�D��0�q#��)�eP���#�B/@��A��)b,O|�X8}�@Hb��������G���":G��i�&+�]� �~C���&�@G����� @��8�(�sj� ~�磌����Vf�:�v%)�$d�ܸ`rUJ��i�`���7٦�l� ��kdCwۖ���0��@z������� ���@9O`�����߃��8醴:�`����/b��v�WiK���8�m�KVT������ջq�JM�H�&������7�4�3k&���򤪼����x�|FY�V���w&��耝�����@8��T�6x�oGlq��������ߺ������J��}�� �~���{c"��w/��Y�~�T���<{g��L
�T*HI��i�{�չv�rA��ǀ{��0���{8�����ߺ��=;Gķ#�Z-\�¯�-V�Gg��rk�3�����wL�����T�ŗ���dPQ]�x���@9O`���W�}�r�zo�^W��F)#dbq��ͬ�X�5X��0�f��J�M����D7q]�j�;��{� �}�aԒT��zq�o-�`�+��wq�Zn�<��U�}Y�����~���{x�9�FY�\���H��`��0�J�o-�?�{� �}�`UR�S�I�b�8�}��33?h����s���Y��:���y*+9e�	&�Y�9��i�囱�7<���E���à�5��Oj�{'3lpf۷0�|��Bxݦ8�]%<e�b1"6��[ ��L��X6�v:2�O�o6lJ��Fnmi����y��1�{@�zm&�;Nm6a��I�)x�P�g�t�t��\hjG�5�Ø��p6sA��Y���$�#ﺕZ��yh�-ȄJ�9nqX���.mF&:r�w]y�>�1m��gZ�8�'����x���:��D�Àw+���VnM,��,-�kX�NTI��U�ݟ���UU$ٽ������f��%M���dm�Q�A�c����|٦�U_R���O����yoծ!4�H��M�XݚX��Kq�U}K}����:��Q���2�sD��}���_ ���;6m�?�ݐ9癞�Hc��9"�����칸���=7;���6ق�[Fy8�=�U��Q�hp�7j�;�4�7�uz���7�OĒ��ߔ��D��n7ifg������8"��b��K��i$���I-o5�I%��yPN�j*i�Bp�Kq��������ߛ�7i$��~9Ē�-ۉ�J#���H����I�狴��{��$�vav�Y�1+I%��Ƶ���D�ʮ˳�I/7�n�Iwr��KrMJ�If�~��ʪ�>����ܻ�N��Խ?Ӯo�bmG$����P��-��p�,�ns��4�j�$�q
8�RIo�_�I-�5+I%����$���ݤ��Ś�I��D�JnC�I-�5+I%����$���ݤ�����$�q��J28B6F'Km�����ͷ�~��7*��cJ��T��P
/]�������癙����+I$���/�Jr�Q�hp�K[�n�Ine��$�䚕������K
)lR�p$t�q�I%���8�^�mߒ�I/{K��$���ݤ��w+P��[�-�;*�i�y�Us��Y�����8�cq�OQJ�d��76H0��o��$�$ԭ$���8�Inl����^ݿ�Ie/z�hR��*q7��[�^����K��-$��o�8�F��ZI.<�kX�NTI����;ԒK��-$�w/Nq~���s´�[�/�8�X�kn$��� �J7$������o<s�%�s¼����\�癙�&�B�`���{rZI-ȶ��&�i)�q$���m����?q獶�oI����sOߛg�����瞮�Ɗ^&:�:��`���WA�}y�� ��8ܱn��N�w{�u��֔�MH.$��i~9ĒKsd��]ܽ?�*^ym�ۜ<m�׽�u�&܄�-I,����o}�3��R��UT��{�������m����~��J�IR�$}h�I�R�p$t6䖒K����In9���]�ӕ�$�[�%�%��)����p���ʪ�_ng7���������Ǿ��m��J���όW�}��D��Y�n�h��T�;��� {�ܫ�P�Qڬ, �:4�zTH|WF�;�Y���Y���:�ᵉlk����A%'���ۚu��9�]������ݎW��m�`�;:���7I� nm��Y�뀡���Tl�����l&� �q�4Y�k lD� �����\eG�z�Lpdr���})��������qۀM]��2�Mm�R��pN���Dƺ��-;g�$+9�y3':����uOV�2�Ľ��f9�`�ʫiU$�Y�Z��B\	p���e�a�u�)�Il��Zv���@�a.��g�����W6���9Lru"��~��XݚXݚX�����[Y�$�DI�Qܘ�l�?���I+����o�|b�76_����#<�לBi��!Q�B����� � v9�ٰ@s��۸�\,�q�v�09UR~�q�`��0|٦ԩWʪ���� ��M����GRFJ��l�3�4�3�4�;��Ձ�����M��4ԍ�U
h�u<l�9�=���j��K�d�ew1�����}ٷjN��#t6����,��,���_y`o���7�/,��j+���3[�W��}��@��H�Xe�=zm�S�o}�Õ^���}�f���܎�q(��H���q`�vY�����`{vx�;ה��)N+.)�ً1~���߾��N0�٦UR~�.��k��m�Q�A�m��@76���**@�j�7���yN�]=q��i�4C��uE��W)qY��ú,��y�Q�����_w�i�CV��� ����**@�j��@w2��R�pdn&�Rwt��RA���ӌ}�i��`�y7]"r�\�-I,� ;��{��0���U"�U��
И�8	~6	� 贒�J��I'��ذZ7D'{,�˴7$��J����}�>07V�X�vX���*9J������ =_?z���������g��)WQX���Y�<uBdC�٭���؃n!���$/&M�������ts���{�b��v`��O����÷g�1�6��)�c�?�.���zg�$ٻӌ�g��qg*��k��$��� �I'%������ɥ�����߾_b������l��.]�HK.C�R}��`�q� 7�ـ��C���t<E|DWz���ʾ���n��.��}�1`*I%�I_����>ߧ���4�5����Ai�ظ�f�a65:�\B5 �������Jrs�{u�.k��q,�<Ӯ�m�;&�'f��{���凧�*@K��!;�dw�hnI�~ݚg�U_$�+����w}� 7�ٟRT�&�w����W�C�`�8�=�׋��Sg{�0;���܎Ӗ(��H�=���`{�0�{��}�~,��my��S���ݫ� {=�`rM�7�@9%�@J��U}������m^k`|��D��G3Ė	By�;���BAI.�`!���=�Ѕ)2UL�0`�X6ac�afxY hv�!��$��/�b���'�l.x7�$	d%��M��ٰ�� ! �gj��.��2&����:��q���
P�J*j�����X~���&i0D��& ���#l�C0!"d�"d�X"	��O��<<B]qe���UK�*P���[�=r�\i����;b֕���Kt�EU��&���������F�����v�r��p�eZ�P�Y�ݚ�ু���;vf�lU��]�9`v3 Z ��u�N 6�ˣvjk-������n�0�4�lSj6�@^��f��ͺJ� $�j���A.slk�o4��t��4��ŝ�I�(��M��<m�����.&;D�r�vT�������a�cT�\�s
�<DU*�Hǥ4���N�xe{/kL;3�sS!�7Ds�ۊ^����U�Yn��5��50it�T��Z��WFDi풳��yղ�h�m�������\]sjb�\^���m,�3,�����)']�gDm�t�,����H���N���L���OIp��:��A��n^D\i�'5��������6ya���𫲵;+N�Z�G�U�t��ā�j�D�W���Ij�e74�T���`����S� �Ӝ�y �-�bP��e��uUUu�r�0^�9pN�� �;��Q�\[Dpl�q��V����2[�m�/-]-Y'u+ζgv�D�ɻ;)�uK��[m�X��eI�͆ճ;v6u����`�A��y���(l��f�kl)AٙUb�������^�E�β�^��DS�58��Vp[���#ƶ��������R��%��,��45R��"��--�9^��۝�UVtRy�Z셒��0�N�)��H�9뜤�%�2�&FFU/�,��]I��݁�d�ƺ��<`Rرq!�=�s\�� �Gmm���5�Tr����ˆ�ˤ��T�nxY���zp�j�3�7����ry.V4+�Ƀ�t�E�Nz]��nq��]��e��eݸ-˨Kb�bj���ų�Y�L@V9Љ�Q�T�vd����K֖)L {V����z�Ӎ�M����T��[��3P+ڂ6ء�ql.��Am#����ZSϦI�:��/Ll���vjٙ�C���.�0���Sފ..(��|�� �����ċ�*�@B�C�=:qOw���w�׷��H�e�[xsr�xp������n�-f�1�ZV�7j��p��v8A
qٟ�y�L�T�����٪�!�;6��Ob�=�q68�щ��yP�e-�n2�Þ#���A����w]�9��.����C�-Fвu�N�΄����X��tu۳���l��0�r#��ۅs���\F���F(��Sv�����?]�ww��{���www޿O���:9����Cyi-Z�s�uǛ���Ws�Z�[o�w|s��	�� �I'' �zx�72i`f�������k���.\�l���C ��Ij�욀�����}UYf�/�7qK�v��r��`}�� od�$� #{Qʻ�n��f��-]�q`r�M��� �q�o��0:�S������qGp�v���٦�*T��s��ow<X�n����4��ڻt���܍��djM��]��S�$�˽''R�t�è��}ݾ~�γsm� ;��;vq�n�X�nϪ�_�w�8�=^�b�Ӗ(��#��7w�ÛAO�]*��:!����������M,��6���S���ݥ\ ���;6�W~�| =�z� Z��۶�����w&�UT���0n��꺰�I{=�`w��q��	M�X�4�=���+��zXݚX[���D�A% ��E\v#�ീ��uXnǷk��|l!�{r������Q�!`n ���{�O߾���� .�k�Er�Id�w-ŀ��ϩ6y�8�;vq�{��|٭��q����`wN0�٦L�$ة�w������|�߷K�!q\p�".����q�ow<X�n����������v���F�)���X�����;��M,;��J�#�T��Ҕ��a�O6x��ػ^&Ƹ�/=K�r��u��.�����|�7&mo���+U����@rM�7�������rލ�h�H;��$�?n�3�I$������w�|�`������oS�8�D���,f�n꺳�K�����O�������[$n˷!��I=���`{�0۳L� �/��$
-��iQڦ��B�&)��������W=���e�#$��R�{�,I�@N���-R�]�VfJ.���;��g3m7*�9�πJ�eK�v��;�gi-A�I����n)DpQ�rXݚ '^� 䖩 Nɨ�Xi�v
Bܸ���7�f��ٽ��`{�,n�,�ͺjR�$��ʑHXIj�욀�o`��rVeˎ��e�?��3�����M��}0{�����=�;��5�[ѷmIq��L�٦���?��b��v`�j�R�}���-� ���q�G/��'���ֶq3�2������
B.Z�;V'�ӥVs�ruH݋`9MZ-���ug��:�v�F�:�q������-[=�Q�lN�Z��sc�gb�v�%���ڹ��#�b9���"[�`�ra.O�"�;(���4�q�K�O@8�b�;v@�I�]n��..R��UM��.��yl�'��^��X�T��%�Iv�#R+�".�r���烬k�N���6�Aͷm��3=�MNZMq��	M�h�<X����7�������7j?&�:N2Fԅ���Y�a��L�����4�T�|�]���M��&�ܶ\Wr�X��� �&������Z��]���.��4=_U\��<��@G%�@����n��RP¤�)V�&����޾W <�&9h��K���k�Ė�!vi
�qtG.��6�g��1h���,��չq�	j��`��ŀ��`n����}]a�}?��������˓���x� y��
U_��1RN�hI����{rZ��U��z���m���*H)��?~~��̚X����9����^'�"8�i����^���@�jLr�n��M�t�d"��su]X^�zpy��K�<�m?S�N8�Q8�9$�l�T��ݔ*���W3����q�0Qkh�'��"i�\N7"���L�ߺ�̚~��3uz���yyQM�0�
7E��91�_����o���;6g$��7����;!n\r\x߿o��^��w�/�)HLQ�% �}q�D2�I��G�*I~�iU{���<���x���N+R(��#����������`���K۷��իW��br���V��W <��@}�l��I�n������>B[\Z�=v����s}��҄��ŵa���m=q�p�,�nSM ��������d��#{[��/�b��=��H������K��n�]�v5��I�^��r�9�/s/t@9/ʐ욀��-�0=��^�&�n�q�*�o���{� �}�`Z��m�0�IW����w�`j:�QM�`��	I,�~��?�RU_UU/��|x�?�`��,F�j�>�
Q�P�*m�HʮƊ��u6vM���3���'�P��3��÷VR8�̚X�[u`j����W��u�<��أ��jE��r�����& 91�@F����=~�_�ԈNT�I�nԺ��������`nd���b۫nlI5D� �IɁ��T��*W���<���y�q`|���_�׀kd�q�		w.<}�i�u}T�os������ ����8f D����}����g=9�;-��
ڻ6˻ ��cq[]�t�6n�WD3��d�E�i/;n{9x��=�n}q�}]�T;<Ò���[l˝"ǅ-��;��d��daz��juȃmQY���=G������g�um�Μ�����y�p�l�֡��;0#�1�h�ݽ�0�\��	����rv�6�)^�F�z���S	mEg���[ �^Mu�W��N{�kf��͛�������Y��I��nS�V��y�q��k1���<�&�:r5�jB���mՀowe��o�$��÷g ��M���ջ��N7"��vg�I&�:��۳��}{�>�T٬;�+��p%��`�OZI :��H	rL@8ᖴ��T����`n��X�[u`���T���Wob�',$Q��ͤ[�� I&�91�@I"����?3���m\�ı�&��j5�[8��q%�����9t���=��D|%n���X�Ut��ߵɎZI :��VUn�I5D� �I�`s^j��AL�$�`���~A�ߗ?s��r�� I&�IQe�������nm�$�R��T�$�P���̭��r�$JF��`w1mՀn���ߺ�?��w~X ��M����w�89 n��������݋ ��V��������i��MȘ�[�:-�]�U9w;��v��mOl2�oY9�+:�E'#�F�JI�;��+wv�������%_��� ���y���{�{����EH��H95ɒ++sn���	*&J�9Vpͺ������� <0� �ȍ��Dң��> ��rP���4�b`���3�,��
Jĝ�8}�ll����H��1M��XjI	��C�H�����H���a�5�X1PcG���f��4F�)� �B��7�v� �C&�@�s@8 ���(:�2�x�;@��D=� �A4*�";z 꾳�E� =^�� ���(8����'�pU������u`bŋSRRNS�I�l�k�}I%M��}0:������<��q`U��$���H$�����`{���p	�H95 �� �n���n�YwN�&s���L���qH(�һ��1���ƈ�H�	�qX��:� ���Xw��ZI^[w��y[��ܒ����,�R�÷�`u�< �ݖ]��o��ӉIJ
J���&Ih95�8� t#(��0nn���}=�`�zX����x=%�����GW��}݁���WRP¤�G�+sv���T�#�P�%�?T�߮����w�Ebz]�c�6�: �/f��6�����cXt�j�v?�ɐq\��GdR����~T�#�P�%�#�R۷r�shw�$��2b���3��:���݋ ��^���I*M���ѷmI ���@w�=h�T��Wnʐ��e���6�#�"l$#q�a�{}�U����X���_U��w� ��}���;�҃Q��X�6��������������U/v��x��-�B�$���t�`w:s�i�*�r6�m�P��!t1�3��\�kN��f�c�KO+p�:�nKbn�:�:m#��\DM�����11�K�e� �fȄ�5pkj�J��W��+�VY���G`�r��i��z����V	�=�ؐ��`x��8�v��M�n���]�am�L<��ի>�7&[#�KqFY{s�i�N2E؛]q`�^������������ߧ�M����������X&�k��]v�z�Ѹ/'8g�]c�,S&+�%�v�7$-�E��t�92K@7"��W,'� �~������73uɒZ� :�`��3��vj��-�
Ed����ŀy�����T��wLξ�j�wq9a"%��ˋ�/����ŀ��ڀ��- ܊�ݻ����Y��,ɋ���0俗�g�? ���Xpͺ�7�ݿ�$�|�L�t�R����&d��[�q�<����7s�-f-��h�T�R	6�9�uX��Vpͺ��Ԓ��{�`���l����$%ܸ�W�w�9��0�1Ha��4��e�op�W~��v5�s+n$�D���Mʰ:� �5��޴��]nVeH�6�JH4)*�;�����`fn���~��`��!>�Zw]�^n�92K@~��=�W p�T�;$�m��oޞߜWn��<[��͑���殒�+]�u�n�tt����99�%�qm�Xn���nEH��H�M�\���u��{q9aQ�Qˋ ��^�@�j��r*^��%˗�����9'�^9����� ��ݼ)*�J��P��Ec5�}�p�^}}�Un�I5D�D�m�a��]~����݋ ��^���UT߽�0]˲�.���HG#���ݺ�=_Vn�r�����Ź������pr%R@I�v�+ŇqX-����Yډ�D@+�;�w-
�R"ŗr'Q��M����u`��`s^j�37n�����H�6��i-�@�j���d��$�� :��K��a��(��'7DnK�{�`flT��]�/ʐ����-V���Vma�fn�� :��H�MAϾ��Ǹ���m!�F�ډ*T�{�z��������osi��*@~�߽���OZ� >���u�9ځV���"n�pv6y��^�\�I���:pK�t��]������鹊����U0j��r*@6ȩ�[�MQ$Q9M9,k�Vf�Ձ���Xwv_>������*i�Cc���OyR�mhz���-3n$�N�JF��`fa�V,�v5���u`��I�N�r)!FY�HnL@rc���R��T�N�E|%(DdI%�J����W]��"�S�$�pU�m�j����ȗ=[v��nj{b ׶����.�o	]��;\gg�['C1�]�y��Gn3�u���6�.��z#' %�e��X���bY�����U��#��Mm��2�dy�Q�n�V���m�lR)Ʌ4e�@��gq��t�smó��!:�⸹̜;S��T�6EU�ʒ�Ȩ��)v��=�y��#�75�67�c-n�hx���p�z$s��g�+ø�=��S��Bo�8���Vwv���b۫n�3u\���F7"�;$T��w �1 �6�]����R�a*A9MI2��n�<�&����ӌƼz��	q\p��L_��T�'��}x��� �vi�w�����݉&��(܉	��͐@vM���� �1��;�~�3/6��]�z��)������κ�Ћ��sv�r���ns�ؠ�fլ��X��얩 �Ɉ�� ��wq܍8[��C ��׋=�����m*���B��y%�;$T�+���+S���5�n�1�=_W���8�=����<h�P�ȭ;��wD��y%�;$T��d�HnL@w����8!�)'��ݺ�;��u`b��`fl�������Ϛ��.p�1�<جO<��ss�6�]�b7QbP�g&���(�T�NTM����1f�36i`wwn���Z��8�S��ݵ\\�� �� ;$T��d�H��ԓTFH�I��͚X��^iT1?�=H�j��b��	�������	�y]X]�vv��Hn&�!�� ;$T�v��y%�a�n'"��Mʰ;��V����� ���`fn�Xה�8�u�*�^.I3�Mi��[���n�Xg9t�F�16�4vy8�II�N�n
HPI*�;����٦ﻸ�Ŀ0���`�{�O����ۻD�� �ݚg�T��7{�`�v, ����UU$fyy��8
!�)7OyR�EH�UUv?{ڀ���&m��J����`wwn���,����r���=1���gsӕU���G)��қ�� g��`w6h�nEH� 9(p��Yw���^�dz�K��-�� �BUx����x�6���R�g�)��q$���""NN�����ݺ�<�w�J����0���w��7M��� ܊�r*@�j�l3��gn�dn�;�-�wq`�v, �wfԪ��w��v, ^y�j'J7$($�`��`w6i`fn���J��%W���,Z7�'�q�m�Q�����@7"�\��d����8�ς����/t����5z�	��ě[�09"ǃ�<6�����g��9�*z#��Wj���H���^.�#0K@��B(�pu�|��wG���Q��8�޾}߀�X��"4H?y��`!����C!0�6 ���P�pNn�HB��%�'n�aD]����ހ�D�'�ˇ���k��%-��aH�:^J�������!�SHk;!������v�;�?������꺪�کl�=�ќJ;��ɹF�<:�EsȀ�+��5#B�nr��3�ZU�!���[��������L��l�)���N�:�F�*��p�#�A��.��e:檩s���[,�j���E`���Vk<u�n�&x����@����B�I��p�D��0��΋�k��nN'[6p�,�T F��\,��n�e����,fcX�=nţ���kb��\�˶�*�UK������YCRܙ����a�6�<�R��D�q+v;�@Ku��Z��k*�85������Ye�b.���sQ��'fwb۱�uI���Λ������;+0\B.�5������/"���;1�2m�n�5n���.��ά������gq����.z�"�a�eM�!a)����n� &鴑l]�W�T�&p�)�ii�%�m��4j��L5U�ciʩmi��yvU�;SU��Nq��6� q�SH���$r��P&C���|��k�0����YA��Ѻ�[�!�͸͸�=. t���δ���Uv���"wW+�ѐ[k0:ԛ�Żb\��f�@%��ȵlܳm@�ez��۔m�r�P��!/\):(��)b�)�U@r�gm�g�y�V�:,F鑅'�/U�+Ht:vr�v���8P=�ka�	�c���������l�`�H8PTl�MczNȻM��Yv�81L� f�m�qT��]v�A�9��YP�s���M"�p�Ԏ��S��䮩�]�u���6ܬ΁85��'�5c�aݢ�S��Z�f��ܔ3%:Ѽ�Աf�
��9AU�f,�&�v�Ǵ��m �,Gj�m�M�d5m.ɭ�0�ۋ=m�=;+=��V��	;vR�h�mYF��h
ڕ�Wl(ۄkN����L&5�su�/5m��̫h��g�V�:�b�������b�dxu�th��>�_uՎ�����t<���z�z�
��6x۫P� ~�@��Cj�M���@���4����=��_=���"�i�T�T�{��{������W?�J�W6���N��9J�ݭ�R��b�:�J�dΦv�&�l��]a��lZ���;����#���ǵ��M$p��P;3�=�[��bw.A&ު�E���2e�t\lmqr�."ڭ����D!n��r'=�l1�$VW�q]*�o5
e��Y�M�us�z�=��xΕ���C�=6��U�Úf��`g.�ڔ�,l�Kr��K�j�U����v��vĖ�r��L����ε&�Mv���nz�ѝDN#�9$
�������*@uȩ vI����僞�z���QF5)%!`w7n�;�,��,�M/�UT�WsW�A������_�;~�`{�L?�*o�����]X��ԓTJr��9,���`��Rﾫ���@GG����8�)	��;�5X�۫ �����K�ޯz�^q�S��P&�eN�]<5�����e��&��Iٻ9����rw���Л��%����o�~����;�uXך����n�t�pRB�IV �&��}\��쪤w`�$sP{�W꤃Cv�^��n17DnK7�� v9�� �5�˙wkM���F7 �����u`��a�O��� �[�Q�,$#���0� ?U}_\~��=�c������ǜw��m\'��&���ٵ�x�V����[�K���B�l����h���������ڀ����U}U�,�b�
�v��227r`{�L �sPr*@�j����#��Wff���$rG����<�w���j��@Ҁc��_y�o�}�w�ʻ�շn6H��7%�殺{��X�,Ǻ�?}UIg���+����'Q����� }�Py%��5�"�ߣ���	)�\-/'Y3�r�n�s3Ys�Ύm�y�����hPVՠwnA�h�T�0!;�eӍ�#��f�yXw6X�ۯ�}U��,�/4��GDH���;���=�H?{Py%��_U��[�Q��ˊ;�0w� {����I�v�� {�� 4��rƇ"�Ϳ쥉W #���䖀;��>�$��UU~�������ݴE$l�ۼ�@s�%��5޸� >ɨ7�ߏ��ۗR۶]�9b���u6UJ�r3�����.�y��#���`�%�լ�ݴ��;� �7�W��,:��V�C�n6H��7%����_�a��L�o������_*���淾�j;N]��[�`o�L�����&���X�� �̢��N%%8�90�^��7ݘ�{��:�$��I+~�ߥ����4��GJR8���M@~n{����@s�%�9_U{꯻�$R��Jdg߿U��foz�����%�KcN�̡,�I�ƒDq�;M˖n�,l��Izm�T�-D�Ugi;9$M��j���V��yգ��걶63s�e�RW����N��F��.�����.�\9{h{;!5��Kecq�՗vݕ'�Q�[�c����6N�:۲���D9�4�vzd��<�51:�b���n��ct�`�߼n�p} �Jt8̅�d��m��������m� ۬�ݑì����1��ṣ.Gw&��b�|ݘ�/u�%U_�����Q�ʑ8�:�w\ ����䖀;�z��vw��w�D�"DDI�`w����,�������]X�,�n�Dq�4�ԑXc���\T�d������޴���$�lQjDܖ{�u`��`s�uXw6X��������n}�C@���{4v�)v%��b�����ླྀ��nJ�NH�D�G%(�I\ �����䖀;��U}�� Qy������h��o|��u��8��
 l~���;�슐욀�2�֛.��r�q�����=�X}UK�M��ߥ���~V�f�)HF5*1ȳ7P느욀�rK@�j �sTi��R/�Q�� 7=�`~���N���ޘ�{��ջ(Z�J�+.\�e�o#�cN��s9��t��㛎9ݘ�J���4��T�""$�9׺���,�6��3�����G�H��G1����yR ���.I��6�M�����`ff�Xwv]��G�2���5�#�,�I
��O_g^�{ذ�kݍ�q9w��[�`}M�� ��u�o�u`ff�X�7��JJr��G%�˒b��H�T�d����?,�������2D.-�VD�I�Ӓu��"Div(��(���/��Sm8�F���ʐ�� >ɨ\�S�E)����`ff�^W�����׀y�O�I6{��ӑ\r_�V�U�����9q�@v8� ��[�n�Er6FF�L����޼���Õ}�������!R�G�ml��;��iƠ�$#�G`wsn��*@>ȩˎb��u�wN����1ڈ�뇭�]r��ӱ��m����?�awn68�5����T�}�R�����r��yR�*{n�J9>Q����M,-�v76�����_�Cv��)�9D��I!`v�=�G \T�}{���BKQ8�ˍ������O�����yR���� $��{�n�nf�y��}qR���� 9T�~��;��~;��PӍ��idv�rY�|�s��P-m	�ɴ�L���(�X�I]oˆ�\<!�y���}j��2�0˂��٪�d�3Es��m�c�\�\9x�L�<���ܜ�|�us��V�X�-Fk�϶᧳u�.y�v�K�ۄՕ	0�<v`n�g�۪�ܥ��;.x2ⱖ���p�6Ѧ^��b��Z���m[��}�����ww{�[������Ė�]��Wl��Q]�,�϶�� ���\rsF��O�,}�kd�e/���}߸}���?=�o ���/�RI%��,;{�X����TJ�$D��8�5���H� ^�~�����Wf����	rIx��� ��w��]����1~��`sL��j�l�PIʰ3� ^�ˎb��H	u�.�3tm�R�Pԕ`gri`z���|��]X�۫:�HƜ�I�rTR?��e�MԒ<�-ŢV#IΥ8�v��˞Cl=���$"�$��Ź�����X�۫;�K��ZJ�#�JRqě���w�8� <�eS0W���@��6ob�;vq�~{��|�l�]��HT�R�piʰ77�Vw&�y.�o^�ob�<�r�"����e�/����O/����@r8� ��S�ZmR�$H��)�Ź�����X�۫:�U�����/�t�GWi벯Y�%	ن�'<v)��Ћ΃�n��D���:���"8�iQ!$�>������}qR��.9�A�[w�t^a�ޗy��}qR��.9�GX�sEM�&�HnQ�`g^j�����rٵ\f ���q	�@��+�� ��������@/}cZl�	M�d	 o���"�$	=���ۈ>����
.�����"l�/TM��V@�jCev�oI�w�`�!��=���=`L��Q�x�*N�l�羽CI�T$"�����L �
V���ς����Z`繊��@�o==E�Ez��6��iT:*>�N�� �t����x��@��]��(`�P�/Q3^wp��۫ �̡=��$�G%8�Vs�*@>���c��g��wkIJR��$�v76�����X��x���R~v��ڀFB�� q ��gH��Z��&�H��9��z-��sP�gdHS�Ԩ�r��������`qnk�Ww�� ��MQ���u�p	n{������{��느wqkM��"DDB��[��nEH���yR[��XH����ܻ�a$�^����� �w�`�=����X���h4#�*��[��r���]�I�Bn*����`gsn�}��}��_����۫��=N6�d�5���{9�V�vku���E�r��;u�[�#���Â��N$7(�J�1w5�[��nmՁ�ͺ�
���NH�rS[��\sꪯك��ʐ��� �f}T����m�$�'r�wr�;{ ��z�[��o�؀��VU�{MJ���*����r�Y�v���u`j��MQ)ʒ������ ՛�@w$�p�yR��H���}�J�ꦗ�����GG���$��.Պ�x_��Kx���4J8(�R��ӗ��kN�Xڣ����Qңv:�r��`BY�<v}L��.��[�O�z�UwBB%�*����[S��m˷n�j�e��IښZ�e��,u�^-��]q�1l�texdXMX���n�F��Nm�a��|v���`��&2�)֖}��m�K���Ѩ�Q����r�������]�2HKF-]����l�pb�V��[�	s�d�೸]K3۔�H��F�{������@r8�������ݴ��Q��BI$v76���f�X���,�v�n$ڡ�EPW�H7 ��@rۘ��qR]nh��ӉʉIV����;�g�����6輛Y�{�w��Y{��[s�*@Nȩ �b;O�ډ�F�M@Q�#��h-Y�jK�״n�nk1��s�qr� V��9gn�7�*@Nȩ �g����=�r��B�e�-�#�`��,��8�� ��D�o5��w;��y�۫Wwbj��RR�~wj]pY�;[s�类ߧ� <��H�̼˖I##���T��z�{{�n�X���a�m�8�e*��I���슐�& %�1:H�ܹ�2[n]��.�Z�x�z�)�қ���q��Ak1���;4
vVz:E��슐�& %�3�r�OyR�^�.��M8�ܧ�`un�UU|���n�b�7��Yʒl���R䑻��.^�w� ���X{IrBUT{T���pD��矸p^��wV���G(�n8�q�{꯾���� <��Hܓۘ���� �Ƣ�ȣ�`own���v��vf�Ձ�0Z1U�HDJJA�6������ml�ؠ��qJ^vD/&�S$MQ*JR/��K����5fk�37n���ՀW3V�ڌ�$DD,�@Knb�_}vI�*@y�ʐ�&/}I&�47��\�,a!$�^�݋ ��R=Wn��b�'���2�⨪4ܫ}_|���*���y��5��P�D�@�A��]�Ժ�5WwP��)4�Cq��X[��	m�@7"�슐�&nf镅��K�Ӂ�Ym����vвZ7W3=�z(8�rs�
D���Ҏ\5���w�O������ 'dT��RIs.�m��Ѹfnm�f�� 'dT��RVf�w�A�Q�E�G*�����<��XuUS|�z���X�7c�FᵻW��+�\��T����c��>UT��{�, ^�ϛv�$����ݤ�� <�=��~�슐�KE^�)WREw��<�v�����@��e�	�wf^�+�����rr|�ݛ�,)�ML�X�r���nq;Y'h�!<njG=vɚ�=�Ļ�t��Y�i�v�)[�.Tm�WkH;p2��u��܏IӔ1Э:v��Q�7]���v��D9��.�C����&��M���=�Mm���\��m�r�69J�v��5��]C� ��P���Vyl
u���m׽w~���޾�����v�˺��Y.Uݱ���"�Ӎz{�i��]�l�i�9��www���;"�슿}\���׀v�vF��n�յ�,|�ŝU_]��ʐ�=�� %�d��/6�N$7nU��ݺ�5fk�;��V�v��+3(OeG$"jJu�`jnb��H	� dT��\˵�r9D�䑦�;��V�v�����X�5��lb[N�R�j�bac�;5�<��u�zת�^,oMv�f�=��fkp����2�i;"�슐ۘ����X��TFJ����R�n{�zx���)"�0��D���˹���*�~�U�{��Ẹ3��&�$�'%X[�vw6����R�EH0q]�i��黻��� 'dT�}�RU}U�_�O;ۡ�6�L���$�X�۫�EH	m�@v8�諭�M��̽4d�@���xh-'n[���s�UϮ�E���q�2�ۗƹ���c��n�m�?���� ;T�ͭ ���j�i�)�RU������Ձ�ݺ�9��V�i[�IRSrH�q���U�{���(!���`cg��}�xr��{�r����8�1��pjJ�7��V3v����xT�$���� ��tv�,�D�o�%i��T��_U}����T������nύm����8�J��2+���͒�ß\[�z8���;QbT�r$k�l��v�ۘ��qRw$���`f�Dq��I#�;��V슐r*@Knb��Wd�<��2���˭.�i��*@qȩ-���mՁ����4�!��7$nU��ݺ�]Ͼ�W�}��Ã"�����Ib�J�ĥR����������"I0ݬ��i-��� 'dT��n�X��:M�D�4�F�*b��l̃Q�e�<P�.�v��L�S8��Nw �7iRIM�`w3n���Ձ�ݺ�}��W�A��`nz�l����'��vEK�}��U]����Ob��H��TFJ����R�w}�Vf�[���*@��]�Y�n�f�������[���*@>ȩ��H�D�2I$vw6�����r���xr���w\��<���#���K=��3�is4��9�C75��15�,>��_^.�<�?2�)�O ��@�TN�x�W�|�3���N��s������������p|FI!(���M�l� ���1P�s��[\���B���"F	M���8	�$�츎�5 �ׂ�<[9�P����J�� 8{�y�k�H����Jh��5�����K܁�t�V�Ea�ڹ�eӢt&F�A��#�I�aҫ۶�K]EseB\��L�zۗ�{@l�I�7%�X0S��ŕ�@)c�fڠ-���˲�f3�Mt���$ѶĻ*Ω�	���Sv6wbnLI�˖ȷL���7a�,�-����z����̲�V��.��LU�P�Q-��pm����Wm�9#X�
�T�J�/hӋm.�H1Z�֔b��$���!*��,P�����a�mѐ-J��%��[���a�ӧ7|�O�2�ԫ*dHհ��J���s�֩������b�&�����g ��k%.��]���Fn�R9�ީ�y���[]d�Y�wO7HȽ�賓EGdͷnNg�l-.͌j�+*�흻m��öʽ��n��s�N�0���v�벵UU�������r��T�y��N�4j�p6xi^e'�I�B�&��J����RZ�ɫ��'t������k!D���M�25Uu����G#�X�k�iӳ�Pz���m�nN6Z����ȍ�tW)� �P9��{o��S���l�"��97�⋢��H��^5��&�������FiD
�f��\�Ī�!�P�$��mU�/Vv�a�sv�r8�A7#��@B]9s�ǜ�h)ݴ�\rی��c[rm����2>�8�lˈe�t�vi4��`����v�����cu����ά�dd�6��ɴ��̰E
1ō8a��U�7U7W]���N�$�sͳ�LiQ�$<�X�\r��켔��7l�n�@�t��x��Rݑ@����T�����i��{���b��Ӳ��G"�;Z2�C+�V�l��ƶ 9�UgU�@^�䫕K���<�<rh9z�2�H�͒E[���5������%��N��a�lg�� ��j��=im#�u�J���6�0�#��U��<�J�]�·4ӺmV�\�:���A��*6Ԅ�~^/U]RR���)Q@8	򯈈�D�Hw\P������(�j 
�HA6�w��V�X���]����%��t���q5S���&���K4�r])��ŷ=w6�]��l9��t�L�dl��[����&�Jh1��q�v�ǈ�>v�{Z:�΢\��n*�{
�q���q�\�uur���p>g�YY$r���V]�=��m�]��-�k�3�k<v/��vnV���3ێ�U9vY31��qǒ�N?=��y���K��/Q�m�Ꭷ��'���[�7.�x��5�n^�l;�f{r��	"M����$�X��;�u`j��`wsn�U���)4�ܛ���}�R[s�*@Nȩ~����n�H�$�Ej9�w� �}�XuR����X�݋ �׶�\r]mn�������;�슐�*@j��`ov��F5N����슐ۘ���- vL�2�����(5٥7KL��[���zpmՔMn�Xȏ�̎�%�\������}� �$�f9h	$T�+��˼�kv6FF�E�k����U^ҥʓ�˥J�5 #���u� /o%h{�R�EK�ctO+�3M���www�=h	$T�}�R\���q&�I�����+wv�����X�ݼ�T�Oޛ� ����i�I�����Ձ�w]��y���ݺ�1n��=�JA�����J<e�Mԝ]H������s���h5�OV����Wm���7k+ov�H�َZIz�����v,�����Ij)%�.[�`m��9*����X�݋ ��Ŝ�Sg{˱Aݩe�w.B���;��`_{�����$Uӵ}�{Õ}�5X��TFJpR/��w\s޺@I"�f9h	$T�+��˼���[q���`�����/zo?�wweX�۫ �j�l�$�ӑ��0���i���n�v))�r/:n�g=3ۜ�v(
n4�Sq�Vu�wv�����X��V��I�Rj*j�����EK�d~��ʐ��9u��M8�7"RU��ݺ�33n���V7v��+3([%
H��)�RU�%Ow{��=��x��Ł⪪�K�iP�(b� x>����~�2�#R�r849*���`swn���Ձ��u`ܭ���"�QT��5�$r�/<�[E�m֮ۡ����cJ����A��r��n�Ձ�ݺ�33n���Vwbj��N
E����o�س�J��ٻ�� ��y��w W{�RN���DI�VfmՁ�y�I*M��ذ����q�]�Ku���w�H�r��*@>ȩ ۗV��T�HMD�AG��ݺ�����ʾ����^�_w9W�W��Q
�ҥC*�w�u˅�A�wq;qɹ1l�q5;bv���64�3vnuf1�7S�Mv幨�-ۭI��0Wn��L5�p�<+����z�tv077/��[�3��3��Z�W!��8��,v�ɺ�6��N�0p�5�N#���=Ta�q1i�h�J[�����?u��N��:���#�sZ�Gf��6��r�CJ����-�4�EF�e�	ڟ���9�~����+��)�.-%�idպ���k��$�C�A�խ�������0�u�n����� qR��$���2��P��l��E%X��W���U&�z���wb�=�wuR��7��W	������V��ݺ�3sn��۫r�n�QԃQ�$$r��*@8�n*A諭���ힴV{�5D�)�8�;�p�����qR�r��*@6�]e�.��h9�-��d�����f�k��ي��]D/nmSmF�D�*%rW ��]Xc���R� ;�We^��u��o3{9W����z��
p��,�|���EH�T���[vfe����Z9q��w���U*M��b�=�Vw~i�7&�JJ�3��Vn*@vc���R ��7h����Z�E�{ﻋ ꤗ�7��<��Vwv���i��k��b`'#c��t�ғ�uŽ�3g8�n7h��i�F���ԥ�J�;�5X�۫;�u�����,�ob��R��$$��I dT�m�H�r��ɷ�D�)�N/�Y�7=�36��UT�!��d_�pO9��|��٥�Ww��R��(ȓ��� ;1�@rM��EH���zf�[��]����$� dT��ͺ�9�7�6HR�'*Ri��O+v^��vk��i�'���Ƴ:�c���vhy36��K��@rM��EH�T��y����o�8�qRnD�,��Հۊ���9&� Sn���^n�xn�V�� qR��$� $ͺ�9��V�8Ԥ��hrU�諭��t�x�ӌw�Ł��T%��P��)�/W������V�{nZ��/owM��@rM�����Ɏ+�}]�E�q)IJJ��p���6;7<��lslP������t���=MBv��+o6�f������� 91�@svi`�ŭ&�NQdJ8X��HLr��`�}{������l'�T���S�))*���XݚXܚX��V�n$�t�q5PQ�`rM������������@uVh{�M8�7"Nw&��������^��?n�0WT�rI-H�U��;��+�U�ꫫa�R�f�*d��b�z�/n�J�I�����7*�u�b���^���m���L�h���78��v�e���_5v�u'5�����۶�q���-�mn+mԜ��͗NY�8-��S�v��WTe�qR���l�ᵰ�ˏ5�����n��g�s)P!�/iӞ�\pt8��Oe*j�D�
�F����ԾI&����%���hr:�Z'�ݥ7f��5�Z��[�a�`�ƻI�b$�\Δt���v����H�ɎZ�l?U}�r�9���5h��JJIC��k�V7f�w&�fmՁ�[)ꎥFG���hI�@>��� 91�@r�ݎ�"��Gq�p������|`�ذ�~����8�ۧ[vȤ�w��� 91�@rM���
�Y����B�q���l��4R엱/lt%�苴��q�6P뵎�c�.s�ٵw�\[��&��׵�w�j��q&ۦۉ�(�9�4���u]��ͯ���[n*@rc��_]���|Ӊ�&�I�������ͺ�9�5XݚXfed�IMIN���T���-�6=W^�z��A���$���V5��W�}�}��G7�� $�^\6̦.��wɳ@gk3]q��[=V�{Xަ�@��lӡ5
�TJ:�$��+��K�����W,;잴m��ytmf�V�m��3Q�#�� ۊ���9�4�
��ZMD9Q(�Dp�33l�^w_w9}�m����L�3,������ ��qS�^	Ȉ�9�'8��Ё�n߇�lSI����#� 6Ը��=z�LR�<N!�n���|5�si����ĵ��1w��h
=��~P�S�T��_m�`J�!�{�x�/��ZŎxz�� C��`Jc6��!��s���xp^ `(:PG��࠺u�X_�W�|PH@�#�|)�^�;Aډ��Ez����{��/s���y���ʽ���J�N��RRU��y����������'���`�dn��]��mA�m�9&� ���T���-����֩8vhѱ4����܌n��[�j׀��]����,���]�#�@�����Ɏ_�a�{| 
�h^��$m5%:�B��ͺ�9�5X�f��{4�I$ٽ˞4B�&�f�H�'��6װ@6����M&�Tdd�8�n�,����_}�xr��d��#��Z��*H��T_��׀z��È��;����W�<����-��L���R��=�H�d�l��l�.�7��e���ι�b�"u�n���f,��v�T�Msv��w�� �yR[s�%��~�,�7�*Pm�u>r���Y���$��_s�;ޜ`����l�t;#wm�m��E�����,�۫Vf�����4�i�I�p��U}U~~^O*@Knb�$�R:�B�6���I!`ff�X�5�w]�r�����Z�R ��.�����v?a�k�ؓ=C����]� ����+a�$h��I14[��E�Vsn�['d�n��K2�u����s��v�y�g�i㎵R��-����	�g*R����m�]�z�|}�7g��R��B��{q��ñ��:���S�5���n��9�*$gv�[b衹���'�Ls
PvyՓ�|g� ���;�������n�;�B�<��ntD`P3�>��w�}�C������s�\X�U��̔OQ�!��C�ݝ͹͂�8��Nt8�EqҔI#m�+@��~v&9h	ٰ���UU\��yR���Yw��FFI#��`s^j�7�4�3��X�}��IR�����Eq\���"��~����H	m�@rc��)�Z�h��D�������X�5�ך���,���(:m:�9B��ۘ���-�6� �X��56x��[�l����=o2�:��蓐�mö�úfg�)����:��&9h9�@>���nb�O~i�ӊ�r&�9�4���_W��2?";N��e��9W����*�^j�
���B�6����B���� ;}s��'^� �j��7��q�ԕ`f��`s^j�3ri`gsn����#QԨ��$NH�kr�=���H�5�꯾����?ĺۯ;�[ �E��T��(p�r�:oI;k�#�m�tiƜ��b�u�e��������o��}qR q�@rc��+��M���DIH��mՀf����U���U��ћb�M�S�(RU�}߻�U�u�s����H
����@m�:����u�+��]X���m���*�wwP���- �� 㚀��ߚq4�܉��ך�W�U}�+��j�� ����WW�Y����-�Z*H��[�u�v��ݮ��tf�*�T��$mԨ�Vw6��\�&9hLr�HZ�4��ڻ�ͼ�7i >��	ܒ���#r����m�:��$��%��{����-��뚀�_d/h����3n�u_ �z��� >��:���E�c$qL FD� P�GC �<_������+��ZM���DIH�� ?US�=�<��ǒZ�}U}���r��'���P�bٮS�S���qPl�΃�m�/L���<���^c^�pr{�%�8�K��UUW,���f��$�i�p��8�3�uXy%�;T���-z�볷O���o��p��`w_���6��U}_}�Y�y�u�< _�P��M˖�KQK��{�I�R̞�&Ih<����Z�5)'N�����V�+ϵ��*��ÕuW�8��2����������$��4�͝���VN`8�����N���͵�D�986�d��գ�۷����4�hsh\"�YӶ�J0�!P�U�nx���Ql��nYN���ţqnUa^�H�jl&�0pr�݁ʡ�UBN������v�����׮�n;v�;sڦ�'\=Ӟ.C,���ݎf�f�(���Nm��fo��G��l#�=���~���޾���JOm�w%=�r�鄢�=/<ۧ[^�f�3�c���C]���k3�.��ݫ��@K�� 8�K@6�^8����J%J�ļ7-�����ۊ�x�9rL@��yf�mm�ٷw�h�T���-ɒZ�$V`nة1��O���Vq����Ih7 'XE�y���Y��mf����Ih7 :���m��{������~�Jz��C/JqCj�D���qSf\%��Ë.�o4[�#����^F�3C3o�vg�h� :��@r<�`��=��q�QԨ�Vw6����@�0�h���$����� 2���N��H�;��{��<�����֫TA���'Q�Vq���Z�$�느���Lܭ��p�ݫ��@rc����- ��^9h����*T�n%�NZ���+s]��y����`~���RU��
\ONF�X���/���&s�D5�\v5��M��r�!{r��RA5��F��������^9hLr�y%�	uyFVZ'�'$vq���U��{�����`op6Țm5NT�V5�ϵ��/CL/U�@6��o��^��Vu惦��ӊ�7Q��c�H}sx�91�@�(�ɵw��T��V.���U��y���=�`~���7��=N1|�4ԍ�PqaBl�%�^t�x��nP�[{Bu�N�6�n��9M2:Q��3^�Xך�f�,]�vw~ۄu)Ԥ�t�����-�6}sx�[p��T��q/�r� ��x�1w5�ǚ�k�V[���Ҕ�D�"Q���Oo���=��x�u�A$��H���E�,	L�B�����zsŁ�z�I���}"rG`wK@rc�������W�Nl�Y�]:.�f�tG1k���S-��y��(��G>�.7K�s�Ns�hES�'\�~���OZ�l��{��X9�ր�%y�T�U�'��٥�#Vo������?=�o:�S`��CW�7����耖�׎Z��� 7�Z�N849R:q�`wj�8��@q͂�sT"�Lܭ����(�1nk�'�������8=׿g*�EQ_��EQ_�@Q�Q��U�TW�DEQ_� ����������ʂ
 ��� ʃ"�4��L��02("�0 #"�0�"�0(0��"�0
,� ª�( !
�2"H��(0�,����DU��U���+�DU�TW�U���+�("����EQ_� ����*���TW�TW���e5�R�אe� �s2}p��                      �   EEE"���� HRTU
*�(@� �*�"B�"Q P �J�P�
��@�)`   )@!T
(��`� 휏NO�&�׵��oJ=���\>�s�|/�y5��w���6��}���}-�粸�� 7ǈ77��uZ�� ����0     �W�v�o
�� �;¯{���ܾ�����{ەfܷ� �>   �P  1� }�j��}�^��__w�=�>[�\`� (�    P1� 
Z� 0  F% ��6   0 � �  ��` �@
l�MD@ ;1J 
 

�P�� h�J� k 6 �6`��7�R緾���:�{Ϸ+��}��{�m����|���ۗ��y=;��+�< Ӿ�i}�>ʽ��W�{:��o}����|*�=}=�}J����}�>�1�� >�  �U �A��
}�����y������/o|^�Wޠ
w{����齯y7޷(r���
�Ҟ�7zV��� a������}� ��[��ީ�������U��=*�|
I�X�r����_}��
�7J�  �<���(  c`
�=}7z���n��k�7g'Tw�J;�֜��s�}>���{9:� �����[�| �}��=|��}�� S�W��ϣӓ\�^ON���}|�<
�8�=���d��%\ =AS{)U(2 h��S�I�3R�SM�ɐ�O���R�4  D�*�)�R� �O�%M�R�(2 h��"$�JR�( �z	߿�����g����w�Ώ{��� z�?� p EO� � U�� V*���  ��?���?ف�������y���4%rIR�Ӓ�����VR
�nNp�~}��\#�ƌF��� �D��.:C`�r�����\�R�X�arֱ���3w�0��a
��,c�2��}'-�ny�8x����i
8���hȱ)��da�	����i$H1�ҡ
ҸFdi�!
���b�$�P��c&9����d���s�O&p��?p8B�P�!YQ��1�Ċ�����dH0L��	L�!XX{�6{��":a�CM79��|�g�粞2�o��/����=��3��z��"@�c�������\���v���t����F,+�$����j��
B��y�cI��%ǅŊ�0adM !Cή���(EH1�!�e�̄n~���?g��~�f�ȱ� @`@�T#�@�)6�9˟�BR5��XH��B6%H$H�XQ����!�J~<��$F�Y�p���2hMΚ{���z��dM�FX�!�	V��%X4%p#D�%	HB Bd��~G�O� �B����R�<�-���ry��_N/�D+��bjD����'�X`���"��@�HC�NYT�e%$��E�I$��!`�BO	C$#	���� ��$��XH0.I,9ṱ��BbAux����������ۚ6�+
�ƒ�J�#1"ZB�@u�8�&G��?$<OX��P`1уC0�#1�FE�p+��1��'����Jp�(V(X�P�!P��\��A���>$Y�t��B6Y���������o����w����d���$)��!e�C���aaT��p#axK(B�+ ń� �̲�2����0��X܅RW�@0Z@���]Iن�����a����6�r�� ad�0M�n^_I�C���}fs��!��S#C��1�#i�'��B��~����*@�����@bR�@$!��	�FD,*��
a�I(K �$�$$HB;\���,(ĲJD�3R�CNC�T�~��P��sw�.sBy3��0�`B�>� G�x¤X, d$�%e!r=��_�r$�a.2��%�cR�p!L!sFsr��-�I���M�K���X�Y#�$d#~��q�IRR�!T���K(BLא�MӖ�3w�H��	2����G�zu����L!R�"ERL�D�b����ݡ=��9�_�?V�.�p!W	!p�a �I6P������3w��i��OZKP�@�Q�@ �2���@�C��f�������c.a�7���"BSܐ���l.���2~���d,bH��R$�!RcHэZI
T��B�KV�fX[Z\�)L%��t&SP��&	�/�=�`��F�� h��ys�=�rI���7���I)밬+B��
!������=��c/���p	8��
��B64 ��{������s�CV'��C=<?	��SbT�"ԍ0���XU!@�_�bP��q��#te�_��g�n~1-H�	�XU�D�-�OҜ`R�o���|���{<�!�n�o,�� f�(J�##�����K�,�!�����)BJ�K)YP�`H�5aB�l ��Ѕ�(A�A�%�YI BY��Io��xL�rt��j��2��#®z SO<	p�#Rd��B�>���D����rK g��H�!%�ƞ���pK�0�L��1H�� 0HJ�:g8K��Yp���[����2BFD��l�,�$4��3��==��*ĉ�F:���5�׈*a�\�,��@a!�)< Ѝ�
P�B��ĂA�R��!�Y	=I����&7��_��U�!BHF�b>��.� x�G���z��y�{��@%�Y�p&��I���3���,G�b$�@�h��jB# ���n"�L0��{��|�=ޠڇ��a���`"j�k �H��T�!�"Z��+B.HF���A�FY �XЁ�Y�H�l�X��(����	 �+%�w�y5�#��#
���h0b`bGD�Ht�@�����N$qܟ�\�C	w����|<ea)�$�J@�B���lf'&9
�X�$�4�Uerd�RGN���)b�<>HG�4� �ģ�J��KCR��Y�Y��$B�� `JRBI�u���3i1y��
$�,#f+�@ ��	���j&DijHFLp�HHE���k "a�j�X@,H�H)�B��"Q! @&�RR��$j0)dd�%FF �+I  ��:���'3g4p�9���`�0����$l� �0�HT�t�p�4��>��
dBN8�
,����ZB,X?�3��g�×5%�Ing�V���9�X�����$�	 F	%�\ i �o���0�7���rX�4%qaq#q�'���t8���Y���k������w�x0d�c�!�́�F�0�lk#�S�@�0i$mŅ�!?P���t��ѮJ"HHB�NE˷�m�7ЗK���KYF$!q!X���=�[?y|0��A�#25$1�B6B>?�7�$���SZHC5�~���/�=����,���4��O�����Y�t��!�?f��o�|�Y�[m����Ip����Ώ:�&a=V1�!CV4�eU:{a�B/�З��sY)@ �W�*d��H��rD�� RI
B2GH�#P�Ec�F�#���(�0!�0�*F^N�á8� RD$bC�M!H�/2sK ���"@|@j2Ejt�P�ؔr$�
�I!$��B����fHaC�ot&�I̦&{�9�����i�L�`���.m��3H�3ܻ�g�kC���Ձ0!�\��I�d}�VB��BՍ ��Q�X��$�����\�i�9=����ü�j����ԌH�H��H @�%s��i#!pu�����#)��=6$d�5-0�W�z,��揞sg
3��M\0b�	ؗ�IwP����<�*f���!X�bH�_H�� \?BB��p�o��7�)+P���!B@ 	# I.F�i4��R�
�4�~�B$�5��<B4�
_ϙ/����K������P�"F�a$A ĊI"ł�J�H�ƒ21H�( �I,�FI!�E���B�	#"B��F,a#@���I@�"��F�V%d����#1$a!!@ ��%�%��zzw�ww�����ϻ�  ���       m��t�        ��  	       �a�                                                                             |�                                                                            ���    6�͘M�@�v��8�g� �2�+S��y� ԫ+��$�:�m�����)�5Y\K$�K(�ݵlm�2]�C�P +E��n[Ki��մ��u�v�e9�Y]�Z�$-�Y%�hk^�^�7dP+�s�R�A
U�Nr�1U��n�Z�V9c���Wl�ȏA�
�� �M�΀�,`m&�*ԩ�V�6�RY	�� �f��;n��� ��km�VFkX HY��D�m�w��V�
�o�ʵT�M2Un��@�qE-��`l�f�l��]��Hǚ�R1��su�d�n�]�VT �UCL�m�ۦ��@ &��lv+2@�P�ݩP%�]����mյ#j�7��[M��h۳m��Fݜ�G]�n�@ �j�U]R���T�T�  R��m���6ۃm���&���s��I�>rۻlm� $ �$ �i,�n�l  �6�m�	 p�t��v�b�gj����D�#2�$ $�ӆp�c��UUR�M�
Ytj�]�[m�6صollrCvؙvU^4k�V� .��AK��8l5*�PVؗq$Z2<�P����QΊ� n�Sr�+U�M@	�vm����A�k$�����^n7+�`ۖ����e�5�� oV���fzKm);��N{
 p�b��j��5�m�@6Z$ m��ۚvŴ-�l��ɑ��]��m[pF˸6������훉 m��[���^����oV���l�G-"Pm��l�6�a�$�-�Kȣ�ݶͶ-���n�b��]�����CSK-��i4�H���sqG`I�5�ڶ8 �p�:Cm�n��k��m�m�` 9�m�,0 l9#���J� 6Ζ1� ;l�吶�lp�d���y�  �Z�m����PȠp5�E+�MU@�=U�R��-[*�
�UUUl�� 8 5���5��շ�v;^���$d�l[F� A����c� �RR��Բ�Z�Z����  ���kpm�5�F�l�	@Ue�5:* 
�^��v嶪�N����-Qk-6���������	�Q������v
�"�i�  �޻lM+8 	�Vv��Mm�$ m�-F��ˍ ��mU�X
�
� �"XbrB$5�&�YF��RZG���q���)5�m�i����m��ڜk/I����x�#��I�f�e�tE�q���6���īUJ��.�5nu����`[m��8�m�c� �ߟ>Y�z�E�kv�Vspm���7[��`-��uZ����8�@ 
Id�\ؑ�BQ�#s�4�<�U+�W
�4] �� �mzrB���r�ܫѓ������\` �f��Sl�v�G5�6�rl4����yv��6�lH�$ȶ�ۂۧD^�����ϛ_�8Xgm���]�X&͊wDjk{VU�a��$� U*�<�C-J�n��i�נ�֮�4W�)@;U� n�	 �:�k@	��7�����UT�}N 3M]AI$ ��m��h�ݱ,���il m��m���8 �-���	e�k6��nݱ�ӠR� l �� Cm�h�j��oD�$[� 5�@ڭ�=f�-�X�Pb&VV�T���õV�P*Ӯv[��s����sQN�J�U�q6�U���ޅ�'j�	 EH �[v�[[v�m�a'�ỳ�� ඀	��Cn�C��m6��`���g#m�*�\�T�U��j��Xm�|$>	  m�p$ k5�m��AH@� 4�Ik�V��ٶ6���6�-�m�n 6Ͱ  ;m� �ඍ� � m����H��E� m���@ 2 m�m��� ��!�i2�H[@Kh �nؽd�V�*k3�r�	��(�۱'m�.�� �� �	�a��  �ɬ� �� �^����hm� � Hm  �  �  [I �#jGt����AS���Cm��t�M)�[A�UU[*s��*� 汤�   � 
��jUꭲ�� ����)����h 	   mtԮ�.���Z�ӑv�Uڥ� ��Uj1� ��6�m�m��e��EH�jؓ[��F6�G[@�nĀ��PE�4�nʠUO*�HMJ��*�lJ��kh ��Vl�ۀ"]n��m����� -�[[����NŽV��[�P�vп������E��T�*յL`M�6M�k9oPhf݀�\i��[AVʼ��s�N�[6������WH͠n�ɗ�.&�8wk]��۝��䮑�b�(I#�m��H�Ȑ�  ��e�m���ڕ`)P��Z���UW���JM����t��$-r�9`.���	 m���-wI��h� 6��np��:[�-����&U�.Aj^(^��m��%���:�[]6v�&ٰ:�#�I�kpl����|�mo�Vն�q����8k��D
C�
�V��*����(
��Ҷ��l �$  �{ vP  [d l�l�rF�am[CZ�r홶�#� �		��$Dmv�E� ۶ ���~�n�YV�vr�5@��"�� 8[@   I�;SD�˶�l�-�-�y�m#m  [Y Ѳ�lH��l�6� N�eH Z�ֻi%�����Um���[s���-�@�8l�$^��4���kM�k�#�  ٶmԺn`p� ||�~o�  m�ڐ H $���e���6UT;��
���������� �f� m� ;e��t���b�W.�t��6����Rv+[��݋hI�� .��&�6�p�����lA�d6l�^��#+TpR�ԫhp   ��` [���u�K� Hh��`тf�-��u2��FG moU���TQ�tMR�ձ�����O�� 	)�,׭��oi�K-݂ۮkp�P�Uz�Y���Է.��\B�ۧ@�4�L9ct����Z��J�P5V[@F�ݭ�啕�T���UUR�s�u�׫h-���ږ�k  �a�K�E��X
��R@vVV�s� [@ ���.-�M�/iV�H��ڛ\ [%�o�> �`-�[%6��3I��`C��@T���C��� m[6ط$�r� 2:@� � ���l]��m[j����[@�J�m���m�-�%,j-l�ki  �( �]��&�n�I���v �		  	�\:tl���I6X"K��Jkn  �Iԣi6p�az�m�m��@[@��EcH�/�2��WJ훦�e��,{T�2���I���ʪL9����^��U���ԄR��q%輐�ڽop����/ml�UUeb4��h֤��l ���>�n�����n]�l<�hV��(z×m4��U@R�2��U#�����|O�*ܜ>&���enVV�l  ��{h
����eͤ�"I.����m[���d 9=���-��$�pA�H��,f�Kn $�׮��ؐ��/F�m�:[m  +����K�\�jU���)o� ��Mڠ6������m��`� $u�[E�K(�S�hp  �^� �m� $��n�Z^��C  ��M�	�l� [mf��ꮥ��VO��m�p a ���Y&� ݶH6��o@�A� *�UUUA X�`m�6�-��]8`nt�i0 $l -���U:⺕��V �@j��5�I'bu�2.u��hu���m� 6݁   $� l� #�Gf�Hm�l�n�5v�  �Z����W���V.;N��mS�����m� [�Jܻ<�Z&b�N]�X���P�[*΅^8��F��6� N����in&�⮪��]�20
�K�v�\K@Ur�k@ m�m�%s���EUE(�*�x�PC�O�(�����Q�P�B�P8��WT��DL���P$E	R�� ��(�%P�ǀ�4DO���S���"����^�/�}�(1�
�z�H���"��A�i�����?'�)��}`��=T5�|��Q���~�lF$T�OP�vz�� ��s��T�A"�P���H�p�� �P�A��z�z'�/D8��F! A��=�z�_QG ���� DE���|EOP��1ʧ��� �/DH`~��~0A�QPG��x�S�A<��A1H��(�^��ʠȈ�D8������/����P��y��$ ���!�ux����t$��A�}:x�=R����蟄^��@����b�DF�E�E�(�{4E�OE��{��D�(j��?>�	�b�P�1E�
��5OLb/�Ŧ �R
����E�� BCT籂�1@C�4O�S���A�> D�PC��
�  ��Q�p �� F�R�@R%�� "'������ ��mAa� m�              �               *�^�l�����/f�*�5��훗fzNڬGG:��u��vR媮L��s�N�&ݺcrե;2�){&K���L�@J�����q��F���^Z �%UV��M�.npzSa8�<���k�8T��gB�[�!sD��.�E��,D�/5�UvQ7v�n�\݇-1�v)����H܍� ]��U�5�����sh 6�탖����*�g=������:Э���	��u�Z�o	���m
�8�D�aH��1'<=qY�ȸ��w8�"�jlW흸L��ǣ9�Bnنn�I�$GOY�m8;t���]*�qJ�M[c˶jVL��\��= I"�$��Prgj�Kҍ���o/+%�����',�ӭ�RNs���۴һ kZ��Z����Ny��ge�5R������@U�+�Vq�ݸB�3�h����ki�f��ΐ"O�-Je*�P�@bl	(fi�d�A���Q�lg�t`H�������Qф[Ch���wtI]SѧnZ���V�G��Y���l!y3u�ٞ8�<�Z�][9����N����]�-�Y��JU��z�!�!�l�:�[h;nW0�"p��O	�]�G F�fJfĔ=�r@]�jۉ�]��z����ӷJLv�x.9P�nmѵ���DL�ۗq/4&_/5�/<���:6M��I2�i1ڡ����R6S���2�]pQ���g2���yZ��[�D��ݯ&�,ŭ���έ�d�h�w���H��m�f�bIF�;"�y�C;nݩ�J�
ݐv��=e���Mxdl��@9*v�Z�����ۻinx-�� �\뗲���5�nF����I��85��7�^�PV���d�y����7ww�Z�ȏ������/�����+�� x�S�C N��U��OGT=uF�'.�Kk`  �`  ڭ�D首Ǣt�M��sUuzݗx�/;��fl��GM�۫s�m ;��f������5�`���6��,"M2l�G&u���s�t	�:S�ힲCq=��GC�)-�J���X�6��)�լ-���̯��p�i���[mT���g"p�Rq��	�f���W����h��7�-�33	���țE�W6NE��l��\�a��x���s������4�� ����Y���~��@>�O#�I��^��*�� �Κm�@�<�\	"YJ�@����:h���Jh�sU����Hm��u�M �٠u�M�k�?pt
�#���i�h���Jh[^�u�M��^�_�I$A �<pi7'F�9Α�&�$']_1&R�: ��3�ԕ�܄�	L���O�_���*�� �Κm�@�|�V`LrdȜ�Н��s�Tb��/��
\t�8 5O�Ph!�C$��_�@?u�@�Қ��!u�LxƜ��q�^t�m�^��*�� ����T�!<�Ȕnm�@�؍RJ�D��Rj٠�u�Y1��ǂrM�Jh[^�u�M �٠}�s��$�I�)������2���<�]�Iȑ������1�$$�9�#�Q������? [��@:�{m�^��;���n7����q&�y�D�٪wb`wC�P�#���i�h�l�:���N�F���X�j5!bUH�Eݛ��y$�����'��mwI )��I�u�M ��4�:h�l�;�6՘E2dNH0݉�l�A�vH�5A�J������Z!�Ra6xR.+j%��5�\f��k���Z�ۛ`�/8�_`7�`�&�P`� ���O��`�%��~����H��� �y0��0�"�ˉ!^d\y��r�F�wr�L�LEP��h�}��:�Q\"��,�%�ܳ@9u�@?$�B\�Ê &$���	�`�� &}��ӒO�k�ؤOĆ�rh^t����٪wb`��D�I}tR\-�p�����h�����S\�.�&��K���N���M���j���4�4޳@�؍�$����G�5l�>�V��2@S"#�ɠu�M� �Κ��hϛi�$�djdNHh�J�.�h�f"j������?R��)�ә�=��<ľ��� ��4�h���q����X'�	�(�4���:����[^�u�NI?!�>����{n�nn����    ꙛE׵����rz���QU�-�og'�+e��Wp��6�%3�/M�`:s��݄v����c��8n�g��#d���n5��@k��[�h�9o$!6��'g���y�pW]���]h���뺊����������2�x��t� p�xc�`�sp�=�wnԛr�iN�������p�ew��v�wu�����`5�Å��bK8�,�\㙵��/n:�WA�;SBd�pSȣMI������>4W�� �Κ���E��didi(7��@:�{�@�Қ����s#OƇ�8��:0�f�02�N0;�ڹg-�1Hb�7��1.ﾚ�ύ��@:��ۑ��#��Q���&rK`e�`w�`6&���������p��%�&��2��+�\��up�.����:;[�"�W�ڈ�3�*��@u�@>\����~�|��@��%��)�ә��{�7��,+"B�Z$rH�"0�"�"BC�d�HH�H�B*@�����bF1�$u��(�O�o$�~�~��?^�~��31 ���ȓ�y0xҍ��M�L	�A�vlLn���p���`�$�y�ff/������`w�`�g,�8�.WJ��q�b`z��I� �<��)�~�u�I&Aᑴ9�ȢŘ����\SŴ��@k��tp����;��[\�:��0�s#OƆ�rh�t����/�S@?^�@�J��j��2
4�4sb`L��b`w�`wv�91�r�J6����h��i2a3�33�:$��w,�;�������ƦE$��~���JhwY�_l����I[��9��ɠ]���0&Eٱ0��D�H�1+�^�����f�J�:te�#�2U�]I��i�u=#ہ�Ά�m�͉�2(0͉�7T���#�0xܒM�e7�3<�ă߯�@ic4���b�N�p����ʻ���0��`M���0&E�>N��s#OƆ�rh�S@;���I;����<*z��Q���tԱ�ơLS ��4��4}U^�? �O&�P`K7bI%@�X5A�0��7i����V�e�;��ŵWk	���y[���(F����S@?^�@�Қ���s\۳�	s���ZI�b`M���0/�S@�z	s��1��iɠ^�F��0&Eٱ0Ҥ�._(ĞL2' �z��e4��4�ՠ~�� �(I��$���9����y������h�b��>�$R@Jò��      t)��#�l���s�<�(�{f=m����5F�nf���kF�ft��3q�'u�xrEӶ��x.*����lG�v���m�N�1]�MY�A7,Q�m�b�/����[��eprf"7d|�)��Uԁ�]Zgj����]��Dɖ*�b�6�����s��������{3�^�m<�v1��-���A_�@�������K�D���%p�l�e�xn���f���p���MuTlJ��"��z�~I'����h��h�����SJ̍<Ɔ�rh��@=�@�e4�[4Ա�ơLR�$Z��0&�ݑ0&�K`wv�9+���ID��@�e4�[4�ՠ�Y�w�sm�H�jdRHhvD���7b`L����$�:Q��r4�d^�Z�ݫXv�g6н���U��u��b��c������uA�f�L	�C���v���&\��pܸK.Mwsg$����y���� ��gy���{�{��^�M����`�&�Ԓh�(�;�&�P`�a���.WB����;�&�P`��e4�:��Vdi�45�@��7b`L��"`HDD�I]���%'\�F������@\u���z{��wXsh2������1[��0&Eݑ0&�����\"rq%nM�e4�[4�)��Y�g����[O�	Ȥ�`=�����w�ڣ��W\���(�L@������R|���2& 8E �0���H70�b�@��/~R ��p ���U�H��"���!*�Q��=|�"H	�x+S�u(�C�1~� ��`��=x�"�������sI�ɠ�e�24o��N/8�¬�X��W���/0�4��|�95��@��� �]�0���*H�#>3�IP�`�1�A�>
���?���U��D �V�c��=�DW��%@�)�<E(�@�W�_a}ߦ��gƁW����Q��Ɯ�11M-f�rO4��hz=3w�����=�upW���w,��L����o4݈�?.��U];s�V0�2ؤ�Ri�C�tl!���9�+I �t�ww���>��]���7u�����rY�.�G�"&#�13������ר��Fe�eA�TV^�%��ff"�ic4�y�/�#}虘���2�VUU_������.�4�{c@>�G11MZu����+	�D�i�����3����B}��גI���y%?����P)���P�"���fs���$��񹞋�˼���
��u��z}3������� �oy�ԒJ�REڳ�J�@[uu�i�nz��v���mHW�7[�S|{�[{<#$O$���޿�@�۱�rX��V�h	�
wysY^"��I�2GO�a��LNO[ ͑?DL��U��˻�� ���#@��o6[ ͑0&H��*��G8q�7U����)�N��y�/����31.�}4�˟<�#!	G"��,�=阈�/{��?{4�ʶI�AJ�  �X3�*�-��`  �A� 
���u���U��n��6N�'h6��#�L�)\��C��s����J.h��]ol�p-��n�M�+�Zs���=um2�&ě��cv�9��'p�\i8�ef`n^Ru�\��vFu��:�9��[�K�X,f�fD�s��0��e�q�����=�[g�I��Pp�������e��?;y���'������t��׭q�F��\X���V�]�{���U�lsع���{��Q���|�Ik�����ݍ �����C�����@ro4è��$R7PM�3@=�f��y�g����M��r��3G�F]����ݒ�ɶ���I������ � � � �{���� �
6=��xpA�6667����A�666>�����Y�n�7sg �`�``�}��o �`�`�`��{�� �`�`�`�}��o �`�b#`������� � � � ���K�f�t�&n��n�A�666=��xpA�666(� �����A������8 ��~�x ��߳<�����\�i�[���T8�KYÓ.�#A�G"%�9�X�X>ӻ��g����w{���~�x ��w�N>A����߾�(>A������>A������7%ٴ�7I�e�����lll}�}8 ����'�� �lo;���� � � � ���xpA�6667����A��� ��A�A��g���s6m&�s7vpA�6667�o �`�`�`��{�� �`�`�`�}��o �`�`�`������� � � � �߹d�.\�sq�n]�����lll{�~����lllo������lll}�}8 �@�A��}��� � � � ����߲Mۻ��7�sN>A����߾�>A���}�}8 �{��|����}��|�����{��g�����Y�s0��04H���4�qQ�`7î�ٍ�+�p��=���˜3.�n�sd�swx �������s�pA�666>��8 ��߼8���lllo������lll�������f��n\4�͞?��`�`�`�߿��8 �@,ll{�~����lllo������lll}�}8 � �A�A�A��������L�.nl���lll{�~����lllo����A�6 ��-�m@@�0O���~�P ��?s�=�|����{�}8 ��ç�nfI-�I��sN>A��A,o����A�666?��>�|������>�|����� ������ � � � ����˥ٴ�7I�e�����lll}�}8 �P=�y����lll{�~����lllo����A�666?�g{������[��)��K�����"�t�tH(����fxՒ�ݙ׈�wlӘnM�ٴ�e��������r{���333��汚O,�-�Ϸ7���ݜ�{����� ��s��@�<�}݈�C��U;	�����s4���@�zSO��ĺ��^�nh�dN�j7#I�D�I����Gၲ/͎�w��VZ1��1����f�����'{������(�Lq�@��S@�2���~ ��&f�0?W�^T��HT��!<�Q�3ÛN��,�;��2q���֚�b�<���SpZ�~(��@q��>�nh�K4˱&PrX� H��.�
�����/#@?rY���DDݝ�4�����Ƹ���9����XeYYyqwYy��c4��V�����L�]��������=狲�5�XD&䆃��X�h���ܖh{�1��h�D	����?��ȴ�����f^Oyt�^��l�tW(�9.��     Ru�c��1�6��P.x��]�3�jE3��������q�`����^v��b�kn˻:��M\Sv*ќ��$g-�켸��m��0n��3�8;e\v�g-�y���eO�m��3<L��]�k����p�:��i{rn�Z�����.�b�e�[V���7<��Z%pvm��w/Q7X�{y�e�Ow��� z����x[�{s���k��Y�=r�b6��+�n�˭N1n����̚jԵ��F�j	��~ ���h�b4��S��������9(ʷ^]f]U�Uy��~]���}317bv�ZO����q1T}\������q�yxh�:�;�[8���>M���|h]�T��FRR-��33�3��Ѡ���?.�h8��X�h�\��`�Ƀ�G3@?u�@�=�?g'�������ȒIQ��'m�v����fYu喍��6uѥ����f��3+)��f)�x�s�I'�=�ύ�}V�����? =�}4�+>Pj7�m�%����'�s���H��� �M
թ�S���2o���$�o4˱�"�i�]Uݼ������g�0�?]�����z�
�U��F�j	��h%�女��|h�h}�~����O�c�H�r
�&f�0=�{��&�:`K�8䟟~����vkCMQ%��{X�-vj�y�Z�պ�0q�۵�7����i_�k�=��Uk��������� �"��Wl3�>4����8�J`� 4��;޻�蘘��݇���y�u�Z�f�2����L$ds4���@�zSe�$D�_�0S��U~���?~�v�����*���_\QWu��"b&f�kY�5mց�r��q3135M7�+�c�/.�.��
���@]iV��f&&W'�? 4�h�Jh��I$�cd�!(�=qt�A��.��%�7vl��)�I��fM�n|��^s�%�4�8�bN&�����^�h�bLLD��jۭ��*��ef]�]aWuy�K7�1����;�<h߼������x����R4��JI4��h֕i�D��O� ��f��{[vxLq�#��4>�<^ۿ��p�y��IOU�Q�+ ��	 �P�����������w�?��\ݒ�*��2���;�[�b#�|߳�;���h��4���I $�ntʾ�pW*����=�F��V&�RlzZF?;�٫xF�$�a##���~��؍�v!���\�ƀ6�VMfVZ��Yē�T���2E�6y� ��f�����򃍸4rC@��f��r���P�<�>k�rYEU�wk/.l����4=3鶟�� ����؍L��D�"���4#Օ^����ˬ��+*�4�r�������9����{���䓇��2@�U"@�Fe<"68$�F���j�"�����!�	T�;�
>�Չ s�)(L#�6�����8��X�!E��G־$`��FT���\�H0 ����ۅ���HF73�"k���(Aq��!c1�3yx�c��w�1���I��)|�x$ȔKN�����&~��$5�!���, L	HL�߃�X~��)�B��GWCR�
� �b�$s#@���w��~I��m���M�,7                                  Νi��н|N�d����۷���JҐ�ۭ�v�q����jx۳N�+���f���JCȋ9�*�}����y�Si��a�N�+-S��H�d�Umm�S�@f�{F�gr�s�v��l��<��qI!�tM�pMg+�r][R��Լ4�_m��1�v{�rJ��f�x�Z nA� ���ҵuV�w>J�[`ͷQ�v%��p���Ҽ��FyU�ȵ�눸�m���bZ��ck��-�<4���:�uϐ��=m�l��s�??|[�N0�=L�rx�<�T�N;��l�H��F�8)��!-M¼��]5+���u�e8�Hm�ZUەg>ě��+���B�U��8+���%ۭv��K�n�v��er��8h1��4'Ó�K�3��@��z�L�ΎA!o���J�ʚf���W���eYeiT�S�l�"�l$֑j�B��eV�1�˚��9����r�-� &S=��:�{�v�)�2w=���3�l[���N�WsZI]�MAq�
���8��g0b�*s�*}w���;�pw;m��v%�Z-��-���*�y�Ij��mh�쭶��kf6����5�-�e�Rn�JxVtG!�yf
��c�n���v��JC���
K6�皂<�]��k�D������O��$�hS����Eڐ�0[;�a֩vz��B�]�S�������V��vv����xS��V�;�ƹ{��.kz��*�d�Cd,/Wer�%�7��yv�d���#�
�%�B\�T�HS$t\%�5�]X�j�e�t�2��6ֲ��rV�;`��>�����JYr;v(���ST�]�1��8x:�����*�k�g-e�	wm�s.�|(=P����o��Q��D>��~V(��T��ѧ����������^��      %�S�+/^��CPb��m4qֻk�RP��Y �fR)�+gY:��܎���m�g�At�.�U�띖y �v���v�:9�ghݦ�OQا<s[cv����V㜫��S��.\k��9g�'A�w�m��r�����\��(�m�*p�0&�UEԛ�ݝ+�v����V�xm!V^�Eac^�{�{�������2�8��1�4�P F�#�����`/���{��t?s����IxO�����sc�}U����4W/���Lq�#��4�؍�"b&}1cO���4˱���#�����S��8h�ۚ��f�"b�汚�c4��pe�K����<��0;������F�6�VMfV^E\Qy��~�����sc��ؘ���$���·=ų�\�yk�bc���8��X�xj�]Rm�:�S6ɬ�.�|�~wb4��ƀ~�Y蘉��A�X���yN)!&��;޻��2��y�
T+E0� �R�!��ү�꯿Uf?u07b�����_~�l���4����Nf�w�M��M>Ľ�|h�ۚ�ȝf8Ԏ�
�$�z���Gၒ/͎�zc�w��4�^���y�F]�U�wuA�ﾛ=��I����of�N�66�mm2ړ��n�ݦ�6н���5�L[�]���}�ݏ��v.Q���:��L��0;5C��UWݰ�gƀ[V<��y0������?�vg�������LIW��A�9���@�zS@��)�b��<�� D1̿��I'����'�p��dq7�ܐ�������^�lh��
=7�Y�6�wYW��qe�8�����H	��}݋�g��0;������~����5kUygh��U�`�5�q0/c�p�k�@�F/���>D�R
&�Ds? {o�@�]�@��(�"'�I�o�*�7W�,��˺��*�34��[蘙�>K�$�ƀ~�S~��<ďUI}����!�@���wr���D�U$�@��u�(�u]"
ȫ3
���C�1鉉�߾� �￷�O;����d:H�5}����?g�y�9$�������%�i7/*�4�r��1舎�����ޭ���}�vI$�(�rl;��Jaն���+�[s�����r�z;}\}�A�9�������h�v�����y����Z�\�ddn@M�+@���[鉘�L]��lhO٠~V�߼�1#ﾈ���'��i��o�9$�}���9��"~�~��<�bX����S�,K�����{��d�.ܤ�sN'�,K>@RD���؜�bX�'��Ȗ%�`����r%�`|�ȝ�~�q<�b]�7{���s���Uow��oq�����'�,K��C�Q�����ı,O���É�Kı/��v�"X�%�"2 Ċ�ޝŰ�     9�Q�I����,{Mֺ㮱�IT�V@R��'�v0�@���C<[]qՏN���9Ӧ
�Oi�c�F��� ������"K����Z������ɓ���l��c���U\K��Gm�n8���h� #�zX�zc��@�fd�;c�GD:;W8�u��΋��d?߾�����ܷ��M��t��=����y�n��!�.D��\�n:5�O]�+m�7m�i���ObA������qj}���w�||�}�kҺt���Kİ~Ͽ��"X�%���É�Kı/��v��"�Dؖ%����^'�,K��3��._�K�ɻ.K�u9ı,O}��O"X�%�}�;�9ı,O;���yı,���ND�Q��,K����.�I2��͹�Ȗ%�b^�>ڜ�bX�'����<�c�ș���Ȗ%�bw��É�Kı,���n�vd��\,�ݩȖ%����}��yı,sﮧ"X�%���É�K���;��jr%�bX��ܛ��Jl�37oȖ%�`����r%�bXʅ~���N'�,KĿ}��S�,K����'�,Kľ���������9��2�@yS�U�scL�����<����lvx����w�o���
�^������ow�}����%�bX��{��,K�������2%�`��}u9ı,O��^[~�s&�r���8�D�,K��wjr+�*�R��D��������%�bX=��u9ı,O}��O"�?ɸ����!�s���Mﷸ��{���?o����%�bX?�����c�C"dN��xq<�bX�%�s�Ȗ%�by���S�L͛3,ܛ����K��@���{���Ȗ%�b}���O"X�%�}�;�9İ:]����Ȗ%�b|gĹr�	t�7e�wn�"X�%���É�Kı/��v�"X�%��w��O"X�%��;۩Ȗ{��Y����~� ꗫ��3�i.wc����L`��]�n�K���Q�-cjU�������&\4�ssN'�,Kľ��ڜ�bX�'����<�bX���n��șı;�����%�bX�{�~ۥ��˹����ڜ�bX�'����<���v&İ{���S�,K��￼8�D�,K��wjr'Õ2%���z}M͹�0��s3v�<�bX����S�,K���{���%�QP8�������b^�>ڜ�bX�'��~�O"X�%����na�nn�ْ\��۩Ȗ%�@ȝ�~�q<�bX�%�s�Ȗ%�by��oȖ%��̃�����Kı>�}ym��̛���K74�yı,K�ݩȖ%�a�1��>��?D�,K���Ȗ%�b{���yı,O�����*����"1�D�;���f:e38ݜ��:�ќ��a�nG����w32�M�sv��,K������yı,���ND�,K�}��'�ı/{�mND�,K�N���M36l̳rnf�'�,K������>c�2%����'�,KĽ�}�9ı,O;���y�?��M�b�K�/�%���.K�u9ı,O���É�Kı/��v�"X�+��?}�}x�D�,K���Ȗ%�b_}���s$�p�m��8�D�,���3�϶�"X�%�������%�bX?�����bX�X�S}U>T2&w�zq<�bX�%���m���e��0�3v�"X�%��w��O"X�%��;۩Ȗ%�b{���yı,K�ݩȖ%�b(����wv��-&���ػ����<=���	�����I��0mڙH��{����w�L-�:��f���ı,K���u9ı,O}��O"X�%�}�;�>Vy"X�'��Ȗ%�b}�ܳnM�sw.̖�\ͺ��bX�'���'��@�L�b^�>ڜ�bX�%���oȖ%�`����r'� ��lK������f�L���K74�yı,K����9ı,K�{��y�� ��}u9ı,N��xq<�w���w��އ��fe�Mﷸ�g��������yı,sﮧ"X�%���É�Kı/��v�"X�%��O{���flٙf廛�O"X�%��;۩Ȗ%�a���~8��X�%�{��jr%�bX������%�bX�
x�EqX�C��}��     �ׯ/M��5�-���v��Ku�i��<ܳ�'s�5�z�{>� z)8�-��P��Kq�;m>׊Z������˓l�k�`��BÙۜ�v���mwlݦP\�^x����.���]+m+���6��*U�+t�sv%�&húW]m�o=7[**�;�ݡ��<�g 2�g6L���f����~ww�����}UZ�:�M<�tF�<9�+bM=�8�u�����J�3lS߽��݈O�b27(���Kı?w��É�Kı/��v�"X�%�|�{��~��,K���Ȗ%�b^��'�]̒e�I�74�yı,K�ݩ�|!��,K���'�~��,K���u9ı,N��xq<���L�bY���n�vd��\,�ݩȖ%�b_�}��<�bX���n�"X� C"dN��xq<�bX�%�s�Ȗ%�b{�Ӵ�ۙ�e6K37w��Kυ��}߾���bX�'{߼8�D�,K��wjr%�`	�
]���oȖ%�b~��htCI�����7���{����q<�bX�($s�϶��,KĿ����yı,���ND�.���=�?��UW��0=<��<s��8�6iC����L��%��/Y-��Kh��.n�r���8�D�,K��wjr%�bX������%�bX?���"�șı;߹��yı,�73����˛�m�ݩȖ%�b_��w��9�V����4�v�� ��H�q"G ��|�G���������"X�%����N'�,Kľ��ڜ��	�2%��N���M36l̳r���'�,K��>��r%�bX���vq<�c� �
4؛��mND�,K����x�D�,K�t��3��d˚\�v�r%�bX���vq<�bX�%�����Kı/�����%�`|�2���S�,KĽ�JO��p�.M�sgȖ%�b_}��ND�,K��{��o�Kİ}Ͼ���bX�'����O"X�%�N�~��x;gA����b,ׂ)Is�4��͆+=k\��ܸ��z>����Y��=ff�O"X�%�}�﷉�Kİg{u9ı,O}�;8O�2%�b^�>ڜ�bX�'}ӹ>�����)�Y���O"X�%��;۩Ȗ%�b{�y���%�bX��s�S�,KĿ���ȟʇ𻉱,O���Y�&ݹ��ܶ�\ͺ��bX�'�s�q<�bX�%�����K��Dz�L[�NE=tR/�("��o��x��&;���t(��H@a��������1F�}��0T�<Gh&���0 A�ؒ0#$b� @Ǆ4���X�	$Z	5��7��My�����ヰ���3��h9@��*�D51Ԫ���lM�O���@�)`Qh��/�~QC��QZx��E`�� ��#N�x�(�!��"����E��@=��|>P�~��/9���<�bX�s�]ND�,K��o,��s&iv�%�6q<�bY����}�9ı,K��}�O"X�%��;۩Ȗ%�b{�y�ǿ'��u��;�~�o��fmq�}܉bX�%���x�D�,K�������%�bX����q<�bX�%�����Kı?�~�n���۷!�e�^��s�JJ�-��婊+sv0�v��sq�ѭѿ|:���kHM�w�����A�]ND�,K�{��'�,Kľ�����_�6%�b^�oȖ!���~����p;#p�����bX���vq<�bX�%�����Kı?g{��yı,���ND�ʙĽ�JO�ܸInM�sgȖ%�b^�>ڜ�bX�'��{�O"X� ?�6&��]ND�,K￹�8�D�,K��/v�wfK�����ڜ�bY�"{�}�q<�bX����S�,K�����K�<�=�;�9ı,N��rv��s7,�	r��q<�bX���n�"X�%���~����ı,K���S�,K����s��Kı?����nff������x�v�<�H��+��m��`��c�u��.�g������%��^����K����N'�,Kľ��ڜ�bX�'��{��~��,K�~�u9ı,O��^�n4͹l�\���%�bX��s�S�,K����s��Kı,���"X�%���g��ߞOs���~~t���fQ���,K��>���yı,K?w��Ȗ?C"dN��}8�D�,K�����Kı?d�r^�L͛.[�.��Ȗ%����؛;�����bX�'�s�q<�bX�%�����Kı?g{��yı,N�I�s�˶eݛ�nn�r%�bX���vq<�bX�+�s��Kı>����yı,K?w��Ȗ%�b+�}��rL���     �qT�Z�j�s������������ş�.�ιS��P"�I<s��8�W�ԃ�:���:x��1\92�Y�������e����Y�ln���`R���y3d�[p6�Si�.'����L�d�){��rAE�bg@��$-�-�$=�mv�����Gk���`G-�����]�r�3���s�K�U[m]�h�D�U�zg/#�V�\Ph�q��6=Kr����w9�)9�ۄ�p�m˛:��X�%����ڜ�bX�'}���<�bX�%�����Kı;�y���%�bX�~�{�K7e�sK����9ı,N����y�9"X�{�۩Ȗ%�b}߹��yı,K�ݩȟ �TȖ'}ӧ�nm�7v.f��yı,K=����Kı;�y���%����blK����9ı,O����<�bX�'{�͹6����2K�37u9ı,N��vq<�bX�%�����Kı;�����K��Q�'�}���bX�'s�������3n�-�6q<�bX�%�����Kİ�V?w�}x��X�%�g�}���bX�'}�;8�D�,K�ݝj���Gj�0Li6*z��nJA�8z����:�nd3�ƷJ�8��kA4'"X�%��w��O"X�%�g��u9ı,N��vp>~��,K�����Kı;�y>ܗa�f͔�ۙ���Kı,���!@�<��1��:<�>S�Z�Nı7����O"X�%�}���Ȗ%�bw��oȖ%�bw�ܹ{M2��͗wS�,K���gȖ%�b_}��ND��!�2'�߾�O"X�%���sS�,KĽ�ғ�]�I�&ܹ���K��2'{~��I���ׂH$���l@��'��ϧȖ%�bY���n�n�.�37jr%�bX��{���%�bX?��59ı,N���q<�bX�%��wjr%�bY�����ߗ��5�m�����u�T���"�>�N�8.X(M�xj�\YZ�߾��ﮘyܲ�%����{ı,���ND�,K���O"X�%�{��O"dK����׉�Kı>����6�ͻ�Y.fnn�"X�%��{�'�,KĿ���ND�,K��{x�D�,K���"|�L�bw=�\���sL۶�f�O"X�%�}�}�9ı,N����<�c�pHB �8�� ���C�R��%����r%�bX����'�,K��M���n�e�٥��ڜ�bX�'o{x�D�,K���u9ı,N��|8�D�,�D�{�mND�,K��'ے�4��e7v�m�yı,K?{���Kİ�#�{���%�bX����S�,K�/�վg��G��1��$� 9�6�	�H�۞�	A�\�;��m�;��[i1nuvb�"۱�JҳU��{��7���}�Ȗ%�b_��v�"X�%�������L�bX�{߷S�,KĿw�'�]�I�&��Ӊ�Kı/�s�S���DȖ'���^'�,Kĳ�����bX�'}��O"X�%�gt�vYw4�\��S�,K����oȖ%�bY���"X�0ș���'�,Kľ�>ڜ�bX�'����76�0�	nf��yĳ�'��u9ı,O�߼8�D�,K��;�9İ5
!��^D��{x�D�,K�{9��ݹ�i$ܙ��jr%�bX����q<�bX��{�mO"X�%����׉�Kİ{���bX�'���w@u���6h��g^�c��d�7\�=�}�8.�%�͕�?�	�iṈ0i���ı,K�s�Ȗ%�bw�����Kİ{�Ȍ�&D�,O�߼8�D�,K�w�̹����9ı,N����<��WblK�p��Kı?���É�Kı/�s�S�?��wbX�}�?�2��L�6Swnf�'�,K����59ı,N��|8�D�,K��;�9ı,N����<�bX�'�ٙs;	f�wf�m��S�,K?��
��8�D�,K���ڜ�bX�'o{x�D�,��P��~59�S"fTș�|Rav�&\4�ssM�y2�D̩����O<��3*d?�����?D̩�3(����yS"fTȗ�{�O"fTș�=����x�Ґ͞���wOzu��u��     �K��3$nX톻rݱ٣5����m���c%Cvݱn��[=��:wգ ���F����n7l���ur)ظ����V=���#r���Շ5�V�F@wK3Q�l�95ؕε����[=�V1�\8���]�ʗeo[���;Y��m��ݺAg7��^�%�5�b6}�4A�\�v��7���8X��;�����{����z���.��\���@l�ԕB�[gT�vM]l��:��r�z�w���WEƠ�n����s��{���~����&eL��G�{��2&eL�}����&eL��S=�;�<�D̩�;�<�sn�
l��n��y2�Ḍ�������� �y���/�xoș�2&eL���ڞyS"fTȗ���x�D�Qwq6&eN���nM�sn�I�37t��ʙ2�D�����&eL��S=�;�<�D̩�/��n�<��S"fQ���jy�L��S"w}���ff�7%���7��Lʙ>�7�϶��Tș�2%�~��ș�2&e��Tș�?��T[ț��ޛ��&eL��S��?�˸n�e�0��ݩ�2&eL�o{w��Lʙ2����S�*dLʙ��|7��Lʙ2�{�wjy�L��S"]��}�q+���a���lrN9є��iΜ��Ȫ֥7`f��n�;��O�~U�\Ѳ���ͻ�~��S"fQ��5<�D̩�/���x�D̩�3*g��v��� _}�ș�2%��]�y2�D�=ߗ�Qwc\�����?����<dK���'��4I
�1]��婑3*g���O<��3*dK��ۼO"fTș�w��yS�ڛ�2&gzS���&\4�ssM�y2�D̩��}�<�D̩�/��n�<��_�v��}��2&eL�{߼7��Lʙ2�Oz^����K�����ڞyS"f_䁱3�}��'�3*dL�>�����Tș�2%���oș�2��yʜ���ڞyS"fTȟ��w�.�y�lE�����{��r����S�*dLʙ��|7��Lʙ2�{�wjy�L��S"_����y5�i����}�g���ح�7*"�'6Ӡ��-vJ����$�͎��{����6�K�fyS"fTȗ�{�O"fTș�3�s�S�*dLʙ����ș�2&e��Tș�29x�pʠ�$�ɾg��my��3*g��v��Tș�2%����'�3*dL�?��O<��3*dK���'��;ܧ���w���'�Q��Z=���L��S"_����y2�Ḍ�����ʙ��Q�A QD1T`<V�����/�y�O"fTș�3ﳻS�*dLʙ���fS�L�6Y�w36�ș�2&e��Tș�2%���oș�2&eL�����ʙ2��bg���O"fTw�Ow���/��J���{�����̩�/���x�D̩�3*g��v��Tș�2%����'�3*dL�?��O<��3*dK�o|����6�4ۛp�t��vsuh��X�b[���ǋb�t���VG-�C�]�=v�n��7�Os��{�}��O<��3*dK�{ۼO"fTș�w��yS"fTȗ�{�O"fTș�2{��n�w)w6�&\ݩ�2&eL�o{w��Lʙ2�g����ʙ2�D����y2�D̩��;�<���ݩ�>���i��ܲ�2�]���y2�D̩����yS"fTȗ���x�D̯�؛�3���S�*dLʙ���7��Lʙ2����s���i$�n���2&eL�{�|7��Lʙ2�w����ʙ2�D��{���&eL��\]mS_Q�`�3��g����ʙ2�D�{9|�nᛳ&�ٹ��<��S"fT���ڞyS"fT�|�����f�?D̩�3*};��'�Tș�2%���'�3*d�m{ۿ��}'Y��u� ���m��1�,��9�N��g2lp��nG��y+��k&i��f�O<��3*dK����O"fTș�;=�'�Tș�2%���'�3*dLʙ�s�S�*dLʙ���)��r�Ɗo����S��r����;����Ȝ�L�~���x�D̩�3*g����<�D̩�.~�sx�D�;��u>�{��o̢�n�d�/C�yS"fTȗ���x�D̩�3*g}��O<���!�Sb\��x�D̩�3*};��'�Tș�2&g����nd�.M����<��S"fT���ڞyS"fTȗ?w��O"fTș�;=�'�Tș�>T�;߿��&eL���ߟ�~EⓉ�xF�w��{��Z����7��Lʙ2�g����ʙ2�D����y2�D̩��;�<�D̩�1v��`�( R@�$t�׺n� @b�A��E�0)�S��`F��UqOq^r�j��&�de	! �6	v�ܶ)�c��|��A(����H��?#��5�O�)<������A�#��]C�єsy����L�D�I��B�0�#�x~�6�8.�4ڂ�$                                 ,�M&��۰����7bvqkg��J�h8�l�z2<8�n�!�q�zA�,��aq���6ݱ�v4j������z,�Xƪ�1�.��^e�ᬀ��]%vv�cEn�����v�:v��U1ɬz�v%2�u���n�r ��.HZt)�M����`[[Q��ĝ�x�����n���ov�Z[\��E������ڦ5�&�6���tM[�"1�e��!3ۀ-�ܼq��ɵ�oe�ܺ�@s�����"�UMuS��K/����cc!���nà��'��]
wP�^�x[�5��a�Z�
u���;n��8S^��rӺ$֒ݬݎ�:�'u�C8�`ڕ����R��ۦ+��K�e��:z^v��ի�Z��Mȣ����۪��hUL`��Y`*ݩlgtXk]e������ �B�ڱ��]���;�i��i^Ujګ����eZU�ˌF۷��e���ʵ�t�dg�	+���k���\d�]t0�#'�P*�JP�V@��%���c����:�E3��&�UK7UeH��3M��9�4.(q��[rg�$�"�\m6��:���l=��'	����5u�9�U��.��EPcr��"�+f�[J�V̛i$��"#��5L�����DlH%1�i�k"��Ab�SmF�-Z�`�'U�1!bI�jt��A��e]lF[6	 ��f���\qF�� �T�]�l�ӄuE9I��[U�v�;f���s$u�L�.�:9��*��Q��l�Yp���.l��K`�nr
,�
�2e������Oc>��T�n�jZ͡�����+�]�5�K��((��꒰��,�I(I�����.'B�[���*�����G���+T囂���.�nn[�%�8:�Q(_1x��N�<�O� @C�T�)�:�����*����w�﻽��~���6�     �ۥ�]n�v9KF��@��;N���'A�[���:����ԻM�;�� yJ�t��A��ض���rV*z ݦ,͎{F6z��A��3�p8�Ў˘�n�s�ok�����U=k������I �O1s�≠U�J�ms��C�qh�Ub���Ş,b�x�� �7]�2�&�n�Sٳ��wy�W���7wwwKs4��˦�F�^��WOgF%���یsVj˺��`�:;�����d�14��w���=��fT���O<��3*dK���'�3*dLʙ�s�C�Q�T/���Lʙ���x�D̩�3*}��囘m�͛M�fn���2&eL�}����&eL��S;�wjy�L��S"\����<��S"fT����yS��W���y��������i�.�`�u�����{�&eL��?���Tș�2%���oș�2&eN�{��2&eL�}��ǿ�ܧ���=�������iK�JОyS"f_�H7߾��y2�D̩����yS"fTȗ�{�O"fT� �ڛ�s�Ȗ%�b}�m�e>�fl�f�ۙ���%�bX����'"X�%��G=��o�Kı/�϶�"X�%�|���Ȗ%�`���A	g���2N�t�4��ɧI6y���]��:����ᶩ�w�wviW�؍Ik0ۚbyı,K��x�D�,K�����Kı/������L�bX�N���,K��;ҟ\&�I2�ۛ��O"X�%�{�wjr��`"�E�"dK���oȖ%�b}>��'"X�%�~����%�bX�w���n�R�ip�sv�"X�%�|���Ȗ%�bv{���c���/����yı,K�s�Ȗ%�bw���w6�M̔ͻw.n�Ȗ%��@ȟN��Ȗ%�b_}����%�bX���v�"X��L������yı,N��,��n�۴�ff��bX�%����Ȗ%�a������%�bX���}�O"X�%���xbr%�bX��o�����7T�ht�����&�H�S����l�C��/Y(��8ݑ]��V�c=ߑ,KĽ�;�9ı,K���x�D�,K�����@���lKĽ�����%�bX�|m��2���t�s3v�"X�%�|����1ș��w���bX�%����O"X�%�{�wjr%�bX�����óL�6Y�v�n�<�bX�}�ND�,K���w��K )"�H������Kı/�{��yı,Os�ffvr�ܻ77ni�Ȗ%�b_߽��<�bX�%�ݩȖ%�b_?w���%�`|� �߼59ı,O��)��nd�.M�����%�bX���v�"X�%�|���Ȗ%�`�����Kı/���x�D�,K��>��X�v�_l���n]t�����5��6�\��2����N&�.\ݩȖ%�b_?w���%�bX=��59ı,K����'�,KĽ�;�9ı,N�Ӿn��3v�n��˛���%�bX=��59��DȖ%����O"X�%�~�}�9ı,K���x�D�*dK�}�70۷6�6��ͻ��"X�%�}��oȖ%�b^��ڜ�c���/�~�x�D�,K���S�,K��ﳗ�Dږ ����7���~w�w;��w>ڜ�bX�%���oȖ%�`�����K���#��H��B��tJ��=I��(��C�"�dK�s��yı,O}73�[�f�e�]��ڜ�bX�%��{�O"X�%��{�S�,K�����q<�bX�%�ݩȖ%��=������뫯	��$�ݛ\����]�FZ�Enm�N4j����n�����wM�mݹ��O"X�%��{�S�,K�����q<�bX�%�ݩȖ%�b_;�w��Kı=Ι���M�wmٹ�sMND�,K���s��>Ac�2%�~�}�9ı,K����O"X�%��{�S�,K��wғ�]�I�4��nnq<�bX�%�ݩȖ%�b_;�w��Kİ{�xjr%�bX���{�O"X�%�gz^���K��˗7jr%�g�2&~��oȖ%�`�߸jr%�bX���{�O"X�%�{�wjr%�bX���m�f����=�{��Y�����Ȗ%�a���8��X�%�~�}�9ı,K�}��<�bX�'�����z~��|�m�      �;^G]'-�q�0&֦jӣ2�n3���+6UC�:k#���6%s�����ă��-ۮ\�^�^�*���.����s���c��8^�0oh�Q��o "vс���ڻvT�3KK��X؆�
w/]U��\.���%l6,M2󍆛h��ٳE�{Vyۂ����t�wu��Ϧ0���ww��}��w��~~_���ia&r%�8����Dӥ������v�ֱ�H��&��nm�m���wMO"X�%����'�����Șf��ɱ�wEp"�84������h��h޻��������cJ<r6�O#nF�<�6:d��6q nH��Y�c�bm6����������4��f���m�a�JȜ� �lLrD�;�&�L	��r%�vڬr4M���J/L墹��5��Z4�stm�l�ν��%�N\��$��H�sb`d��w6&$���ִ�]ݗ.\��y���(���@�3E.[��Y��Y�"f&j��}�2<r$�yi�4������4��h�z��DV�(�QdI6��SU�l�`}��;�&�L��T"�7HH�M �m��މ��c��ؘ���y$�J��.'Gi��Di8y�/V�-�h[�������g��bncJ<r6�O#nO���h޻���W��@��6�R2L�.�*�3@�Kc\�Uܞh6�@?{�o��bE_b�������#$s4����$���y=r���+,A8�D���m���o$�~���v����b��4��M ��4��f��n�~�����b�)1�RA4ӓ@;�vGL��0�&�q���x�mٺL<U�f�W֗Ի��Х� ��:��/ph݉v9v��0���2H�sb`l�eo"��D�c�f�ﯪ�m�@?{l�=�w7�"ѯ��I�bBĸ��&�ɀf�L�0;y���u�iG�F���mɠ��4o]�	���s�~
@�T �;���I�yF��FI�CR'$�=�w4�<������y0���˓�$�E���t�l!ѭ��؜�e��t2�W��9s�Q�s�9&(�~#L�D�h��^�w�f�wܳ����{�qP;�2⋮*)s���rD�76&M��fٿx�}�ؾ�x�ƱI�NM �~�M��f��7$L	6�K����̋��������O�ן�� �����4?��<K�~���|�E�,�&ھ*`݉����ˠ'�&�L�#8!��s��Knn����� �  %�
`��ց�nza9��ipd�s�7n9Ƙְd�h�1͝�
6���{'^���7k۩J�'j�Ł���Ů����8�؁��ݣ.n�NZi!s�n�۶��6X�W(�8�q�Ny�����\����@�W��%��jQͥe���k(=Z�N���<]��x�uh�m�U��XX�@����Ny?n���i�v�لu���BWV3�X�N'��=�m��]Ө�zR��"G�D☐���^�4�u�������M���iG�����m�h}�7�33T>oc@��w��f�3>�D��ǎL�"�I&��}��~�@/u������[��`�i��I���^�^�4�u�y�����˾Ň�O�0Ȣrhd�0&H�nȘ�9ƒI*�B\�ծ��R릔Tn��Ugf���g �h����������\�TM_̓}�&�0� ��0;6�K�O$rdM���/��l�?y��f$�B��Va"� � ���p^s�-^��=���2H�5Y9�V���Ȓn
L��f�^�4�<�H��hw�nh�Pu��D�bBQ�4w,��Y�/���s1T�y�%��iG���L�ۓ@=���ϻ�g�~�h�@�<�uI$�$Jbw7^���;H�:s)6�ۣ��:z.I��t kt̟�g�wSoLx�D�I=��nhrY��g�"bPsy�*qN�ܙ�]Y�efF�}�,�L�I�}���n���XW�'�ӘdQ94$��y$�~�w����{�3��*@�S4��#� ��  \�����9������sp&paLA��O8&"��7��#dӉ) ���H�x�&�H�D� 1"� /᧊Z l#�s=졦�א Hā'/�\�/��!�S�S�:�)�tG�:(���(����C� =��␬_��8rI<�{��O;�ݺ���.�ۛw7w�"/������?~t�76&7b`vmF�o$rdQ���/��h{�h�@?^�@/R�$�y��k�d�A���Nm����[C�nHI�k�6��r�̽(�QdI1�ɟ�/_��^�4��?� ���s@�;����"n4��rM ]�7��������4��t_;�(�ərh�m��w4�z� ���;�&�1�dR
H��c���0	6&_|V}_]�_%(E�
��B"T�O�f��I?^����4�#L��&h���oY��Y�[�s@�}�裸BdJrc�L�$��{r�:4�N���[����qlQ����+��{J/��V��tޞL�"`L�� �޳@?Z�S��7�H��9&�~����#���0	��}��fzW�\�<�mɑ7�@���s@=����f�~�٠u�V�(�QdI1�ɚ��0	� �H�{������i��;���� �i!(�{�����$�����~��w�N��#�%?5FB0p"�fP�D���}��     G7T��^��:]4mjjW��;];ljNӨ���
��Q۵�<�\�#�.λ.�<���d�s �=��
�,lY�7����hR҉,n
�X��Pj�!��豭��f��@s�赌j�^6✶0nx/f뗩.eܗ:Ȇ�����Ůy�b�d:;s�sl� ����=7��,.d�Lٕ8�����/������;5��͵��\�Kը�<�m��V� ��)�V�(cM�cJ<m&ərh[f��Kc@>��9��@4�h	,��d]��#���I0&H�flLn����W�r��u�L�26)3@?^�@r��DMR�N���hWtT���i���ɡ���fx���4
���������b�G1�I���3@����ff7�? |�� ]�_$�����[���T�8��t��3��餺�[laԃ�Ns�YoS�B�����rdQ9#�/��h��h��<�����=��I�D�"I�LГ����TT�D`#�VQ� �4�1h8.�7�QmUVW�m] �L��0&H��9��M�A��BQ�4�Y���h�w4�z��;�%�n#�ۑ����y0=����0	�wbm�$d��h�w4����<��<�rD���$��er�&��[j��v^�c=��2����[���n�jtJ�L���6��9dlRf�{�Y��f�~�,������h
�����nbĢrh�@?{l�/��h������A��/��G1�G"�I�sy�/���f����f&���� ���?^˲2'�92(�rh}�b���i�n�&7b`�a�8�Z�YLprf�{�Y�fy�/��~ ���h��hg���I&@h��9:TKu��y�c�"���$vM��{a=:Ѯ-��������69�I	G$��}����4�w4�z��q���Pncr'9ĘrD�UvzO:`�ɀL�0;�6�2c�dR
I�^빠��4uC��@>��@�QJ�\�Y�V.q_0͉�L�0䉆�������:"k��o�ÒO�~))3�B.�"����4|�h����I�hf���U_U֞�I$�9K�$���*K�nJ�^��e�F���l��懑�[ڔ��]�w.���#��.�f�Ɂ7c���~��>ﾚ�\�ddl��ȣ�ɠ^屠}�4|�h��7�}>���ɃM��X�O �������wnh�>��lrƒ�I�$L�"`M�釮�g�v�s�m,I�r#nM ��@��s@=��w�I����ID����� fN���o�m�     �ת�e�Vk�l]Ht�家��wi_4r�.�N-ڷV�g&�|$��Ԝ9�`����'�F�	yegr,����nptp:�P�Ʀ����le[=cm�0��!�n;e3��-e��8���@iT-�5M��Gj��	�q:R9�e��G:܉�·��j�ng����L�؊Nu��26�F[�d����� t�z���X7�mtF���\M����N�Ik�!n�X���E�m����dR
I�{�WL3b`$L�"`mʹ�N|Z�B�%�|T�36&2D�;6&}��9�"��������$33J[�7X���`�f�Lsb`�\�Ⱥ��Ȭ���3C�>����f�����36&3b`vmF��
�%J�8�f�L3b`6&ܑ0�����_��vmwXI�Ȼ���N�x�SN�����!�7���r�ZZ�6Hb9]�!%] ݞLf��;�&ͻ����:����	G$��Y�?�ꪗ�Xw$L͎�f��̮.�ڏ��dmɠ��h��i�bGu�h���@��t��C�&ݎ�f��&H�rD��qV��S"��'3@=����@;�&ݎ����^�<�I"�Ic��v\n��X��s\N����Z�j�M���,Sq������p#_Ͷ��??/�?^�@��s@;޳@:���Y�!qY�Z�I�w$L	�0͉�Om��՗b�9�����/u�䓷�{���H�)���"��3�V�L�\�<�� m��ťyuYw��UV^efF���vӽ }Mր[�h��h�����8�$,Q���%Z�������4�ƀ�r��?g���\��iuu]A�d��[�..�� ��<�g�փ��	幤S#iŠ��W���h�bM�9BI4�w7鈘���N��7Z �,�T*qN���LP�8�������Z�޳@��s@�[����s(㍀L�-�I�0&�t�+��W�类�}z����sDq
5"�z&ݎ���0	�%�2I|i$����.���إ�Rk�R�6N�r��;���n��.�d��������#_m���s@��z}V� ���/��Ɣn74�r)3@��z}V� ���/u��;��'SmH(�$,QǠ�J�.Y�����i=��N�}���J<rH�FӋC�<ľ��4���.W��)�ց���Q���,I	$����\���ۃ	;�{��S�B�R�M�q��3���'�O�d$%
3��7��燄�2҅�s
3���z��ׁ�	��u-D�x<ދ�瀧 �>��«0���� �2�E��JEc??���,H�z���<<�V0�����0`�=^�Җ�|p"S@��c��Hy;�������6٦�                                 ���v�p��C�<�*�u��fa��`���r&���)�6��p�f�4��W;����;n
N�'(f�����F��wbl�dN��1]����gf�JJ�l�z&L�<�<\L�x���V����۪q��.YW���R��u���N�L5r璹�����aG�@���6��"6�֧v:��H�����p�\6絻j��ݥ�^` ���hm��{vkK�Gky)_/���q]���\<ai�lѮ8 *�&�M��gw7 F.���'Z��Y�Q��\r�۲�ۑ�Aר��L�&�λ�WF��l�na|�U�v��֫���:7i���$T��&����UK\P؀^T�J�gD�Ϝ� �cn�1F�p��,f��a�i^��j�� T�Kɓh��-K��e���F%1�]�8 tj)�ڶ6�}l��t��U�pʵI�<­���i��4�n&��ø��yk��#�ʙ;4�]��u���,����t<�a�ԨAD��.���u:R� ���I! ^�^�7[��u��v��p]�)pザ^e�h(�,WGe���86�X�14V��ɶ���n�]��T9�7A��d:L���6:�Ã	�+{n�H�������κyB{u�����^��v<d�!!Y\����b2gt�ёB\�W�r2��K=��ʡJ���ŷ�yμh�ftuY�[��9���.���=����Yu��m=r�ۮ�+�s2S��b:F놴��Kg\KM$�A�m�����MI��l$HuMT�qUI2�@�!�jd(��tm�`)Nf�qT
��n�i�5��Q�d��bg(���C�	@�Ti�)l)s\�m������'QOP5P:������Oc����N1D_T\T_�.t �K��OrL����     	8��9"q����L1������ێq���b�9m���M�ֲ��F�O�����]��k�g�Ʊ�u����+�������6�a��9Bw9ov��.v^��a���]��9:5��:�ҦY�9�Kd!�&nuA���;���C�P)$��n.�����b9��;Y[��v�	�U�>lҷ��w��w�ް� �N��B�Qƍmͮ��[��g��;ax+��[i1nbC�I�7���$ds4U���9V�%�����������Ŋ8��*��h�٠^빠U�^�u9��s�8��"��Y�.屣����t���ց�*����̈o#M�4�w4
���*��h�٠_Gk�(�iA�ۑfF���^��bb��~ |�h�o|�{��{�������X�i�g0vn�M]qK�gC=�odƻ�-���a�0���ą�8���_m�{��*�@��|�4�� �b�qi$���y��v�	6N�;��v��s�U�j�=�ě�&H̍A�4��hwW�U��h�٠r��u�F(E	����
�:� ��4�]��a���a���qǠ*��Z������'��*�W�}�m�5�Ї
GM&�yN�kȵ���S�[=F�;s�kV-�S�Ӥ}79��rĭ�L�0&lt���9諭��z��-߾Y�lS#�2!��6��/�w4
���*���l�/��ƔN54�p�f�Wuz^�V�����+EQų���'}��9$��/��ۙ/"��*�����s1N�N��y�/��hwW�w������)�1ŠlL	�0%͜`K�e�2�s�@��U��1�I�#�1�O79&kٴ��K�t��-�:�iła�/�lh
���
�9S���i怗ؾo��1�D�����ؑ����怾屠ut(-E�]�EEe���
�9V�/���>Oc@t�� ����yC�$Z}�h��xrI���I���EQE��1>�i����q�YqyE�e���h6:`Kݜ`K�e�	�&$����}�RZ[��.ʵ6���uڋ���y8�w[]A���(�d�A[IW@���0%��������L��71�1!b�=�N�Ǟg�@���'��*�W����tZ��X��LQ�- ����/�w4
�W�U��h�bM��#$D��M}�c@T�^���hz&bg�w�?f���������"d��f�o]��NU�	r�}�c@�D�D6���     D�/kSd�g��'7c�\��/T��!�[��I�r􊹧o�~�?N�{X���K�v��9N�Q��N8�����V��0V8�r�y�6.�n�b�\EQ�%+Փ��-��m�s*��j�q���b��g����wf����N�	�<k���B�][��]�N���ۭ�#�z��L�WtX�̶V]�W��{�_� �Z��n�u �^n���U��-�l�x�X)Ŋ��+b���0�9����8���|w���@_r��&c�I�h1]\�Ȳ�/(�%��2D����n�L	xl�� -����ۦ�m������I'��.屧�j�p�h��@_��(�j<i6�$��]��N�@/�����_�f��;�����8�$*V�0%���f�L	�0߽��������;��[���uؓ�8
�x��Y�k�]��J��7�^f�'�͙Y�^W���}�c@K�É��Ǟ�?���h�D��1Ȣ$D�%$Н��xs=IDTEj�D�c�L��s@/���z���[��1B(H��h�������<�c�3vy{٠r~��:��ົ��*`��ld�����7c� �Ni�\�<�!�F�Z}�h��6{��='�0��s�ȒIQkq����Iݫ�n��s�Ѡ�6b��z]U�\ZU&��Qt�te��������n�L�{-�L�0&������Ɠo�4�w7�y_��}�}4����;�'��6�9����O?_{y$����%/'�B�
$��h
�s�p�y����w�:�4�$����qhx����@��ۚ{��ޮ�@��7R(��|I����Mؘr�[ �"`g�}�'Y�͚�D�'iۮVX�Asȗ��Ӻ�0��p9)"���w]�z4��R���Mؘr�[ �"`w6:`r�0�<x4�8��ޮ�}Ă�p�w4^���O���8�J��V�76&͎�݉�L���[�sb�D8G��ܚ{���hy|�3ɞ��@�;\iF�q�I�"�4�Y��j��@��s@;���$� <Pcd��X��z��\S��Pf�y����'�����jطSQp�M��F&�Drh�Z��l�/u������ߦ�ݎ����$NH�FӋ@-�4�w4޳@/�ՠ{퉷Lr)��E!�oY��j��Y�r��u�F(E	��y"��y�����,�r��9{�qG��'�}V� ��0&lt�&lL	�}[s��q      :�s���m�{�	!0�X$˴'��\�W<o&zw7h��c��5.�=8��sNƽ�7`c�\�j7�r7n�^IӶ���%9�h�s�D���;\��0d^(7(ض͒si���z�n�R3j �!Nu���۫��
K�(�\��M��hg%�n0f�ٝx�\���D^�<^�C;����l�:;2�L�{w���������N��W��[�9�/F�6y��,�m�*�Np�e�����Dq"�H��M��c@ܳ�3��}Iրڇ��\\�5F��h޻�}�4��� ����y�G�?�pj7�M�I3@'� ��U���'���4�؝m��7HH�M ���@/�f�}빠޳@�q�ҏ$����|V�&lLU{g�] ��&2�[�~������j�s���抱!\�n�^�JAn�m�0^-��g�ktp������L	�0	� �{-�Lؘ�*�~�BFG3@�ޯo�y�3ё3s Պ�rY�/�lh����ǃN�= ���@/�f�}빠U�W�Ӛ~+1�G1\e�Veh9�����=�Wܯ@˪�-칲8�9"j<�7$�/�w�g��lf�����~�I$��\���%����qs<�t��%�3;�׆z�V9R--b�$�O �����׳�`/e�	�f�L�ͫ�m��7HX��@/����Y�_z�h{���>w���d�8�qh��h�liq��3 L0��:p0=/3tMj	��
i �][�"DN�<S���@�	A)��aF�$�$!!�HI##�܏� �=(��=� ���Ŏ.��#+B+@ I ������P_H4��Uz~ ����BF��Ԫ��P<�`U��I�5BH�RA?*z!��@GU��Q���j~ �^�W�U=PN�(hht�g D����� 꺭�lM�cd�d��RM�]��z� ��V�_z���[��1H�#q9�^�z}V� ����������[�I$�D��c�y�-s�umѣLF��@�]�yk��WVx�-r�\`�(��ӀF��ܯ�@/�f�}빠U�W�Ӛx�1$G1<�UfV�/�f����'��:��@��h�\�8�j,�7$�/�w4
������ ����v�5�G�&�$�������r�- ���O��"6�a?�Nw��I=�Ε��r6�Iq��uZ�����~�W��;�$�I�Nc�R[9���[]	YiH�э;��:[<�g�օ���Q�q2H�m8�޳@/�f�W�� ���@�lM��d�d��]�h��k����sw��:�ܳ\EP�û��e���y��:��@�ʴqT4�h��@��9EcǃNRM ���@/u�}�4�l�i�<E��(�&E�h݉�Lؘ�N0	�������@��`��{=����     ۜ���n�O*L���o|���<��unwYu�l3����GMl�ڻ�S�.Ona��]P:�g���3�'�z4��sзkd�@���2��6{F�Xf�6{h��gv@�]�[5�u2Qãdv�E��/B�U��S���#Y�qn�S/=�:�f�ˢ���hB��I�<9:��c�#�v)�^{���v�����^�e�v�A5��R�U�9�aKcu㞛 GSWY$dx㍨�4ӓ�>��4�l����Y�_Gk�Q��x�ڂJ�� �{-�Mؘ6:`o��N��q�ؐ���}]V�^�4�]� ��4�뉢��⼻�����U4�h����Y����ě�&H�H����/�w4d��L���&�L�9I*AL`�I,P��nmv%�/^wC=���]�<�Q�d$��m����s4�l��r� ]��D~�|�ƁԠ�8̘a2�n]��w�����V��kg�^빠�f�{Ni�,ı.++Wi[ ��0&lt�&H��uZ�칲2<r(�X�ܚ/����=��`/e�	�a�8�Zn516�$� ��4��� ��h޻�"��$�x�#��΍Ƭ��n��^7O3���;z��9�C/.'��BĤz}]V�^�4�]��mz{�u��	"d�8�qh�Y�&bf�|�ƀ뛽 _W*���{��H�dcrhu�s@����'�R� �R  DddA0I�"b""�������E+�re���U��h9��w�ހ>����f�}빠z�:�c`4�����&^�`g�r�&͎��}�$��w�~��~ �+�s)7M�`��7+T-f,���nf{[\Z�l����#ƕ]ծ++Wi_@='�f�L	y#���U]�$���)1��4�-�qT:��@Ru��f����G�?�pj7��P�f���z~�U�������@|�Ɓ��}��*�q<HII&��g��b_r�- �ߦ�����$�X�;��7��'��}�r�����iŠ���/�w4�u�}]V�{�vI$Ɂ�7���m7Y�D�@�ް�&��E�M��ۭ��Y$r21�4�]� ��Y���h�z���[T�(D��;� �{-�w6&͎�{Fr1�s	�p�����f�y�%�_�4zύ�S�x�1,I�b�v����������=��}W~�~Z.W>�##�"�LbnM��i����t�s��;��U���: Eu�Jh��7n�n      ^�?����D�:�p:���3�aS�����Yi3�͒\g���؊|�tk��!�u��ݣ����F��k�$�:�c1���3[`+�ht=YEBvN-�։jzס㭓d��n���f��}�y�[M.��:p`&���h��H-<v�R��T��\�˰��3��N�ۧ9�N7_h�쳳�,Š�I��˽�����> {��|��u�Q�Ll�+�]�m=�v�i���kk�����S�F�Q�jL����@/�������<���nh8wѸ�n.U�gC �{-�w6&͎�͔�;�k�&�����iŠ��4�]���)���h�Ct��Er��s�0&lt��j� �{-�~���9Z6�cp�dN9��zQ�L���;�f�LeȒI��<��M���][V�U2�f�E� X�5��etsv��FxA�=��m��/e���������![��\��6��I��{����Q��*���|��035A�L���_Uٷ�s�2<r(��&��>�>4����_WU���4��pj7���q�0	���sba��������.p�?�q8�O䆀_WU�͉�3T�P`z������IW��@:�j�x��]�鎕�L�C��I��J�r��C�[qnE�P˦F?�m�?��f�0;����m�&��rnDc�ܚz��o�gޮ�@?{�h�*ڦLnL�������N����~}��"�B#<<�3��ݳ@�Қ��î)��⫾P���l��0&j�V/z�ƀw�V�#�bN"�H��ܳ@s12�k?�,f�/��h�o�v�9�!�4��ie�i�KԐ�����˪�뛒���.5�w8h݊�i|�L	����j� �{-�w6&�v�5�G�M�G��)���h�z��қ��fy�9����N7Ą9!�r�- ��Y�_zS@��Jh�>w�����iŠ�ؘ5A����ꤾ��*����U�y�����}�D����CȠF7&�3T�P`/e������A	��\m���dM��\g��"V��L㋷f���M�-�䵇CV��0	���sb�}�}�v���+��Q�s�I ���~�̫�͞Ll^�P`
�_*Ȫ���J��V�;�f�0;���/���=^���q��#Rdrh�P`w5A�L���;�a�S��ƣƒPn�zS@/�����w�N��{9$����# �z@CMH�B ɺ:�p�����b�F �A�~R�$�����'��TL�:(�4�A��b@"Ł��Dg��x@ A'�Q*g���?fE"�B�M� ��bB)#��!��D������H�VO�`��Kse44Z�*� 2��Q"��G��H�)9����>O�R�u��JJ�*�$'9�0�$H�m��S���!R�?�_�<9秱�8c�F��D�u/ �V�8����X	�R$H����,B# �	�Y* ��x}��E$ H                     ��         UQ���
����^p\ٞ�)\VaB등n����g��d�Naz�5�u-l-&SH<�v�v20�P9ќ`���C�%�R���1�<�l��BQ�v- l\L���Yn	��<>�9uCxr�7}��	���a]۳i�Ī��H9ce�e�cfu-G�Mk7gvO3κst��nS�YiS�8n��vwA4��U�ʅ<�춋Wj�v�dǚ��Sk��r�lpq@[mۦ^K�ೖ��!����^[n*UZs�`'�1�Y�Ydu�jA�:���h������Kw`c����P��j��I��Ș8tD�ۥR�ӝZ4�.��h�Y,��f�l����1��7U��rUJ�����6�L&ԛe����#R�l��,��ݔ�v랪�� ��u�x7uBMN�	(
�%��T��ٕ�)T Us �Q�$�nʖt��@v�Hl5�m��J���X6<��F^R�h����Z��s%�m�d�t�n�u�L��y8iBß����1�2���D�lJC�n��^�r�`�q�v��'oWA[�ں�`���V�)�v�ki��+;�[HK<�$���`�`�1����[Tk�Y6��)ڴmQ��(UZ��zpc��`�qr%[/cmGdi+Ĩ6Ť��9x�]�ѓ-��sl���֍�خ6I�z��]'��ۭ�����-�64�H+��	�]���
�Bz�jn\B�ַ���P��㶸��[r�1�&�f���m�[�q��=:y��=gŹZ�m��k6�m�/}��O��X��F:{$�y�und��삼�pڍ�i�n��'����9�/ P1U�j����p*�vƫB쁬PhO;{����ۄΰ�J��Eǋ\pslݠ+�nK��(���<my�j.������# �o�
׃��:��|�<?'��D4��@C@=�
��~S�P��N ���띳w7@     Sˣ��׎��쉣�i��C��Ba��g�$���`��6��6�G�;��)tV����HvM��]t�k)�uC�+�3�	�<�~}Q��խ8]t�D��n�u������,��۞�Z4��+�x�nX݂�f�ű����֦U,KhI��1/dq�Gn��zu�d�xA��8�]���3���%ik~�w�w��/���7^��s�z�On{sW3H�a������FBĘ�/��6�n���n)�x��8p�+����f�}�M��)�w�>��$R6I���l��0&j���e��}�y�G�X�܈q(���>�>4�v#G15C�N��O4�J��A1�A�����M ���@?^�@������0�c�4�% �4��ٱ0&j�sT�{J�v��hwTs�p/F��/e�T�����F/^a�Y��Q�Wk�
>�vlL	�����2�[^^�r8�ܑ�2	�4�Jo��<ϳ3̞���K�4B�<�<"���N{��9$��_�$������G�?���q����zύ ���@?^�@������]���q����}]V�~�f�}�M�������٠^�߱4�R6L�8�r��f�0$��L����3��:L��M,�d��F�8.��f�a�;����mA�V3�5�8�BܴfՕ&�P`I�� �{/��v������i��	�B	�9!�[�s~�<��N���@_v#\LL��QԠ�}�c�4�%Nf�}����f���}j'�������NI>����{L�"�Kp�JE��4�ՠ[n�^V��G\�L���2
���ZU�:���� �7Z ��@��l�I!�S Ld	���j��	�l�Ŝͨ��=b�ʑikM�Y��nE�[n�^V� �٠^v���ƫN'm��(���ՠ�4�ՠ�4����iH�l�"q���m��j�m�yZ�}�T��C�DH9&��ҭ I,�ԕhTL}S�+[�0 c��;����y�:a1�A2(�Zm�@/+V�[l�/;V���ݒI �sWm=�t�1/i�k��m;U�ql��\�OWW<u�LN)&9�0cNbQ����ՠ�4ץ4�f�{�sOf%E^�e�ehIf����汚 �s@;��h��Ȕ�ܑ�2`��@���	%�:�u'Z �y�/�Q\�G�$�7 �٠���f�yڴ��q��lƁG&�^V� �٠^v� �٠?>>H2AR�߿g�ff�����    .ۧm�t@�v�K�[��P��eɜ�q�d�[6�r�	e�u�:��ɉ�������/v�)�1#�y,�]���>>��rW�]խu�M��m��&7m�9l����H�	C�	�θ���<�����gF%��f�Gl��[�AiS�ٔ��2I�V�e�Y�g /3��g<�L�a��|��5ٵl�wL��������d'���lS2��te�<��VX�C�k�F��N�Kg��x��;�J)t�2�}�߿�����ՠ�4�h�Hڦ7"Ue��f��ҭ��D�Um�5O��7��1"��O�	�B	�Fհ{�Lm�lIo$�opî%0`�ƣqɠ��@-�h�*�q3T�y�	��(yTU��R- �٠^v� �٠��@���$�dx,�<��<OрK5�c)k�^�l#�W<n�s0tFG2�l]-I���j�m�yZ��f�}��8�j<i%�h��"g�bb$�J�V�$�h�*�;�����f4
94�h����LU5mր6�h���EXfe226�Zm�@��Zm�@/+V�ﴍ�c��DH9&�y�lI �r[ �D�˓�$���1�u S"n -���Q*��K=��p[��͵qS�a�mrtv��El�$�o�^�^V� �٠^v���0�L71��rh�j�m��j�m�����T�X�jE�'{��$��;�ɊX��Z�@�1�y�/<�3[M ����]q�L�Ȣ�	�4�ՠ�4�h9��������Ayu�TeUV]�V�[l��ՠ�4�ՠx���va�'h��i�:���v��}�b7�Q�ӛ�K,�+�25f�.��@K4�l9���@6�h���jD���N- �٠��m�@/+V�ﴍ�c��DH9&�yڴ�f�^V� �٠Z�mY�1�A2(�Zy癉}��4�n�$�C�dA3=D��È��EN��"}y痒OoHN�˥��E#�@/+V�[l�/;V�[l�;�[�$�b��2I��q�M�]LFf�n±P:��k�kV.�t���;�8(ԋ@-�h��@�����ʮ��F�D�	�4��V�$�9��ST�Sn��D��Q~k�|�8�"ȒQ��W�|��������Z��tn'���ے=򼩠r���}V��%~��{�;�!�I#��(h��@k�:�����u#@�s1�7��'�m�      xѺ/.��q';���3ײu�nCPs��[�gYú7'\�N84M�h�J]�;z76�mڃ��k�;�Ŏ��l����zL�![��L9�G �;��N��n�D�t�دӜ����W�[�{d�WIW<nP���Qѣ�Q��9���j�����ɏ@��\d��&w%��e�;D�+���:��y�l�/{���7�#Xkeѳ�v�<mu�U���mg�u6�Js:��U�!�uN�Dr�S$�����������u#�3��Sn���ݼ�� �n-�����M �٠w���?.�:�9��s	q���M �٠w���*�� �e;���1F���4��ZVנ~W�4޸৑�$łrM�}V�U����M �٠L]�j����Ϙ�rn�0#��$��챺t��R�ms8��	�ْ���^��� =�h�7w��3m��9���qȟ��#�ם6��a�y�9��If��_*�$�}3T}Ы)���28�6�4��h��
��@?^t�=�,�rh���$�;��Z����֍13T�y�Z�m�<&57�F��*���Ş���{�Lsb`��I$�J�X�9�%��W����Fe�Y�)��p=r�c��n�9�&�$qǠ�:h�� �z��k��Qc��,A�J7 �٠z��k����8)�nDI1`��@:���v���N�=�%Q%٠8�
QZ?�o8p�B*l8��)�P�S4A?:AHc�5́��p(��.����"<W@'�I*��5�6�H�~���	��J_ b:!���b�0�I���OE^T��!���2#Q�B8�)�xs��θtB�3"O�����B0I�p��G��+É!��X� @��x�Q>+�h���_���h�O��"#�Q���(�P��<��?23��M �٠uj��5�*�����s4�z ��hIf���<�+��h����N9�$z�y$��lؘ�`e�>���f�'ln�u�#�&�0X�e.Cج��ؓYw�<�N��앝f�.��톀$�h.Y�*I[��@7Mր����#�#DmF9&�[l�*�� �Z��f��sJ����27���`z��q�Ir[ �D�$�0?.��
b`��Gzj�h���I;��y$@=`�E�H� �*$Tk��%���g$�ϡ�L�r`�y�(�Zm�@:�4
��@:�V��y�y�{ҿ��Li�28�q!�4�iץ�m歖�=�)���uu�8�TH2H8FdnE��NI����@��zʒ���m���T;����*1$���VנU�@-�h[f��>N��qȟ��#��ՠ�4��@������5	"�3*2��5M�� �y�*I^�u�M�dn��@�DیrM ��h[^�u�M �٠fvfa�U��*�ܜ�Knn������    ��l������`�����'m۵�Z�n�n�ٳ�Ы��lܷ���F�휎%��n;sأf�� �\c^]~�;�7X�lFL]f�"틱��pm6 v��mq]�I��e*xN^�Wk	��hq�.7>�[c��m/�ڸ(�ZndJ�ck9��s�t@���u���i�h��H����{����w��g������SVM>��M�ss��	�1Kչ�61�۵kcf�-ёg�c� �A9&������:h��c� �y�}J��*�� ̼�� �Κm�@:��V׿fbĀT[������*�� m��\�@-�h^t�m#29!��$�͉�I"`7�`H�Z.Y0q�E�$���Vנy�@-�h^�@=;��I2,���zT�I����:n���kCnVv������������q��CNI4�:h�� ��h����QT5	"s6m6�f�I'{��:�=G�Q��y�K4޳@-�M�dn��@�DیrM ���m�o:h���K���cP�<�rM �D�$�A�I"`lL��Fϋ��70�'3@:�[l��f�m��ٞb����I$�	&��F�������1��3YǗF]�⦡gs�m�KH�;���0'�y����}���f�m��ם4ڪ�3#�I��Lf���GLf�IcE��8ԉdi"'&�m��ם����F�� ~H���W
A��OT���}��7�I��~�I=��tn'����nf�u�M �٠z� �٠w��*��$Lx�Ww��$�hbf"�O? 6�h^t�9�$�`23"�A�5V�t� ]uF�<�k<��/�nm�v��t9�g��4F�c�h^�@-�h^t�m�sK���cPDy	$�m��l�A�I"`6&oh�gŬL�E#�@:�[l��f�[l�i�,uL��D�p��� ��4$�Bf&T�:DĒLJk MSЗ�w99$����r빻�n�x'$��f�[l�����$���ߠ9:nB�軒oWb��e�zu������W�@���]6̔H�ɠ�4�:h�ϼ�3<����_��kU���q���9$���0	$Lf��$�07+m\CP�&7����4�Y��dD��� ��h�2�E�^a�q�u�^fh9�M<��� �֍ I,�;��ݞ�#�I$�m�˭ �Y��f�S11�&'詉�w>���|��     M^�M�Vv�ݽt�+i,�|����kZ鰖�]l����y�Np��!�}��.�*iŦ�so�k�-���Ŷ�al������ݘ�e#{*a����Q��Vܑn[]%)���7b�Z�&S^�X�WciÑ���5���g�mzsN^��t��:5Z&��.{X;i�i���%��ۖuC::�:�����y�{�w���߀$�-A�S�i�uȽ+��[��.�V�m�=��g��v:�\1Wn��9��r~ �|��4�Y�Umz�3�����<�Ȕnm�@:��Vנy�@-���29!��NI�z��k����4�ʠH�F�"rh[^�u�M �٠z��|���q����#����4�Y�Umz�y��i��I&%��MH���;\ga�d����Ʊ�vyw �t�z�CD�P�&'<Q�����h^�@-�}������r'�<�@P���&�I=��b��E"��<T>X��,A�@��<�o�@;F�$�h��wK 2.�Q<�rM�k����4�Y�~]�_�1�25zם4�f�u�4
��@=�p��0HO �%��[l��f�U��^t�>�33����I2<F
y#Px{v��.�-�n���+����H�O#�I�䟀/��Umzם4�f�բ�p$d�#I94
��@:�[l��f���:��q����#����4�DA�U@ 1R��\���{4��W�~�UB8���F���[l��f�U��^t�/vD�0�A(�"$�@:��Vנy�@-�hٞg��_�I'��fK�R�@[uu�qN�.�ݦ;r=v�F+��vn�6�IjL	��D��?��u�M �٠z������4�F��@:�[l��f�U����:�y	�(�4�f�u�4
��@:�[kQ)�nE��NI�z��k���3�b�t"�(��0X��0?��^}���'�L>>p$d�#I94
��@:�$�h.Y�zb&&�C���̚3ɖ���Ѽ�73\6&�=i�[<�"�Եڣg����n68�n'�CnH� _���j��bDO�M��>B���a��e^Me�� �Y�b"�Mc4M����y�[�?���	H5$��ύ�k����4�͵r"�
ʸ̼�4��LE;mހ&��@-�hzS@��.�)�ә.����Z4sm�� ճ ���$�� ��Ҫ���� *�� *�UAW�� E_� �UT�A��@H#@1�E a@@�@����DP*�@�,E `
1��@�, `"�P(@,E b*@*���*�
��  ��� *���*�UAW� U�� W�� E_� � U�� W�  ��� E_��PVI��\�4�h��` �����Zo�h   T�      � @+Mj����         �EB�)P)PJ����
     �*	BB� �(EB�R(
 `    ((��  �P4���s�RŸ��:��,��ǀU9ʽ͋�q�֜ڧ��'�>8��T�}�t�Y� i��1S�PN�R�7{���5���  �  ��V� ;��s��sj�w ��<> �  
� c�7Y�T�O c��9��M�x� �}<{��La��T}�s�/���F-�i{������k���mUgTnwה�o��͐�s�><'����*�\�˛t�=��>� |  
 ��� �}Yq���WuW�|ϾgҾ��;�H� ;0(��;@� �� �� 	�  � � 1AL�X�� f  � 0�   "z �@� � ` �@*�  � � {��@16�ك�� �*� ����y���w>Y*ũ_��}��޷�o���� &����{����B�t�/9�ͺ�g^����{��y�[�����rw}t���_y�+� � �  �P )�O>���=�}��*��i}��xO� }<����[ޭ���ɮmOy�N����\��'�K�W ��������|xNzzr}�����֜�w�����<(�%�����-�s��}�u�� zB��J�  �)�����J�  �=U*�C@  ��U*M��� *�Jx�)P  !�)" ��>�?���i��������;;��w���dTW���E@UuQO�E@U슀���*�T�"����,;����܌��}/��0�<��,�k!FdH@�d3$�)pi�
�
�
�@�]�4��'9�_��a$𘒒�0�21�Q�1V,C_em�yw���s����׫s�{����=��3}�쎄��@��CHs���(]�חc�#T�#L�ǁ���I#���w���$_�fB1&{�<�=�bFYW8�k�sώ��IF�� ���θw��p�������O>�<З���u�<J���%2V�S A���QHA2	H%	Yy�.��<�d;�(L�������3�yI}>�#~C��EhF����
4�s<�V$|e0b�`�"�p#C�p`Q�P�� ����LH\aL!P�=E
��|���}!L��7YsMe�6\�apH00ЍHT�Is���\Xԅ1�p#R�)���F�i�.BᱬB81�)�.p%��.�!�	LIL!L�PGӌL
�R�R�����!X�P�I#YBH�FH�(�XR�#F�Sr�;!w���<$
��م�;���0`q�$�&�%(FҖ�aL��\��XҘa
��3	q�	k�XG�z0���i�A�BI {y�O�s�6K����f���<�7	�g8���V��d�=t����d
)(�
2�	p�����C�W�41��|BS��4 C� �;�~��a��"@���!
�	$���D�ԃW���!~C�P9��yot� 	��"ōee�NN|�|�2ß}���&T���*��V�R���UQo�����xL��sxp�/3�q����x����)���w6oq
�_�^>�G��E%�P�&��62f�B&�}g�==��5����20����sB����v�d�yD�(Hh@g��E�$�����*�^���	q>�=�]Ð�\�������o��	�C6\	y�򞙃 D��b@��H@`F!B@��0��}�M�Ys��]�� �@�Z0�b�YK���M	����B����_d��J���+(Fp#bD����[��i��{�;��hRS�L;�f�HCHP�FVXؐC@�$�/��sy�=�w�ad�>�H��R�fʵ����W�0 B-*QH�s�3lߏ��s�^p���!��5aX@�b�CQ����S=7�}�^��t�7d!q`P��@�B4H	�"�"�1 �"T�ЍIsy�.�y-�u����#���߼<7�48�F�4�F�1h8��'�		�F�B*HZV�R�n���0�4P��t�30���,�'���4������ 1$
$B,� �,B#����J�4Ӟz.�$�}*�0R#`	�� �X�bRR���J�+����q�P���c� ��-L$X$#Q c A�ĂD�b(��0>M�!\%Y��^��{���! �0`�q��H�Q!B��D`j: 415xF�)��������⑤K�c�c�+���4%�
Ƙh�J��̦��@�[���ir^{�����0�rn2��'7��=SB�qH��)_�JF�m��<��M!	o�x{�c�3M9<��y��U����=�i��W�n��/-��t�/L#�hE��h�n�����3�i�i�}�=%���Fʰna�����5�F�H�%
D�E�=l���y���#10��e�@�%p �XW���h@�*F�=�����^�_#I7ФqaV]氦I�����o�.o��!-����ϩ�H�"D�xh�&��0�G�e�b,b�21�+Ba���}����w�i�B0!�
�)��,��fsc�Ӈ�!�Y�2�C, ŁHЍH�H��Č��wR�g��_�܅�5!q�\I�CsHsxÚ�%p�RO3Ͼ���c��L~���"@`��tjKW*����Br�s�Y�A��],��{�	&�x�b����K=�1�N�NO-�O=�3|\���4��s�c3���!��u��HQ�BD�˖f������dr�/}��'̓�C�}�J0<p�=�䦑��}���5�B��.2�)�A��,�@l$Hː�L������7��<��哜�'�)�$L��M��ݷ��F���D`)��L����OY@�F4���9�F��&�<��Y������D0# �0��%*X�b�GNE��FZ�#�  �0JO�R���D�I#�%bB,dY�$ D! �F,D�E�V,h|F�@�D �X�DE ��HMa�	~�𙛙�� ?�Bʨ�uN*^X,w0$�`�0�!��0H11(gIxN���!i�� �b�%H$B%.s�s�3�# z�u!���4������$�,))
��bF@.1#,�$i
B�"��D�B��\�&��{�=�zcșJY�H��H�Ƅ��HԀT��D�,d���
�0�F-?kCaP$X�։�D̯��hK�]�e���<WjS^�l�*�,�o�_]{��_́E$..��,����.�0��g��<�9��9BR\Ќ���L��B��  V�˫P2�!�We�[<���f�3R�$��1�|�����|,+}��V��^��e���z�+B�ۮ� m�Y��y�������a^7�z�s+�0un��n��v���y!4��C')�3�|wt8t���Ͻ�对7نO<HS�Iwi���!��!�,�'\�N�!e}���g�9������}#�������7N�u���{❺���t���G�%Xf~-_�a^^��ɩ�&����f��g�փ���__:�ֽ��w�_K|�y�<�39N��>}����_R�3��$!�_<8�0hJK�p%3aYR%3|��"Ny2��)��\�͔��$a3fn��D�D�̼��#��L��c�ɐ6�@���SR���1�&aM���uA�B8԰k�}�)���`e��ܮ����$s��e��[��_Yr�RYXKn$�f��ý8����x}�OR�$"če�/���<�BN�P�ёX\��Ǐ��������,3xN:���fp������i�4N.j�^��/�*�MNg�y��|�,)<�<!k)I$$a �)�!
a��IZ����k/�y�xy�d!�,�#+s��Y ��� G�\vf�_<�a�/��+F�XF��E�]�Lݞ��eo��7�>����<�)�9�{��o��                       �                                                    �e�                  �|              6�                                        ���                         �   [@               ��                   6�                              	�                        ��      ��                                                                             |                                    :�ft�N99#k9����s�U%Ӵ�c����l*��U*�Q���s��\�l�u�x1�Z�{X����u��̵m��!p�Ӥ[��%2R�A�D�%	���
v��'��ﾏ����m�jUe��η��lD�x8)�X6ѫ�WX�V���yP%u<nĄ���b"gX�
��n1� �����S`+>��^�N-N�1Ӝ-uuk�G�l!r�3��s���[�+sq�I�p�b�k=9��;�KZ�dz�p�Uk � ]<�N�
� ��뤋-�[%�  @�sk�m�V��eU��[�����6�;�� �6�kn�� l ��7m�Z Ik�t[h��bAtؐ m�  �+Z��m� �yj�r������mp     ��  k6A�m�';m�m p2 'iĩ�5����J�\�!�ix��%Z��3��ej�Bk�nu�n�Xv��5���c�B��6�UV�X�6�S�Y��m��+K$6�@�m��a:$   	t���� -���K!��ڐ��5����2�U�U٪��m ۶ j[cl���  ۤ�t�\UT�*5UJ�!¡�a��%�[p����������q:�UV���n<f��n�����^�l[(��e�B�Jp\a�����j�3��YL�t�=�����  �.��ݹ��RF*V�l��Z�.�  >_�� ����E� �%pm��͒-ΒI�l@��I�n�����X�hpyĞ�:�mp��� ����   H ��ū��_�~t�d����u���۴�(j��-�l�IZ��Z ���e�����ѩZ���8`����md��Z̫�u�]���^Xx+�e۰� A���$�ՠ�n��U\�:�ĩ���1�i��gÞg�ݨ
�G��U�i+�U��C�;�7*������*�]l���m��]�崻��ŖM���s���+�ZUP R�������K�` �K"�k'P�zd0M+	��$X[t�l%� [[l 8�a����  �ݮm���f��[\� 8m�` yËl�mr����[�$����Uf<�"j�U   ��B��` �b�v6ڻn 5V��j���a��'�69:�m�$�E:��Bm��!+�V�uU��F��&B�`��mm�$�e7kn�V�A�b�l����}erU!J�6ܚV�UQ�gcq�sMe��[6��o�lN��6lNn�a]&�]�eeK-HM]Z�n�؝Q�U�ei�wM&���Ŭ5�I,��OM��i�Ŵ�J��PPJPur�no;$�8Ͳ(���6H��l��h<��@I�m�nٶ� YD� �  >�N�}�� �m���R�WK�N��lsd��IL鳝6�i0 ��`6�m�f��\� ��`��V����j�p  �` n^�vݶ�d�l�:ې��m�   h��t�`��$  H��6Ӭ́mK�i�@���m�XA�#̫�
�UR� ��m�m,��kR ���lN��mҶ6���@-�J6Z      [@7p [}%� p m� e��� �� m�    H  p�� �`    	l�`-�-���ۀ��  ��l 	     l    	��`�s  [[ֵ�lݺŒM�m���  ZM�c���m���Ym�O���l h���kq��� �M)k8�F�6֬�$%q39�Z����mT���W-.��8���n�   �` @ml�tU���[W$$�&�L���gI-�h  ��9!��$6ZH�	�,�Xm�e���@$m�  &�&ٷ    �  ��  -��:md��oͶ��� '@�    ����    @  �`�`   8 l   �� �  p 	�  m�      ����   ���6ٶ�kn p^��R�,����];9�[y�[A $�V]�i8 m�[-��M��� ڶI,�e��m���m	-�Z�6vy�e�e����C�r�U�  ����hN�I�pll ��G����̍d�-͝�D� �  a1�m%l[du�kk�-�[@   ��(��  [d  �� [@�  6ݤN� �  a�    �~�>�� ��� �ڀ�yB�����
���~�e��b����6 keYm 
^�a��`�c#P*�j�ҭ�t��E4��.�d� -�p�  J�@ �m6ۀm&m�p^��� -��m%�af`	�	�9�A8 �k�VIm�(�������;&�t�K*�А�Hm&�[R�m]UT��Y�m���[�*�U[[J�� T�1���R���mJ���TQ�A��*��l vۧLm�kѣ��M�Q�RNK5���G#�����;A\9q�[�7�n%L�S�s�M+�c�@]�\�����U�&�j��j��(�6[`A��a� l��i�`*ꭠ�Tݥ%�yn�am����͵�/6�^����3e��`�Ŵ㞓E��^� ����m������޲� 	 �:ۄ� Hky�  �ְ9!m  ������۵l$ru�� m 2-�@OA ��6�Ĝ-���mKz�[8�r�M��m`�5�8ݬ�ֲM6�l��:,�Nu�#�hwg]���  [N�M,֝��� P}���@�6&�+��  �o�m��H�-6�l�NI�� IͶ�n#Zan��;@��U�mA����ڶ�-*�Zm,�%	�e�I)��u��|5��kz�&��.���R�V��m���;:�j�As<J�S��sô�ݍ���U�����xN�x�	���m�۳����� #�6��d��4�1)*�[�v�ҭ���-sbͽX���:Ѷ���':�[m�M�S��m�� h  ��h��2�ʶÖ^Z��FVm����mH@8�ܲ�B��RK��i�V�j�sS�2�]M��Z��q$���ʫh
ڪ�L(n�M���a\�\�Zl˲�[v{�w�[����j��ݐB��մ���$8=m۬�!)���jČ�2ql�ƋВFh�l�L�[@ ����1E������' ;��nmnU�-0� �:M�h   8m�F��0-� ol�gk�l'F�  -�-�ŕ��@   i'g-Ųe�p���=�D1�,lu�k��X�3` �+qwK:��5׵�[4̀H%�R886=6����X��Y�Z�s#�:�9W��w�C�|�V�هa٬������Y�viσv�p�������/hKEq���-�����JՌ`��7;kQm��p�iKsff��\͹$���DDES��G� p���� VŊ@"Q�5�
����G��w�N�� :�`����p�C��H�� _@T��	��Ղ'��N!�<q�)8�h tU:x!<|F!�x��) _EwB�j�s� �TC���8��<b�#T�<�W_|��
�S�*��P�)P9D�CQ�Q�=5D�C���A�P�"d �G�@�C���+h��4Ԃz��_N
zO�� = �P/� ���A�?!�;p�O�CP�DA��z�C�4
���Q���x�)
V��T���0$HT,��T�ԉ��z� ���≀�Fb��� | �T2�`!�x�!�����/��P^��"���Z���H��D�� ��`Ab�U~Ab(,�z{���{׽���` � l          �   m� �  � 8  ��   ��8 m�         ]6    ���              l      B��&Hn��I'k��8��.����0[ғ�_3Odd��*��{$�5wE���k�A� ƒG��kkiV��	ڮ�[A��Z��iۛЏn0���^\�e��e1�l8*]l��h�u�̍Yxt��\���3퇧ˏ-<����9�8�4��:�7M"���l�n.
E"ݚ4�#A�M��I�[�l2ֽ�m�����;�|��e�ųǶ���qՍvg�3���S���\iې�s3��v!��k n��g��F��4k�װ]�{(b��/��GOomR5�˧��!d��md9��Oom�g�a�ɭ����*�v�r�%J�6�bUj�)y�ۢ�����n�go]��m�
!�%�l�<HT���#���"Y��DURa�r69�,��L��UU���e^����i�ThYH.V��$.�k5�ծǉ  ��m�ˌm*�VvͶ ��)vA�Y��ɨ1k��g�x����jdi�X��d��l]���@��J��Tki��UT��lt���k	��'�Zb��g[A�C�KnP�i1<1<���$)�9���ҹݠ�ɱ�@��h�������$�w<����5�e
�ΰ�p��Í�e2Q2�ڛh���#�	L&t�g\��tV,l�e�7�kr9�kX�M���g�	��5ǧ�;s&8�W�sb��b8b��E�)]Se�����t�yc#�̈́�hp0ʫۮn& �5���.�)'���mX��4�-ښ�ۨg�R�����D�\�yҒ����[��m˙��p�wl�����bE*�g���5�W����銝N�����᧊�� <������$$ J6�m��Ն.���  I�� ��#�tۭ��շa�-t&�U�g��mr�J�Q��19}�az#u����q��n�g�ɤlvS�j��33��8_2P�-��4v4�d��RvK�V��XՎc-����kn�<�Љ���.mf$h�a�������k���5�8+[�v[���L���"��Y9��m�W��W	�{�9ݓl`Exܢ���pv9�p���ST��P��C��ŀf�_ٷVs�V.Grd��tۅ8&�`�1�����r&���]>XXJp��ے��7���ܬ��U~K7�� �w����c9�D��U��r&�����0=�0=���ʉy��ĳ/��� ��ލX��vD(ջsΩҐm�UUKuf�L=�E�]���z��̡n&���Uێ�iS7B� ��ʂi9�7��`}��V��Vٳ���IQ�B�R�fc�#���}R���Va%�&����,F����b�rU��r&�dΘ���t��6B�T�T8ґXf�,;zXf�Ձ����ˑܙ$�Tc�8'%XΘ���t���������~��5��5BNv�r�LH�'/���ri�]e��օ��3m�h���O/"��x�����LoGLgL`ym6��7
���`n>�`}��V�s]��ٶ��(I6{`�M�UT��L��v�zՁ��g���	@�@�	!B<�J��6Ձ�9�����$�E���X�yXf�Ձ�����o]X���J�JT�!x0=�0;nD���t���M���-�1���\9��hW��ҽ�{6湲�lAŴ�&{�3�N�=���A��\b32��"`{z:`l�����gqNH��T8ґXf�����~H�t�`f����ܬ\���%
�˦��5J���i`~�m�:!(or{���޺�5oTi*�$�餓����I>�;��'�����T�=U<S���,A�M��m�D��%%X��`n�t�������2��YW�R�v������������/�q���ܔd��3�ν����Q┘�m�������07z:�y���0:�s�@�H���mG�������u`n>�`}��X���J�9N���"�3z:`v܉��e�L#C�R�ө�&GL��a�
�w;�=���{���޺�>Fw�H��%C�)�r&���:`v܉��U�����I  m� i�a�I����H    ��ip�&�����e�Yݹ�L\�kp���պم�獙2f܎1�qD��n�\izG����ɃD��5��ֻg8ݬ��8b 6]*�h�xր��TR==O�-� Vx��Dю.���ͱ�p�sp�L���[s�7�-7��rɭ�+.,q32�-���GVx5�b)ߝ��;Ͻ=��_�Ѷ��Hq%(�t�ӭ�r6�)V<��[5�V��s�q=�ê��dT���@���VguՁ��������i�z5NAJN�I����mȘ� ���>H�r�iS��03BK2��"`n�遳������P� ���F�qX�06vA��#�mȘ�/�@�I8�m7*���Ł�w]X��X�m��D.���SU)�uUT�2�=��U�eh����R�5j�4ӽ����=*�fܒ�NS���p��z���}����mtD(��;k�����M:��B�������y���Tʄ�	)/$�Rb����֬ݵŁ�۶��D6y��朦��Ɣ����]X�8�=�:`v܉�GEffR���5JÔ$�v���Ձ���`{ٷV���:�FJ��4�p�>��q�+ջ�}_�����׽�J`UX'���ܝ���k��9�Gj��R�I�6:�L�!���� ��m��.D�ݑ�gd�:`{��*@)ff]��Lގ�; ���選����h��%B�*��nU������۶�I(��JҊ�ɽvfuՁ�Mo��Ӕ�I��G�7�&&�GL��`j4:�,T�7!��ݝ���u`gl���;���T裍2R �H��!%�܉��j��-<�J��CsrWt�;F�1���+�*�E⻼����遳�l��ݝ�ˑ��$��H'%X; ���遽�107z:`r�'Q�NT�餓����u`f���06vA��j괪R�XX�	fS{�b`n�遳��꯯W���"Q/��NI>�ۤ��fwc���j�����B��?��j��l�A��( �IL���Fu�ﮏ�8Z,��/fܝ�n{YK�'�Lg��L$q6�nW�o�x�3;��ݝ���u`b�[�*5H����VgGL�ɉ���e�LEo\���RnA���VnΊ��;��缬���gqN~I�b��ۑX�06_D�ݑ�{�b`r��$���N	�Vv�,��7gE`fw]Xm~��w@�$�I$� m5�.�v�8 �    5��[_�h����sN�^k� ���$u��Ѯ�qT��C<cnE��ܞ�St;�m�-"u;�f�p�m���쮌J�&R��٥,8U;S��أ���	5j�d-���
�2)�,�FG�I��j��ݱ�v����qܾ�9�����&9n��P����t ڮ��\۹�3v|�� x ���ۻt�ej�ͷ�^�s��-�@7g1�z|խ�dv��*��'#�R�'dq�T��p�>��Ձ��107dt�������JWk+!,�`ovLL�06vA���u`}��J �~r4ܑX� ���쎘ݓ�� �@�D�m�X�8�37��ݝ�}���Ŧ��Ti(�pi�R+{���d��=�ce�Lik�-6y���##nygq�/=���v���;gMx�<3��2[��d�Z��%���옘�L`l�����U�'�L3;�5��Nfj��(o��W�Y� �8"A�����~��{�������X�ɒ9�ӧIBrX/�`ott��옘�L`E"W�uc�)��Vn�Ձ������X�yX#�Ԥ�������d���[�1���&�6���'Z�!�UZ�CB�z�SI�V;:��dw[�ڱՄ�6���{m���U�f&�&06_D��#��d����� I#��I$�3��3;��ݝ�fwK�RF�9�IQ�FS.SuN���`{2����]��Rhf���B&���5����p���|n(�� }��0`��>8:�c8@nt�5�G� >��#�<<6�K1m)��)���$
�ڡ�!(0
n�"A�}��0G��!e,��7�ў����<R��b��	
/.��ЀY�ǌ�1��="B�r�m�`)HE�(Y��d#"��x�'=�HcIYR������OS}("@F��p�C�$ �A$!��z X~T=OA �` �����y$���m������t�I�2R�U�����{v�?f͇BJ?����V���SQ-�1P�mȬ3�X����y��u`nl��7�R)��OҜ�#�F�I�4��ݳ�8A���tn�v�uS~��_"�2G?:t�(NO�ս�`fw]X쭧�|��߾�������:��)T�n�l{v��Pٹ���3��,�w��_��QS��$�(�qʰ76���~��Y�"Ǜ�`foZ�=��Hi���"����S��
o��V_��9$�߻Òp�$�dHq0]	(�B�_(J"=������0uUJu5SUUU`}����^�DB������zE`f�R�؈ȝ0I9$�/Ccd紓� ���^;��&{u:[vsűp�w~�_���Q��I����?����Ձ������z�������Eo?Sq��I���L�+=���"guX�zl{6���I)�W}�MSsNQT�f��o�U���ٳ�7��j����\���R��T�	�aꥯ{����`g����&�;������5N ��R;3���������|��O|�V����^���J�I$�I$���m� ��p �   ��E��;u�I�p�����,��7^�<�uH�0�:�v��	�=��	�	f�[ctH�+ƫs���:����]m�V�Q���XwjF�J����0{v�d�G��IN-b��0X�׳izb��#��Jņ�8Y�����V1�v��N���+�=j�F�ö��7TʣTM�w�w&�6�6�U͂
��h.A���c\��P�]�.��	��YjS�ӒR�P5%h�����7d������OΘ�E�*@��?GnH�ΜX�y���V�Ί�I^y �F�G#m�X�~�Ύ����d��R�iH��I���ug��oy�X��,Y��Ef���m6�c%I%0;{&&�w����~�쎘�������PvYV	c��u�s�u��N���B3P�ƶu�p=v���8]�ᠡ�1]�b`ñV���GL�����ܙ#��t��,Y���A��=�Az��%���'�wv���6��P�I���ܵL�i��-��~t��옘�`jޖ�����uE%9ERU���p�3fA��z[gGL߹e
�]��X����ِ`jޖ�������������߽����(�����&i��놹&�\۩^��G�ͪ��v;p5+��1�"DI#m�|��;;z���޸X�8�1s|JM�#O�$vΎ��ِ`jޖ��V��n66ӌd�$�sz�`ft��uG�v�TE�$ck��,P
�`�x��~��2�����R'D��"�=�,������,�VӰ5��ɒH:8��7o;��Ł����7vq`{�/��FD�HʍHm�眚\�;��ri����V	筥��3m�#�Cc*J[��
��7{���p� � ������Ȁؠ� � �����>A�����?N>A���������A�A�A�A�'צK%�m�3HCwvpA�666=������A�A�A�A�������lll~ϻ�8 ��~���� � � � ����Rɗ3�n�\�ݼ|�������� �`�`�`��}���� � � � ���?N>A����w���A�666?M��$�m��n��fn�>A���������A�A�A�A���~�|����~�?m���ll>h�QH!"|n`t=Px�>A|�?N>A����v���!�K�n�\&�� �`�`�`�����8 ���~��� � � � ������ � � � ��w�pA�666?�~�����r�1����f�=�9z7J�c�lv1u� �^N۷��M]�r�&y�骞>�����s�o �`�`�`����� �`�`�`��}���� � � � ���?N>A���㿿C<6fi��	�s3v�A�666=�y�pA�666?g���|������s����lll{����>A����}g\��]��f˙���A�A�A�A�>��8 �~���� ؃� ��A���?��A�666?�~�����lll{��럩s-���4������lll}���� �`�`�`������A�666=�y�pA�66
� �����pA�666?d��d����!2n����lll{����>A����*������� � � � �;���|������s����lll~��	����  m�m6��ְ�� m�H    	�����J����)[��q�}Ab{=�����w݇R�Sja�[fqn��9��9,�I�bY�I쌎�n[e�������v�ѪV��.5F&�����Pk��R*]u�����2�i(eqd���/Lp�ݥ�n�r�ޓv������`�fz�Ľh��3e�i����&M�\��)���\�T��ڣ��o���ca�ц�6���v%κ��';=E:����8�+w4����� � � � ���?��� � � � ��~��|�����s��#�lll{����>A������d�M��7ss37g �`�`�`��}��pA�
666?���ӂ�A�A�A�A�{��x ���?N>E�����_ٟ�2�s%ݷ	���� � � � ���?N>A�����?m���lllw��8 ���߳��A�A�A�5���M�N�7!	$��?����/{�G`}�_��fá(��:��1op�����(�nf���ZX�������`n��Ӕ�#l���$���i7W��@���!u�8�j�
X6�v.'���w��ʚ�u\hzN�M��o��`o���32��D%��n��9�5.]L�14������\b��^P��A�H" E,B�4�$"TR� 8~E=�{������������(M�f=R0�ԈR��wOE`v���RZ��v��V���&�N��S���v��1�t��v�9=ݾ�`b�w�%DB�R�&�,Y��/o�>����;vq`nNQ�I$�E����uKv�F2�&�֯#���i�ݷ�q��V����f�K�jUL�EUO���>�����,Y��Ef�����
(���36辅L�wWŁ�~�l��_�$mw�S��28��D���=ݿ�$��{���?�@Ҁ��
��	(�������`w��E����rUUAөH(�a�}�`�zX�:;I���`k��r��B�@�԰	�c�W�$�x�gၫd�����
.v�����nN�t�c5�k8��O4Gh��un͜0c��o���ӵs���(�P�$����Ł�;��TB�ÞwM��ݤ4�Z��EK�5T�̭/�BPُ;��;;�����w��f,'y�hT�)9�s5E��;��7۵g�(_(���������u|X�{3���l�U.QUSaС%�wU�����̭,�'�".��RӈKTB�_(�^�w���.�yLԩ���(����̭�`|�B_DB_w~���������S��6� 	$����1�ny���A�45ַ��$k�����pݟ�w���e\*FGtH�r/��t�`b��`k���J��]N�׌�rT�D�UMU���۳~�
S'=��`n�u;s+K�ID6k��tRe54�sN���`fem;9(�M��q`fOs�?0�)$��UR�U5Sa�_$�%=���v���`{Ӻ�>��СDL��}VGu!���T�K�3TX�ZX(P���o>߾�36�%s}
��Cp�F`Ed��c�F{�i7�R�J^�Cꄐ�KO��f�30Z��>�6>��p���BR�k˻�~����  ���          $      �� $ �      6݅�            	��    �                       ՜��ٚ���'��u���c��(��p����{HcD��v]�c���{=�ug�nn���C�� ��k��+u�*�^
8؞3gcd��.�b0j㌹�6V�g+�'W�]Q�R�����rk����z۬n3պ71���:���&�oe@u:ۍL�OOW	f\�Z�;�ł᪤��8���z�\��m�2���!�7T��3�uŜ�݃r���M�\\�p�:�(}}�}���۫��¬��ī�i��"�K�\�gn=��O5ra�*g�{k�n�������&y�`X6�5�m��	yTݕe�4(<�@R���&~H�@��5;p	�15Pc�Sb����rn@A�y庪��� .Ӗ��SʫU��m�@���Um<���U���2��6�c;3�ej}`�iXr���@�GJQ���2�T9u��«�wϾ�[']��p���
��*�Ulce.Y�u]����:�	��r����)Vz{E����	 �!�����ڶ��� �6��uM�ɞ�Ulͤ�=�����G�X�D�V�Ҽn���Y%�e��j�rk^l�vڕ�"�7��n�gʹk��B�v���#L7
��Wg;���bF[�C865��u��R�;p��������H�"�s��Og�ob��͎���Jz�Ƃt�Cm�|p��ƥ��nY�g2���6Y���ZȐ	Q�E��;��
�e3����v5�1�kz呣;�Z�[�^`*XT���	UU�-�=��@B�(t����J�n�ڢn�N���qcd�.���ڌP��� :Ap<8 TC�� �~@O�H����l�������` �Z�v�`  �    	���������&Km��˰\etz��t��;�]�g�:)��2V�t��n7\Fy�n�p�s�X�
��\�ۦ�� �(�H��(�[m�v���G��+��+vy�(��\i^�n�Cn�m��7&�r��`u�y�Rk���ؒ�mS;v��Җә��,�,3���!����<���3qRI$�Ӗr�����G�u�9�9];�#rA�����y�fN9ژ������O��ب�Xf��3���`�ڰ32��$��÷k� ���)�I�i�R+ ���I&�ݮ�`v�q`y�vo�"f1f�Sq���c!$�����ݜY�&��t�guXY�YNQSN[�U73T�9%	���`c����XtUU.�E`r�{ɑ����T����f��$�;���]N������ߏ��
.q���o{u��8����:��[�C��
�,S~�w{6���VƙSH�����`fem;s+O�%脣������I>N@�)��w�O��{���\��E�P���h�� AC�+r~���9!��`�ھ��Cg�v�c	rDT���vn���fΈ�P���Vd�'`f,*u�hs534�j�P�C̮�`s��=��N��DB���|Xƿ�~.�d��r��;_�f�脣3o��n��;��i/�)��)���5Mؙ��rc���v��D8�V0�Ɇt׎2j1v%?{��۾��eL�kZI&���X�8�3r�UU|��������Y��6�ȋ�g�ICfd�; ���Ͷ_(����&F�*@d$p�7_����Yǁ P��{�|��O{��9$��K��4�$�3d�79'�������������s+K.ID$�L���a�����*���*��̦P�([�z~�w��o�j����J+l��U͂T�S���O
�mv������;�b�p�f�ͳ���ǜ�Rɔ�m��-U7�ݮ,l� �n�B�J��\��	Cgr����Q33Nf��3�y��B����76��s+K�IW�Ư7থ*nH�8�`�zX�n�Q	&�v��3���<��S52J��N�UUa�%�BJ{{���wWӒO{��rO��S�!J�L:�%
����ޫ��r��"j��H�&f��72��>Q�Q�w� }�}V��J�+��H�1	�'�"D�&N3�ςi\�#ͻn{FC��tm���M��ݬ��tnB�������;;������$�0��������)M�SA.h���_B��ͮn�������i}
<�5I#] ��B$���76��s+K:o;k� ���{)0��i���UM�rP�v��3����t��R���Vuq�$	����nQ`{r��9'��_�����̭,��߫��������` �m� ��l��    .��+�QMû2�NyB�5udҍZ���{0�t�;�I�r�H��4J̯^���ٹ�O�gm��vl��WmUJ�������iVR[��V��n��rk1J�7�#��=���\�i��a�n��Ͱ\����ټm��.Y'�� [�Wg-Ic�1�vu�;����{�߽�|��i��T����4���f�) ��K[TrާKc�Mv���/�r\9RD��;sg%`v�����Ł�����lt۔��I����`N�T�l�K�H���32�ܦԢA��=�<X�����yo��ޞJ��v��܄""�GI�����zl�V�aГ������9�4&ꐦT�9��^�́�J!�G���}/�}�WŁ��ٰ1���h�:�&d��I��-G��5h�1�Ӯ�IK��%��ms�����������ծ�j���].�����������������҅H
^�2�Dr5`wl��
!(]	(��_oM�Ϸ�����w��""ɼ����`�U-�D�Q`o��;^�͜�D7�����,O=��R�9��ʗT�>��������M�����w+KBQ�%/�y���~��%Q9J)Q9�����;�q`g=�`r��`�*B�JpĥDo��y�v�Fw&v���#:ɹ��m=�k������9��VO���������ٰ5�l�_�n�t��ĕ3QUCj��u4X{�7�Cg<�wk���Z_(�ٯ�s�hM�!L��s56<�3+e�h�!b�$A��)���NI=�oM���x�c�9T�'USa�!$�v�]�۵Ł繳a�%	��t���I��$��j���Ł*�{�K+���s��32�]��{ju�:S�Qqzz��=�7\5��p�	l�g
���U۱�Mg������.�͖��o��l���6fV��	B�÷k� �W��SJSc��C����߫�~�H���vn��������P��5�y�Sj�NR�E$v���Ձ۳�=
7������`b�j��IsIˤUf��rP����`c��5�vl
��IGD(�����foT�D�I�ŉe���:[-��ݒ�wd,��.�Q�"R rH��A���2��^�x���P�q�����A��D��w���~!88����������X�Zt%���v��T��%9���UM���r_(�I��k�:w�������"� .d���%,��fe�Kf�l����`{g5��$���`n�\�b¶�C�KsC��áBP�}�v������l�;vq`b���6��r; ����~���|π������ٰ)$����Ve�U  
P��[MkN�      $�����m*GH�&����mwAԝ6'I�h'C��x�����/���Ѻe���o0�]�$�����v��y��#��c����g	Hm2���0�^��j�Hq6w��Ů��<���6�x��-��V,d�.�--��ۦ�Yp6Ij��{��j��x�*��i��iGN�6��{v}
A�N�<;{q��������������X���Z����72��<�6yD$�0;;�����Y#�MJ$q��g���!�oM�vwU����X��$��PM!QT:�,=͛ �ͫ:(ow|��{��W�6@n"��7�BJ�ޫwyڰ7r���(QD%;_w�`c5�))�DЄ�l��j��;v��>ޛ_�f��(�_�ϟҋ��j���)��N�|vh8Iu�s5v��Q�Vye����_#������ʪ���u|X{�6�n��!G���n��'�BT���r.�|�@à#"�SZB�5Q� ��P?��f��g$�l��6�V�С��L�H�L��e�&�ly�6d����%�IL��_?+Y����ڔ��I���fl̭,l��I>��VN�eT˙�S�R*jf�������:���<��v��n��9N�26�He���8�t�,�m�%
�����V�
X6�v.�g����]��t���֮������ޛ_�f�̜ٞI(�÷k�_rOђ�j~r��v.�v��n�������ٿ��(��oI"�&�����M��=�́�����0��$��t����`�}�$�Z��"�`� ����b� A�1"��#�"�zL�=x�����F*TU�+`A#�c�z�.��H|�j�!!|QQ�e%� ��|A<��R$�Kh[C�a �������00��;�w�{���>8�����({�}�"��z'}ؐ�.�
��'�� ���t=:
x	���/����q�!Ǌ���Q"��qbB���.�&����?G���[��&�5U3a�>�,}�6��V��n�ͭ'D��)Q�MA9o;߫����ϼ݁ݳ�p:r��t�s��rr�j�2��L�&��E�X�{X�7v7g��?��d�~�Ģ��f������O�7gzf��͵В��!���v"����Q�6�F�$���{��tt��:[ ��?�RD������K�S�R*jf��޵`y�l���ݽVs�7`b;xd��1�*
IV;o� �ޫ2sfl%B���$U�A(D���w��}{�O�H4���88X����]Ӽ��{��Vv�,��Jw�R)LBr5�ru7=��2�sP���<.�u���r	��7?�F1�l�9�B�RG�{�������nV����`z3i0��x*I��l	�06vA�M��y��RGuq=��G5ܫ;k�_�f΄�ݝ��zՀi���1Jm�#N�p����y�ϼ݁۽u`b��`b+5�6��7 �G$�7^�v�����W���;���?����_�~�  �` �Z�{l 6�$    m��I/,1�ap�5���Oe��#u��͞����vԝ��]��a뷈mc���sM��/��K�O[����n8�N#��#��l[aʶַX:p�,#Q�U�JOE�nA�����i���+��n��t(6���㎮.������Llũt�.N�:){Q՞8j$J���ww������Kn�
�Nn�F�.�����N��N���W9��z�Y3��:���au5�(�G�3���.�]���zX�y���%7?7(�H)%X�yߒl;���ݝ�w6մ�.S&��ߥE%	�H	��/w�������7ݽj����`~a�E�*�������y��z����������`g��I<�u#������V�_���;ϼ�׼݁�0�q� Pi�9\Ӊ��>��v.�t��Y��`ܓ�=`����9ژ˹�
g�an�m��������v�sf~I~a��j�8��<.��.��77o$�����O`��]��BSe���ݽj�����<��m!dc$���{����V}������V�w����z�"jF�JR������DOo~Tv��ɠ؈Ovo7`j=�)���EBAI*��}�������{����V�Y^�蔅�0��q\��-�L�d�5�ۛ�H�ۣ[S�.�ctDU���a��+e���uO�}�����Nĺ���B��3'���y��S�O�AȬ׼݁��ۑ0$������L��	~��ɪ���k�ޝ�c��Q��*������~�vmi:$%I4�SPW�07nD�$���i�'GL�\��Ƥ#��Vݽ,͑&�07nD����b2�I]SpL�G��F�ړ���c<W�IP�3���+�ٍ��ڤD�D1�I,͜��'GLۑ0�1���ґ��-,K2�RY�0:tt�ݹ ���9+��%7?7(�H)%X�8�?�{�>w���7�����r��nF�@#��woK3g%`wo]Xg����Ł��2��Ԏ�(C�X��&�07fA�I��)"u��5W=u��X7/g��6�n�\S���6�f���<،6xL�Z`I��gd�3���W�I3��5i]M*�s4�nV��BI��ޫwk������DBl;��br�"�'QH��ޖn�j��޺�3r�1���_�(�1ɘ��얘::`n܉��J~����'y2�9��擤:�vnm��%�]����X̭�`~K���K�z����N��~��  � m5�.�I�  p    ��ɱ���XݴVcv�Z�O8�:M�D�b�'b�v܋Ag���8uq��5�m�:���;���6�F^���)���	�uԁԥ��S`�L[(< ,�f��;T.���/!n������u�t��6�"�pՓcrh�[������c�+y.�^$���}]��5Y��ߞ�w��]�Yp{e�e�gok&��Ob�8�힚�rm����M�+:張E�AI+@�����zX�9��z���|�G(�:��8��zXݒ�N���"`y��TE\��(��n�j��޺�3r��(M�oU��ͤ1�}$�Jrɚ�vN���"`:c������L�q=/��P���`f>�`������X��VR��ȝ0I9*B�]'@�u�jn%�e	ٺ�Ǣ8ps:[ ����DF�19M�R4�)�ooK3+e����"#���v1f�)��U-�%UUX̭�w�aE�D�m��{��;��������H���c��7T݁ݽj������P�;������Go�ܦ9EA�I*��Ͽ��ŀ}�}VfV˰�O�{�7���9Dp�Ԕ�4�`������X��Vv�,Z������I#L�Y7[X�����)��ӹ�5#�:;��M�։�FT�(����j��޺`l���t�}ݔ!S1f*�E�e�N��/�`:c��Z`gV���B�
r�]��{v��#�B�BrU]�W.��޵`�7���7)H7I���zX���N���K`j+z�+_],�Uf^f0;�%��05l��$�,�;�HB�I�@��%RP-s�H�wgk���CDOU=�k��27�N�������u��e��05N��$韾�	$�V��ᒛ��(�8)%X�y�nmX�[.�3sj�DCf�󞩪jHGN�; �w����������7ϼ���X�~�F��Ia�{�}.�;�����k�Ģ��b=Uv�zX��P��$N�Cr5`����o�y|�w������>���Qs�Qqzz��=�[����Ͳ�Cl�P�X�e.�:t�sad�ɋ%���җ����1���-0	:c �F��c����V��/��<ՀooU���ٿ�D$ٌY��e�S�F!�I,�j�7����;��ooK+�"FA���9���`b��`����ou��Q�ᒛ��(�9B�X������36rVI>���I<WxD�eVЅp��
�A������!��"H�	 	 		��I##1�@�B�a�4�"%
R`�
@W(4���Y�)�I)[7�	�B�e��IY
X�l#|�9�*��ﯯI���'���~�v�����  ���                -�  $ �  	    n�m�            	��    [@                       1<[�p��l�gix��u.��ۍ�.�u��l0l�)�`���s��3gj�K���A�YL��l`���.��	����W.�*�6��eٞ�f�0���r�7��v;x0���+G �e6�b��T
i��^^��������F�u�h�u�ǶL#�m���I�z���)L�R�X 
�we��Z��mel\�;	�n��e,�=�����;�5�\i�w��;R��:ۃi^b�����hr���q���;v���c�^h�ƽD��9^�s1���l\�[��ų<;����r�/(n`d��!^�* �u+%�)%ΉU���)Z��t�+�� �Nɹh�mi����*�[��n$kn��l� ��
��Z���@��Vqۊ�e��e�
�`+��qU.X5v�; ��1�Z,@F�N�(M����%A���v�j�t ��J�U[�.
j,v�C�/�S�2vI�[Hy-֓&0@2�
A�j���E*@&�S:�sp��Gh�<��qdu��M�{��S�e�<��ٍ��M����8�'��ݫY���ûk��P;D[F24݌��VF��t��i��[[%R�'�87H&�����ʇ�܋R�0/I����S=D{g����8n;t6��b����=nLM��Dq�-ӻ(	�ڪ�j���1�7�4��Ÿ��\5kn�x���n���'b�v�\孧^�.����e%!�*�Ss��o[��t��9|��]�"�[�(.r��.ûmr�e4�΂<Db��T�G�B	�:��"���Q=ׁ�@�]��d�wwwt  m�m��;` p    ��6�����"j��n���ڠ3�x��n�h�f�eĻ{j�cv8�����^l/v����wP�����h�i9k�8�+iL�%�eGv�BV�s�+��uٽ��=�P�$����՗v�%dK��1�0-b�/<p�׺��)�lu�I�����Un^��+9ie��{�`���k��j�qq��}���W=3�t�Fuv9��2�ɍv�N$NFJBp*:pq���,͜��f���B��wM��c�n��Q8�E�cw�$�$�[%�	:U�DD&�Fm&�9�*�UK�7`��05l��$��ȓz�ˉ�q���,Y���zX�9+ �ޟ|�G3��bq�S�n��;I$�t�y$�H��K�$��?g��Z�E �Ϳ�~O�T\u�7����ҦN��p��:ⓖg<oo	���ek��ܡ�#$�|�[�r�i$���������ꪪ����w��$�W9�D��%E)�+I$����]UU6�'ܝ��]���K^�t�$�3��F8�r�9B��y$�\��I%'L��K��]&�IwoO�I-���d�9QF��JD�%�}wrOg��]}��4�JN��$���]���������R
*RO�I-{9�i$�N��$���[I$�t�y$�ve�\�T��hgd�h�h��%rK�8͟)�R�	��\�_#�6nkI��v�m����ͷ�;�m���ͮ�����a��_� ��G�c���&f����I(Jf[{����m��>��y���H�s|Q	�(7JH���]:g��]}�	��_]���=��r+i$�����J!6F"
I>�$��\�I$�t���r+i$�N��$�W^JD���QJPV�IooO�I,O�[I$�t�y$��I%8��Yf]�q��W؎�c���[ �ìB� n��V���d5s�6t�77k7b���n�i$��3�I.���I):g��[ϓ�S�J6�@��I%ݽ>�$��I$���Imܗm$����"����4�MI>�$��\+I$����/W�޷�7i$�{�>�$���BAȎUR�d�:��BQ3��_�6�L�L�n��~��嶾ʪ5�L��B���Pa
�:���n��^[m���!��Q��|�X�sv�IooO�I-{
�I-����%�:r�F
A�:)"'Z6tZ�:��̂�\�u��������p��MZv4�ܒ��t�P� ������%�b�ZI%��>�%�{��I-eo?Sj4:rE)$��ױp�$���=��r+i$�N��$���H̰n2TR���[���K�N�I-����%�b�ZI,f��d��r����Ij���K�L��K��A4�K{z}�Io>N�FB(�7NN'i$�nm~��|�([[o�����ޯߛo�w�ﭶ�{ӻ���~??8� �`6�mm��a��  H    �9Ȏ.3(q���&ؠ̀J��en��:�(LcN�jkn���/N�qhݞ�ă.�� JkY��ղ;ve���c�ҭV����ls������P�N�R�D�e�v�u�'8jenP�n厺.�NK[; <�k��n��t���=�sgk�kۮWk%c2�l'�%8���һK.�V��{^M�1˃�:�Cr`7D����z{tS�+�Q��A5BjI��]�p�$����D�yS"fTȞ���8�D̩�3*g���O<��3*dO]���N�t�7,��/ș�2&eL��ݩ�2&eL��o{s��Lʙ2�}����ʙ2�D���e�y󻉱3*}���e��]�˹���S�*dLʙ���]�y2�D̩�w��<�G�Dȟ}����bX���ݣȖ%�b_��͹r[�fY����bX�ʞ�{��*dLʙ﷝������L��S;���<�D̩�/����'�3*dLN��������4�w��{��Q2'�o;/ș�2&eL�����ʙ2�D��{w��Lʙ2���w"y��w�Os����|}�k��j���Q�]����<���<mp���j!�lW`�K�n��n䙗tۦnl�O"fTș�=���S�*dLʙ����'�3*dLʞ��܉�2&eL�������&eL��S�>�̛�݆i2f�wmO<��3*dK���x�C���M��S����<�D̩�;���O"fTș�=���S�*~v��L�����seݒf�n��ۼO"fTș�>��܉�2&eL�����x�D̬D!�3*{�3���Tș�2%�{ۼO"fTș�=�/�2�&��2�ssr'�Tș���؝�|���y2�D̩�y��O<��3*dK���x�D̩�3*{�wr'�Tș�2'���['l��t�ffݗ��Lʙ2��s;jy�L��M�M�1ϳ��O"fTș�>��܉�2&eL�����x�D̩�3*wd����I$�Ӗr��g�Ͼ�]����Lq��lr�p��f4�z�˼H��wbF`�{�L��S"_���O"fTș�=߻��*dLʙ�����<��S"fT��gmO<��3*dKݝ��\�۷7r䛻w��Lʙ2���w"y�?�c�7jdN�����y2�D̩�y����ڛ2�D�o��x�D̩�3�����y�4�w��{��S�D��rv^'�3*dLʞ����2?*"� TdUY�j�=���.��.�<��S"fT����O<��{��;��{���Ƨe�t\����"fTș�=���S�*dLʙ����'�3*dLʞ��܉�2&eL�̻4w�
e˅�d�%IE54���.��2&eL�}���ș�2&eOw��D�ʙ2�D��rv^'�3*dLʞ����2&eL��w��Qs�5F�fn69۷=m2gdw'V��ey��d��N�$����Y)әkqm�w��Lʙ2����D�ʙ2�D��rv^'�3*dLʟ}���2&eL�}���ș�2&eOvK�L�L&�e&��ȞyS"\��>�y;/ș�2&eO��v��ʙ2�D��{w��Lʙ2����D�ʙ2�D������ᆋ��k{��ܧ���﹝�<�D̩�/����y2�D̩����<�D̩�>������Lʙ2�~yܲ�K.hK�ssmO<��3*dK���x�D̩�3*{���O<��3*dO��'e�y2�@��! $`H0�� �yʟs�����;ܧ����ߋ��#Q#�E��&eL��S��w"y�L��S!��{���ObfTș�;�g�S�*dLʙ����'�3*dLʞɷ�훛3��j��CD��L�B�����K�0Κ�nL�=�B�-�Y��IS�����2�D����x�D̩�3*}�3���Tș�2%�{ۼO"fTș�=��r'�Tș�2&|}��f�I��4ۦn/ș�2&eO��v��ʙ"X������Kı=��r'"X�%������%�bX����ɹ��搹�.m�Ȗ%�b{�����Kı=��r'"X�%������%�bX�}���,K��;��͹�n\�7�nm�yĳ�������,K����?N'�,K����؜�bX�O �v'�y���yı,V��H��B��)���9�d&Bd&'����'�,K����؜�bX�'��{x�D�,Kٝ���Kı=Q�H�*�� ���  m� i�a��   �  *���\d�d�;u�j<W������jݧv4�:ݫo0�!�b�]��5�!۵��������m���ql���c� # =��n��V�a  "^�.\�:y���k�TZn�&�[zB�vc�鹹'xz\��;[3��6�h�Y�u�:9��tXfԍ��e����3�{�04N���b��k��}YywV��r�4�\�'��m��[�M!�{ҍW)�������{��7�����Ȗ%�by�����Kı=���ND�,K�t����Kı;��l�Yt�K�swlND�,K�w��O"X�%�����r%�bX���ݼO"X�%���ݱ9ı,O:v�\�ݗ6e�7v�<�bX�'�;ۉȖ%�b{�v�<�bX�'�ov��Kı<�{���%�bX6��3.�0�ٛv��Ȝ��DȖ'�i�׉�Kı;��֧"X�%����'�,K��;�Ȝ�bX�%�����ܙsl�n�M���%�bX�}��S�,K����oȖ%�b{���ND�,K�w����K7�������.q���ש�F��r`��WM�p�Df��/8��\3�l�c�DW9���搹�.�Ȗ%�b{�����Kı=��r'"X�%������%�bX�}��S�,K��w���sL���v�����%�bX��{���Q�Є �g§D�%��4�Kı>�s��"X�%���oȖ%�b{��㶙�L�f�n]܉Ȗ%�by���yı,O���Ȗ%�b{�����%�bX��{��,K���zKd�˛��2[���yı,O���Ȗ%�b{�����%�bX��{��,K���>��yı,N����K�.�]˛�jr%�bX�{�v�<�bX��#����Ȗ%�b{���x�D�,K�;jr%�bX��N�w��7&�2`�f�N��{1���:���m<�lLc���qۓ4���ӵ×"��{�s�bX�'����ND�,K�t����Kı>�s���y"X�'�o^'�,K�����̴ۅܙ�m�܉Ȗ%�by�v�<�bX�'�ov��Kı<�~��yı,Os�܉Ȗ%�b_O{�,�ɗ6�6�Jf�'�,K����ڜ�bX�'��ݼO"X�g��a!�Ƅ��1�$�(-N2�3����!�d��&�L���(`eHfb c��P�̒�F�F��p1 �(�)��L�,�,H`�	�\�
�	�(�jr�H2ư�����X0�o ��E}Ʉ�妐^n�GT�u�OC������u}\@]�=E�Obӱ;���Ȝ�bX�'�i�oȖ%�bw's�&攛�B�̻��"X�%���oȖ%�b{���ND�,K�t����Kı>�s��"X�%���ݻ��neܻ��nm�yı,Os�܉Ȗ%�by�v�<�bX�'�nv��Kı_�Y��~!2!2K{��Jl��&��=�+@u�뜼n��[UӤ�<�9��oJtr4F�C�sL����w��oq�X�{�{x�D�,K߷;jr%�bX���v�<�bX�'���D�Kı<sޖ�'n\��fKsf�'�,K����ڜ��Q�DȖ'�o^'�,K��?~܉Ȗ%�by��vq<�bX�'~�N��s6�\��S�,K�������Kı=ϻ��,K������yı,O~��Ȗ%�b{����swM��nI����Kı=��r'"X�%��w���Kı>�s��"X�SȲ����lO�y���%�bX6��3-6�w2��ww"r%�bX�{�ݼO"X�%��۝�9ı,O=߻x�D�,K��w"r%�bX��������e��SX��"ny�9����3�[N<>nPMy�6�۲�㉸�쳮��ͼO"X�%��۝�9ı,O=߻x�D�,K��w"r%�bX�{�ݼO"X�%�ܝ�̛�Y74�n�wmND�,K�w��'�,K��;�Ȝ�bX�'���oȖ%�b}��mND���L�b~���w70�˹w6�����%�bX�gnD�Kı<�O�x�D�,K߷�br%�bX�{�v��bdK��!oK��ɛm&f��ND�,Kߴ����%�bX�����,K�������Kı=ϻ��,K���z[,���wr̖�x�D�,K߷�br%�bX�{�v�<�bX�'���D�Kı<�{�q<�bX�'A��P"`�(�5�u��7�od�  m�m��Z���� 8     �OI7�9w#l�GI����^z�|V��8����Tێ1��>�ڱM�8�i�#�ծ�ձgrNm��]��N�n�'H:@J�ؗ��X�̞5L�[�u[2��1;j��T
��;S��]�ף��9^.��j��.��`�(xY�s�mQ��˸�6�ixK].�?}���|o�]��ஷ��M��"�4��	��&ɡ��K��4�mh��#w.f�]˛�b{ı,O����<�bX�'���D�Kı<�{�p?*ؙı;���'"X�%��Oן���s3M�$����%�bX��{��,K����i��%�bX�}���,K�������Kİl=�:fZK�neٶ��D�Kı<�{�q<�bX�'�ov��KȤ2&D������%�bX�g�ۑ9�L�����8���*�&jJT�GT�'�,K��w�؜�bX�'��ݼO"X�%��w��9ı,O=߻N'�,K��N�fM�,ۚL�����,K�������Kİ����ȞD�,K߷���yı,O���
�L��L��Lw��Jl��&���\mQ�K��9}VCxP���k��sk�v�N�,�K^`�����{��7�s��D�Kı<�~��O"X�%���ݰ?"�șı=�{��<�b�	��D���5DҚm���I
�LK����vq<�ϊ�*P�vԋ#ec �>���!�9��wݱ9ı,O�߻x�D�,K�[L�d&Bd&B��M�6d��l��ͧȖ%�b{��lND�,K�w��'�,K����؜�bX�'��ݧȖ%�bw�	�#w.f����ݱ9ĳ��Ȟ����O"X�%��w�؜�bX�'��ݧȖ%�b{��lND�,Kώ�v%�˗4�rMݼO"X�%���ݱ9ı,O=���O"X�%���ݱ9ı,O}߻x�D�,K���m���1����cs��ćC�5�&��ț7/N������ J67r�b�Rдow�,K����i��%�bX�����,K�������Kı=�{�'"X�%�}=�t�w$�ܚmܗv�O"X�%���ݱ9ı,O}߻x�D�,K߷�br%�bX�{��8�D�,K�>�̛�Y�4�7e��'"X�%���oȖ%�b{��lND��W��i�6'�o|�Ȗ%�b{��lND�,K�߻v�f�]˦�mͼO"X�%���ݱ9ı,O=���O"X�%���ݱ9ı,O}߻x�D�,K܅�vXK�n�I���'"X�%���Ӊ�Kİ�����byı,O����O"X�%���ݱ9ı,M���H�0I9$d��) ������ѹ8\�L����WY��4ek��ci�H�e��Oؖ%�b}���'"X�%���oȖ%�b{��lND�,K�w�Ӊ�Kı;݄�I�su�s3wlND�,K�w��'�,K����؜�bX�'��ݧȖ%�b{��lND�,Kώ�v%�0����7v�<�bX�'�ov��Kı<�~�8�D�,K߷�br%�bX�{�v�<�bX����7w,�$ݙ�nn�Ȗ%�H'��ݧȖ%�b}��lND�,K�w��'�,K+��	E(��F��� h�`��`2
���PdK��dND�,K�{��f�%�ɦ]�si��%�bX�}��ND�,K�w��'�,K���ݱ9ı,O=߻N'�,K��G����}E��j��t�n��.��`V�[d�iRi]��N���`�6tޖ���yı,O~���O"X�%��w�br%�bX�{�v�'�2%�b}�s�9ı,N��۷s7$��]�n��yı,O{���,K����i��%�bX�}��ND�,K�w��'�"��"zΝ��3&Bf\�H'��{N	 �'����I�=�~��yı,O~��Ȗ%�bx�%,��37-�-��q<�bX�'�w9�,K�������Kı=�{�'"X�%���Ӊ�Kı;�{��]˛��nff��Kı=�~��yı,O~��Ȗ%�by����yı,O~�r��"X�''N��������r8 �m����b�� � @    *[/�մ�ټ�����W�L�49�\6Z�"r��]r���i��7spɹ^-�\��֦^�m�.s�{f�*�L�����a�%�fyݠ�*�h�,ݽX�VSmD�XU[8.��/9���ඎ�������v�\�9�xSZ��6����7']��[�8��}���LV4�%�褜^���!%��xhlkf���m���ɶ��70�'.N�Wc�7.ɻ���Kı;����,K����i��%�bX�����,K�������Kİl��黹d�&�ͻs7lND�,K�w��Ȗ%�b{��lND�,K�w��'�,K����؜�bX�%����ͺK��L���Ӊ�Kı=�{�'"X�%���oȖ%�b{�y�'"X�%���i��%�bX���vd��p�!��.m�Ȗ%��D��w��yı,O���"r%�bX�{�v�O"X�%���ݱ9ı,N�{۷d��&d���woȖ%�b{�y�'"X�%���i��%�bX�����,K�������Kı:}��
.q���bz[��.���ɸ��v�0+�N��\g�n�e��I��2Gj7dND�,K�w�Ӊ�Kı=�{�'"X�%���oȖ%�b{�y�'"X�%�����S�3s,�nfӉ�Kı=�{�'!��؛��w��'�,K����dND�,K�w��Ȗ%�bw��-��.n�.\�ݱ9ı,O}߻x�D�,K߻͑9ı,O=���O"X�%���ݱ9ı,O~;y�L�4��wm�7v�<�bX�'�w�"r%�bX�{��8�D�,K߷�br%�bX���v�<�bX����7w).I�3n����,K����i��%�bX�����,K�������Kı=�{�'"X�%��O~���0\lT�(s��	y�`P���5�ew�gg76�b5ٷSq��3�M�wi�{ı,N�m�Ȗ%�b{�����%�bX��{��y"X�B�WsW�	��	��M�$��SsD77-ͱ9ı,O}߻x�D�?(�S"}�m�Ȗ%�b{���N'�,K����؜�bX�'s��77m�n�5Ͷ��'�,K���ݱ9ı,O=���O"X��_�5" H)�������țy����Kı>�{��<�bX�'�	z^��K�.�n�m�Ȗ%����=���S��Kı;���'"X�%���oȖ%�b{��؜�bX�'�������wwL�nfӉ�Kı>�{�'"X�%���oȖ%�b{��؜�bX�'��ݧȖ%�g��I?+DI$���G%μ����f[y�3Fv�e�n.֎#��\�1�x�7�\�7v��Kı<�~��yı,O{���,K������yı,O���Ȗ%�by����d���˻nI����Kı=�y�'!�)k�2%������yı,N�m�Ȗ%�by�����'�ʙ�3��K�jUQ4��U+!2!8����N'�,K����؜�bX�'��{x�D�,K���"r%�bX����K6�.nM&nLͧȖ%�b}��lND�,K�w��O"X�%��{͑9ıq�A�*%~������yı,N��;2nm�ni��slND�,K�w��O"X�%��{͑9ı,O}߻N'�,K����؜�bX�%>���Gj�ͷj��s�&ѦM���mL�Hg\"�p)ӈ�����vY�m����ı,O{�l�Ȗ%�b{���q<�bX�'�ov��Kı<�{���%�bX��%�{KM.�I�wdND�,K�w�Ӊ�Kı>�{�'"X�%���s���Kı=�y�'"X�%������w2�n�m���yı,O���Ȗ%�by����yı,O{�l�Ȗ%�by���8�D�,K�w�m����e�swlND�,�	Ͼ�gȖ%�b{��dND�,KϾ�a��%�bX�}[L�d&Bd&B����D�5Tə*�����Kı=�y�'"X�%���s��yı,O���Ȗ%�by����yı,O|OO�
}�}�f)�i���	��<�|@�ϏT(�y��z`w��LD�W�,���.�ED���<i4B�D�J�����.R�>	�TfE�ـK
�h
W�<�qH�%R"A ƨu<�C�2����ψH���D��(A�D����hq|%Z)����  h [@               �  � 8   8   �l6�	            ��   m                        SG���S�0s���,���ρ���1����"u���;�������ܔ[p��kp�s�䴅mU@v]�7gSd�vQ��4+Ulֺu��7m��>������gp��Mɑ�`�	�8ݎ�e���v��{[=��,s1�g9�v�8�ٺ�
�P�;���Ű�%�e��⮊�\�݉8�/j�,� �5��s"�7A�Wur�N���۲g�LkѺuݮhδ>�V+b���t�&�ٵ���R�g�u��]��m��;2	�7]Jݷ3lb�%��d���O=�=9`�c��*wl�C.�2@ڶ���R�hX��dS8�U�(0ii]��Z;Z�XĻP��h�I"z�ۮ�<D;E�� ��[��egUUϕ8.2���Y����U�0u�`��#�*�P��g��c��L�E�Q��U�&FRy�&ڪ�U��8nd�`At ʂ�UU�s$젰�uh�a��uZ�Y��o[(y��nt9/h`q[@*�����UmN���헗<�����]a�g6�[�+���n)SSP]&1�<D��]M;�{d%���h���|�Źڝãcsɥx��q�h�@bv-
f�F�����/��T�t��ڦ�2g̬ԅ�Kּqz�Fy.ڀ^g����W���j�ϖɮqO<�Wu=@܋P.�Q88��w*��8��n�����)���
��uQ:�̸��]�u1�d,=���69�DI�+��]ӗ�E��� ���*�KR�����r2���\��0��u�����N��5w-��@�DC�?!�׽�uC�� Ph�C��U�w������w�_�$ ��mm��a���l    \[u�>9�lC�Exӧ[��.<���u�����c�V�q�'j����,���L�ή�A�-�v�s���ɶ�sR��;@,XqC) ���3{P��ᑶ�&�j������ކ�2-�k������b���Վ^ɨ.[�<�0���-L��Y�w��:/�M�v�k)-0nz:i�IU���-J�
�p5���nz�b��i�K�=dͻswdNı,K����Ȗ%!2em2��	���e�ir<B�!2uu2��	��	�ΞL�H��4��.l8�D�,Kﷻbr%�bX�}�;8�D�,K��v��Kı<�~�8�D�,K�>�̛�fۚCsr���,K������%�bX��{�'"X�%����i��%�bX�}���,K��w��st�͛���s6q<�bX�'��6D�Kı<�~�8�D�,Kﷻbr%�bX�}�;8�D�,K܄�/iw	we�Mۻ"r%�bX�}�v�O"X�%��A�{��byı,O{�~�O"X�%��{͑9ı,OUw�/z(Ȕ �$��r	��4��)�l���ktg�*)��kk۩�<������nf���%�bX�����,K������%�bX�����<��	�������Bd&Bd.讖��k�幻�'"X�%���s���: ���blK�w�"r%�bX���v�O"X�%���ݱ9ı,W�w�Ks5E9���T\/�&Bd&'{���,K������yı,N�{�'"X�%���s���Kİo�w:n]-�nL۹ww"r%�bX�}�v�O"X�%���v��Kı<��vq<�bX�'s�܉Ȗ%�b}����ͺK��I���É�Kı;��؜�bX�>���'�,K��w��9ı,O>���Ȗ<oq��o���R�j��z�v�g��W������b ����3�2�悺�gM$۶���؜�bX�'�}��'�,K��w��9ı,O>����<B�!2uu2��	�������l��b[}��oq������~DND�,KϾ�a��%�bX���lND�,KϾ�gȖ%�b{����.�.�I�7lND�,KϾ�a��%�bX���lND��`�C��"r'��=�O"X�%��w��9ı,O���;�wst�m���yĳ� �2'����'"X�%��{�Ӊ�Kı;���ND�,KϷ�Ӊ�Kı=��Kl%�r\�7v��Kı<��vq<�bX�'s�܉Ȗ%�by���q<�bX�'{���,K���ogrm�$��I�m�]\f�ػ���\q�"�X�t0�� V�[dQ�WNJ�{���oq���w��9ı,O>߻N'�,K��w�br%�bX�}�;8�D�,K�gs���.rnݷwr'"X�%����i���9"X��o�9ı,O{�~�O"X�%���w"Y	��	��E�L�HsRR&����<�bX�'{���,K������%�bX���r'"X�%����i��%�bX���;3nn�4��̹�'"X�%���s���Kİ~���r%�bX�}�v�O"X����2'{��Ȗ%�bw;��sn��3sK3n�l�yı,�{u9ı,O>߻N'�,K��w�br%�bX�}�;8�D�,K�o{�rm��m����6u�뜼�{��������Y���r2�H�'Z��f�+��Kı<��vO"X�%���v��Kı<��vq<�bX�s����bX�'���̻֝��m���q<�bX�'{���,K��s���Kİ{����Kı>��vO"X�%��]�Z[a76�.[��br%�bX�{�vq<�bX�s����bX�'���É�Kı;��؜�bX�'�����e�sK��vLݜO"X�%���n�"X�%��s��yı,N�{�'"X�%���gȖ%�`�l�tܻ&a7f���۩Ȗ%�b{���q<�bX�'{���,K�����Kİ{�����Y��g���~~H� �  ���I$�  8    	e˫���h��s�%d��I������,��<v��F!��e�ql	 pzt �z���ӡ����.V�n�r�ԥ� .�68fP�Ʋ�A�擇���#�UF��m�c���q�Lsm��r�9jm���}{r��Mv�M���m#��GW�}����0�Y��w�I��jn��6���HY��Nw;8#��[6���d�k�/nRhv�MƋ��M&i��N'�,K���m�Ȗ%�by�y���%�bX=���r%�bX���v�O"X�%��O��v���!��nm�Ȗ%�by�y���%�bX=���r%�bX���v�O"X�%���v��O�ʙ��~��74��74�6�͜O"X�%��?~���bX�'��ݧȖ?C"dN��lND�,K�{��'�,K��$����6鹙�I��u9ı,O}߻N'���G"dK����'"X�%��߹�q<�bX�s����bX�'���̻֝��m��m8�D�,K���Ȗ%�by�y���%�d&(��t����5��BK˺�S�; �N�Ԧ��9n��=h�lb��ׅ.�#��MGh�(p���A��m����~�"`n�B���0=,�]�3L�ɻ&n�I<�w��|I�BE!	,P�'�wZ+vw]���ZX,G>��N�$R��X�+���&�d�"`j+e�F,�^Y�^U����0=� ���w�q`|��$T㔩£�N+��Ł�w���޾���9dŖbE��5]s�T<a���O/<�p����:벚�e9�����L��fu�k'�O��H�����Ll�05�!D"�q�F�37��������t���_r�>���*Aͩ�D�����gݼ�y}�s��vu�|���B"#�w7���͸�?dNKi�-������b`yl���\��������r�T7(���H���+3z�X�yX,�vpt����$�8�cvMmĘ��mt�}ڍ���㎩wv�Y�g�$��F�*u!"�����޿���L-���"`j+e�F,�^Y�k*��u�OԐl��z\�����h�t�S�R�
�4�V,�v��������7^�5v�8�D�/�-��r&�d)��}������U_�I��A��(�)R7N��S��&��lI�`um���`���!�������w�����v�Ĝ�ź�����^6���a+¼�?&��lI��U}��A�3�Xߟ4*A^r?�m9"�>Y��I�`n�B���0=R,�Z�Y�D���G`}�8�36qV��V�;����s�T�N�$R�p�36qL��[%�=&A����)���$��*��{��RX��v{���'������I??���G   ��m� ��l��    3o\6���nî8�tW�͵Ԇ����s����YS�rN���t���}ѵ�}�v�5ˀ�Gq�x ݳg�l�e� ���V�tV��'N�����u�����gm*��$�n�3v��xqt7!71��g��y��=�m�g��i8)T��Ĺ�]s\:�Y��j'(	�# @͛y�w7.M,�n��:5���Yx+v�{�����E�:�Kj�Ɲp�GA�)2*�4�X�����t����n>J~a�;����Ή����,ʲ�2�� ����`w_D����`b�qD�2F㠍�`fo_�u�L-���"`{�IR	v�31b��g���[%�=.D����`{���*AR�/�]������-��r&�G���& �^,�����մgN��/6�bس���n�`���n�bg��^St4h��I��ߟ��������[�Q.VZ��-ݛ�L���O}��y���1�D�uA|y��g|��}}�;�}���Vs�D��8)I�����[��L��S��
�%M'E5SR�Ӱ�	�s�lt�;3g`n��`j�����ǈY����w����[6������
.q��ιݪ�k˸4Cی=Ϝ\�@�zuַ�1��gl='Uөr�1^�e~��0<�K`zL����}IRm)$�RI�,׼�-��� ���0=�_Z �y�B�W����[�d�궨��2��RA�V� �-\	QH
�N ĀB�Ԯ�F���B�q�9�@�@H�H�|�*�Pr*�*�V"�H1Ho� ��80 E���
!��8�T���: �DcAdR'P"|81	a11pɂ1}��  @��	IKkX�H�!I[d�f}x��)r�N_)B BiKmR�Ik-�,�*HW��hE9~��$'�@�� ���N�>*���T�>P5@���3���QO}�}��eA���LT�!E�ff],Fa�2�� ���0;��`yl���b9�F�m7 ┣������;��`yl������&,�K)����:��r�6�d��[ewp[�s0`������k�c6.�����z&��lI�`n�TF�f+ND��GN+���I�O�J�`n��`j��r�E%1�)��2�ʃ��&��lA��$I)I��'3eq`n��`y}�s�`ӥ �TS�������!�RI"���X�yX,�lI�`n�TA$Yf ��I�4�]������ۛ�[V��M(�ݺN�#d�s�ɦ�(Щ)P�NH������A���P`w_D��H�YFfeҦU����Z_�ٙ���7gy�,�w��U��F-G��5i�	��+����[�d��}H��N!�JM�,׼��w;�}����\X#;�NP9EGW���[��L�ʃ��&����t߿��  �l�A�����l� 	    m�zo+���`��)�8l��K�F���c�����Nѱ�i['[e�CakY��r�{Y�t9�E��6�UHMl�+ԚUI2t���l�C^��
�_�8����8� ��yz��5rP��qº�疁GE�͸�mƉ�7h��`n�A�I�V�����-+����3�Q^�rmq5��٣Xt=�N��R��.I&r�pT6h	%"D)���yX�+�u�+����ԫ�#dr9("p�37*��[%�=.D���q�iI$��N�`n��`|���s�Vf����=hT���FӒ+�[��L�ʃ��&ʯ�������R'J)�G`g���͕Ł�������`fwDGLNI$�&D7=T�jr��2���o"L�U���@r\.�ʍD�NB5)������5n����g�I/�=���bΞL��:�u#��U<͛��D_�(E�����d����e��^QYyb����lI�`n�T���5v��)��������q`f�T���<�K`r��au�yv��1^�ʃ�����lN�X�.�"D@ �S�TQ�>�	wFS���w�m�2�¸�wkh��2��1�br�eڤ��[��[%�=; ���\Xo�
�1�B�m�#�>Y��(l�mq`fm.,~͛䡳˹׊J�DG#Q���Of���C�`�B$F�D	F�H]�	�S���1��l�������)�S�����������`|���wN,Eg>�H�H�b�Wx09wK`w�W�}2�� ���ŀWwu6�1	�%8�u#���?WA��\g�3�z��.!y":Z�:]*L[�1�d�����yl-��� �����;Wo(8���RT$B��wN/�I�3k�^�M���vo�BI�o��j6���������ջ����-��2}��
Yw��j�SE�=�ޛ�;����ZXbK�
""�d�;�3�>hT���n9���-����GL[������W; �[7�]C�=���D�[��	���l'��+E�L�͝	���g\Kq2�O�=; �����z[�d��"\��JL��,��Vo;�����q`b+9�"F
F����f����6t$��mq`foZ�?#;�r%NQQ�'����`}�8�=��V	%gw����Ή�UEHI
q
G`}�8�=��{�W�r��>Y���VW�+��@�I$�I#m� �kXn�l 6�$    ���a0���s>�AS��b�=cq�:2h+�pS/��If���wi�e7Gn.1;t��,a�'&-x�];�cz��ŷLE��}!���-���'Q�96�*�㛉�O(ĵ�y�v�uu��ݛ�S��Րp��l���qp�0C�A���e�+mP����'�^G=Hⴿ���w}������$�:�u�& ^����e h�]��N�K�IN�ѕbF�m�(�j:�0��Ձ�w������IB����Ł�����I���F��`c�پ�J<�lt�;�����)*@��
��$���gs�>�ܬ͜X�y�Wr�P�J7*7��^e�=.D����t���z���,G>��JT��qJjE`fl����-��[��L	�bX]!b��R#Q��t'SώpG�
86l��cn6�q��q��r&(�(��#��,[��[%�=.D������w����������f�6��?B��d��������Ǚ�B��}��r�R�T�����zx�36q`j��`|������7Nf�,y�6��ٰ�BO��Ł����y��lbI��ջ���gs�>�X�8�:���"��$�9C$����hn��@���e�v;7^�,�l�-Gh��c�A�
I�$���gs�>�X�8�����w)�5?I"JD�r;�|`���K`yl��ը�+

S%)�*jh�=�,y�6dDD@X*
�Ta��$%������	��$�5�{�`{���<�흥`�j1JM�«��5os�>Y���w_��O3o������6���jGU6��ٰ9B��w_�����ջ���MS�����J��
5Rns�[l.�ղ2��9ۨFC�^.*#���%7%1�H���f�,[���w;g#�P�ܔ8X��`r�-��[d�?�_|����La�FD�T�p�9wy�,�v��07{ ��|vRT��%wyUSa�1�vl۵���eiaТ�$����B_CI/�{�M���u�K�U�,Yy�����d���<�KrO��?���Y@Һl:��4���bهm��㱴ӻ��z�=(�7I����t�b`n�A�nɌ-���W�U}^A���`j+|�J(�rE�&�`���I��v��������gq"nTM�U�I,�w;1�+3g��,U��
J��qJc"���"`n�A�nɌ-����%H�A����ŀfwK=�����3'����yE��9P�_�@�$	O��vJ�ZƢ��L �G" �`�}�ш�c	��F���7����$�/��C�<a	�s�Ѐ�d
�N�p�
�\ib�� oO
�))�! � �� + ��R,#`�:��&j)I) @bVV���!��/������c�)�#�A'�$���,5G�U�'d/ �"_�����)�eUi<� �����"����M�r9,%��3I� '����{�]��ˮd�߫�;{t���{�  [@��         	�      $       p8   �l6���}��     �`     .�    �                     � (��Y4H��dj�i��X4�8�z�h\l!�n��mx�z�-s�[a�k#�s��ь��@��&I[@c�;)���'[��ʵPV�v�g�&y7n���g9g�e�@4��P�����3��N��bR����Ph�qZ��[<�#�W��M�sи\�Wl�/q��:�l��tR�ݜ\���`��y��a=����(�N��+��g�J'�w�9���γ� ԛ���۶��[�'��7�@촻 c�l���,v땦Vڝt�u�� �e5�<U��&v_<Q; qz:9vUNn2���է�bM��b�J�Ҭ�[.�2ʪ�j�N�]Z���*���57Q,$�UP-�֧jZ  ���+<Hڀ��ɐΘ�v�T�����UB�OI%� 4�6�d�����kh�t�;Um@�,	Rz���W`6n,dkiP�MD�*�UҮ([H49�ö�R��A;G��m���tqF��'0�	�b�a�h�KUl,�du ��%Ip��l&;Q.{gvs�������<��5��Ĳl)��z��D�q
ؓXg4v�q�p�v�qխ�X]�g�;�Q\ƀ*��Tjr1�p@OLnܼv�p0�����P�OԨqhSy��-�՜m�)s�$jB��T�K]�lhTt��,s՗����`��R��63 ��z��3U،qUl��ݻF㖫�(ٺ'��Y�@�L�v�a�L�3�x6�!��
iܯ/J�Ž)���n�zm�ul4�Δ�:Fv]��9�κ�v'iz��.�%)���H��ϐG�(	��"�Q}D����G�3�@�@���������"@ l �kX^Ӷ�     �f��� ��t.�vy��\�'���8����]����s��nQz'��B�l)9��8]�,n�-�x�z݌��:I1����h4�as:]��'-�U�ِ�;ZP�r�^��k]�G� ���팺�a�k��dƋHr��� ���*�	l;iݹ%�v�������#骩AHn��ۻt�-�����^
���������G,v$S��=�8#�Յ6(�r�fxlI��J��p� ��K����}����Ł��6RT���(m�w����-��2��0�1���S�jB���qG#�3:q`fl��3;�����`b�k�J:�t��`n�A�nɌ-��� ��Vs�QGC�(Ҕ7 �ޖ�;���Ӌ7g�tQƙ) J�9���m�^&89{3˯VN֨l2<� 8�i%$"8H��&JUbq�-�v�Ӌ7g��v*���Tt��Y�n�rI�{�����&F��B��BK�BHJ�^�>���ٿ�%	6c�p�P�f�9���3����-���[�d��k��y�*RD�>�w�����`~ݭ,:y�|X�6�i�>T"�o32�]%�=&A���.�lݓ���YRN��đI;/J�������m�۞y��w�%i�n��g3�I&����SU6�����ei`c���
!%����b�y���Q�B%F�(�`fl��UT��{��ž�>�X��}J)N��F���X�y�,�:r_%��,Q�U�|X�_���D܉2R�����gs�3����y�֬{�6���SS4����EY�2�&A������l.�vՏz%"��'$�d�P��T����W�nkps�d�+Tc��pF�jZ�4^���GLRK`yt���Ӌ����tsj@H��`j�����-�Ӳ��J��|e��̶�Il� ����˻���v��5*�F�)��ӎI=������{�������
x%������l��]!�:UN��������z[ˤ��d�Ԙ��; �Wb��X�K�5ik���8�Y�e�L���.�Sq�I!rW09oK`yt����{����&�M�Ucq�-�w���F{��{�u`j��`b��RF�8�$Ȝvݳ�7z��%�{�����5��IR��n+7z��՛����-��}Զ!]��f��2����<�K`z_D���	��{������   m���l� 	     �$���O����,X��W%�a���̂Ui������|;�r�\n���8�l��yn<T��h/]	��7=Y����:�kkuL8�88v�ZjU�[qg��z�*�v�\ ���[*���ӽ��Y���vjy�����Z�fL�c�� ,�m�\��vn�����zբ7�����!sd�yw&͒e�f���� l����_q�M<Upi�qӞ4��q��X۞5�S|GIR R�ۍ��yw��;9�+7g��v�ڧ ԥ��������k��J3v��5����n��l׬��R�AҪt��vn�)��]%�:vA����)b���ҔӅ��������`ol��ߢ!(P�n����3Rܔ���*j�]%�:L�{�S��
�?��Ypz��q^�ע�ˍ���nLƺA�Iao^��C��
6t�̖e���; �����n����-�f��1�)���#qX�8���U}	(#�D"��]�1�t������RM:9��(��,Y����;>�P�t�;7zՁ� �M��N
����`yt���}{��-��Wj�R�Q�����{���$�3{���������n�*h�; �V%��/��C���;�2���ۑ&{�-���%�r�4�%�v.�����09l����-���&��\��0r5R���Y����;9�+7z����B7Q�$���#�<�w��'�ϻy>� �ŀ� )! "/�T=n��~��'��g j��RF�SN*q	�`o=�`fo]X�y�~X��v���2IC�wYtw�������l-��/�X�.�"D@ �S	Q��v՝ќ�r��m�,��6Ñ�+��:���O�\���bB̦)��]%�:_E�����Ձ����R�qQq8��Io�D�s�`wOΘ�K`z�Y �J�HܐQH�缬��Wo;���պ�IQ�Ba*4�)��BQ3{�5�����f�5"!DP"�G��$��HFA�I2�?����}��גO����v�#Q�(rU��������`o=�`fo]XwwB
��$��Q�RA��(i5f�ӵ�gGD�{j�Nwa�t�R6�Z��J�%M�I����`o=�`fo]X�y����ܧ)&A�'��9����m}��}�6�wM�M�r^��#����7��޺�5v�`yl���}ԶP�������16ꕁ�sf����6l�J"P��{�3�r�*@z�����`}����%�[���֬{�6+TB�w�ޟ���ߤ� 6���[nkXd� 6�$    �][��ax�����m8�=A��(����G�뭶���"�lE:=su�=9�ib��W��$6Ǧ�v��ІԶ]�N��jW�b��V^ں�y�R@:JgtM�R8�T��,R3՞ڶ��տ��o��6��y��(QvnϚnj`�8�>9����q�[N�l�\�7e��w��{���~���Kn��Lnu������s�ۖۥ�5oW2�&�̚4���&�3��%$\?+3z����������+�s^��R��A���X��LS��=�"`t������)bX\�F���V��v����������u`|��!�)��7$v�����Lގ��K`r��^]�U�%f�+���}w��mȘc�V�z������DԤ�%;(`'Y9x���Fn�%h9�sօ����)���BJQTT��7�@3纬�� �^j�9u��D�9A�������O/�>
��UO}��=�x�����7���񲒤Sq�#k/�}e�LoGLۑ0=[�pP���qD����{���7���ܬ��+�]%F�	��S������;?~^z����}��o��Kg�b��2�k�@�N���x �*뱳)��gn��He퍦�4�/2��"`{o�`l����W�������F2R��jE`}�y[��/�`n�t������$W�w��%N'N+�{���7�������0�sb�tW�3�B8pH x�XG�B�"P4�}���.��q>F��L��|`�uh!��E1#t$4�9R�h	���d:t�������Q�L�xp�y��F_:�H�d� N�R�Ĳ��r�e0�e332���T�@͇(ՀF`�%�(Ry3$�KY�0�$���xS|N��zӎ<8�'��V� �GQqU:�B��^|)�S�>E:�'�(�����!���9��������]�*H���qXf�Ձ���`~���%	�V�<�9��E"r����q�+�{���{���7�����H�0I9$N1RRLs��uP�g�K�Z�����Y�e�Գ�ּ�b����Q�`}�yX�yXf��������;�y� HL�K��M�b`l�������r&��&��J�D�RST�)���u`n>�`}��X�yX�}J%#Q�(��`g�u��;���Ӽ�.�D��<"��y����$���C7%)L��8ґXc�Vs�V�����������(��% 	$�*M�UF�6:��{:��eX밧!�C+�v๮��q7)JJ�N$�_�}�`}�yX��|�Q�{'y��}j�MP����v�Nk�P�"lܞ�`{'y��yX�\�3�R:���n+v�Lm�L��0=��0=��� 9�*$mG��>�`g=�`f=�`n>�`}]�ps�Q��+'d��0;nD��܉���}G����  �` �Z��l�     �Ҭ���\ۜX]j�����4%:G���_g�LH+��ٵu��D@\�^�6�pH\m�IڞP%eU@]qn�$@m9vM��ff IƲ���!'H��0)��i963�Q`C�tޒ�f�k��k;�������[���GS�H����SLl>^�R�{������>����(�]Y�n��	qa|[��$�����gi�{mκ��Ҭ�t��WE0RL������>���}ޖ�C�ԢPr5R��7r�>�� ��Ձ�Ӛ�(���gqEL���*N4�Vk�+ �ޖ����������ܙ��%N'R+ �ٌm�Lۑ0=��0�U�,$�ST�m�`}�yX��Xc�V��,�{�)�	'$�	GQ���O�;q�;���71��g��g������I&D�tDnP�M����V����goK�{���)/ʎc��Q�`}��o8�@ $ ��H�"C�(U@�6�d�=;���ˊ�l9Pj8�RE���,Ǽ��ܬ�Wꤳ_��]�zJ�F�**`�cv�&mȘۑ0�1����ԢT��6)I8��ܬ��+ �ޖc�V���v���Gd�]#V��i��M� �a��s�%k����1��*TB#�H�%!B��JE���V��07o�`v܉��#��2��Vax��LgL`n�D������n��Hj�$5M6ܖc�Vzw]����FD$�5�~��=��?v�X �3���$�V��LmȘΘ�ݾ����줾TKTHڎ+�}��3������������8�q�  RI?9A�N.f���!�ca���r�۬\%�9ڛ��m�I�%$V��,Ǽ��ܬ��+��IQ��5%D�I,Ǳ0;nD���D�6t���.RĩI"lR�qX��Xc�V��,͜X#;���JTIƔ���f���6�zs]��D
!!(	xU1��-�~�/$�_��n9I�N*q	�`����{���}���gs�=_��+�z%"��'$����׷^]��&�s=l9���u�N�j[�)(HcNR���ۓ�7_yX��X,�~�����1��"9)�J���L-��Θ�ݾ���!%��6�p��JU2�i�y�6��07o�`v܉��ȀB���MF��UU~K}ޖk�+q�+���Ŧ��TjP�ԍ0RKw�ۑ0<�K`:c ��}�ߒ�~H� l m� ��p�8    �,�On3�E�U����֗iL�k�&�0#�/ur�۶�����[n�Rl^����J��8��nw\��	őJ���[$u��D�M�)^ۚ9��:l�JҪO�s���ܢ��!L�M`�s��s��7�c�
L�SN,��w��K�gi���P�������{���>�M�v�lOH�۞A/N�8���c��!��؁��n��ڴ�"Fu[�Dآ��{�`|���v��36qa����#UP'R+���6t��d�"`E�Y�yJ�7
q)%Xv��36q`n>�`}��V���	rDST�m�`fl��r&�GLgL`j�e�3)eZI+���r&�GLgL`fl���w(�@@�8��n	�����nJR۪��r��zU�K�V\�1��x<p�8���_��]Xv��36q`n>�`}Z>��DEI9V����"z����ܛ��e������w]X���J�JIQ�3��`v܉��� ��#�R�R�Dآ�������w:`:cw�#d+2�e����b`{dt�6t���Lۑ0��{����~�E�0�z����>Nщ��5v������"��η:M\�at3���)Ĥ����,Ǽ��ܬ����4ս�U!?5M6ܖf�,ۑ0=�:`:cPl,�Y��)m��vzw]��۶��$�G�(QC�ڰ?zs]�� �M�C�4�U2��0=�:`:cv�&mȘ�r
D�TQ4��`����{���N�?{vՁС(�;�L�)ʐ����7=�C�g�;��7#�c*OOn�Kc��G��r����]���ث����_����vGLgL`yr�%K31]����L�0�1������3��TӔ�4�Vgs���07nD��(�����N�p�$� �ޖc�V��VM��)	��C�nV�|��|X��
��I��i��3:q`v܉��2gL`g��ĤŖbB�$��Ƥ�s�ʼӶd��\����Y9һ�]u�a5���F*�q�m��?ˑ07dt�6t���0=���ʅ3�̼L�0�1��2�ܬ�G܀Ct�D�F�r�;f07z:`v܉���Ww3+-R�TL��U�B�y�ߕ��=����� �ޖ���ԢT��6(�%X�"`g�OW�:K�=��L�W�}@���������*��"�*�U��TW�AP_��P_�UQW���@�E `�@�����P_��P_�@U"�*��
����*��
����*�� �
����*��
����*��*����
�2��;���:�����9�>�j�    �:         $P    @  �� �P ��(B�HIP���J����AE ��R�$�H� ��AQIT�%@`   �QR�    
Z�5�R�n��y5�Wz�-:_x �{�}z��jU�nW������|�n�����<  _O'ӽo'�>�	ҙ,f��qeu�O�_pN�| �  =� ��Ǭ�,*�@     X ���Uͯm�UV��QdԬ ts�ҹaWsr��ﻪ',` 6�Y��YW\ \YUf��� �B�n�����ۓ�N�=�� =����;��Ω�Jw�� @� � ������qjU�'��YK� rS&���<��7+ӓ��� �"tq�  !�bt����}�9>.��w=i��)��� ��n-v��ξ��ͻk����}���J� *� �� ϕ�����u�<[�ks��{ހ��}�2��,e4"��} `D�����v  )ف��;: �f�4iفE)���b {� ΀  "4��% �  �UR��  UY�()H�(n�J �E1�p����ħ��y]_y������� �*Y=t��� ���ӽ�N�/� ,���Zw����uK� ^�=Jͻ�uy��M;ۼ�Q� z�)=�*�@��������U4�# �=UI6��&  �"{J�e%F�  ��(ޥ)P  	�)M" <S�O���������?��|�==�{��9��*�5���*���E?�@U��*�����TQS���N��O��܋��	���r��"Hp{��L5�S\��P������)�*J1!
a�>&��j�:�Q�I	e���r�d���^kp�p0���ŀ��C����i!ql�$�z�L�ȷ1��˚%{��w��L�Ip�BBP�(��H����5�.o�|O�@����t���˶P�D�MVT�J B�Co
R4�7����]�oZ&�r�y��ˆ��&�(S���)(F`@�!!H�H��\H��
�l%��u�^�wD���	��.�B�w�%	xK��o8^>@]3CA$
a�;ŀV%1!L�S��Ğ5
Җ5 � ċ3y �{�p�\�����0�pĆ�����.��;N�i
C$#H���s�������@4��-0��f�i%�\��˵�HHp#����B�L*������V�)]Ń�l�)��ߴ�[���ё) �ߓ�)���J��� CT���%�0�����6oh�gn����`j=vl�nh R7F� P#H}�æo{Ð���T��53�S/y��M��!M�h�z|@����	��I��}
�S����=��hJJl�ǈ^y�IXV��Ł�:K�籙�H�a� D��� o��n���3����>&k�ߐ�K��I	n�I]�0�C$&�le�!BY4I)��0���B�J�,�����Xf�ϵ�F���0��|oA�����E��R%#P �	b4�<����-���~�k�/�n{�cd�����xކ��� ����\�%!X �F��g.��s5�3:�d���̹�٧����,`A�æ��G�h]o�%���~<jV}
g���^��M������뒮����e�g4K,!y݄����C����ݽ:[��|ߡ���}��)�e����5Γ7���d2, 0H�b����F$H�`�!Hk�4܅f��P BK��i��k�[�7��������sa�:�)���H�H\��c���m C�
�HK�$�JF$o�&��dֶk���7���'!��iYa��B��B6%H��!1#qH�)�3F�F1ٽ쐗\��88@�) BC���Inkz� Y��� ����I�Y�l�-l!B@���7ԡ�) T��Q�5�B)0B$`B��b�$ۯ�cHH4LLM l��ăd0���#��4ɢ�f�	�0R����!�Ie�C��n�a(��XDj0#=�%�޷�s�\�g����J�(��B�)7s-�|����h�j���$��b�B:�&�5�ЯŅ�')�̇Ғa[w�ː��{Y�����F�X8<֝f���S
p����f��37��͛�)�f�RVr^롛%	��)
J���i@��ٽ]��3W"I#���y��t-���}t��5���˝��{"H�u����U�v�j\�۰֦�0�&[��R�Ĉ2d&3��%��9�<��!H��bF#� �64 ��$X� @�Q�0R��D�1"D!$J)H$��1
�"H�T(`��"0`A��
�Ep+ELh��I @�E�E�D#�X�D�Q"@bҤ�)FV���`i@)$J%H���`T�DaX�A�VJ� �L!$�`P���!���c�!FH[�ې�MI��#$a"NrNe&�!J]�6䕌!���A���Dq$I��M��D�B����0�)I�K�B��HJ��+��2�I	a�0 ؘG��F��X�5�IIrJ��hDkH��%�4Lo�6LO"��=9��ۚ�&<3!)�a5{w� :�36������lI�Ww�I�%	�``iaVb�@�9�$�04ofr�5�����v��
B2��HhHD�3Z>�F# �`F$�cï��Dng��a�xp��&BE��+�$���~H���\�vh�� Ire�y�o����}�}S��n@*˼14~0`�0��rs\��v��h%�D)������S���\��̝��5Ӽ�}��
-��	�����P�T����\5��h�i�sl��+�4l�04�*�@����Cq�0 S$x�{��%o3�}
���w���o_mԸ�s�k�r$�*N�%C!X��P���! ��dH��E����9�܄��9�8�9u7�k6m�5���H��a�lJA�p\D5y~��HX3+c	bF�
$�BB2$cK2\���"+�C�	�bH��֠F%�{�L�X�B- �swz�y�K�����&�7�p�͵ ��R$$�$j�B�����jv����9vc`��<%Q��#��2a���1,t��_��H�Xbܳ7�	��FkSwF�sF����
�y�oC9�5f��pd$$�Md5oщv�6t�LsFa32Z�hB!1�I<y�Fᙲf�'��90e�f��6��hÌn[�roE`� ,
%�.���xH��2R)�1%�bD�Lյ������]�)��`bX�"ƌ��C��R��YK3E���r�����)/0ӌB1R�D DH���x��4a�R0�d���6H�%��!njJJ�	\$��Ddd�C3�D&�H��XXF�F!*�X��R��=w7�ܜ��<s�8c7�2j%�IrI��`�qz�!:0â�!)1#XTԤ
��D�.o>ɽ��٢S�9rܼ�e�����v��5�$eނ\Ѡ֖4�ZA"@"@�#Zѩtm��!̈́+�J8m�$���GI�BF�24�.�˚�5��,Oj�b&&}����;�	͚��k���L�0�Xh���[��|��'ݐ��.IFė>�Iu���q޾.C<�!��x�h��|�9�_��o�&d�HWm!�ČC�!�ϋ$.���;���6m���o����%)�Mĉ��H�d�s^�2j�V[�5e��Jl��5��)��j�!�2BK��Z ���1�)#r�G��̸S}),Ӕ�Y\��ibحa�M�~0�����$ �Lf ���a.�1��S&4�9��q!�%K�0028i�3p����z8r H�-aB��75ÿl�ׂOfB$��![%d�#iIK��C4L�Jj����%a\%3S�v�3�&�m
��5��3�w��,�a�H��Y�2ˌJ�F8�D%�)p�	rSeaiIZ�Id%)!H�˒�K�Z4�$ F3�\�O{�:E{���Ӝt���J�$���D)�Be,i	���iC5��85	4̒�-!i�Camr%4��3E��S;�&��C�D8s�
Cw�d�0,�!0�Z0�(`¹ "V A"��a�h�H�feΐ���h�2��X�!�!u���S
SH�j��%��
IR5
HFH�V@�V! ��"ZM��+�%�i��@H�R@��Ԉ�(l�#WVi"F� X�IW�,5����"hb��E(P�@�AĈ¡$Z)4I
A�Jl��00%0��p\�!p�j��1+)d�2KjB����\)	$$-L\�)��"B�fC5q4D����1���JbH�+��
VD��ef���� E"�l%�5y�B�i����߹!��a����٫���o���s�޸�.�����6a�h�M�0!�%"\�Jh�K��9�g��ӟp���G���s��Y�9�_t�db���l�����t%�p!L}y�h  X|                                     6�-�      ��                �K��          �   � m�            m���        [@     ��h 8� 	"m��M٭�k�D��u��F�Zŧu���K�2[�i���v��)6溕fy:��2�9�p7 ��.Q�9��p�[S� ��)-)<�u��ij�Iڴ��%�Vڮ�m�88�U2`١�j���  ��۷m�llp m�$�����-��(   6ٶ��`�h6رv����ݶ ۰�m���8���I����6:��RՑu�h�R�\c�¢�i�	   �f�R	l�J�UV�pvCgm�Y%�n����H   �  m�$ ��m�m��`    �-���25��$H�  H�gԖ�   � �� m���Ɠl�m��4pA���&�%� m�:��o]�Z��`mH  [x�4� ���lpW����**M��$5R� 	m�h � �ŶG  m�m����@R�t]c"�*�ԖہmH  -�l p�� �p �6� 6�    �H  8   6� Hp       H -�l [C���h,3�m����`�[@�h��eYV�۫j��-�H� I4��m�m�    � �Ӭ�`�� �   ]6�ڲۍ��I�  zwf�n��  �ׂB@@l�    %��6� ��� m�X[%�m�   A�k���򲲵*��-�l� h 6� -�   $      $	5�  �.�0�Iz����ݠ*�U;�n�� ���6��/�rH�u��  7m��� ��[v�RG 7m��    	  6� @�h��  -��$H d��l $8 ��l�[v�m�
V[B�ҿ}W�UVƅj�+ER��A�o�W�N � #m��K�͹�C$$dsV���χ� -�$ m�  -h����� XbCi.mk/BI0'Rɂ@ր ���"rf�v���I!���-7kH��M��۰�-�e�/m�����"�3��;0�L��a� ���Um֑U[uǷSm��n���Gv����].sv��*��3�k8ŵ�- $:�E�v�a��:�  ۮ��Q���m��N���$�;���ܐ�3vm���@�eڥ�I��o  pk;%�6��>6ˤ������O�v�
ڧD�YWj���ِK#gf�Mn�  R���J��Uc9��[�Úۯi�0]�$ש%�l[Rcm� 5[�'@�Hn�0:A �[n�A �j-�n�2;s*�X��S��8F]�v�	��:��BX���&�[lc��z��v�b� q�i6�ĆٷaӖ%ZTᗀ��&��j���{^ݎ�Ie�]�
��Kjҕ�& ���� p��:��^�Ie�  ؛j��� 6�ݗ��mm�6z��w�^��[RN�`m����A�Æ�X�p ��m��6 $ [I�	 ,� 'V�b6�6�����@+n��NbZ�TI�z��2�m�H���:	����zi�b��.[�vq�\�S�g�il"�`�8[V+Ә�']eiYN���%����`q%����2��x*�w�O��<�F�S�g������7S�����m�ȭ�;�j-���y�D�k�-��sK�Ӥ<,�vZt��;�dTB��v��V���~������8����t�:�9�j�m�6�j�f* ۶,;�M��W�]��R �v&�{b�;V�UR�Ί{j��m��w��/횮�` l�p͖��u�j��5�"\0L�&�Wc��:RN[�7�&��k��m�m�:Mk �� -���&�t��"�)��k����]�8��L�;���-8  [I +��]���|�a��`<�*�gq�%�m���pZ���lKd���	j�ɵ���Nv];V�   G8	��  d�f-���ޠn��k[eg� �GUm�U�+�ŝu��I@-�hsZ��xa� 	m�mM�F��� m�uuUW<�F�� v@� �`p  pv�[��vKh�m�m$H^��m� sm�mN�m%��tN�֭� �Ä��-�y����[��UP    �󭣅�pm�m�	�["m�m n�U��M��N�d�����6�    jؒB��P��W�
�+n��j[N6ۃ��צ�դ�^�m��PڶI,�I0�f�8����G�f��   I::�{`��.�v�Zl�I6�m���-��EMw��8�8嫅�M&h  v�t�N�ٺ��T.uq���7,8ʹ�V� �鎱�6۰UM�Uc�Tq� ktݭ5�ٹx�`¥�� �����sn�K�&�����N&ڣ��K�cm�5N�4�ʩgh�nAb�s�� �-PV�u<��Gvwt'c5ՉM]�����F�n���B�� ��	��k��>��Jv^ � \�]Ft3�	;:�:ݔfI��2�[�j�v��~/���I��.8�Ij���譪�,��פ��ĕ����Ɓ���'R�S�m��vˬm��S"�76��� 6����]r恖UU�.�ꀥ-�@�o�WԒ�+H��D�� *�9ZU�9�;4Y�j��*qH� *��V6�u�RHx ���	-�B[V�+��4\�91{l0�Z����b� 	�E*�TI�@;Y��n�ծn�l�[ b�}+�zڬ�d�mY0,7��$�Iŝ-�A� ��M�8smm�v�_9C[��[YnXl�Ix�` ��u*��d�e`�iVږ
�ڪPI3����˰6�V1m�@	e�nH�	�p-;I���/q���Ͳ@I�;v�/V^q���c�IF|#�1\�f�V�͌�#t��8�����eo;��4�W�����Й���#�`V�n��W�>Ә&1fl��H�TZ��ne���6  �v�kI�H8   �6�  � h�m� �gI��cI���6��/J	-��ӡ�۫6��I�]$kh[@8 �[D�R��W[TH�km��h:�,5�m� 8 ��1m�cF��m�m�� m%��h�*�jm�fs
�L��! -�#�'ϟ�   ���f�Z$ͺ��vP�j���h6-k�p��l�np���V���6�Ė�A�l:,�VT�hJ�{l敊 ��sЬÜ�&�7f' ���] K) ��c:�x�  �6 m�ԝn�q�J���P�U��+(��U������!8�v�n��n�6�`qmm�)۝ �l���.ݵ�ݤu�dq� �'m� ��JKR���UT�^1����@�V�Y1�]��Uڦ%��8�*A�+�WQڶ��)�u]"�E���Z�I�m-��l$ @�g��l��#�8���ph�����]��Sv� ,�0i��qm��r}�����k�j����J�i^�_c��V�����VV�T" 9���m6��q"G �M�N��.M#v�x7\��T��a�m���ni��NZګv���9x���	m���m�   m�6�H-�-�!�ӥ��qm ����sm7h'-+uN�ڠ	庫�H���ֵ�䛭cZ��-��cm�e&�j%\:�1����VV�UM�IZu n����y�hl����a�p���Ř]c�M��8�|��:k=�- ��gmt2�H
��m��L��;R�T�t2��5I�rsr�تU���8v�;<ˍKU]��7�eTܡUV�^{YC! ��:()ـ���pn�{Y-�Z�HM�-��]F׫ڞvu����62   Nˮ�jڑ&R��|�'ͻ[w����� j�S�.�USq�����v�f��z0���M�m����� �`   m�ԲP-��	i$Ymx[v� ��  �a Hm[ 8m�o]�΍�j��V�R�U+Y[����;@�V����{`H��m�d�h�B�^b[�{�hS�y�m 6�$R�㈜��6��H8X�� �ϋ�|8�,5�����V��p1j�Z$�qg�/6��H�5����    6�m�m�p6�E�^�u{�}�
"*P�D�NT6�T��*����iERD!�!�@!b�~�u^�cX
QM��[J� �P��!�PQ(D�:@��D4������t�� �l"��> ���)�G�/X��Az/�>Qx���0v'��"E�C�+D5:*����pD���b 4����'@ �8�������@�
�
y؎��"���5:��ч"#�C�OPS��1���N��$��@��ދP�u^!�8��P�A��E�PW@0
�8#�T�*1v���ʏ�>>����*K[HʔR ZBZ�e��6 	$!"P� 	# � �@��bZ�5ёda����@�@ �� ���4��� S��Q<�l�>"�������D�B , �!Th@�+�b(�b�R�(����}׻���ӻޞ�����      �@l� 	e m�I�  m�  $�kS���ݎ�v�w��`�t���a4��0��7lj���\y ��j8�$){�a���Lq��UPY"u��T�ʩt�8T�6ώ��[R�Z�ڲ;X�� �-F�	&�@R�3�N��PK*@�j�S^G9+���RY ��V�mE�r�)�b��!*��6�;FB��+I��m�6y�w%	0竁�e�(:��y�j�%y��j��X��n֛"�)���nـ ��ZE��֫6���͐����õ��˛��"ҹڛ
�u&t�/��-�k4dC���b�+9�����\�4Y��˸��a:d.�f�Gu��I���{Z�x�x���7m r�ۧq=s��*��9Kd�4Y�|��9�-��v���6��`A�s�1ŕ{\�;l��sY��y�I����Iƞq��!��W7/0��ٓ`�\��
�$�z'�x�N��V������v�1C��Q�łT�ۖ������v
خ���+��7.�kp��U!�Cam��v���3�ԯd�:��:��ջ5JwR'YF\���Y6��e�D�=E������ۢ��h|-�m�6����\E�1��Qm�zDm�F[;m�Y+=T��U�r�Q@%����`�-�mr�g��A�[��h���5���Vw`���جq�=#���K�v��q�qP*1N��͘�ܻ@�+��ִ�g��C&4��6��%ˠ�F��2�m��:$���9�"Fgז#0T�K�G���۔"cD��8I�R�M�B�����W�Y��ͮ��7$�ev��Q����>�y�V��"�˺�̤�n�.ng���b������TnT�kۣ�du���	%�ɶ�j�0�8��I�N�Ʋ��U���w�4S�Dv3g��\�&qo<�����M̓K�m�\˶���^�����q<"�5E��@¤����CʏPZ�ER��P��`i4��"���җl��|��] �α��5�H�@r�WKD��p��۶
Z��aA筻wX�F�fM�n6�34�ݳ�u�λrq�p�\�I��Ҍ���)<j��g����7nT5��9ۄ^�X�nC�'Q��*�����N������mx�b�gf(ܢ�7j��÷e.��S%C�S��(n�q��(�|�l�,��2Ie�iv�9�v�>;r�ۼ/����<M�o��$}#�!�n��>���s�3=A޾�hgz׉�${��f^����s��b��[��{m�7�A�c�Š^r��ط ��T�[�u{��ͭ.�4�wsj �-�>y� {�����,�Ԍ��x�E�{yv�b�y�P�n���Wꪧ:�)ߵ�z�l�ыFժ\���ڹ�>9�H��θ�
S�VQ���0�|��� ^rT�[�{�*��uF⍼��1�H�s��m��Ϗ<~`�q"�v�����������ڴ��,k��N!2�1h�n�ϯV��]��/@����
ܤ�85�JŠ}yw4�n �l�ط �{¯��6��3wv�b�W%@�`6�h��3>�w��cIG@Stn�[F��x3�����u�q��c�r�pY���&�icx�&8�^����s@/-�����ڴg9����"H�h˰�� {�
�*~�����>�$�G`�����w4�ʴ�R"�"��H	��H�y�%���4�h�x�m��I��ᙵ {9��J��`+��s��T���d�	�
E�[k���`+* �-�=}t~n��9-����{N��dv�Wb������7�9z�-F��=Q��/i)8��b����o�����b�[e@-ma�҃M	���>��o�3�3<H�}��;ޮ�h�٠}�;Fbd�NdM��Z{��@o��i*�]��f�����b�cx�&8�ZW�� ����^��!�K�J�]�w�|�uB��HbL�H����@����9�j�8��|�+⭝���1t���,Mg<\�V�8a����kϓ�p^����$�q8dRx��`�RO@���9�Jh�י*�$��?I3@j�n�b��Ȧ4�h�%4+�&�{m���s@�r'cn$�ɒ$��Uy݀W`+*ܲ�y����1��Q�$���\�{4���h廚V�4����A&���`+*ܲ��� <��9������,��uN+B����A��UV�>��<���^h�j�m�B�<�ڹ�n��V�R��M�#�m�q��l@:�V�,��OFq��7��X�ܜ��v��%M�u�\��ҕڄe��hv�p��a�y�ќ�x�g֚���"CUcu��Z1��mؘ�t�\�e�Mv6k`.-Z�v3�c���v�2k�	���{Ͼ�/��s�xRbⶳ�)�����ǳ�8���1� F3 =C��Z��ա����m��~߻�:�݀W`�T��aW�u�NA�c�L�8��o䃝�f��w��9n�s��V��M�X�I&�}W`�T�e@:�݀�Ĭ���晁y����*ܲ�j����@�*.Q7�i4I�9�:ޭ����ͼ���h�UR���o�g{����S���T؋0��

��Z�p�O=�t�T��z��r��_ �I���y�?��$�����ܹ��щ�(Ӓh��[���E?�8:"�kP������74��w4+l�@�*����*�6�v�,�j���4s�h�L��q�$��癋���K�fh�y�|�ՠ|�^������6�qɚV�4�٠{m��/-��|�T��L#d��lR����cd�x�S9<nȽq-��Di}.�۲�/r�3wv <� �YP�T�l��T��'��l�@�,��*֮� yv�t�%�'D�1�3@��s@�ɢ�0�03�y癍��4���/2�8Gu�y[X]��@:�݀.�,�廚�s"uD�1��Q�$��`�T� �Wv '�.����q��`�q��v�M���`/�&�"0�d�4욥���>I>VT� m]� ����._�d��G#�L�/-����]�d���h�w4|��bmcx�nD� �� ]�|���*�ݦV�#@�D��h�@�۹�>��B�%�I*�������h�v���R�c�h�w4��ow��uw��@/9f�yņX4�<�3Z6L��pY��ͳ������77g����;GJ)�q�4I����/�S@��&�^r��n��k�$qF�	��+�� ڻ��v��T߬�����B�9&�^r��YP�* ڻ�ܛ�n�^�yWy����� |���� �h��ј�Bcy#��&h�w4m�� }���ޭ?R�]UJ��� *�Vb��+���֪�W��[���\K��*ەi�F��&vڨ�)E�RB�t�:A���啒�ܡH�F8���������t׮M��s���y-嫢=��8���cc���5�ݯ6ǡ�-��a�����H8�m=�z����n�N�W!ʗG=�\P�����n���8�7`����z��8�vݘ��l�Rn �p`m�n�Ns:ڠ�g���g��KC/n(�]/�qC�+���W��n�a�<e\Z��y$16���nD�>���y�4�� |��]գ�^�]��e�� >y��ʀw�� m]��9f��H6	���=��h��s@��&�{yf��Yx�Q���3wj��T�w`�; �YP�[R���c�f�U�M �]�|��Τ��k2��2�f�)�<k�ۙ�=Ol6��ݻH��|�5ֳX'�m�cF'�NI����ޭ��<���w$��dY�2�f��e�]k[�{����JC���^森�@����`W�L*�t�3M���ݨΤ�]� ���w4xe�16��N7��&�<� |��:���wp�ܺ3+n�7wv <� WR � �[d�;�mXof<md�&�6�ȈH\�vɷ]�k�x/��z8��엦��Wd�Odd���A0LrO@�{:h�S@�[d��f��T�7 �r"H�@�����&�}m��S{�Gs�w�5�2d�˽���i̙��e��~M��(h%��"A��bn�F�T�YsHl��K���J�0ąJ�7� fD���Zca(�٥��	D�5)�1�Ŋ1H�H�����6���Е<�a!0X�1��H�Q�k��Ig���V?'�ta�*x����vd��G/�xl���^�	z�bxzT���H��,bx�����8�fB�P-��ۄ�1iC{ٱ!E���x�����Rq�B���{H��&d-���x��Ft�����V1�cHBB�hC6Γ{.��#`=:2�D�ϕ �����tTC`<8&�*��������@���<�S���ߵ�nI����}�A�6�1��Q�$��%���I��^3C�U+��&f�@;"�H��I�N)&�m��/,���ɠ��︨��f�1�4G�:���ùĽ�&���ѓ��Y�9��GU�9��d���4�)�z��h峾z����}�l�&�M(�r7֮� yv ���R]����� �o�$a$�@;{٠[e4�)�z��h3��s�H&	�fh�f�����hb*�U	
� l�Y�k�ܓ��ٙ�.�.���Y�a�>�f��)%ܗ9�rf�ϟ��F�2)�d!�'���Ş9ջ�x�n�'��m_�m�q�6~�p�=i��j)�d�Q��>\����f��YM��hs�n���~$�i�4�����R��; <�P�'�8�����O@���z�vh�@��!�L�)��p�u Z�������k�blQ��N-�k�@�y���������@�v���O<�b�$�H��H��8YB�u�3F�zqζ1��h�x :@����i���,&��ۗ��b����_|���S���`�`7"���ˤ����d[�;�ò3���<��=�n;]D�v�'��ݶ�ω�ď%��t\>�I����Y���N���1�D��@<XoK�m��nӦ��O";6�B���1:���u���9�8��9W���~q�}m�a0vV�f(ۉ���vz��k��hm���#��A�!w:�o�$a#�����-䦁x�Z��f�s8�PӞ0lrM�j@Ÿָ� yv�g7��'1
4H�h�ՠz�vh�@����v��`� ��h_�v <� �u b���f#o#�8��rM ��h���O@�}��=V�4���.l$�Ĥ1L"k�asg�����k�H�s�l��l�ph�ћ��l�����x���o%4�j�=V�;�y������s�w�x�D�L��ۆ�x�[�fy�nfcg����-䦁o%7�����u��LM�B)�͸���?� � ^Ԁ=�pꤲH�F�#	���-䦁x�Z��f��ĹQ�EL-� ڐ�n����H���{����\��߶I7��\Y]��k�"�+ί�N��rm��V�)O�����!=���@�[^�ye4s��|���D��S��^���z��Hwj@Ÿ�:�3+p��8��q��S@�9)���<30�3�"�A�PZ���������U���߳3H�\��G�q$�9�䦁ye4U���S@�5iR"F�F�m�@yԀ}j��R�ڐ�v�~�:��:zض$�ո��u9:nZ���F{&�`�i�:�x�=he���_���@u ݩ yԀwRk�Ol�9�ye4s����=Vנqp\���"�&��;�R � ���Τ�tخ)�4HD7��h�k�/.�7'�"�b�ł$��g�y��g�m���Uk�'$"�0pݳsH֮@u ݩ WR���2��<.7�v(� ��8�h�
:������8���U��n^W��]��踙Yӟ$�i���~���䦁m��=Vנ�q�2�I��rS}UWd�!�~�'4�������|��s"n6�[e4W-zw31.���@峦��+ˍ�Cǐ����������3BURW$�h�Κۑ�ҍ9�k�h����}����Ɓ����u*I~���ffc�!m�É7m�E���臫��kS�+�dJ�9�];�^��%��sA��v�v̈́���u�5﷮��v�Cg8^�$�y��q=�������B�>kn����ܝu5�.[2��W-��-�6ؼ��u��d��t\�9۞7PF�uf��n����&y�h�.�����AK�vl�Q�m�`�W�m�:�����rWl��[ՙ;�0�^�w{��V��KѲD�դ���zrH�b�s�^vE��o'�c�r�=��_��E'�E�ȸ���h�M���_XI�/@�,��y�+�Y�e��o��]��I�NIz{�f��<�"�W�r(�L$Q8h+޽�7zD�*��y9��"��מɟ��5�.jˬ��lA�ll_�������y~����A�A�A�A����6 �66* ��s߿f�A��������Y��I�2�f�6 �666?{��6 �666
�~���A�A�A�A�{��؃� � � � �����y��~�Lɐ��k0�jK]�ī���Q�myw;tm�J�����0�����{�w���j&�jf�\�ff��A�����o�؃� � � � ����6 �666?�����lll}�o�؃� � � � ����e�fjj�5�֦�A��������Db?���#� �
�����¬h�E� � 
uڪr<���s}�y���6 �666?����@�A�A�A����ִIs.��Z֍�<�����k���A�A�A�A�����A� ,l{��M�<����~��b �`�`�`����_ڗZr���\֮�A��@�A����b �`�`�`��߷�lA�lll{���y�����؃� � � � �a��߳WSM��f�VfjlA�lll{��M�<�����A����{�����y{��6 �666?g�O���ػnڭ�����T������V��8y�1;�^�V9���x��.�4HsX�M�<�����W����{�����y{��6*�����~���A�A�A�A���L�.a��,��.�֍�<�����k���Q,ll}�o�؃� � � � �����y�����E�A�A�A��/��ѓ52�k���M�<��������y����b �b�,*� �Z(Q +�*� �Ҩ�;�����6 �666?{�b �`�`�X�*�2C|1e��39��0�IW¤66X �����y�����A�����o�؃� � �(`��{��A����~��e�fjj�5�֦�A�����~��A�A�A�_����b �`�`�`��{��A�����o�؃� � � � �޷���&���[2Mj���j�|���]��6��ϩ ��nK�I�#�"4�ww����ۻ��kD�2�,3Zѱ�A�A�A�A��~�v �666>���lA�lll{��M� r6"����7$���_ڗZr��.+�e��q�*�U+�I��?I5h�ؒT���h�Nb�2���0�4	&C@���O$�%�IUs��=��;��Ɓ���I# 9���4;IRUrI��$䗠6��IH@��[	$� �B���(�������nI������a��)|�-�Z|n�R��T��}����~4m��
g˅f0X���Lӆ6�n��/�4�����qnx�&�1x.
���L���ݞ'�H���P�/@�{:h�f��z�IR_XI2X_Yfb��g9�4�3e*UUWd�!�I2o��U%Wg�nK�9b���/3��fa�I2o���%WrL����t�=�jNH�j49��y�%rM��$�h��ꪤ��J������� �R���E<x���m��<���^�����x���ƀ��
q0'�%>�`��)+ ��%P�QM���E.zV3���E�D���}��	��kDQ��4T����j�A^R����.��Cr\��:�jI�A,���	�:zON����߿�       �  � ����6�$  m��!N+WOg���N�ƌnÆ�m�dE!��ݱ���ZtA�)--z� 
�ݩ6,�/cI+�����Af� 5Jtڮ�u� m��[Î�ûmJ��9üV�UW��gd9��T0��jڸ	`���fݪ���d�m�1k; R��fUZ�8{GS�Z�ʪ�b�Ud�v����9~'���*�^j	��e:ٮ;	V˵�!�jU�m�[B���K�z���CѪ\]����0 q䇷mlj�9�C���m5�K�5ێ�#��p��݈�δ�1�##^�з:9xq���#��8q��٧ql9l�=�8�g�m�M���8f���}����ֶ�m�h�EKә�nSzM	��Mԫ��c�ܷ �Zs\v�A�Ԉ��*��wb���dB��y��/8b�ک��v���5��f+��c�<�qٝ��msd&B�jSB�Ϧ���Qy:\rR�{-M��X9⺝���؅Ħ�MJ��ӳ��pԀ�ZڪL�ʋ�ظ\4�eUN7� �d��]�;�//}n�_Vy��q�j�e8�ۓ+ոv�#f��_e���8�m�It/�n��Vgk��f���<��v�XY�΢���[`Ъ:�q�u���ײ�l�l*�`��²5;f2ck���. &үS��v����R�p���jI9����_o�
��=��k��J�v���C�����Yn��Շk�;�Ӷ����7lۮ�=]���H6�3� t��֛Ny���<�ņ�V]�1�srpR�����d�����˝v�G��6�V�K��v�^=	�H�aE�@��u9S ���W�E�.��ȵ��5c��h���'�;n�a�f7l��q��s���l&�c9#F�Jܚ�Wt��νK�4�Z۶�j���]a,�]����s�9�Ռv����ƞ�m���C-�]�ݣ��RB:7S��|.���Dx/�C�
W�D��;Ϲ�kZ������]2u�;T��'s�W*uA��n+ON6,[6C�����mTeu�x�
3+cS���i������G�;K�5�üu�F�tOOGmAOYW<�l];s�EtE��	�kwt�ױ�g���l,��N��ݰn}u�5\ۑ�.a�o[1��4K���Z���������]�7��r��=	0�f��e�qO�P��!9��̽���𽵞x`�N��&M˻k}�7��G�������盋��1�!� �8���u��@}x�J�}`��h��a1�$d	�4[w7��f$v�K����6U*Wg[��/���Ç0�f->Iz[�i*��������q�1���hP�-Ҫ�&�@�d4��hJ�J��/@���2	�"$�#��h�S@NI���C@�x� n�j��[��Qے�f����]ʼQq���/;m۲��2(P(��fnn��1��H�RI@��uh��u�g�U^J�����@�3RrG��Q�H�h�S_�<�0�0xP�P�hA�P�$T�R�%�IR�R��Ɍ�;C@�ws{��$��r'<ȱ��$4��h�f��+�$ՠI2V�˯���,�r��/0Љ%rM��$���3C�U\����C��333�#0ŗ��4�ՠD��a�L��۔�>����a��A����m�>�X5ti�v��\��g��L�q2_�����F<Q85��=���[e4l���$������Z�9�8p/(3�/�4�3bUJ�d4	$ՠ6��<�<H�8��� ��$q��솀�z����*��D�$�d���?NΚ��kx��d$q�䆇��3����.{���{���@m�4?(�RT�&�}oLԜ��q �I�8�@T�&޳����Z}�gā���
Ý�k�&���M�i89,8�/]9��6
#�}�����}�+y.�y������:��*�}a$�h�\����$Hh�M�y��䚴	&C@�x͕Uv4�����f�����$���3H������}�D�i��x�pk&hwĕ�6�!�6�J�v�J�RR��*^T���Z��C9�E�s��y����hT�W�{����=�{V�m��>��K1��CmH��<Q��쯛N�5ѳ����F�H��/8:�/�c���8d�On6���gM�)�[e;�������W޷���d$�����7��s����O{<h��U��L�$P1�#�����@岚J��d4&C@:�ݶ���sZ���4%+rl4�C@�x��9��;�9Nɑ�	4�Hh�S@����?���u�f�w޷�����յҭ��k��h�nu�]t�D@,��͌C�7�/ ,;��%�Ղ�j�:r�"�C����t��G�������T�Jmq�1�׶��Z�p�q
x)��M�	g�<��i%�s;!�l�{qu�M��6P�ŻlW*�r��ձ��1�(wH[o�o����܇'��iS��X�P	�κu�7i3t5H$�4�F�� �{��}�>��?t�k.:q]�����V�&	��2�=����G�d�o��Ȩ��y�6f�$���ƈ��?��?��ye4[)�3���4[}i��ei���ni yԀr�@u �Mv��dm`����$�h����&C@�d4�w8�bd��4�m�C��{�4����ye4l���q��7�Ő�FG$4�3@�䪼�^����=�g���4xŖ���7�d�dq`�G��K�F��k�x�&����qr4\�����(菱�q��8zogM�)�^YN�$��L��4vN]�2�b�\\W�����k�]��*�U�fL��$�h����K�I$��U���1s0��y���@��x�x�%RUJ�9��$��@�r��$�"s&DG�����&�@�d4�3B$���6[���F<�p��[e4l����]H{��k&������.����q��C]̫��m����.�:��z5e��{ݚ�[�&6�<ؠ�=���[c4�2$���I��'Sɕ��e����.���ؕU�$�hL��m���y�G�_z�7�Ő�Ƥ��!�6�]*IeP�T��H��E HAB� c	��7UI|�$�~��d4��4�tg7����8_3-fg0Д�$�I��$���ЕJ�+�l4���˾e�Z���4�3@�T�%$�/��d4l�����ck�²!#��?����A.����q^p95�ti9/����1{���/K��b/0�[ՠ6���EJ���{��@��k��	2H�ɑL�x͊��%vG2�!�>��}K�?g�fy�e����ǐna4���@m�4��*��MZ�!��׋9e�s��y���J�I��$�V���hb�J�ꪕT�d���?5���&DLoq)�w4l��m��-���>�Y޼M)���6���"��E����t��`���qdni��}�ssw7�H�F�RG3�?~�?�S@m�%U}a$��ͨsy���#��2�fs���T��$�hI�@m�[�UKԩ.p���9̣0�\\W����{<h��H�*��MZ�!�uX�\\�9�3 ��BR��$�h�{��[e4l���kW�QL�s,��Š6ޭR�$�|�!�^[��?<�>��$�I$�dIJ��6:0e�P��m�0�u�}�<l��vѷeX�v�����uGE�[C�h�Ivۅ���sn+sݻ%���C��]l&W�8��1��n뗌�g�:��!dw���{Z�r�3���s�����v�;�<��=/6��.B��d�'�"����VN���Y�MWe���`쪅*��v��u�nH��.[��o�|4uS6�!�.�~�w�{��;{|����l�;�y�1��n��|�i�����H]�n�����|�?V^����ќ� ��o�>��R_XI3��v��d�<S�����-���*�M_������h̆��.7��1�iĤ4m��-�sO�x�{��@�{:h�ˋƒS�jH�hw̫�O��$�h�f���y*��~Z;��=NH�'"�$��[e4������MZm��?_��8.	��qR/`n����m=6���n�9]w<�-�}͠2�]M�q�$�<RC@��h�f��z�*��I���r`p��Q̺��]jnI�{^��8Dk����D�!B(@�"�E� �D���$H@� �XD" I�$!E �� Y�a!iD�I!"�#	�)ā!" �!H�	0�����*��~�ՠw�<h�f�I]�_d����Lx�N{��h�M?y����<o����~��~4��u���~(�E�9����h�f���hEUrI�hz*�F0S�����-����&��$�V���h?[���
	j[r#��)��f8�x�,]i�m�wf��=cM߾�_t_�茼���o�ِ�oV���J���$����1���7�Hh���)�[e4l������6r��ֵ�'�334{��@}x�5jԭRFWP��/����h�"��6�_��4
B��zt�U6px���GV�A�""���' q��8q_�}�^�A���
���đ~�5�t� ls{	��$�A�0���� 2	USPM��+�dc�#���M*9���!*i��Ha5�(��:+B2CZnI��Ad �@�!�,Bb�� �ؖ! ���b�� |� !���U<� x�� ` ����%T��J���^�~rf�~���3+//-qq^f�9��%�9���ye4b�����BR\o���π�d4׌�?[�2�k�ӻnH�2SnTD��푀z���l2^ݜ<�ͯ=��]8߾�o�&Xk\�?ͱ��6���z�}a.I�����M��G�@��h�S@����٠����#0#Ơ���h�|�+�93@�d4��Հ�Cxӂ�����޽���@m�4:�VURB@*T�R�y��>��&4��G#"r=�Z��l�|s!�;�|�=T�K��� ]K�M�Z�'��Pk�㛵�=Qʏ�on�['�"4NH��j9'�I�v�t�/:��H|� 8�.������ʽ� :��r �.@u ŕ[�'�ȈĤ4
��@���O�%��t�;�Κ3�K��Ƥ&LiG�|]v���gM�e4
��@�.q���Lx�8%�8�l��'f��%�9�;�_4:T��330p$-�k��I-Z�M��7P�<h��:�獮m��r�Z�ڻ;���&9�d-��^�'��k�[>z#qƞ�^�*͋;<g,Wo[mq�b��\m��@�S-k��0�k���E�wYּ'fC��շs*��l��n��Xs�s����v�	jq��m�)]��#�ՠZ�[����>���;=S�Ȇ�:�������w����t���ϗ�0�[o<�kS�����C�b��ć��T���f�����1�F`(5!@����4
��@���@��h�V�������h�|�Wd�'4	&C@}x��{�6���91�#���{נs��Ӿy�v�t�>��V��8Scq���X�#�9�Jh�S@��V�|�]�^�|opny#O)!�^<f�*_��|�'4������c��:��:M]�������s"�����������;]\g�Y^Z4ୠ|�3@w���w��EUK��C@�]�$�dD�ے\����<��*,*���9=���ܓ���@��V���1�c�1�,JG�w��h��J�W�$�[s�ޖ�,\�˻���UU%�͆�rK�߻��*��{��#�rXb�D@��4m��*�+�9�Jh�)��,Af64�$Xc���lå��%��7ŧ�ݻ ګ��(�Eė����ŋ�f�$��7@귯@�9)�_��|������}h��$� n+�77 ݩ |�@>]H}�O�<�#�^v��B1���$4󳦁��]��4�UJK3�����U���4�F4�Q�Hh�ʴ
�����3B*������.�ŗ�,�#2�v��9 �v�� ��n<�}V���((�& do�׎"-�lE�Z���3��gh�+b�rD��ӄ�Ŕ��$��~䦁~�����f~Ϙ~]���z/ߦLm�
4�R��h>uހ����א�'x\��B(�6҂��=��hrנs�Jh�S@��X��\$��D��*��{� :�.��g�ˀ}�9zԒ<��2H�}�M�ow��}�z�
�k�9ʰ��x�eM9��!�)��M�1�8��շ\9��V�4��+$KӲ�"3x�I��h�ʴ
�k��y��/,�\Y���i��i��/0�>|뽊�*�s��{��#��@}���<��e��Q~�I�H$��"�?.���}�M��h�ʴ/��bhSi8%�8�}�M��h�JhyR^\�O{�!~�,�-e��^r�.���4U*���>[s�w�' ~@��@l�H�{��m�6�ͶqΎ�'S�i�6�Y3`�s�v���3�H�:���:eum�r�j��ա��[����q��Ɍk��N��-l�0��v���'r�Pz�@9�6��.�Si���Tj�ӁNu��v�M��Tn��	{��3T��7>�!e�x۶�V��l���"v�sӶw#�x��<�o���h81�vcݮ\�kt��"뗀���{���ێ��e�:�]=�u ���y6�z7Kv��Hb.�@񃡹MG���OE7�D���� ��N�}�@;ݩ |�@Z��̲�G�7�r��x�ygM���{_*��x������$xq,dq�;�@:�����9 ���������Hhw<��wzhuޭ�z���UW��ϼhZ��yr��v�q_0�� 9����{� :����%��H�B�;���	b�����g8��3����v�}�WL�����s����nE��~z>䦁ye?��y�>a�Ͽ���z?ͦ
b�'�'�Ϲ��N����9׌�:�����6+��]����3F�JC@���{_��I+�nNh�!�?�-�uxe��&�!��}�z��޽�rSC��{�4��Xǋ;��5�N-�Z�*}{��d4�:�@�_����;��ջjKW8�N�X��:���q��/7`y�vV�1n?����m�]�����Τ� ���zڴF('"0rC@����>�4�޽�rS@�,���8I��Ԇ���3@w����	B�D��V�B��BJ��993�@�d4˧k�b��M�6䆇�]w�z�4�)�{y)�q}��&�b�'�7����hI����4m�h�m	�?$���L��u���857�m��u#�ٵ���2��G+�z3r��|���;N�+0o� ��Hj��ڐ�_4�P�%��AHh�Jo���6~]��������h�b��E�G�7�[����i��K���x�;9�^��2��G#��c#�C��b��@�d4���B�!	��Uqe�[��,���C�C�"���;�g������޽�rS@��q���l	уF�A�۪_-�T⛶;W��<�5�m�=\�c�x��LLs����;V���@���"�I}a���r@�$q&�nE�U�^���1"�Κo{��{_*�ٞbE�����1A�j�3���h���ʩ]��r�	nu�8.Y��
4�R廚���Z�;⼻�@���^(E.�3.��ڀ|�7 o� �Ԁ=�lܓ�40���U �]Qh��Q�AV)w�:��H(F$22�;Ic5�R@бĖU(�Mk���6*�,����YJ���{���N�{�zw{�v����       /Z  -� ��  �  �@��If��%�2�����ؒ�I���"5�vl5"^��2�c����I � fx������2��Ӯ`:��q�Q�]�TVU]L݁ݶ��2� 	k[��"�v�����FQ�B��&f��F�ٶ�eU���������::uT�ţm�vY{vؕV���7(�;�M�^�7���gf��A;EV��n�f�.6� �R�K�j��ۥ�Um:9I0����غ�R���!� �U�x�f�pn�bv1��o7���v޶I+^��O4�lv�p�m�v�[�QHnm���jm�9���Oizv/FӤZ+msL6�v��O.f�i���qx����c-�%�t�6�gh a9- �]�0�g��/2d���K��:Ƿh�m���t�Ȕ��ܝ�,�W�=�lCX��N֋d��akOmIٹ$�VQ�����x��懕a�P1)����	���=L�<�,S��[�Ȼ`�H8�1���Ggg{s�J[]KF�,�a��W����掺y%���Sz+k�ļ�(�Sꮺ��5r�2�T��=�۠��x��í��q���i-���O��p��޴s��n#����WmRT�uu�I��!.��#N��rgms��B�HW��N�hȚ3g���r����㎪��:7N�n��.볳=h��\v5����8;p�<��tٮ�GUñ4�KFsm�;:��^;m�fBw%@���k	>v�#���0����9�5�<�����\��US�n]�])�(܈'G���v�X4K�]��0�ܮ��.J�<ͩ D)��n�Th�q�]����+i{ ��֤A�8{Mn�n/l'<z�g��9�s� ��S�70�8j�pF�C�͎Sq1�tq52��V^Е{n�q�`ek��X�Z��ظ��Ľ��`���C��]Nڭ���M��Mp25�fKs^E�E�ߐ3J���z���vx<�>D"�B����
mݿsZֵ�k30ֶ�U��15����#l-&,P����	k���l��4��+���V�p<�$]�Xr�ͻgwn�Y���0�$�eM��3���W:��;m���g�nɶ��vyD��vt[j�RY��讗v� ���Q��<����3��i��ighw.��M��p��ZF�3�c6u��vw-nH��pD�O<�JJ�=�����|���lE�'LǛ/�꺌��y�N�:�cOn�2Q�������n9���H�̍��z�}�M��^UUT���}3Ɓإ��y�g �u����ڐ�T� ���rU�\��l���30������@���@>{R �.@;ݩ �ͭ^��\Il�f�q}۽4
�z�}�M�n��p|�ԙ#�'�$4.W �ԀyYP�e@=}t~;2����dq[�s��4W����<����=��Ew^�f�9���%^�z��8��m�?���r��<ʀu����W ���]�[z��J�K��vO�hw�z>䦁~b�^(E�6<��@>y� �W �Ԁr����\"�3#�4+k�9�%4[w4:��﹠}����P�	�cg4��3@��/��C@���|~�۝��Ba�u�����h`�5�E�6���ܮ棗�z�͝ĝrb�s�Y�hm��>}�h��?�����p#��h_�dn4��(�$���V�*I%v;rs@}y�oV���n���I�8��&ۋ@���@�9)�x�y�|v�hWj�*�8�M���	8]��g4"J�{�5h>7zm���%�1����(����n�)/�$��w$�����}������l&�fE���$q۱��X�裮�z��{i��B���sa�����w�;m�@�{��K�	$ՠIȋ4��"�3$p�*���x�m�4����=�S@���Q�F	51H������iW�$�\���>�5ww��k������J��~�_�䞾��r���1P�@@�g�����M�����#pc�I3@�Ÿj��� 
��mЗ����K\��|�=�����sG<��k�;A�����k��Y̬}��r�ڐYP�[�u��M�C�4��(��9�Jh۹��1/��ՠu^��>K�cMa1��J%�@YP�� o� ݩ |r:�D���"s4m��8�k�9�Jh��h���E�)2L� �.@;�R �ʀ|��~�}�>�� �[C�,�}6[�m� x�$�±�tm�eʯWm�`�q������g�ˡD�2]�]�6�y�[�J��s�$y��g�ۇ���:�m۝��!q���૮���8p��kn3.�����8��v���a�M�f�V_k�۱� =Z.��&��������GO]���ύj���s�a �Ӎ̗�V0�-I��ӊ��?��X�;�5�f����^�63�b����]�m۲S��v4F����S�ME��?���Jh�*�p�r y�o,͢��v�wt�<��8� o� ݩ �,9]Ȝ1E�I��ڴ
�kӞx�8� ��s@�9�Pm���.���wd�Ԁ<��+*��㩷�� ӂX��@�9)�^[��{m��*�@9ŕ��#��]�7nw[�]�㲼�pl�qgv�3gOmt�2m�i�	O#k	�Q)����˹�U�^�Ϲ)�_���x�I��'2�̩�U�Vawː�j@YS��T��'"�r�Ȍ��೙�@���{� ,�˩ ��RK�����-a��hD�RI+m�4�5h�)�qrנ|�\iL1c�I4�yYP�R�ː�Ԁ=���(�*��ɧk��{OJ�68�v�g�-j�y�x����$j�Ι�C� �u |� ��H�� �wR���Lj)�4�qr׽��<�1"�:h�{��{l��~gm��y��ڻ�����~m�ЪPUT	U%eX�R�#�䗠;rs@;��._k ���.�H�� �Ÿ_.@�+n��;ʣ�(EF6<���=]H_.@;�R �ʀZ]YS��	e9ٻe��X�,3g�F8�z{k݅������[n9pN�C�(�l�.@;�R �ʀ|���u[r��&E��=���H\�s@��V�W-z��˂�F%�8�I!�<�����\�/j@:�8챥"~L�*��@����Fhb�I"�B�$�����:����RcQLI)�W-z|�����O@��w4
�+�9�Q�p	 ��LEn��rkcFJ��s�Ţ�燝��vƮ͵�Y�8�y!28%�H�y)�^[��Uy^�W-z~\vcX�c0q)��� ye@��Y����9s����I%~��_�B&��c�s=�$��Y�$���RJۺ�J��s�P����H����W��}I+l�5$��群�V�=I%�8*�S� ��9=�$��pԒW�����U[�n�m�����m�bAE! V��{������!,���ph��	�
��*��Y�uMը4�Ț���N-��Me���2̋ugtkk���GYƙv�c<�7]Y]�����My�Z��v��Hopim����{^4gY�����ۋ��6�S��[�y�����֍+���!�����b�f��j�b��2��\�u�{1wQ�Mʖ��8]O��؎K��d���i{YǑ�eלuι�q�tp/VK�z nm4C�&
4`�ƲI0ԒW�����U[��$���{�I[f�$��8s,iDH��9���U[���cm%���}I.��pԒW�����_c�)qI�b�bI9�RI+�g����n�J��s�RJ�w�����7� ӂHRO}I+l�5$��群�V�=I$�-���E��kLf%��jI+�}�}I*��z�I^[=�$��pԒ_}�ۏ�	v����p�<��6����={=On���WR^]&6:3vY�L��Dc˛�}I*��z�I^[=�$��pԒW�����V��&1-A��I1�I%y}�s���	�Z����nڕ�群�V�=I%�8*�S�(E�O}I+l�5$��群�V�=I$�-���G8�pp�%���$�RI^[�{�IUn�ԒJ���%m�����0��\mL�,�s=�$��q�I(�U���߮�䙨ۻ�}o���wr�R��|���Ke��k�Xі4gj* @���4d^S���>{�:~�&|�7j���.I'1��I~����RJ�7I%yo�������w��������%N	!9=�$��pԒW�����U[��$���{�I�;1����F%&�J��s���_{fn� �'�i�0iT�H"@��l�HK�,�$B D����,T�
�� ���%!�,i����3+�l��	$06��Q�"ư�(A���"D��R @ � �-f�w(͑4P��e	HP��I�����ы"oc#M�5�`�=���AS}��H$I%*�B`�L�eiH�G7�$&�rH��,��L%%�X�P\n��jMf8�"A�+
0jB�@����*J��Ah��YV2E32�`e��0D������ |��TʚG�q@y��o��9m����7RJ�Ů���Q���{�K�y��w�Z�Iv���RK���RI^[�{�IZ��ĵR&8�ũ$���RK���RI^[�{�Ir���$��Ae���K��s�V�,��!q���o(ӫ�b��p<�Z�@ ����'$0P�����\�n�J��s�RK��ũ$���RH�P�8,X�ƲI0ԒW�����<�m���ũ$�o{=�$�l�5$�1�̸ڙ"X?�{�Ir���$���{�IrٸjI+�}�}I/��2�RajcĜũ$���RK���RI^[�{�J�#�Hc�@̗�Z�J�%jm�q,SB�{�IrٸjI+�}�}I.Ww��W��}I/�÷�2;� �2lj�f�w��H)�n9���<�9:yy�Wf國\.v̓��I%yo��%���ԒJ���%�f�%~�R�!��1��h�����@o�V��ޭ��*�#�ō��'�7&ho{4yw4�w4yw4yʙ�bds�2,�ɠ/2�,��* <� ��GE���Y$��^[��[˹��{[�{�{f�>:� ��>1, �(`�V�P��5�kZֳ3h�U���s�n�@� \�0��mN�7h6w�ܙ#'An�u�;7j�5��"G(�^lm�:�p;�c���x�76_��u�������ry�.���.�gRV�2��7l�6#G]˷ uӀ��wQ�+��m�N7R��l�rwni;m�njq� �`x8^�!�H]��x�[z�}��[c�INv�E֬4����_�{����|���%8�mm�4tv�b�L�a���w<��s1; ��$�l�sYv�Q�����V�>��}z�R�_ ��w4e��	���ncBs4���* �ʀ/2����3"�b����@��s@��sN����ho{4�v`�1��SMɠ<��̨ �� ^v ����!��1��9�����[4�Y�}m��|�׉�� (�$�Do:�3�S��5w ;�K�&:�N�*74��.1�(ț��7&h9l�yf���s�z�����>��Ǯb�pęH�$������i	
�@#`A

��!�
L��T(T�BP �&��lܓ���7 ^[4s�@�c`�A$�岠̨ �� ^v߬������2�9W�š*�Ur9���� o�h��hg8�B����ncBs4���"�π�MZ}z���w������闍.�m�nJ[��~^��v>�wn���&,��̃6���U������Ty� ]�y�ܳ9�1�ܚ����]� �-�o,�/�Q�1E�yѹ'���nI>������V�$+���s@��q1���M�an� �]���<���*�ʙ�bbpęH��yf��3�w��=����r٠s�q0�"I�9��:��8�Œ�N�ؼ��[x9^kY�� ��\Y18E�$I�}m��-�ڀ˰y�U_��okv�2��ڀ/2�r� ^v�e@=�9+I�ȚjcBs4��h�� �̨�Ļ��/h��n��� ���ʀ/2�}��U_�W�K!D^��	Q�L"���a����h���0�� j'+.�7`,��* <� ��߽���o���9ˡ�N��[�
�s����v�f��<��l��N�׶-WM^-��������T yv /; ye@�\Li%"nܙ��� ���YP�T��볹��ʼ/(/
����`���;�Ҡ{��w��q85�$I�^[��[˹��� ��h�_��)�,O��y� ]���YP
�߂�O{����� $-���5�ۓŶՒt;Cx���uFt<n����v� v&�ɍ��,�e�!pj��D��DMnW�M]��GQeރ�����3�-�۶n�(
tl�K�n�qf�K������ۯ%]��nh�m�ǥn%B�וu�\���s̕�u��}�<�����<��kvͻGBP!���b:�x�1�Y�ti�����\��t�j��ܬ����]'EK��Lp�X��&ud��q��7H"bSI���jcBs= �[4y��* �ʀw���t��3M�/w`��Ty� �h^
Y�$�D�4��@��s@^e@�`��n9���M.�/�/��"UI*��hrf�7�4���mˉ�	H��0Qɚܻ 9�`VTy� ����8�~�GVݨ�l�ܕ��Ũ8��T��n�N<y���t�8la�������`VTy� ;�`ԫZp��hq rM�n���s33.k* w.��`U~3�����9�@o�V���|�+�G3@�s@�8rV,����Ƅ�h\���+*�k��~��̻�/h��n��r /; �̨.Z��g��;՚ٝ�'�I7�rND������k�k[H<�#o6�6�qZiے�a�]���Q9�&����s@��s@��� ��h�F�~,��I�8'3@^e@�� ��� ��)���I���U�^�[�4���>�$`6"���=<X�]���r�h�lNd��@�W�39��Wr9�rj��ՠ;�@�8d��I6$�@�廚�* �.@�`u��eM���D\�-�F�J��9�ǎM Г�mi��w����B`L��<���f�o.�o� ��T��je�홻�|�\���@w����%v9�rj�-����g�q����0nbR= ��� �ʀ/2������8әnM��h���_{ٹ4���+[k *���r��U�ŒI�i�Hh����� 着<�@>z����	�ݫ�e���m��T�QĒ��+Gmc۰��kyG��mI6�-��ѱ�$�o�߹ 9�`:�y� �����mf��W�w��� 着<�@9�T�Z��Ԝ$lbN$I�^YH<ʀ7ː�v�W^[���7K�?^�y� o� <��)�}�92�n%$m51�Nf�W-z�ך��h}z�
J�ʥ�ROC��p�I�6���"��v���;��B�#C�|}&�Co�D�tj%C4���-	J��^�%s@L"P,H���ϥ !���7�n�4��� ���>x3�X�"�#6� �_��@6�^��<_Y�ܮ�!�Q�w�K�q����g�H�@ �4�R�`]���"���h�2����;���       -�� �  �M�  �  �  �8�=�Ǟ��ZW��Xbg���+ۙ:򮡩+Xॕ�R�9%��A���Zv�`��8���ӡ�n*�X@y�4� �,�B�:,���d���g�n=@6�B�TF��m��V���n�nuI��l�e%��T�1��u�JBP�9���efь^Ӑ�3/]@�&�w���GK[�U��2��I8�ԚÚ�Ym�7l{.�P��1��` ��R�9�+3c�Z��y'ŞK8ӻv��o-�%�y���k�;mK��{^��&��u�S�Q��.1ї'cCdf"v�ar(�QhJ�u�l�C��ab�h�k+��Azs�a6÷�7=4 ��N%�js�wY�cq��Z�<�R��W�z5͓CÍ��Q���v�=������=�"�<7\�Y��^��-d��)�vX�W���ҹ�lgg�OWB��rncI4���]�[�*.e�$�zt�� ��=T�дj�stK`�έ#��ay��f��b[zI�V8�nF�J��\�ɼ��\�%�خ�n��I�v���en�>��:�Z��;Fe�}�m�ay׸ˠ��g���Fl���N9�A��]�ص˦��H��	[�{l�!6mv�'�=����[G ��P u��V�8����ٺ.(�#�79QF�Y��ꃢ؉��ZX��Kn;7X�m�V&^1P��g18z�N�9؁ڧ�`{�<Z�Λ[Tֺ�Yg�������rjzr�mV���{I!$�sDd�4�T���JD�\E
��H�jT�l<:��c�:u�|�wD�`�EQ������\�v��XCG�vws�ѻz3��W8L[ngA�Mٺ�
F�t �Z�CL��=W��u�kd	j���f�DLU�z�^�㱒Ȑ��g&���ݚ'��Xbx�u�.�
��i���{����㪇0U�S�/����  �"	U�� ⡱;�ߞ���w��� 8յëb��TQ���sg�EC�ә6��9�\і-�Z�T�[�S�0;(�6'���Ч9zL�F�b=�z Ѻ뎎��,"��G�Q�!ۺ`"���h�U�֮\㲻��n9w6���q�!�p��يUj�M�!cq��;lٷm,U��`YC�ݯ/c]s&l�Û�{������xx\�gm�[R����P���;��{������֬eذV�By�M`��[y0�".�xyч�/4�rD����JFĤ~�_����9yw;�����9h���9� �Q�ܚ��9�T�\���n9���M�����H<ʀ7ː�v ��h�Q&4��)�7&hrנ��Ty� �����mf��g/�fs@>m�*�U(��|nj���h*T�w-K�-+/�9�.F�koK9{��u���67�z��t@��,C�&F�$lbN$5$���s@�9w4
�k�y�����.�wy�Kf��>��l�(�M� ̞��f�זh��h,��	�`��|� >W`,�w2�~�u	��Pi�,JG��h��h�s@�����'RP# q���v �ʀ}�ʀ7ː��`����Qm�cKt�s�6����n��٣]��ً�'vt�����g��uh�b��@��z�}o��z�%I}a�����4��(�B�L�*�@>�v �ʀ}�ʀ}�sov��wBԍ2H��r����3�Ϗ3��1@h'U�(��s9훒v����=ﯛ�6Ić$�����]�﹠|�Ҡ�� ���UZ�Y�[��eѹ� ��� o� ���YSm���s�2Qғm<]��agFz���6�qZ�E݋/W'q���ȓ>\W+%F�ͨ|� >�v �ʀ}�ʀq}�u&��Q���$��y�7���+�95h�j���h��/��3L�3r�3/w`,��e@��~��|uOHD�Ɯ��_��h��4���ԒiP�R�UIVdv_s@�}i��H��D7&hr� }��YP�ʀ}�.�h׷$�9��⃪ۂ5�6�I���瑦�����k�P��d���a%���I��ڐ�T�2����jf��Qww�w���� }̨|� �rS@�#-wy1Ɠ��h�e@y��Ԁ/j@:�;���	��9�W���������g����4�2���m� �Ĝz��f�)G'��?G5h��4}��UR�ԫp]v� tm��n׶u�W��l7'!�91�th:��� 8wm�]j�R�J���iJ�v���B��j,Y�K�:S�{ug���Z9�n��I����϶yx#�*��;�(�NE6�x�vN8���E��Wg;0�����&�ѣa��@t�Zw;Ӧ֞�m�5iи,�׍ƫ��Wb��ü�j�ac �n�M���N�\&#�����x>;w���n͝ȡh��Α��Sd���\��<�c�����	18�7&F�F��$>��v�<ʀ7ː�j@���o��n��3Kͨ�e@���Ԁ^[����3�ď�{����BF�nL�?�����Ԁ<���� ����1�	)"d���Jh��h�]��Z�ysH9�1'�Hh,��2���C�Y���V~��Fm9ı,O����2~�Z�挳m"Nk��$h�+�v�(v�Wv��2;d�WD��M���i��7���{����~��Kı=���Mı,K���M�"X�%��_l���%�by�����J�\n�����{��7��}���0�:	EB �>�A�9���ߦӑ,K�｛"n%�bX�����Kı>ό�[����֥�L�����Kı>����r%�bX���dMı,K���6��bX�'�Zߙ���1b<ϯvdm��n55�M�"X�%��{6D�Kı9��iȖ%�b{/����bX�'��~�ND�,K���<i��5m��534D�Kı9��iȖ%�b{/����bX�'��~�ND�,Kֽ����G��1b�Y���q�J6�yy��E�/j��K���<%ؓq�
�kT�b+<�Ve�F��w�{��7���̾�bn%�bX�w��m9ı,O{ٲ&�X�%��}�ND�,K����6j�T:��}����ow��o�iȖ%�b{�͑7ı,N{�p�r%�bX���f&�X�%��˞�p�DƜJI!�g���1b<��fț�bX�'=��m9������{�^" 
�@ GoTJ}�̿�f&�X�%��}��iȖ%�b����j�ֳ0��Z"n%�bX����ӑ,K��_{17ı,Ow��m9ı,O{ٲ&�X��������NY�A�0�{���oq��_{17ı,O���m9ı,O{ٲ&�X�%��}�m9ĳ�n��w����	�m˦_�n���2��4�'��{m��	�;C������}��?ʫu�L�����Kı?{��iȖ%�b{�͑7ı,N���ӑ,K��_{17ı,O{�w���Y$�W5�5�M�"X�%��{6D� �J�D��ߴ��H'�~�BE$Nsﴛ��%�b_O���M5��nd���"n%�bX��ͧ"X�%���bn%�bX����Kı=�=����G��1g��֞F�R%s[ND�,�"~���17ı,O����iȖ%�b{�͑7İ<�"}���iȖ%�bw����	֚����{��Y����}���Kı=�fț�bX�'{�p�r%�bX���f&�X�%�{�Gcs��ۢ��*�hn�]sbͱ��Q/���vN��Ǝ{$F�������h!A��Y���Kı?~��"n%�bX���iȖ%�b{/����L�bX�}�߮ӑ,Kž����eѭ\��]h���%�bw���"X�%���bn%�bX����Kĥ&�5���\�\)YI�vrf��˷F[.h�r%�bX�������bX�'���6��bX�'���q,K����"X�%��|fz�ˬ˙��R��bn%�bX�w���r%�bX���dMı,K���m9ı,Oe��q,K��}w���Y2ܺ��ɭjm9ı,O{ٲ&�X�%����6��bX�'��ى��%�bw�ߦӑ,K��g��kZֳ1���V����l�<���0Tt85[�`�"�T�n���K^�ڍv:J퓪� {=gÒ��.(���ۍ�	4�_3�a�n�m�р:�9�LͿ�?g�v���,l�\���ڃ��uuk�gm�/��x���h�Ȼ�b=�gd�\�pzṌ�6�t�*1�c�x�V�fPt�f�)�v�8�-���Z���ͭ��ѣ-Պ
&� �DP̛�mِ:�r8$I�P�i�ۀݖ:z[/,Y����m�fJ����V�\Yn���x�,K����"X�%���bn%�bX����ؙı?~������G��1e�{�l�	��4܆ӑ,K��_{17ı,N����r%�bX���dMı,K����=ߓ�g��u�������tؽ)j��Kı;�o�iȖ%�b{�͑7ı,N����Kı=��_w��oq��������a"$@l4�iȖ%�b{�͑7ı,N����Kı=���Mı,K���6��bX��~�̖eѬ�kE���q,K��}�ND�,K�}���Kı;�o�iȖ%�b{�͑7ı,O}�'��պ�!55��#9mɎ3�
훞Mx�{c`ub3H�����Սv��l��w�����oq�߉���7ı,N����r%�bX���dMı,K���m9ı,O��g��[���.je-�f&�X�%���~�NCțAXYD	T�#�1�7��{6D�Kı;����Kı=���Mı,K�U�dQ(Ɛ��d��3��G��1g���q,K��}�ND�,K�}���Kı;�o�iȖ%�b_O���kSV��u34D�K��"}���6��bX�'쿿f&�X�%���~�ND�,K��l���"<�y��[#�$������=<�y�%�����Kı;�o�iȖ%�b{�͑7ı,N����Kı?��ԥ�JkXCD՚̰��N�=q�h��vcc�Z�/i$�L�9�Sv��uLu:�kT�Z�SZ�br%�bX�}��ӑ,K����"n%�bX���iȖ%�b{/����bX�'{�~�.���̳5.kY���Kı=�fț�bX�'{�p�r%�bX���\Mı,K���6��bX����l�d�kZ�).�D�Kı;�{�ӑ,K���z�n%�C�}�0�1p��C
$�r7d����R% TB�a	��p���)HP�D%$�bT�e%G��
�gk��\v�����OQ��R�K��#!!K:��!Y"X�$Xie%l	�VI5�����uf�*[Z\%���+(ҕ!IdXHЕ�XBV���H2�\u!2�#)�^ W �lP^ !�
�>At��]�F*���"���;"f���ӑ,K���fț�oq���y�?�V�@5��{��ŉbX���f&�X�%���~�ND�,K��l���%�bw���#���ow�?��"�,f�����x�,K�׽v��bX�'���q,K��}�ND�,K�}���qb<�y�խ��bqL�(%��6KE��\���W�V�C���F�L]�!R���ɖ��]e��]�"X�%��{6D�Kı;�{�ӑ,K��_{0?�2%�b}��~�ND�,K��������nd���"n%�bX���i�~c�2%��/�ى��%�b}��~�ND�,K��l���%�b}߷�20$������=<�y���V��Mı,K�׽v��bX�'���q,K��}�ND�,K�Oc����ؠ�K��{��7�n�{�����v��bX�'�߳dMı,K���m9İ1v�"���?�K���bn%�bX���~�.����&j\�֮ӑ,K����"n%�bX~#�߹�m;ı,O�~�Mı,K�׽v��bX�'��M�Y�u!�����˒��,�§Fg����3֞#ήt#�+ukfh����OwȖ%�bw�ߦӑ,K��_{17ı,N�^��r%�bX���dM�1b<�y��N:�prD��bN�{ı,Oe��p���r&D�>�_�]�"X�%�����q,K��}�M�"~EAʙ����~�̶�3E�L�����Kı>���M�"X�%��{6D�Kı;�o�iȖ%�b{/����bX�'�5�h�V�&��kV�f����Kı=�fț�bX�'{��m9ı,Oe��q,K��}�M�"X�%�}�x��˫nd���"n%�bX���iȖ%�a���_߳�,K�����6��bX�'���q,K�؁�f��� �����If��M�4��Td,�u�S`;j�妍Pq4�a�z�U�"�6�e�n4��׷;�Ȃ�ڔ�,ɐ�q��&��ن�H�úޝ᧝��n�b�{3*0�v�FcDn��6�+�ls�jL8��p�P�Eq��ϱK���}��Z���zM���ܜ�&�J�B��m�k+�[x@��ܝ,�0�EC�R޼�Zݐ=�w������9���u��K��۳ۚrp�sՈi'n!��i��w8{h���h�8�]����=�{�K�~�Mı,K���6��bX�'���q,K��}�ND�.���M���S٠�K��{��"X����Kı=�J��bX�'{�p�r%�bX���f&�X���_���)��p�3��G��X��ץMı,K���m9ı,Oe��q,K��}�M�"X�{�������!Q��ǻ��7��bw���"X�%���bn%�bX�����Kı=�J��bX�'��z�3S5�[s4d�Z6��bX�'��ى��%�bw�{�ӑ,K����*n%�bX���iȖ%��{�����/kV2�1��T�ƍ����4g���o]#�v��V�D�G"�١LL�52��q,K��~��"X�%��]zT�Kı9��a�"(��Ȗ%��/�ى��%�b~�kߴR	Ա-���w�{��7������Ǎ�
y^b&�j%����ND�,K�}���Kı=߽�iȖ%�b_C�.C5&j[�.�֥Mı,K���6��bX�'��ى��%�b{�{�ӑ,K����*n%�O1gܷ��!"�NL�3��G��X���f&�X�%����ND�,K޺����%�b{�{�ӑ,K�����?>��Y;�}�oq��K���6��bX�'�u�Sq,K��~��"X�%���bn%�g��w�����螶�W�ήT,I��r����!�O�=`V�@����D;�m��ɚ�5�Ѵ�Kı=�J��bX�'���m9ı,Oe��q,K��~��"X�%��}�K��Yn��h�ֵ*n%�bX�����? ș�������Kı?}��6��bX�'�u�Sq?&TȖ'������B5��w�����oq�ߩ����X�%����ND����d HFB���dND��]�7ı,N{߸m9ı,O�����.�h��}����������߻fӑ,K��������%�b{�{�ӑ,K��_{17Ļ�ow��k��؉V%�}��oq�X�'�u�Sq,K��~��"X�%���bn%�bX���6��g���{�����Ǿ�0㱢�Zl�nq���Y��]�v����rOn:3vY���;�52�K�u�Sq,K��~��"X�%���bn%�bX���6��bX�'�u�Sq,K���\֮kRMkZ�L�h�r%�bX���f&�(��R���Y��)YJ�VR��F�X�%����ND�.TȖ'�/���e��Aj�����oq�߿���Y��Kı=�J��c�"~�߸m9ı,O�~�Mı,K����n,I(�)��3��G���a�D�������%�b~�߸m9ı,Oe��q,Kʁ��P �C� %SI7>��ND�,K�a�<f���Z��MkR��X�%����"X�%���bn%�bX���m9ı,O{ٲ&�X�%����s��ͱ�oWC�]�ٻF�Ҙg���+��K���n���"��,��n��Z8��bX�'쿿f&�X�%���ߦӑ,K����"n%�bX���iȖ%�b}3�=5�e��355Ku���Kı;�zp�r%�bX���dMı,K���m9ı,r�k~f�b<�y��9�8�F�M��S0��Ѵ�Kı=�fț�bX�';�p�r%��C"dO�~�Mı,K�~�6��bX�%�>��1�52�K���&�X�%����6��bX�'��ى��%�bw����K���ȟ��8D�Kı;���kZ�a�I5�k5��Ѵ�Kı=��f&�X�%��#�߿N�Nı,K��fț�bX�';�p�r%�bX�|��ݷ������Ŗ�'ln��U�m���--�i	�*c�}�}R��8�KP�wSFR֬�<�RA��Հ���5���%�3��`�#WSZ&��Pkf;m�ohgI�KeQ�HnM��t�ez�;��ˬe�^������חm�k<����ewPGS���mC���u�.ݺ���mM�N���Q�X��(v��OK��r6L.�����w�~�_7.y'��[]�c�;�7\kE�Ś����\��g�w`l�u�l斻,��T��ı,K�~�8m9ı,O}��q,K��}��'bdK�:��~f�b<�y��+�CME�J"Z�MND�,K�{6D�?�"dK�~��iȖ%�b~��ى��%�bw����İ~�>-�5�.��aKu�&�X�%����6��bX�'�����Kı/{�Mm9ı,O}��q,K����잳R�r�d�Z6��bX�'�����Kı/{�Mm9ı,O}��q,K��}�ND�,K��L��a�WD���-ֳq,K��}�{[ND�,K�{6D�Kı;�{�ӑ,K��_����bX�'3����Z�6�.��B�M���6�����=�{5��,;��$V��HV%�k�w�%�bX��ٲ&�X�%����6��bX�'�����Kı=�}��ӑ,Kľ��ڙ�h���2]e�7ı,N����"H�ș������Kı=��=��"X�%�｛"n'�ʙ������4kF��kZ��h�r%�bX���oq,K��}�{[ND�,K�{6D�Kı;�{�ӑ,K���=7��Iu�a.�u��bn%�bX�Ͼ�kiȖ%�b{�fț�bX�'{�p�r%�`~T&D�=����bX�'����5fj۬��Mk5��"X�%�｛"n%�bX���iȖ%�bz}��n%�bX�ϯ��ӑ,K���fOA�]�at="�Z9�w]10��Qls'��j9�1������0tFi�O<pWov�X�%��}�ND�,K��oq,K��}~��B�H���u�N���}fK��˚5�]hؒ	"}>���z%�b{=~����bX�'���q,K���{�ӑ,K���:F��,$����G��1e�_���"X�%��{6D�K�q���j'��m9ı,N���'��oq����������`Z�9ı,O{ٲ&�X�%����6��bX�'�{�q,K�ȟ��g�m9ı,K���3ԙ�nYu34D�Kı;�{�ӑ,K����_�\ND�,K�{��[ND�,K��l���%�b_v�찙sZ�]=��a܉�ӵƢ���ȯ�1�b�r�$:��O5r��VB�V��w�{��7��=뉸�%�b{>�=��"X�%��{6D�Kı;�{�ӑ,K=������LT�(-2����{��'����r%�bX��ٲ&�X�%����6��bX�'�����O�y���^EN�C�K#j$ro���bX�'�~͑7ı,N����Kı=��f&�X�%��������bX�����fMf���Z"n%�bX���iȖ%�b{/��Mı,K����m9İ?Q(�j'�~Α7ı,O����W0�ֳ.h�Ku�iȖ%�b{/��Mı,K����m9ı,O}��q,K��}�ND�,K��_C3XɗV�ӵ4�UvAzx2�aq���m����pY�g5�-�K�e�p2����{��2{>�=��"X�%�｛"n%�bX���a�Rv&D�,O�}�17Ǎ�7�������F[K�����,K�{6D�Kı;��iȖ%�bzg޸��bX�'��g���Kı/�>���5&jۖ]L�7ı,N��p�r%�bX����q,K��{�����bX�'��l���%�bt��0��jL�֮e�h�r%�bX����q,K��{�����bX�'��l���%�bw���'���{���7�義0�٠����x�,K����m9ı,O}��q,K��}�ND�,K�~�bn%�bX���]�4 d���"D���
�\�3@<5�)�#��:&a�pvl*�Ҝ&���`?1�8 �S�vҐ���\! ��C������1V3M�@�|,��!�"��o��$I�1����wAB
� �X
AH0`�b�/n �� ��"��E�l��cdSH}� 	xg����o�`��W�G�W"��1��R��[����	)]i	"���2����c�F�2���H0v�z��'e%e�j�g^���ڵ��B/#`���]��$C���wâ\5�_�"'�����f��9"����E�e�&����%6J&��BR^ˌ3�G�!��� �SB�
�XS���Ya�S�]3����`sV^�Sr��[F���+bAA����`E(��H�"E�	D�5��4�r���zM�׿;�����       [%  h � ��  m�  �����N<ì`3V�Xb�l=��v8�r�iI��,[T�$�8)�+�l��t�\�EZ�Ύ�8QUۤ�R���5�� jUU�A��͖Y6�M�njA�9ŞB�=W`��CS����tJ��U ��������r���f�`{N�[B��컧Ps��}�*�I�m�^w�<eɵ�iV�W��[pu�!��[a��T���U��ɪI�ی��k��q��vAi�����\P��lȾg��k(s\������n�����3iD��/`9u[��6�Q�m�S��#��f�k�(Cq.�97k�\��9��C��.���;-g�^9V*ð0,��m�6��sl��*r�"KoJ�r8t����+w8���u�jm���IϷns���X��n/U�/;%��j��9��.�+ъ��4-�06����s�ʯS��/e�U��˸^�j�2�t�Ye�^�Ni�V%)�]�Q	��5׭!-T�y�=}�|�s4�=J��������[dM�·$\�s���k��
�Ɠz%���v�q�a���%#���n; IǷF�鷬�Ly��5y�hΰq�x6�q�6+e��ܬ��1Y���v
�:�EPKٍ��a$�:9,��D����'u;h���X�s]<e�r�vz��7�qͦ�]�p9B�����fGQ�f�m��,=��ںW�T��l��݀�h�K:�8�苪��C{�Z�Im@��3�B��ؚ۠]�\m�m��}?;�]S�Nm�9C�c `b��*����Ԝ���z,qt�m&�+knz�6�Hc�R��q*'s�:Gj��|geg;������YV��C�l��"ŵ�D�;r�Z�����=��TR�E6Z�}y����&tn�z�oWj��nCu<���C&�SLY|��]Ku�V���X���)��_� ~4"<0����(t�w_kZ�R�PJ�W]��8xK6���Ȭ���I9]4�0�L�;߯��2�ӌZ�nf�HLWW<�{k��]��7]��ђ�'�k��.v�h�d6��c������գ-���8.lgۮ4���iћ�����ү.4 k#�i�W\�*�7Rk;r܎�w���z�%F�ٓ��[����&�.t�D덊�6���!��w�wx�ccl��eё)�r7
qqh�#mا��Du�p/�n�����Ғ:�̀�KS_{�w���%��߳dMı,K���m9ı,Oe�ى��%�b{>�=��"X�%�{i�|f�&�Z�
K�7ı,N����Kı=��f&�X�%��������bX�'��l����_s���~sߟ��5�J5�+��7��bX����bn%�bX�Ͼ�kiȖ%�b{�fț�bX�'{�p�r!��������
�\]���K��x�,K����m9ı,O{�ԉ��%�bw���"X�%�����7=���ow����ߝ$+�����,K����H��bX�'{�p�r%�bX��{Yq,K��}�{[{�����oq�����S*��.6d^l�
�僃�G&�܃��/Cr5�$���U3!��շ,���H��bX�'{�p�r%�bX��{Yq,K��}�{[ND�,K���"n%�bX�;�s/u�%B�w�����oq�ߏ����#�	 b� J�ΡE@�MD�=��=��"X�%��{z�7ı,N����O�(eL��{�����U�9�4�ﷸ��x�?g�����Kı>��ԉ��%�bw���"X�%��kڱ7ı,O����3R�k3XY5�ֶ��bX�'�{z�7ı,N����Kı;�J��bX��?k����r%�bX�a�L�f�&�Z�
K��7ı,N����Kı;�J��bX�'����r%�bX�}��D�K<�y��/�XQz�X�	�CDm�� ;ub�lGc��8G��2e�Ͷs_N�I�K�ֵ���2ۭND�,K������%�b{��6��bX�'�{z�?"�L�bX�}���"X�%��k�W���l�ﷸ��{�����n�6����L�b{߷�q,K���߸m9ı,N��Ҧ�~Q=��������/�����w�%�bX����D�Kı;�{�ӑ,A:	���a�����Ҧ�X�%������r%�bX��O���ԙ�nYu3Z�7ı,N����Kı=3�\Mı,K�O���Kı=���q,K�����2�ѣY.��33Z6��bX�'�}뉸�%�a�>���m9ı,O{�ԉ��%�b}�{�ӑ,KĿ�����p�i5ў܍�#�8�Y|�c]�0Yy�l�W�Q�qf�[�ѳJRU�\Mı,K�O���Kı=�oR&�X�%��}�ND�,K�=뉸�%�bs�}O�5fe��f��SiȖ%�b{�ޤMı,K���6��bX�'�{�q,K�����m9ı,^��=�u���֌)njD�Kı>��iȖ%�bzg�q7ı,O}>ߦӑ,KĶ�3O1b<�y�c୎I$I�e�Z6��bX�'�{�q,K�����m9ı,O{�ԉ��%�D�U,O��t�r%�bX�{Y���0��8�����1b<�ÛM�"X�%��{z�7ı,O��p�r%�bX���\Mı,K�z��ہ۸l�mm�8��M�0��:n�S�r9�Ѭ��A$Y�^�x�p$�˩��Kı=�oR&�X�%��}�ND�,K�=뉸�%�b{���6��bX�%�'��̆jLշ,���H��bX�'���m9���,O�?~���bX�'�Oo��r%�bX����q,K�������5�Feֲ�fkFӑ,K���z�n%�bR���f���eJT��R�JI���q,K�~��iȖ%�bv{�浩�kY����֮�q7ı,O}>ߦӑ,K����H��bX�'���m9ı,OL��&�X�%��u~�5f�jf[u��Mf�ӑ,K����H��bX�'���m9ı,OL��&�X�%�����r%�bX�"�{z� p���ykGTI&ΐ:8���U�t�+���ڎ԰�9���Խ�����:��ӱ�[n�\���`�[Ǝ{9�o`��6�G��c{��@���V�5��۷k;e�ܢ��9#���* {j8�4[u�؞:#�a.	XhH)�ʸ��N�Τ�fe�7���Cՙ!�4C�Q�Iw[�H��YL,ȷM���k%ԙt[o�Ҩ4� z�޵��ע7�i���;(qqۃ�!�\�٢����n���9U��X�p�^�$�'�ı,O����"X�%�����Kı=��~�ND�,K���"n!�����s��ʪ�hg W}��o%�bzg�q7�DȖ'�Oo��r%�bX��~ޤMı,K���6���r�D�=�̿�fI�&��je%֮&�X�%�����6��bX�'���D�Kı>��iȖ%�bzg�q7ı,O�j�����%-�ff��jm9ı,O{�ԉ��%�b}�{�ӑ,K���z�n%�`~E*G
Q��m/�VR����&^p\�3Vܲ�.�"n%�bX�w���Kı=3޸��bX�'��o�iȖ%�b{�ޤMı,K�}})�-�δ�y�\Vv�{s�/�	Y�na#�q���K1����ܺ����sL*��{���D�,OL��&�X�%�����r%�bX����q,K�����"�oq������Eh�c,0����ı=��~�NC��Dr&D�=�oR&�X�%����"X�%��ڟ����1b<�yR�� �JLF�6��+��1ށ����UR�������4g�9H�Q��b�ȴ�ʀ=�p�Ԁ=�pU���b��M�&h�ՠw�3;jޞ���ՠ}���>�7q�dRqXU��5�ɳ:�'C�8�=��9��v��q�7�i��5l�a$ȰR-�S@�v����y��ޭ�/1���(ŉ8ۄNk�V����h�ՠ^qJh�R1�$�#�@��vnI�޻��FB3�Y �x�登g���|�@���P�2c���37j �-��Ԁ=�p?��U_w{�hs�͊H��F'#q8��)H�[�{�* �sp�u�~
�H]�������\k�xNd����u�W];R�@��H�%�F���\j}������?~oV��λ��/�#w��y�x�ddN8"�>����x���V��T�_��@�.%l�LR@P��{� {�u�@Ÿ�����U6�&L�"��fy���zh�K�?~oV�ԅH��*�*]Ig�����׽�h�ǝ��)�q���i {��ʀ=�p�� ������%cSOn]s��h���b��׎�Jv�y��\�	�ћ��l֜�s ��͸���b��Hط ���P�2c�A�ܙ�^>U�^qJh�j�>����$}��b�&䍤�N'��T�_��@��w4�ʴ��Y&A��LC��@�;V���z��uބJ�*W����.a��Ȝy1`�Z�[��^;V�y�=7$���]�8hP�	1t�t������@8յÖ������X7=��B�KJU�m(G&�>m��bSk��]�u��7n�`�t��ώ�[b܇����۫�����u���;���ln��ї��;���½+D�����*n��N�k1�676�:���6f	�)�;�cn)g�<�ю�m�W*u�Nv��0�.�;�7���}�]�~�.p6v���v�	T���ww������>\�+e�$�vv��`�#U���	<F�x]�z�sg}Ŵ!O���VšCv������z��n�,�_2�����ȰR-�S@�v����/�@��q�o��'��� b��YP���=ש (|�\��1ēB�qh}n�y���H�[�z��[06���ot��ݨ����Ԁ>Ÿ��4	�����Ls��0l�h�8�k�M�]Hވm�q��/�f�j:��QP�*ND�qz�L�s��-�rd�?��|�rDI���LC��@�;V�<|���7��s�7$�s�]�=��S@��\m�@��&,�@��w4���wu�@b�����spې"cRf�x�V��qJh�j�=������Sr@ncrdX'��r� �n��T���_���u�v����}�\S����l�m�U糸v�ͣ���#գK3p��`m����Ÿ�YP���wu�@=|��h��I�B8�~�s@�|�@�8��~v���%m &9�')&hO}�z�I��_l�採҉����9�8�/P���D7nU�j#����D'GdޗA̮J�R%X:އd0��$1!��U6���᳟Q�HT`�[�UX�ų���?|F@��~��h�tU����� ��Hܨb�H�7"�i��8I@
��kaӯ�� u'�?@)��1	�X���j��B�D��� O�	���u<*���UЩ�J�ׁ|(�6|��Ȉ�!��p S�4���5�k�'}��n��[�nH�ND�qh���/�n�ߛա�IU%q㗠~��g.�����Y�y��-�=� {9��������a0�����y"���oV�N,�`̜�-��n��ͥ���#�&,�@��w4�ʴs�S�y�y�;�ޭ�u�8��CdPjm@�n�ש }�p���ع�7#�7&E�qh���~v��˹�^>U�_���B��'O�a�?�n��^���w���T�@b�J��߯�M�'d��Rch��I�B8���s@�|�@�⻚�ڴ��Wz��Y"q%�b�ʎz6��W9�8�<%ڳŲ�JkQ7T�p�mb	�c#�Iɞ���V�y�w4�w3<�=A�w����lNA�#w|�_2�/@}�[)%J��;�/@�d��/*���y��gV8��1F��I{� ��������g7 {�R �����#��ȴ��s@�|�@���/�ՠsV����e������u�@b��YP�{�ߛ����Hk�u�Ü����^���*�oU�i *k˹��z�:��9H���\#,�ѵQ��v���Â�vtp���q�ܗ�m����m�ۗF��d�]�gGe{qlD��#�據�5����>������y����Mό�N�'	�;]�N[�X����$�(�\�g<.W:N؁��3��3�Cr�v'����܂�wBp-�'l��vLF���;��|v���l[;kV�M�B�N�t�nx����[��q�p>�M<���u��R�r�G$����?�ڴ��s@���@��;27�LX��'�4�h}n�W9^�y�)��3ă�[�ch��M
Šs���W9^�y�w4�hg9+kLsNL�*�+�=�ʀ>Ÿ���r����3wp����sr �[* ���ʀ^>U�qp@�*SƘF4��!�:��qwl��3��s�7B�b6�+Tu��{��Vn��@b��YP���^q]� ���na�D�,�@��{f� �$�)"ŀ���Uᙜ���Pط �_���1G�D�4�ʴ[^�~v��n��5�(�&72H�D)���J�=�pye@�n ��w#x�ŉ��pQ��/�ՠ}�����Z9��4��.�u.��b�����8t���cn<6;�rnzq�[��ѭZl�k�HLmD�hP�/@����x���rT�-�>�bх��ma���� {9�w9* ��ye@=�b��i��R-��h��]��͢��_����߻��r|�uh��eȇb�("H�h� ��* �sp��P����2ԍ0X9����h��^�@���h�j�/8��'X���D5$Vrm�8�+nƶ68nA����)�r�/$��hKm �H܈�)3@�|�@��{��ڴ~�s@��UƦ(� {�� }�p����9 �7Y%1bMF8(�h�j�=����r���h����MA6��sn��T�� s��?��~��"��u_Ȩ<߻��rO�gߦK&��dr(ԓ4
����W��_��@��w4��x���b���ț�����FwD��+���7nma�m��HW;�E.,�$$�#�4�Q2H����h�j�=������귯@�����%�DA��Pط ��T�� �J�߳�<��t�#q������Z��w �9 {�� }�p������9#�B�4
���y^�~v��˹�s���7#m�p�ФZ��ط ��T�[�5��EUV�N���=;��=���} m�:U���WM�ո',k�s6VwR��9���kgt�u�?�{���R�'�{Y#��ux�c�ӟm������q<��gPs��Ugi� ���T�
�<�ڦ�I�9l�v8�x�#.�Nݵ=���,�ղ����MM�m�j�U�X�\��u(tI�#�K�MK.؋r�ۍ�;"Tˊ�)c����RvH�ku��O�#���Ε�$����Xj@vx3�h�b��S���E�{4��]1"E�G�E�`�8�pQ̠}����=����h�� �s��҉�&ҽ76�<ʀ=�p�%@Ÿ���B	�c#�G��^;V�o� {�ye@>�n�n���������rT�[�}� o�4x���'�,"H�h�ՠ{�* �-�;��P���r�ͬ��!_N�D���M�����pE�v��+�v�pQ5���Ʋ7���Z�[��^Ÿw9* �-�:���:fћ��֤ԷZ7$���]�h@c� 
U:���>�ՠG�/@���h�;��܍��cB�hs��h�ՠ}yw4�j�/�Q�bɍ	�ӂ�� {�y� {��rT @�����M��Z�.�x�P<�ط ����0��@m�z�K�N��ns�x�,�9:�7m�5�1n�Qd�A1̑�ۊI��h^\� {�s*�-ͼ�r�p�v�o6�y�P�n �2�b��cY`�Ȑ�AG3@�v���էꪤ��T��D�39%�9�Z�Yr�n5���"�=����ڴ�W��^;V��_V�c�I"����@Ÿ��ط ��+@�y�yyխ��d1H
46�dbvq�5�"��=g���@]���p-�afxd�jW�cB�zm���/�@��w4�j�9�Q�bɏĜBb�f�x��ye@Ÿ�� ��M��6҄qh}n�x�Z9�w4�j�>���1c����䙠>��;��ՠ>��Ǵ�RM]���1b��hQLH*��+{���h��bp�x�&8�Z9�w4�n��T�[�w��+6�Č���B�gq8�˫=lޔ�J�z�+�8��d�mcP�� �"E&h�ՠ}� {��l��L���p��x�E�{����;_z�o^�x�Z1}[u�a$�HJL�/���� {��ʀwv巹�n�ƅ"�ff+o_��s��Z�[��s�ՠ_��,�L~$�s4��h�3��~π�_H�}ǹ�'���P�EPh��*�슠*�UW��T_�P�EP���� �Ab("�0 "( EX* �"(X� �@��
�0B"�0 ��R"�1X* �X� �B"�1 "(
�0A"�0� �U"( Q`��#ET�"�
����
��*�*�EPj*���@U��UW��T_�P�U@U��UW�"�
�EP�1AY&SY��-�tـhP��3'� aj��_`�  Ƞ 4      h @  v�   ކB�$
�H� �@*��   �R�P �P�  �   RB�(AH�)J��  �
A@)@ l�@ �@ft �R�w0 �� ��馌@�M,�Gon w���#���yoo  6����[k���� �����e��W6�vrw֫炅8u^��W�7K�N��  s h   ��P
H ���t(�y����5֯��ޏ������
p�ݏJ����޼]Uv��.�x װ�o�k���׀ v�瞃�����V-z��9����ܷZo|�'ϫ��:��N�ͧV���� �� �T� ���{�}��`�wjۋK�\�h_8 �������i��x����|� ��f·�����������>|� :�Dt�vb��f)��@��o�;����y7g�}�:�����( �A@� c0 ;�/�۰����g���Y�
w(�}o#��6�㻔��}}+�7�e^����/{/o�o����
`����}>��z�޽�՞#���O{�9�齷����ɻm����| ��( P%AJ (��Q�C�۴���yw�}���{��{������JD�bSJQ� :�A�(Ħ� 
b 
D4�0L��� "i�M;0 Sf 5 �� J()� PG`��   ORdm)R&@�T��1SmT�P  �z�Q�J� hت�mE)   D�	Lʔ� ��h�IJ")��?������tE����.L�̧�NڇN�/�%Tt�
�*�QEO��
��ET�PU���*���O�����a��g��ͤ���'ܼ�W䃣Q�3�rk�Ö��H����](D��X�Rk](<]f�%�(��j|a���xH�Y���GFs1��6ān�7R5�o\����	���ct�W+�Pv���V�Z�ϔ��J80B�嫅'I�JEt[��]9>��6K�a6d߶s��$It�3\�P��4��R���)� �I����f������Y�P4��ֵ����$��0H°�Z���RA�
D�_<�18�ц����5�#[��
$ 1J�pH]c.�V=���s��3���F1�f��%0�20����xpٴ�ͽ�g3���׌������@�wNz�<O/�PU���%|�Dב|UR�)����)��)�4�B�Ț]��E,�u_�npB�;/�PB�Ȍ�k�a��dXK��[�o���d���t�WWZ!V5���d	Hi��k����j8\tq kS.�u���4.�`:R)�FnǄvwxe��5�j����l���1�Y��3)&��ǻџ}{�{~b�a5�K@�.��B���Ѳt��Y$��M2���]%���7
GIF$"�!�p۩�Md�ܦ��EF �@� ؑ�R1[#HH�F0t���]@��HE4&��Ԑ��.��֜�jB�!�	i[.M:�&�0p%!��E$R��P-%�$��ߍ��M�ɭa��6��h�� �D,�bD�������`c���������)�1��#��O�q��˦�] B˽8	[�mq;�\�[�Pr��(���AN�R*��T+���B.�n�����$0�&�R�l����]нQPy�}�I�v���]n��Y|K�gH ��M��2i��P!lkwJ�%ծ�k�64/��V%(m!U���'�#����fs��N 	F���(KyI�6L�y��nc�.���,X0�VS;�54a��%0���Fl S�zH@oM��\���<��_g	{Ņ����E���:} I�Y%)�HG|>�	t��AI4�neb�"Բ��$�o�m#�]k���d�ﺑ�1�.��D�f�&h#�F���u�]1��sWl޵���c�&�I��$f��{���!�JU�R�5I)@�n����w���s�f�u	n�e�|g^���!�ưH1���������>>>,��i�M&i�#]+�
�XY	�)!I-%�j��,$�Ku�|O��fh�Ǒ���ª�O�:lO��	�Y���t�]�9�y$#Ͼ��(���}ބ�
In��\�!���XB[���滁
1!�f�˭�$w�	MK����i��$Ix�>��h�BA�]o�}�ʤE �ħ���~�K�]���kwG���ňD ��@b��D`�
$���������o�<��357���}��k5�����w�H@*i:B�@ :�#���)ll	�s$!�w��,̈́��!(�
�5#@�H1��04��SL���!R1�$#��F�ŉ�pX]f��l���d��͘p�5���7͚8�bK�o��X��������lk|�>7��ooxj_������ӡgHXP�	"E"ł�)$ �"-xm��g��������~9!Ņ,�B�P���ƚ6��3f�y���!t2����t�h, �B.��$V(E(B�����$�S���6YC8i!�6a#���d���͵#�k{։w��!nI��x�aM����(�lA�D$@��"F)�C�	���߽)8p���3{�oiO�p�C=�����0$�M:B(�E�1
@�D!K���};�!�x���)�.�)���H�m;��T�D�d"� ����>�<��>�=�n����/#����.�c@��H�R*��� T�BB_j���4�
�_H��w�7���ܤ!-��Ӂ�hh��B�A�Mf��%�z��9H`JŁBM\p��5�]f�sv ��5��{�-�!"o�)�$3�[Y��4K��4"��DHƑ#&�!SLi��ц��|a>щ�#9��{������I!�)��Č)Rj�$$It��G{޲�a��2���FT�
2$R�+��gI�]�*Fk3�za�K�f��	ϻ�ɮ��;�F`�� Q",7�c7��	�FIl.��\1v��&F��AB�"�@���.��	�Ԑ��֢q	$X�]�HI!&wz�.�����$,"���X� �1 ��0N&��5�^���SR�+����r�cx�gRRS�0
E
��p�5�ss��Tn�Rq6�;���%���eX�Q%���+��9�����8]�\����
D�k� �`A`�Nޘw����5�]I�o;���c�v�H%��ӛ6m٭�B�k��+�a�r�BE�B20`H@��(�H����O����t$H0��HN��h���.��4�%,jD�"Hf���"I�$Fm�jt�٬5�c4d5�&��o�̖jb���s�$"�"F1	ֱ�H�1	a7��՗�V3e"��p5���9×}�k�0%�]�X��(JbE�$b��"E�Si �H���S%1H�WJ&+��
��� �T�1b-*E��7�f�0�7���vK����O�5t��7*��B���*J���}Es��n��h�9��L�)`ń	,�HHicaZ��ۉ�@�5�hH)�HH0B)(Q!(D�) @�H�21(Q"5hH0"Ԉt$�AB*� �F	�F�Q"�H�$B,b�H�b�H�j��F�R ��H$$F��	�t�l֢�e֋
�-R���P5�X$J$P����11��D#M	���l$R#�P�
,D�B��Lk� ��������:(b���IGY	��.�a+	R��RjC����.�Y!��F$)�� L�-���!
j�E�%�!� R���! �!	w�}�H&(Fta�}�t#~i��B@��}�zYIe�9����%�%��k}�w�e�meXMa�]f�n��t������K��>����v0�1a��f��,~J�_��n(�5$`�f�8t��!���c��]8�9ϰ�|�����B�3T���7Revp��L�;3'>J?atIlfk����.QD�
Gr�ʺ"��1��]u%Ҏc�<�������3��������c$�e�`�� �t�˧&]�[	�^HjO�]I���5	0�h���4@�4+
��4H�HāT�T��,,������CP���b}���������gs�9��u��]jݓ��E�\4K�%�
³��rvI�e����s��                                                                 �`z                                                                    �           �@                                                                  � rv�u�l8muSi���l:0UNH$t�.����Q�('��Wm<ݺ .���['�Z��w�e�2�p�.���V�T�Y"�ŀ�� �[\�XԵlM��/F �L`6��:��� �M*�5����g2���\�x87\*�\\�T�R�Dg�m�q�n�F�zBWe�[3��5:)T�rtUUZ�*P鴒u�i�F��H,��ص��ѷM/<iV�v3:�AD vE�z�.G�Nʩd�rH�⮺��k�\ �7m���*Z4�u�䎑����m�� �Ė�!n���l H���o���d��ز`�m�,�a�mVQ�5N_���[UT���Yn��J�(꫕eX
�N�@ m���ipZη��u�am���K(  �'mo����,#[n9��        l�p 	 q��d7+�T6���[j�mUV�N6��ڶ[@���q mIsS(�u�Sl��Pkq����ճ��.�/���ʠU���nA��6���+
��,g94%UWU�{R�T�b�y����\��i@�gj ܼd�:t۶��
ZH*�iT�tJ��j�W�/��'Gn�`FWq��n�F6֛[@%MY�M��G����i�7Un���vYf��a�l 6�u��Ttܐ|~?>.L���	t�%���㪩�i
�J�R۵R���Z�mlL�[qm-�  ���5�m� ��M�n�Cv։#�MoB]m[@e� pnBI%��qv��m  p Zl      ���%v��  @h��i��mHZ����vjU�n��t�v䊪�[�z�T� � 	5��  ���i-l-6 � [W]� 	p�nkv�����m�M��J8Z�����X⫪�T.���;:]�hV������7C��_%�ԫU@Uʧ�;dv�A�Uy�p��8될�nL� l���UmJ��n�˜��P;j�ڈ�N���7`��J[,��N�;l�UU*ҭ۶�ތy&��l��և�ܲ-�u��-�p�XI�l�6ؙ1ve����@�*�BUS� �����
���klְH,�p��T��Y\� ��*�T�6Ҡ�nXC��yj���� �:�5�ٳv���NǶN����
'wYs�H��U�l�iY�  ���)���am  6� �� H H I 
R�� � ���۝� �~� p k �`    $m�    7n�� $    )m׮$ �� ڶx�L��ݶp���l��*m�۶s,;c���� ��l  [@  m��ۀ  -� 8jF�T�mm �`h   ���kXm���  � [Kh    ��l �   5�m ���	m��  �e�e���4�m��H��#��ʺ�]�*��v�lrmp lm[m]5�   ��nٰu�n�  �   n�H   �`���h��86ݖI�N��$K��C��� 'A�M�[��Il����WlX/.^�,ÓK������j���p�]�H�$	ӂ���kY6�8�ʽ�UT�����auCUU*�UF�@��� �۳���Z�/P mn�����k��:�+r��54$����ֶ��-���Q  �f�$ �  p�Ú鄜A��N0�
��[mnղ�( ��i4�������m� h�    �m����@H  ��t���v��i$���/Y/[@  A�v��a%�8 �]�� m� /Ze��UUU`%YUV�� ���  m� [@      H  �   [@ ��沷6^^���K���q�( -� l�  �.��e� Z�i0��I�9����� 	      6�ph   �E3I�&Դ�[�+8ewc��U p  @    ֱ��wQ֑�   Vԙ�D��;b��5sP�u�(��� �-W)AT���)���z  �8m�`tڗv�K=<Q�@UQ[4�
�U��9�]�YC����%ՙ�o�[M[Z�7Bڗ2�n�����ZͶ�,�jp�u��!������:�Y��  �$7^ץ�yr�۴�;nl$u�Kd�	d%�;\ ޽�֖���H ��%.����ٲ�M� �^Tܤ��`ݶ��D�$ ֵ����q6�&�� .�@  �   8#n�`ڶ�W��[x6���%)oT�m]��P6�[n�l�L   ;vڦۄ��8 8�b�n � �  l��            �z�M�m�m  �  $   ��[@� lH m��i0 � ���VB�+YF��@m�l�p��e �Y�4���!'l�m� J�kh�F�  �ݮ "@  km��@p   8  �  p    h     m� �         l     -��h[[l    �[@H ���v�  {=��@ q�l�-�mn���KM�ޠ%�m���mk�	eH��`n�l B@��sm�m���gI"L�G��۶��m� p  �$�Iq���[n� 8 m  m�  ��� А H[M��` �    �@�� h��m�6ݒ@ ��  �I�[\  �8u����~zm�l�V��p4��j����k� �.�Y���I�O&�N�  $���V���gT*ʡ4*����#���5��@WUE��m����� � �`�n��l:���U���f�t�����h!5�b�sjͰ�Z���K���������W���Ν�܋ƶ��m���mH���&�-�d0  �A�ccekHܜN�m���W�L�rY�-:E��ͺ�� H���Mΐ  -��e�kh�w-�d�T�m� H�� �V��U��8�'ׁm-��I$#��`���M/3� � �m��5��P .�IbP�2����=�A<�Q��Vl����W㷾�6�nɚK"@84V��*�U��n2�:�K���+��gj�Z�55WOS��7"ʰ� �:WT�UsڢBj'2U��q!�����{[�)v9�-RT��gn�F��9�ݐ�K�Kn�T�����A�t �8�̍��\۳��֢\b��K*��u�phM7�6�q&tq�lW��":]�-����s� Sn�Lp�l�m�4P6��y'[�̶i|��wm�:I5*�mU��xř�9��!�4�Z-�86���T�Қ�����(�ͳ��ؤ�i����qӹH��
&����{Um�)�-F�2��%Yɲ��n�dh0�u͎&�fK�ګ�gd�Eɦ-�H�W��M�+l��m�	&��M,�D��H[@���N	Z�P0ռ�Ud�L�0�[D�m�۰��E� ]�v݊0��8����0 �:�b@s��'YI �d�ڛ^	��n
��U<e�;ZY۝�<�Hg��}v�k��n�I qm   �ݨu܅���`�X�eY��Y4Iv�$�b� d�!�ַf�V^����]��ΐ���������ҼP�Q��lpҧfB�m� [Mkm��\$ pj�@n�%l�@  ��lm��"D�k�� zq�  �s� H  -��� �h-��@ G\hMRt7]esi*tێ64Jes m�6�ֳ2ff��TTQSh�Ch��!US�A���� �@H� @P��*��+�>G��AK���Wt��E�z!Q\
��Dq� Q8.΂�"��W�D6&�
�)S�@��GDBU~� k�h�N�p
� 0 ��*>��z�8��_�O�Q��0|�D::��1	��=�l�Q��AS`�x��6"T��|�G�	�x��ʛ��&�*���^�K�E�v�!��b;U
�h 6� �t(u�b��A7hw��4�Tt� ~P4y%
��ޯ�V"@�} u���^�	��z
�(l 4	�Sj'�.��ʉ��#��R���@�E
��Lx� q��R#�?"�� �` RF(�b� �b�~U`�P6�tp�+DځD�����UAWb�$�?�@�US�YӼ�y�y׻��            m�      p      �` 6�           UUUPl�Gt.�u[���E�j��9�;v��̖�,[�4bLd�ѹm�L�4�5�L��Y�L��|��xɴ�f|&] �z2ꪪ�T�y/T�A�'E��;w-��JYks�*�2qzN$r0NL�v��,-(:�s��ث�E� x��L�/������*h�ֶ^�n8�YEX�=��#m�
&Ӳ:3\�q��zM��v��ۙ�=�M]�Ԫ��r�Z�Ӗ����۴�lE�����5)�]�x�I��Q��(�jj��H��� ��Up
���3��2�ն� �i���n��� ��@m�dv�m
����Bl2��R�]�Tg�类y � �mb�U�:F;*T��ƖZ��+�]��8��Y�*�b��5��`Hֱ�iml�g�u�6��K���U�
��yX
ڎZ�dt��,�ۙB�j�1Mx5�J��UN4��c�lrލ��|�'\k�n�n��I��Y'�ط5dײ�$�'��{��$�"R�W�a�U�i�.��\���l�u�ඁ[T�v�s���,��
�{#]ע6�[�"i�� [M��ΝeMU��Y` eB� �Pkj�M�v��hrR`�m�������iPIL�sOh�k��u�8�IJu*��6���/aR���ˣ5P �m���8�	�@n�n��87OUu�D@<�`6��<��4����ͧ�1kA��r��,���k���"kh$5�t��2�i��uU�A\�eB�-yd��KǦ�W6VV�[��x瘌�=�^wW҆�N���A�A<A�\�՜��u�nn`B����4�a�VFx;:,�nj���ѱm�u�-�HK��;i#��U������*uWH$Wb�T?��O��¡��lAZ A>E��W�fffff`6��۶� �D���%�x4��r�gC��%S���th��w�;\��fE�Cgi�	=W[#���i�6�&z9^*��b�;&d685�8
ݦM�A�N�۞qo14l�Y�<cZЮa@t�k�)]�a�ު<<�J�N�RN�Ý5��a3�\��㋗]��`�ɒ\�K�֮d��%�K.���j�_~w�����UTP�g�aNW��ܪ��g���ϰv pll��n"nP���wuOw[��~��͉ �'>���I�}�si�%�`��oq,K������f��f��5��ӑ,KĿw^ʛ�bX�%�{��r%�bX?w���Kı9�{�ӑ,K��v�y�k4Lɬ��KL�fT�Kı/{�fӑ,K����&�X�%��{�6��bX�%�u쩸�%�b}�o��̙�f�f�eѬ�ͧ"X�%����Mı,K���m9ı,K���Sq,KĽ�}�ND�,K�z��j��.�ff&�X�%��{�6��bX�%�u쩸�%�b^��fӑ,K����&�X�%��� �����ѭfK.y���e�7)iGVq�ެ���K�SZ緳u�n�;]j4<6.d�/w�����,K�k�T�Kı/~�iȖ%�`��oq,K���ND�,C{���~���.*=�7���{�K߻��r}b?+����ND�}϶bn%�bX��}�iȖ%�b^�^ʛ�bX�'���e��f�2f���ND�,K�{f&�X�%��w�6��bX�%�u쩸�%�b^��fӑ,K���=��Y�f[u����a���%�bs���!���j%�}�~ʛ�bX�%�}�6��bX�&������bX�'�g�f�Y�8f��5��ӑ,KĽ7ı,K߻��r%�bX?{=17ı,N{���Kı?"�����
:��Yd�����[ �Fqm�]���F�q:t	;��ҳڳ�뙙S�,Kľ�fӑ,K���鉸�%�bs���"X�%�{�r��#��R9]�&��tFH9�ffm9ı,�����bX�'=�p�r%�bX��ײ��X�%�{�}�ND�&�j%��[����\u�e�L�LMı,K����iȖ%�b^�^ʛ�cENa"Z�P�!bj%�wٴ�Kİ~�zbn%�bX��l��u�p�j�5��0�r%�bX��ײ��X�%�{�}�ND�,K�g�&�X�%��w�6��bX�%�����̹�na&�.fT�Kı/~�iȖ%�`�����Kı9���ӑ,KĽ7ı,Ow=����̶�֌�Q�[u����K���x�m�
3�)��V���Δ/U�j�����x�,�����bX�'=�p�r%�bX��ײ��X�%�{��6��b#��V?Ȝc '�G!9Vr�ʱ,N{���?"�MD�/���Sq,Kľ��fӑ,K���鉹�G)�r�'����G��}ı,K���Sq,KĽ�}�ND�����MA���17ı,O�~ߪ�_�r��G+��\m�D�F����Sq,KĽ�}�ND�,K�g�&�X�%��{�6��bX(�!"*;x!��Ȝ�5�T�K�r��#��tHHԉӒK�|r��İ~�zbn%�bX����iȖ%�b^�^ʛ�bX�%�{��r%�g�g������Fr�YQ�\u.�'�'�=�+6#�ľ�d^͡�d!3y'Y�]d�d��Kı9�{�ӑ,KĽ7ı,K��ٰ��>���%����bn%�bX�׬����s&�TɭY�ӑ,KĽ7ı,K��ٴ�Kİ~�zbn%�bX����iȖ%�b_[�[�L�m�I3R�eMı,K���m9ı,�����c����~���ӑ,Kľ��eMı,K�dX�Ը�j�ffӑ,K?(05���bn%�bX�~���ӑ,KĽ7ı,K��ٴ�Kı=��i�e@R"�C���9H�#��Wٙ�iȖ%�b^�^ʛ�bX�%�{��r%�bX?{=17ı,LC�~��  ��  �o3K�ҒvŲc�tNn;NT�ӫ�k���ڨ�76X5��J�Wj��Y��8��j�ɍ���W Q\$�h�72k�����?��`+$��[y�kn�=������7<a@ݗ��ˌ�M:IR��ܲ�ݹ�t��r��[�{�g�ا9�k��2�5�䈍�:*n���5�M���?{�����w��b'
�v�1�׃��P�ć6��獧�%��F|��ɇ��e�k=;L�������bX���쩸�%�b^��ͧ"X�%����q,K���ND��7���O�%g�$������{��ı/{�fӐ�H�&�X=���&�X�%���߸m9ı,K���Sq�G)������F��%�8X�%����q,K���ND�,K���T�Kı/{�fӑ�7����>�}c�z���k��{��~ ���~���iȖ%�b_{_���X�%�{��6��bX���LK9H�#��W_���X���7I�W��Kı/{�eMı,K���m9ı,�����bX�'=�p�r%�bX��E{�������L�3Ylp�.��b�kF��d������r9�c�\�OkQ�@��\침�~oq����}�~ͧ"X�%����q,K�����&�X�%���*n%�bX���ߌ�X�ո�j�ffӑ,K���鉸@��X) H|�J�D �	�Hv���,M����Kı/{�eMı,K����W�)�r���X���T	��17ı,N{���Kı/{�eMı,K���m9ı,���������ow߷�}���CӴ��ND�,��5^��eMı,K����ND�,K�g�&�X�%�}��U�9H�#��WO,�ێ��Fj�32��X�%�{��6��bX���LMı,K���m9ı,i{�"�Y�G)�r���I$�n6��WY�'\�� �S[�ϰ��Z�ґ���'bm��BK�=�'u���}��� �k��\�-�eOp���Ɠd�l��Z�wW �����v�[u�5�ĳSy =�]�fc�&�!AP���Ι`{�`v껩n�`��p���{����d ��p��E?��_�kpM��] [f@z� ;��m��^Z��O<��`�+�ܙ9�:�����js,��	�t��M��a^M	:��F[>߿~� =�\ ����t�Z�mi����li� ��p���{����d��cI���ַX�Fۀ�\ޮ��� �k�{ݥJb�M&n6ۀ{����+ ����P�#�za%yv���8��:����n���3.��U�W7������{�� ^��m�٭�SU���k�w[s!�\�]8Q�U�[�7#�.���勞m��m��}�| ����t�}m� :��u%�n�`��p���{����d ��p��E?��^7�a���] [f@z� ;���.][P�֓�kD� ��2 {ָ���=�� �r��M7��X�4���Z�����ZXmڰ=)(J�"y���wO�/�   [@[@  Y+��O'\�*�m��R�js�2��d����O��3��Ƥ��n$�i^9]��]�LM�V�nK�*�upJ���\�X����m�l�@�$�4�qQ�&�1�����\]� keZ��Z�%��̆�|7�nհ�`�V���=�g���]�%�-!�O4v�y.�m�Qm��,��<�4�v�������w��Fm,�Z�[���7^�{[���0�J[\�+�շE<�ZF��)$,�F������t�}m� =�\��*S�x6�Y��n�WH�ِ޵���Ԩ�ǫq��&4��ِ޵���WH���X�hX��5f�� {ָ���=�� ��2 u۪�KS��L��6�wW ����l��Z�������yjP��y91v�G�v�Jn��[�v�e[U��n�]]p�/W&oi�y(���=�L�:۵`�u�	.�����F֦��T��iB��3,߃��ti	SA����~rL��}k�{��j嵦�o5���6���Z�wW ����l�׶Ɠk5����m����=�� ��2 {ָ��T�5���7m�=�� ��2 {ָ��,��)nf�$�@CM�6�`ᶶ7����θ�ݸwC�$�Ƈg8ml�٨D�H�G	!��۫ �s%�{ޮ�WH���X�ih��5f�� {�Հfc��t���W������m�8��8)%�ff��Ʌ���a�C�q���l���7 �V\oY�i�gX�N'|��D��F1"1a2:� �"�����d	�O���o�8k�\�!�i@���r�6즈�0�%%���eO���F�����&��i�ą�*2���MS*�"��,���:Ic�z�L ��l���CƳd�J2�jJ1fR�$�K���!��!���`�"F ��#*��F�@`�������*��IBP%aFV	F��F�Hz&8�b��Mb�5&����I˦+2F*L��A��)�o��<��"� ���|(���4�K!B���
ʯk�`^Հ���C��*D�	�a�����~�۳K ����"У����>�|��}�MJ2q�G*��d��ڥ�nπ37e�~����{$����\.����Y�%=Y��ؒ��.4���ooRIfx�*M�#�u����z�6�� [�� wZ���7�ݚX�[q�SR�D�Xf:��37mXݭ,�n�fL�&���D�U$����n��&�Z�wW �jTZǫq���j��t� ��� ��V]����]K*���&����16=jr	�n�7VV��@�ݵ`w2��̺�������^ݻ,I2r#����Sn�����N99�<�n��9DaQ��lU�`��W ��� ��2 {ָ�uŢ��[�԰��޶d�l��Z�wW ��*U-f�?�i���w����`������`7���&��z�<m�� {ָ���=�f@>�̀}{li&�o�� 31Ձ�3w��{wmX��X�����   ���  ջ\k4��9��Vg���<j½.���Ŷ�:����YZ�" t�G�>�n,b�h0�JX�M��NnPt[9��䮉��B1�Ճ���Fy��<���;�<\Z�d�5�D�]�s�wlRj�h9�˲E����|�?;o���`v'�*�e[ݳ7��<B[�kD]�<A[����f�����w~���|_�*���k��N�C��,�sJ�uF�\�l�s�ݓ^����2�Kkf��~���d�l��Z�wW �q���U#�#�`}��W�H=��`����s.�i#����E9�&� w~��wW ��� ��2 v,L�ҐBp	$�Գ3e��n�XfeՆ��n�}Y��W�R�M�5U`{�ڰ?	{wz���V�����ϟ} 6'RsK��Z���y7Kj�ׂu�p�w��Ƃ�'`���;:�e,qsG	�R���V�7V���J#���V�ƶ8䒔N��RG*�;��q
D��B�Q�W@��X��V[v���Gw�m�D�R��D�Xfl�=��YB���ڰ�ڰ=������CQ�$�UT��ߪ����X{�,6�\K36X��oGD���
�+��V�S��] l{V�ݫ�*��ݛ��nA
Sn"��"MЛ��gV�����RU]���!�.�غ�[����x���ݹ"jr�rW@3?~��yd�;��j]��nڰ>��;��<>�ITI<�G*���ڿ�BS&f�ٻj�=��{ʪ���f�M_iJ�7B�K���f���ٹ�b��A��x����H��������Oߧ�ٰ1t���j
��Pb�U�򫋹��Xf�Xa��6D�n�Xx�;\�I%(��J�9V��Kj��f��37mX��X(Ku��U*���j�KN&6Z�s��v���k�;G]]l�iAӶ�n�O�s��.7#�ԧ(�tI'@7M�,y�Vq�Z�.���`f97�G"%5�X�e���s�W=��]Xg���=��/yʮ${�=N:��G*��R�<�mX��Y�%
dl{,{v����y	�'*)�7I�Xo"&s7j�Ձ�7j�Q脠HW*0��E�P}�o��rI��՚�%D��)$�x�Kk������K �s%���ʭɻ$�IN�Wb)7k�n�0�e.3��a�F:B���类sz���%	u��N)ⓠf~�u`}ܘX{�7� 31l�5x���j��*8Mr���:e���8��X���pzٓۧUVƚi0i	���e�{�Հf�ϔG�s����7���>�,�܎�Q�(�	$��K0͖f���(K������O�t5����I,�2�����9����ǀ���XQ���<㪪��  6��  �8M�ҮY�-�o$�smvܻ�Ds�#��]ہ�)͞2^��,Wn���vGk#t��9�I�[Y^ ÷ Z
�;����X��/8r3��q�'��9�����$񋺈�wMn'S�pF�ed�ʪ��ϟ>h���˭ۦ�*�0s�-^3�C7%�j���ųՉx�ͬ��ds��N�9��rwwy��<�=�8:�����;���s��牔�iᨎk��Н�3?r�Ei�q�NH���`�'��;��`���|��ݺ�<��kS��i��,�̗�ă0͖��u`}�^�9ă5jf��Q)!JA�,��X�v��
&|����ڰ�쨇8G⑌�X*�r��y��v�߫��=���TD(Je��X+V�ڂQ�#�`}�XU\����_���{�̀]���&�楂O��q�\c��D�Ť9�Cչ��7U�
�y��N�����wq��L���s�?$���ڰ�X�v�K�{ZX�;q�G��M�X�{%��sܬ�HW��1��]1��#�*��Vk�,�n�R�2f9��-R�CqGD$���u`}�Y��G��,0͖|<i�JIȘ�t�6'�oK �ݫ �1Ն����<��kT�S��Cp��2X���w�� ut�w�V�m���"��4��h{a��+�\r��=���tQ�rn�I��զZh�$)89'�~�-�O��ݵ`w3��3v��UO&�G⑌�X�e���ʦ�o����ߥ�{ǲ^�+��k[��T"Er��絥�{�Օ��(JI$К�� ��*���M����rO������?5�G��ӕ*I!a���%��V ���y�V�%>{zX�;q�E�8�D�X�{%���9�n�_�٥�w������I$�D�-۬�X�'������%�ц$E�_3��H���v���{ڏ���z����~m�wmX�L�y�Ԕ.�%(J/�=�6 �666=��ں�s3u�Mk3S5��A����~���T,llo{��lA�lllo�=�6 �666=���6 �(%���u��]]_�2e�5tMk&�A������f�A�����߳b �b�! PA�}���M�<����o�lA�lllo�_�S�՘d�����͈<����`�}��ٱ�A�A�A�A�o�؃� � � � ����6 �66
<����J�)� ������w6 �666?����,�35�f\�˓3b �`�`�`������A�A�A�C�D��~��؃�lllo����y�z�͈<��U�W*���W1��n��I7j*:WcV�d�$�z�ح(�#p����bl1;�ݘa�kz��.L.\�fd؃�lll{���M�<�����~͈<������f��A�A�A�A�o�؃� � � � ��{W���\�2��ffd؃� � � � ����؃�
6667����y���M�<��������b �� � ҹU��-�7#�@��Iuʮ|W*��z�͈<����{���A�Q�A�A����lA�lllo{��lA�lll{�_�Zᙢf�sR\�3W3b �`�b��Qu{���b �`�`�`��o�lA�lllo{��lA�ll?�`��~���b �`�`�`���?�u?�3E�ɓY���ɱ�A�A�A�A�߷�lA�lllP�D��{��6 ������y���M�<����
�cЀ� ���:2~��`
�i�~������k�D��YI�u1�]��u�Z�HP��Ym���`B�R@5$~� F!
PD+d�a	�`�XMH�A����(aFNAɥX7D%�a�[�"	!"�2���GD��&���Y==��h��h�]K��I���<��N�>t�~~�                   p      ݶ            �� -�jK.u�.�Vi���R�9����+�n�3d�i��a��h3)���e�l�y�n[a��o1����B�w]D�sp�1��ir�h�֤����S#[�j��=SX���;�mn'��ctk���"{��GS���s,SE8ċ8�@r��kv����3�;*�YA�R�(��8�÷=s�h�M�&YRN�^�z!;H�K;;g*+v΂������7�@%����v���q��iP�����SU;�m���k���,e��@%�%�6�m@4�I6 vU�Z.5���(�-U�͵��V �$���T���T�LYM8��4���mTUI Q��FӇ9;x;Mp��9���c����s�^�x�岰�
�@#` �c��X��j�YYT�H5���qĆL$��R�UT�O�{Sԩ�[s/\�em�ԥ�}�)��'
���3D�]�Z�z�� �k:�q�Rmۥ���\'g��݉`�����YN�͇���b�p��e%U�m��̴�]E/:Olʲ�EU �&���m��F�d�v<���{10��.�m�6j�֛5VI�$$i����f$�*�l�lĝm�:\�5�c:��\`9�27��V�U�檀�S6��y՜X#�*��\�:3+Ҧ����[�gi�[��X��d70�Zʈ�l�v��]G:w�5We�{2YC�����I�Ke�Z�7"����u���/V�I��qɧl���7mr��ͳ�u��nsbM	��(���8*�q��"GCy���n�rs@�=<��f��݊tR�������`���#��<:)�5��"0u�2|N��
��׫g@������λt�j�^U��n,�B��7["�t���=����w�{��~@�������u?^�|U� N�'P<�`���}��   [@[@  X�۬͆�����ϑ��C�ee��nd�kY��>(�%�]&�P�����4�N��Md��G��{-�gm�A:
�Q�{�����̤��F������g�k�X��U� 4�A��u���� 8ob�SJ��7e�*cAO��1���q�歮ܼh�ΰ�'Z��\�� Ӡ(�M�+��������w�}�� I��2��6�^�ү��y;sՒ�NY!*�=���u��|��қ���˄ֳkb�����ٱ�A�A�A�A����؃� � � � ����m@9����A�ʮ"�UŚ�0����'$��S� � � � �z{�lA�G�U�.��� � �����y����؃� � � � ����؃Ȁ66;�f�C�rG �%�*��\��+�66=����y����A� �A�A���ٱ�A�A�A�A����؃� � � � �����~֮I�0�rٙ�b �`�`X ����6 �6667���6 �
Q"������:�)����{�����"'NT�$��w�����9\Y�l���� ��������m��փ4A=R=�*������q\X�g�3c�:7E<�{��#Wq�E�#$���6X�X�L�D/�Q���X��<wR:%78胒��rao���9�
*Q�"� � 	 �����i`�Հf��$��1�֘��$�T䌎sf���K7��q#0ݖ��K��lxㄦJ�G9E��P�s7j�7j���2��J#�ǿw��7��x�*�\�8r��� ��b�ͽ:=�,�n�m��~����G<Lry9t���N:�U&�ѭ�r����&ru����n����S�|��`�'#�C��=�X�L,�̟�����s�����?*�_�_���"4J���t�؈�2��`��X�^�Uq#����H8���J�Ȭ��ٹ$�}}��AχH�'�Ns^�<X�5Xg�\m�QG*H�JI,>J|�"!%�n�?U����`fq��ky\�Ur��� ��jn�GD��MU���JBY����ڰ�?^�'ߟ>�%���[�m&^�����������E&
{q���9������|t|��7V6�m�3�-��޵��6���{f�V�Sc�%2E(n� ���Ԣd�ڰ36��38���A�k�HTrpRK �ղ��raf�,Ǻ��ݖu��C�D�6G��_�g����X{��#^�P������f���=��2�Q�$���<�`~�9T�������}�� ����m��Sc��l�bxX�'c�/4k�������ƾo{|K��g�;��,]��1$��ϿǲI��,��ɇ�A��U��ŷq�$����i��v�ޮ��n�{��{ݷR����OE�`ַ ������b�i#�͖��e�������r&I!,5fM�`�l�{8ޮ���ubU�ǌo^��{X����v��kK3�́�<�>�  �H  �n�r�N��cm�òJ�i�WR��r��vL�2�u�u�m���dٱj8�g�\���֏0�2�S�r@>�U��j�uG'n�lEr��vT-�w��vv���&�]�^٠�1�[*�xq�ù֦ؕq�=:5:��N�@ӻ8N/6�nfX�+u¥�-��4��g��a-��h�N)��d����~w��{�n�0�����ۮ�I9lk]��յ=#�W˃���w���C�G#v��ș�� �~������[�h�W /gQh�����4���ޮ��n�{���k�]˜��37^�1=d�[����u��z�,�Ʋ5 �"t�J�Ȭ?�I{ٲ�35l�>�L,7��&�;���n:#��JQ�`�,����\��ߎ���~V��%��zd�T�I�ہz�@��ӎ�I�U����;&�B#�<k%s����Ҹ��wj&�tIM��I���,y�+ �}�y�|��ղ��jz���r&I!,{&|�Ur��9v��ݝ��t��K䣜2~����>��rH���37��{K7��]��,͚X�bco%I ����Is��O�`c��,�L��3���}[�MH�H��$RXw&��@{���k�_u���m��j�X�l	<�On��n'��x�om<����m��p��&�W(P�#q�����I!�7Oŀ{���3�ԔvCٵ����9;�T�NHX{���W�W)����K��~,{&��U$wqm��tF�"�8Mr���ڰ;�L���I""�U+H�)G�?|��~�>��fn������:#�&�tF��ڈP�ٷ���֖�c����2�θ��-_�m���Ɠd��@6DBS��� ��Ձ�:e��I=����X��Ƶt��3���ѧZ�Q��8���=��cK�{[��Z�--�Tݖ� �{V��Ձ�:gД%����թ���%G ��{K��P�Of֖{ZX�����Q
8��V�i��H�GP�I`{?OŁ�:e��""d�{V ��Հ���+�	(�"HXmUUqfm�`�l�c�V�V�GcTD%���,���q�ŉ���� �����>�t�=�X�\�ܽ�ӌmH��L�����>�դqNS�b��ݶ5mV�:��l�����TmK��茐Rrtw��,��g���cڰ3��Eq4�tF��>�L/y�UU$f=�`�j�3������DD$��4��<����#��#����~V��%�ʮW9T���e��l���b1:o#t�G�T�j��B��ǵ`��X�X�݀v�5V&��&jn wYu`jID(^ͽ:|ݛ ��Հ���~~��   �h  8c^ܗdײ�{X��3�1|�Ήj��tv��H��W��!;&i�0�
mt�`��U�t�ݧ�"3ks'j�z.������gB�f{�vK�y\�p�,��۰��x��UVdA��;����v��Yg(9O���i;�4:,�^��S�q���p�|ћ{s�,q��f7-����+�UU+Ө�،�A�h�Gp����δ���ٮ�1����V�O����{�������6�� ���,�76�c���$� 7���Ն���QʍBI�y���D$�C1�~]�7~����mi`y�NKkщ,I���W ;���U�W�i`f=�`}�Yq���HM�a��*���ղ��i`{�1X~��W?s��Sy��X��'r(萑���5%��ra`mUUVd�_ {ٲ�;�� �+[om���'�&�3n�m�{zW=�|0T�a���c#؝�b�n�!�owq7��cL�w+v {�\ �f�\�}�K�Q������Q�˹$���7���0Q�#bFaaE#!  D�M:"�A-O�Ą�_�����}V������sz���թ���rpNK �ղ���0��Q�D(\��>�l�����y'+��Bm��p�] �݀�Wa���U%��e���7�������t�RQ9�k���X�������^Z�-M��9c���K1ôn[���p�\l�bt��7��x��{��M�O���Hx�bm� w_� w]����j���f�,�-�ێ��J���V��Ձ�:e����c��D~��Sff��܊:#$Q����~��rN��鹣K�%C# = V,XL�{J@�$�!� @�, ��D"��ա}��Ev�I�Pt|�P�l4s���HŐ�ȄJ.�YU�B0%IX�@��P��4���D�)�������I�YP��H��M$i� H�+xv���T&�� �d�/HA$X�`� ���h[)+ ���j@�)
	$(,`+(�+$,b��,F��©(B�j�*B�
2�B	���X��:Z�I��[KBZ��2_��*�����C�H�W�'ʠ|��y��N�1��"��6�TDB\����v"=�|�V ��Ձ�8��(�NEQ�G��Y�zX���u��z�@>ۥբۭ&b֩�,��V�J[���ͭ,��=�|��>�:]��γu�`���c�>�cUq9��34�t1��6&���t���~vQG!M��> �ղ���0�=�~�9UU�������?g��hr��(�$#��z�@;�� ����v��3Q��7�����f�,��K?s���l���K��~,�Ʋ5!"Pn"SrB�j���e�fj�`}ܘX}�U}�r��?{>���|��n:#�D!G%�{زXU�m���4��ߟ^�?������� ��M��jT��(j뫶�hR��	䪮w=v���/�wv��w"����tF�����`{�0���6�� 35l�;�֞ҎAS�SI�2�] �����>�t��q#�Q��z(�)�%$�`�l�{K6�Ļ�X�uX�bt7��Q�SpnK��K3V��٥��V� ���}K�D�kOZlo]X�X�n�g��j�3��?���~��?@  m�[@  Y5��6����wl��;b�ю3�[v�
�mt]����oWR6�C�-E#�;q��H����z�kH]��W�k9Y�>�sEU�{%m-m�fUi���s:��ջ��sֻaLfKK��&��v�JG�YrL��r�5�ƣX�
�'����s��s'\��n��;]���# E�y�v����~���{��~|�~K�W����/	�WcV�`�j��:;5 ��Ny��]ca���N���W��4�UG�~_�>�l��V��Ձ�:e��x�GR%�%6�V��%�q �ղ��i`{�1^��[q����B�K �ղ���0���U\�\�ou���3K����E���W&���2���s`�:�ԔL�����Z{JI��#p�����Nc��{;V|��c������30�2���a;�r��d.����@a��w�a;�s�^��x�V>m������3��;�L��d����7���I��)�7%�{ز]Ԫ��W
��!TDBH�ձ	{�3kK�7f�=� _R��<Z��i�7��>�t�38�ٰ�L��j��ڰ��8�JJj8�$,2���*��ސ�͖�p3��s����`{^��G�1'�ē{ =� w]���������I�~� :�6��d'T���`9T.�U����s�G�觇��w��j>|��Dc��(��3V�������b�UUs���,{�lr�RD���z�@;�� =� w]�~�Uq#�=i�)$J����8X�u\�}�}������(+��W��L����f����u�I)���V��%�{زXw&Uř7U�f�N��9#)�7%�{زX�w�z|c�V��KR8{��7M�(牎O'&|^�i�Z�3�f�p��Saۨf5����G'r:7$��E~m�]2���s`�u��d�v��7Hܧn!�$,y�+ԃ�ݖ��e������<k�'�q�r��=���3��T�f֖|ݛ��q���)$�ڤ�5l�=�X��V�Iw����|�;�GD�!M�{�s&���ݖ�v�{�m�m�$�lz�@�۶���F�"����dl���3۞���2CqS[�?�d�[�޵������W�=�XZ�N����
�SN+ �����d�ڰ36��38����$�S���$ख��\ޮ��n�z� /�uh�-�(�$$RXo���Ł��~V��K�K3V�W��7)��R(9!`z^>X�DD�n�@7\�X�X�X5"�E`��=�g333   ����  ����煉���I�V	�ڥX�L��X*�sup�k��g�f��͂�Q ��v���,�D�����bZ�����E���Jcv�d�u1�6�9F�����t�βWf�keX�ö\Pʨ[��{>Py� /h\ok��h���������y��m�mm���v��ܥ=vTJ�	vuͯi�w;���'������ 휎ƪ��ݪ�&�:q�I�:wO\���f���W�6����0IY����~�8ompz�@=���}{lkSX6!�馶� ����] ��v��K�$fj��:$%D�(�G ���m��k��� �	bx�#J59$�p��繮�=��`亰�$�#����Ł���O8��ʧ����ڀ�� [�\ޮ�m��Ɩ�[m6�4Onjś����qkX��m`�s�m���u������$;/�(I �$�w��Ʌ�՞���ʯ�]`f~�,�������1�	SU`{ΙdBQԜ$�{�dվXf9`�Y/k�H��t��q4�ʄ��2u�,�n��Dɺ�j������4y<qH�d��Ӓ;ܪ���e�n��`w�0��UU/=�vw�i�D��(�)$��,��罷��ynk�<��vj����$�$�H�7��a�v�m��xҔx���]Ar˵�l��s��{���Zw	��Ӆ�>��K�z�ouP���x\�]ku��I!,��;ڮr�1fk��[,�&�UĎ�F���S�T*Hӓ���� �K�+�BNRIM������X���ر<RB8I Ƣq�~�%��e��٥�՞�`y{���ቡ�j8���I`}�0�7������ ���z��m��uaՇ''�����k�'\/^�Uո̝���?>X�OJ�M�IB��21)P�������omp�t�z�;UO\�21�i����c��+�q���W�`{����:�����.5#�*H�T��Xy.��L��8������ܰ=�X���JT�p�5%�󔻻zX:��Nc�� P�Q��UN�ۀ}�r�tm���X�cL�{oU �D}	F�����l�V[�X��s�j�9�����'l����61q<����n	|엮k��הɞJ殷T�?62s,��V[�jQ��׼��׮HG	$)�'�fyd��s�H��i`d��X��_�$�C٦�$�&��1�	���K�=����q#�ݖ��e���a��NT!$��z��Z����=�� �Zv�X�Z���jm��Z����=�L�=/,�u(�$��$�$��.��5i�����Ēm��t=F@�tA\Yڎ$ �`�
5@t(�� ���-��#�R��*s��b�d��b�M�P��11GH�$�0�p
�,O{o�y�$���֑7;9)@��.������                        m�               [b���\����/h�3ɧ;t���m	͹=l�͋m]�K8�l7=\	�����F�7[�U�d�y�i�]%�\X��qځ[;������ɤ�Zd�Րxۜ�l���m�rp�����3����ۆ���V�]v��j�S��ͭ�KR=��L�1ٖ�[p )#"v�[���m1l�M��U��X(�6��v�ۏ\������Hs��ʹ��.�B�9�V��_u��/+���m]n�u�\�� ��i�-��N�d+c4�x���%@�J� r�m��m�m��z�&]�L�r��5VƆ6*�`����)U�HL�)`�ְd����R�յWU($�vu�˻ܛx�`mӬ�slv��,��n]R񗮙ᣐ���C[���s�O�i yj�eYYXr�ʵ��X�Y��U`8m��m�I*Ӟ� �Y^�
H�.���iג�6�Bj�CKs>"9����&V����[�l<�L�\mحm٪��L-��Kk��h'�V�gF�s�뫬�sm��6��X=�m@J�@[V�I�d�����6\�ʺN�]s����n�&�������b[��Xm&��[E��kh,T���ԝP�<�#�l�q���/=�mE66JӶ�6Q�e�䗫����̂vH�5%��#�[�l�e��ɮ�v�vɮ'l�'[�G.l���n4h[�uu0��[�u2tJhWh
�^=U��`���Y	�m��mm��ѵ7D��l��d�x��Ƀ�S`�&;7E�Ŏ/nw�h{On�����rVuι�n0��m.-��g�;���`v��73�n��U�+�;cKˡ^�o2"��P�9�s��V��/Y��<�cFgev�v��MR� h�B��m�� ���C Q� zP^��/�T'���=O�Ezj'ύ�mh�p@�o�fffffff` -�$   J�b�����@�u����ºE���i��fa�*xxz�z�K��չ2%��۰�S6��-)DD�OA6l��5K�Vs��ʽ��O���%ɪ���մ݂��R�Vֹ̛i�-�Hm��@���kjv[e�Sf�;���n��]�Yͱ�L:�y��T�X^�*�Fk3��c�ʽ�'5�s5�Z���D�:Ll���m�A���M�[W\��n�'k��Y��:�'Q6 ��m����Ձ�:e��x��DGd�ڰ���К�x�5��5��=�� �ު {���3<�^�*��RG�-M�D���m��@;_� {ָompz�@>ۥա[������ڀ�� [�\ޮ�m�]*��4��1&&� ����] ��@~���I��}� m��ҺX����F�;����*Z�y�] ڷ�src��HZ7$�hM��n�WH��P޵������e���F�4H�R�$���x�s�
�(�κ�ܺ�=�L�=U[u��ѫG��5 =�\ ����] ��@>��5��ք��7w[n [�\ޮ�m��k�w]��Z�'��I=��n�WH��P޵�{k�{��m�m�T���.����	\�eᕞ���݈�`5���f\�,Sl4�S��6�����{�Հ7��a$�!������6Z68��5QƜ��;��{U�U$������@=���t����l�r�UU�7�����2�!vM(��ku@�\ �Ժ�Mؘ&��U`{Ι`d�|�y���J&wG�`j�S{"#�dh��{�w��i��=�� �z��&��"��n^X�kn�r�n^�e�=I�bH�{%;un�e�E"j'9���Ͷ�>��`-:��] ���}{lk[Y�(��RI`��^�#�٥��s\ ��p�TkZ��z�X17 �����P޵�N���)rG	�,6�\��s]�{۲�1Ճ���P�@��C%(�D��! `�? �*� F) ����� �a`�!B�
�"m�����M�ei�4���6��k��\ޮ���@;˫m���R{���,*k����m��d})@�͑���U�l[��1W i6�cm��n [�\ޮ�m�@z� =�]Z&�M���y�/b"&G;��;
d�ݫ �7\�.�Z���Ƶ�d�ڠ�k����] U[u�޵�n�ǋSj {ָik�{���mP�m�kk5�=z�tm�imX�X-�X��X�PBHo�   � �� u'�v���.�L;k^��v\��l�ND�u݌<�V�e/B1q�uƳ8��J/Z�ԭ��!��B��α�4���]h��dgeP��J�k�l\t���Uй�ۜBONi!�A底�#��R�9��E�u��\y�U#c��M=o%��m�Qz�:���G4d�N����-���{+UUP��Λ�I�Ss�I��llZظm���BW�|��Y��)$�ut,��_�o�߷��mP޵�K\��u+�6�[z��� �� =z�ik�{�0��$uj1�����Gn; �{V ��Y艜�J��m��=�bZ��$�P�`�s�{�� ��Z��K�D��z���ۀ{���mP޵�K\���ū�=S�&\��\[s��O\Ge�aMi��r<]^����*�ZMp�j�������P޵�K\ޮ����&��SZ�5u���'�{ٸ�p:�@�e���������\���-�Ԏ�mH(��$��vX�L,,�P޵�;�j��X�7�Rx�bn��(�ͽ,;�� ��� ln�omԮ4��m��Г ����� w�ޮ��um��lƚST�4���nw�r���Ŷ���٠�4�(k���H�tԌL�Tq�#��2X^���t�{oU :�Ui�M�m����3<�^��U${�4�<�5�{�,�ቦ�j��'$RX���'����:�~ܨ��H������7��X���F����D�,K�� ��� o%Ն�B�ͽ,kֶ7#Q�n$�4�v��K ����] ��@>�Z�m��jNu��6�#����drnU�mN�@��O0�gYz�*Jx�n"���}��}�`����z��Z��j�mf�I����t�{oU =�\ ������WmcHI�m��k��� ����]-�	1�Z�P޵�{k�{����F!@G�HQBJ��w� �#�"r)$)�9%�f�`mr��m���5�{�,���tܑ6�BR��sϞ����n��I�������`O,h碑t��Tz�kKq6�SLcn�WHm��k��\�.�Zצ�x-{�l�vު {ָi��=�� ���mkZ�[��Ԛ��� Zupz�@;oU ���ֶ�Z�O5���ۀ�\ޮ���@�����ݖf�v�)M�"l�K�Ʌ�����=���1ՀBIG"Ȑ"D ��D��UW�|�   hh  
��77�C����m-IVㅳʚ�VU��vi�WKC��Rm)rָ�p�n��4�Ձ���@��Q����8-sْ�B�������j�=Z��J�v.m��
6����`s�3�S�M�ز�
����h�yBvyGrGl#��7M�0g�s���76�XB�\\�s�rd�m����Xa�{���㽽�y���p5��UmI��E�'���[p����ŸG�6�3����R���D��]� {ָi��=�� �n��B�	c[�5�� =�\ ����t�vު uҪ�z�i�13[pӫ�{���z��Z�ޥիZ[�5������] ����� Zup�h��{���պ6�m��k��\ޯ��'�ߟ} 6r8k9��u�ۈ���-Y	���Nԛ���|J3y���ʵK�0OM��w�� Zupz�@;oU ���֦�b��V���p��͈Y�l �v��̙߳�rO_�T ��p�D&�x���#6��t�v�T ��p�� �u+��{�����L�v�T ��p�� �s��t�Ii^4��i�U\��u`}	B��v��ZX-�X�sۻ�mH㑶"@i4�`�N�Zŭc
����qg�\��9o��[�J�n��9$Q���,w��3� ;���;�54�mSq����ΐ�j�^� ZZ�ܴZ������ �� >�\.fo�	$�F4P7�6�1�����0HXX��*j�<Db���7F@��ډjQ�5��*�O�QѤѡ�YE ��J�]@��B���h_��P�
�hiƂ&ڒ4A �t��F*A� �@%E�	���4��V6�Q�B0��Z!E���M(:E:� W�yU��ǁ'RP�HQWC²���,|���'�'��ڀ^� ZZ��t�v�T��cZ�ưկ4{�������Hm�@z� ����]�f�f�X�*t�JQ�ˎ]X�[S�)2�'\�&s=�
Uݘۀ{���mP޵�K\��x�#I�H��,,�w��+���,tݖ{�����c1��6��k����] U� :���kRm�z��m�J����2����ð���!Aޮ%wθޥիZ[��i�M�=�� �] �k����t�GV0L����`K�z�zu�][��9�7�8���.�ա�`͵�U�6������� Zupz�@W�$�H���S�$r|�K�˅��Y�d���Ƀ��^̼>��s��k۪\i�QP�R���B�I-�v}�Iud��I/f^|�K�˅����c��:#iH6�r}�Iud��I/g��I%�e��[\�ot͟|�^x�7h�4��ԑ��I/g��I%�e��I,��>�$�}��ݶ�	��A�R���J��GA���(Q��}�   �m  6��-�nyVq9��&׊MP�Rƞ^g�R5C���D��L��7�<M�����R©:�u��HN�ɬ��@�
�"�)�n���M�r�yedP��':�ݞq�حcX����U�ݢ�Hjm�rn�����λ���z`$=����6f[�]���p��Շ1�j���v��6�7r��������/-3i8��e�N�qI�GL`�Q�s����`�=��sN���L��]�Z?@�.�If���%Փ��U|�K6f����?���r�Q�f�� >�߹>�$��`�$��{�$����i$����D�ᜳkU���>�s� ��{�-�6��ߡ�I%�fϾI,l�"q�IҐ�' �$��{�$����i$�a�|�]Y0v�K���I8�Jr��E��%�e�ZI-{�l�RK�f������~~ }?o���4\��Mx9�P����'������C�ݯn�G�"���EB%B$����K0̟|�]Y0v�K�3��ZIfm��Ifj��umH6��}�Iud��W9*��������	@Bؽq9�}�sלI%��I$����%�剻���#�"���^ɘ��$���I$�����}����~��T�n��D�/�Ims��oд�Ktݟ|�]Y0v�K��ߟw�� }>�j�j(�V� ,�2}�Iud��I/f^|�K�˅������ �;f����D��K�q{l8&�(�ˍˠ9z���CM��T�L%˖�r}�Iud��I/f^|�K�˅��Y�d�����'�ԨB9i$��x}�I/{.�If��K�&�߷�}����6�� ?~����z{��^�O������դ��z����deƜu���B�I,�2}�Iud��I/f^|�K�˷������s=
��{Z�����`�$��Vn��z�K7n�If���m�~>��v�e�IO+��c�ڧ<1^V�u3v���`|s�k����I���Z��H7i$��>�$��.�Ig����%�h����N�����PMI!$��e��I,�>�$��-�K�ϟw�� }7ߴȵu:�| ��d���L�ZI/f^|�KٗI$��5�&�6')��'�$��e��I{�ߧ9m����n�� ����GIa-Q�T��`ԀFTF�i �\��[�����֧�H�dC�R�E���e���$��p��K0̟|�^ɖ�I%�U�l���7�Ŵ�sɣ[`;]�����uE�$���*i���,<(閷v��?����-$��3'�$��e��I{2����}���v5։f�� ��}�~~ {&Z-$��f/�I%�˅�Uo$�n���SI'I*m���͛h��^~�I%�z�i$��>�$���n��r6�I#��K�3�$��e��I,�2}�I{&Z-$�^#͍Ӥ7��i��I%�˅��Y�d���L�ZI/f^|����>���   �   �65�r��^Գ����Ҥ�jLOm=�cf���m��ŋ�Nz]F���J����5S�4��P�ivj'���P��Q�)��3���Q�vz�7�W5�,������0m��f���ٷ/;d��Br�Xq��۩�Uy�>9e�0������9���a��/J���ߝ�������s�H�oh�i�#��u2��ɥx@g<���bMj@�L�u5ԒHu$��=��K�2�i$��x}��̀{n�z��[���Lbn�d�t�{�� --p��=Z��i��t�{�� --pu� W-�$��B@��Z���(Jq��X�V��Vs���+Z�ǸcC�� w���d��2�d�ffy[���m�Ԟ�V]�$����Af�z�k�)	�<�]V���dg�%6��q�Ԅm�	'�{7n�����ِ�up^۩Lm6�z�6�M���2m����g_���Z��f@>ۧ$%���K5��cv�<7Vj�ǻj���K��T�4��6��@�k�{�� �s���l�{n�ik�[���Lcn�d�ΐu� x��6�\�����)(�A��EFƊ���]<E"���kys��z��J��ϖ�hK�
�U4Mr��{��`{�`Ằ=�̀uUmi&�! l���ِ�Z��f@=�� �֊֦���ǻ����� �[2�����EPz���7�Ϧ��}��>�;c��Ƥ#n�9,?s��R���1����7j�3�u`y��-6��m&�y �s��l��-pu� {�m���ki����ݗf7my��;=\[���"n�烴����@k�$�1��ĳZd�l��-pu� �t�{n���-Om�lm� ��ꈈIL��mX�i`{�z��� �Z��JM')(�$�=��Pw:@=�̀�� ꎣկ���z�i��ΐu� x���𑐉 ��E�V! � �$�"=
��7��y��u�r�P��<Xަ@=�̀�� �[2�g�O�ߟ} :�h6���4/;��5�D���u�� q��O:�r]e�u3=<1��w[y ;Ů�d�ΐu� {����	��%�pяw��y����7j�3�:�<�\�3Sz���M���H�ِ���T��3e��ݺ�:����2��Q�M2�d �\�l��}l�@<��9�G$�!$� �Od�;�ڰ;�L�=�v�.DB��\��m%�l��	�V!�~�L/�D�d^ۤ� Q��rzQ�bA�3�A*�j�&��v��R2��ОwOq-�J��ک�+�Gt�Z���J�*@(!(�J���v��=,�A��QV�U�@�'0ؿf��6�]Ih�p�AipC7�}(��Z�H@�,��~�{�                   �     �               Jrs��h\�������B�\X0��u� �6��	�%��u�k��6�����\m�ztU$l�Vysn�vs�6l4�Բ�nl�f� ��#�5��[bx���=�@g����m:��(����,9��v��G�1�I�p�{ �&�R��5�5�I�f`�Ԅ>cX8��uBp��7'����,�m�S����^|�[-6(Ká��{�v;f[m�O;f�8���Nƀ']d��ѵ�ev���4�i+b�� �m���&��i"���b5���R�mUUK�Z �j�������j��d����`�:x�`	��Tn�{EUQZ�V]�LA�C���͵jy��Ń�>8�vڷ{sm ��v���Z�Nʶ����VV۞�5�֤�j��v�[J�p�b��)V��q7TH;lj�0չ���l-폃�fUY	�q�h��f�h�܌��=�.�X�>7Z��]u��Y�ħe�M�d���ppF٪s����Jd�k����0km��'��P�^��z�SnI˸��v�V�3���;J�Q�Z�WT@T�P/�j��9����^�^ق{^(���ɷ(��A��-)�Wr�T�B���m�9,�&�̆�v�q�4��y�E�vz2[�l�im�Z�gI����eh�ɱ�v��T���v��I����>��R�	�:q�v���8�\�ِ�m��z3���<vw*�q��}��,is�l�#)m�lN�QM������a����n-Vj9yќ.����Rrv<\2�V�9d4v�K`@
��ٹZ���h&t�l^B�c���{X'���&�4�i%8�Uv�A���ۭkVq pC��&�qT�6�?���*UD��v,F;CH�7�P~�B�=&��   l�  �n�+�nr�9�v{��]^�6ݩѷ6����<�NӸx"�欦v�Z���6Iz��N�Ca�B��sr���,���y�m1	��77j۲VԦ�=�畩�{pu��Ւ�O�v�gf�j
"iV��jyj��I�A�s��1�W��Dc�SGX�T�Mv�m	��.���;b�U7I�w�u��m������w{�ϒ��19�:�sϞ�ӝ�'�.�,���͍��4�A��Cu���p�pCc5��`w2�`{��j���{Vo�=Z�-x޳Zy ����u� ;�W ��̀u\���F1$7�����ڰ��Jgٻj��u������ưĆ=ԛ��:�޶d��H��d�v����4��"���;��X
#�ޝ1� �Od�6�U[�{$�$��n�uJ2]��`㱭�b��ca�$*�s���ؠp�ԛ����i7��L�{�f@t̛�|��ݺ�:�M��eI*���U+��j�$�,�Q
�P6v����̀{�̀{n�.��Om�mky >�\�[2��2�u� /m�mך�S�ש��zِwY�{���Z���z�!���f�R�=��X�z��V|ݫ	����@������7nr1�pqT����9���o�"g�ӯ�CtIJ��+�8���tǶ���X�v��K���Vwc68�dEFB$ܕ`{1�>�� � �Y���TBk�Q�Q9,��u`w�˫/��.s��Q
U�p�P���ڰx���r眺#�2(�$nJ��W+�T���U��f�@���}�f@=�NĄ��$��o �Y����>�� u� �_߲�*P�S .�lյ�(4��LM`��ٺ����qֺ��B������Z�@wW ��̀}�̀{�f@��5�Ri9ID�NK��]^�V�����u�2 {���-��in�oY�<�}�̀{�f@wW ��̀u\���F1$=6����e�{1Ձ�7jð���Y
"!+�w�@=��ZM�{��{�7����>�� u� �Y��:�x�o[+�Ӟ�3�n�i(�=(�]]g���N�d��';K��4���*�ܣ�'��߾��}�̀{�f@wW �ݺ�cX4=z��M��d���w_� [��>�� ۧ!jU�y�V$�@=� ���}�f@>�f@=�P��u%�[x�Z�@u���� �u�W���X��5�Ri9ID�RK��2��2�u� >�\����[`  ��  [���z���F4���ns��)®k�Â�嶌<PU��XiNՑ�@�I�UV^gn+��c���Wa�b�� �t+����͕�Ϲ��6@ ��[�e�x�	�8���l����X��"CCVһ˻pm.˷���{j�Q��d��(��k�+���sl��[�nN�rK��FF��2��t߽�y6���rF�*wgj��'�/]{F3mŉ��s|��u�C`2B'8�IJ�AG+�{3n�����Z�zِ���I����MXާ�{���Z�zِw:Oܪ�H��f�n$�2&� �n�޶d�ΐ{����!5�����,z��}�f@=�� ��̀u���u(�^�^���y �u2���ڰ�u`w�ڰ5(�Y��K�L�N�rA.�V��\��nzv���vz.k��h�n��{&���s]��r����Հw��n֮�cu���5��z�u���IV��%�W+�PGA8��"��Ͻ훒{��M�w�˫ �,CX�&���N$�>�e����5(��{j�<�Ձ������5��޳Zy ����u� >���� �U�M�-z$7��{���up�l��ΐ���ĩ��X�ci�=���F=Y��,lW��ݺ��2*����Z����wW ��̀}�� ��̀}�ڢX<i�=K��zِ�����d �����ԣ��c�6�o Nw�ٹ'�w�74N ��Q"<�㯬Y6X{v���ŋ��)�N=X�y ��̀wW ��̀}�f@=�P�Uh�m�6ַ����zِ�����d�Z�m��բz����pv��3��{c���q�.G���r��H��QE)4���q'%��s.������d ����-�����޳Zy ��̝��ux�>��s��f�Ի�6���z�@=�f@���}�f@>� Z�Z����iʩ�r�XsX�7���ՃJG%Ur����������D��M�Q���T��2�u� >����	l	�JyIft��!T�_%Z%�x^�䃤�����9ּ5Ѯ��8�A6�X�v�{� �c�������,-Z��n���N�����u`{��}��@>� ިY��%�Zcmky >���� ��� ��̀ՈxԦ�r��Ĝ��]���`z�� �Y�����h�O�ůF��M��}�f@=� ���>��=�|�<������O���   [@t�  /M�8�פ㮣7>Q�e6�9�J�.���5��l�f��.g�]WS]����k���P�ZSn�b"Z����v,��j))�F��),���%����0)ХJ��L��S���ԩ-u�s]�a�UCn6ݍ<jA涧��c%��΍��>M�&u�sƜ0�k��|%~x+8wf�L�丸I��oh����V���֍k3)u�Y3&H�&փ���H����vM�Jp-�q�n�3�a�w5�I�1�В׏S�o�2 }�]��7k�Q�7��n��O*�D����ky >���� ��̀{ݗW��U$wص�tJ�BD�E$�;߿L�}�f@=� ���>�n��61��y ��̀{�̀wY`uw1�X�'K!)�ND��`w�̀wW ��� ��̀{�m��*�GlVӝzv��i��U;6�DbyZ�.�C��.�d=���M�6����>�Z�wY�{��{n����n��.��fnI�����R�Ă!�K!$��J%.Q��j��nՀw���Z-S�0LִM��l���d �up�l�U�V��1:���ҩ�+IB�ǽV�����P���ִmo[c�Zְo sX�v��v�{�a,�{@��&ӱR�V��Җ�r69"&���,��n��$��u#]�f�L��+�{7mX�v�{� �c���ԣ{���z�j�u� ��̀{�,�s�Ո���#)Iȟ�X�;V��VJ�QP�N�!*H*����"B0��&��	h�µ�>�~�iu�$�%!(u-�-#H��ˌ4���TZA.�iN�c�t�aHn����#$��h��F��P�;h��6/�Q�P�&�Aъ�v >�����P�����z�� ���e��Տ[lou��wW =z���d�l�{n�n�պٺ�=�� ���>� �̀wW �libM�kh5���4����[/�h`�d[���kr��n�X�� ��|����&	�z�&��[�d�ِ����W�n�1V�I�)�ӃMJ�ʰ3�z��y�� �ݫ��Ձ�:ᵽm�kZ�M��wW =mp���u� {������m%�j��aD�n�XomX�ڰ�
-%����7�w=��w��]ky3Ymц�������d�ِ�����O�>} %�uW^ڶ�,�Σ�X�Z�n�ny� �.��솽���hyn�E�ɷ��f@�������d˨�F9Cu�%%X��K�s�n�XomX�ڽIDL���9;4��"J7rX�vX{�uf���u`��z���1D�m5���wY��f@�����o���l��jbխ�y �d ����k�}�f@7?����`YUm��m��m�h��= q�LȽ���Sq���o<�2�j�;b�ܽ�dg�v��^(f�rn�]n�m�0��*��a���öӏlg;A����#TB\�5�3��q/%a�'5�Ϯ�뎭pn����qn�6Ԯ`��	׀\����^�i�����=khL�lS;���l\6ܐ�]��!��.R�صKm�ld��<����z u��mn�by�y����&'+1�q�	���8z���.�srN)�lxkZ�m� ��8�k�}�f@;�� �ݵD&�lOi,zۀ����d�ِ���[�R���Zz7���n�u� �d ����k�{n�V%q�[F4��o,>���z���Xmڰ;��X>Ҭ*x%�[x�Z�@���z�2�u� �d���ě4ijǈxY{v�s����q�u���,�8&�/;)9:���"kuE�^j�owZOu7 ��d��2��[	Dv@�{V�6y<�
��
�f���7$�{���*b�{���@wW :���*���I[���l��up�� ��̀w�Q�r���I*�j��f� ��~p���[f@>�mQ-k��M$����� ��̀u�d ����'߿C�����]�V���-�!��5�6A0����!� "��y���m���2�l��up[f@=��Z�Sƍm����[f^�	L��ڰ�ڰ;��X>��@n��T�rU�}�d�=��V}��.$�	%��S�_n�Xuڰ�rrZ��R$�q'%���ݖsv���l����iuj���lMbi��l�[f@wW :���c l�!j�����5��f��TJhӲ+�uѲ��4{�܏X��F[��m�MM�]�� �c� ��X��X�Ɗ֦��Z�m��� u��>�eՁ�̺��H��k��t�jR��5U`wj��7j͈S/wmX7���<�7u�B"Hकa�K���XwmX�Xu(I.�DBJ��d��*��4kh�o���f@wW ��d�d�uih���%Ƭ��Xe�sk`�ָ�:�k��c{X�7F��W7�˩�n�<�W|�o�����[f@>�f@:�2 _m�mך�[�֓�M����l�[f@wW �K�V��ִ6���p�ِ{2�ͤ�fl�n�<��x�r��64��ِ�������sw�=�͍9
%�U�w�����v���v���B���N����   mm  d��U�e�uZ���z��h�v!����ub:�;���3����`�	K����'-N�єw\�ҹF��j�[�Y{A6�6���\D�)�բVzK�aKj�eF�`��/m 4���c+N��u������:m۞y%�ϳ���۞���RU��������N4�&n�z�LMd���g��ڬV3ǽ�~���y�uo}R��4�Yp3�k�*�]��7[\M�n�O&��.4d�@Y���k�i$=m���\�d��?r����ٛ,�-M�EBRrID�U��n��J"d{�j�1�� ��Of�yU�z��F&�ky �l����[\�d��TV٩��16&� {��׫�}�̀w�� /����[���S�M�=�f@>�f@=�f@wW ��V�m���1�4�Q�[P'лKp/B=s�k��r����T �i��$j2GrJ�����] ���wu� �mZ��=]jfI��XnI�{=7�i�Dw�:�8��d��2�V�ֶ��Z5��� ����\��2}],����(���6E$��X�v�x�X|�L�����g��&���Sm᩸��d�Y������,�wf�n���Л���}�j9v������/�������mu� \�%	���17���_� ���:���}��^0;{J�[�OCbo �Ɂ��L�^�2׬�{n�qJM)rX�eՁ���V��>�A�`)�5��=�rI�{�ܓ�-�ͭhM4�y ��̀u�2�>��Xmq,��`b��޲�i���T�x�X	B�J|��@����2��V�$��I I�i��x�8��Ԇ�Z:=1�M\O�:�v���
����5��� }�\ �up���ם {���K5�ףZ��� 3����c�`u�2�;���$��35jn�FJNI(NK��u`}��X����W ��Ukbi���M�&�XyL�f:��:�����P�\�eUr��v����Fܩ)6�����W ��� ��H�~�%�Lm�,n�淯B�z�6����ܸ�9A��A]V:�rd�{5��� ~�Vq�V�S5D.��Ձ�f�S�21��K�{.�R7�4����\��jU��M����}ΐ����W ��̀}��Z�ްkF�x�d ���}��>� �� �ݵD�Y�V�z����}��>� �� >�I"�EH@0>���|M��`K���u����H�C���h��@/�1D�Y����9�F˫��gD:���+�!ִ�#"a)F�)��ɺ���*K�尚%(@$�KYy~�o�ύ�s��y�p�h�@)X�iH�U��JV%.�?i�bmJ)�,P���� 1ҫnڐ`��TӠKt�H�\4		Y���"Q�(*!	U�pC!��r!d��hI��-�@���~�ٙ������                  �                      �I���yn��{�8尘ys�s�`�n�\;YŔJ�ks�у�l%�[���W'5��n��N�����X��%�Y�C��AJ�K�@��]d[�4�0�A�{w��-`��;���b.Y7W1�qu���]�d��"%�LXy7%'ka�lUAPM�Q(t%�W�]d��Q����ig��(ؙYZ�%6�%vgm�z�Σj�fm��&D`,���l[vK��9;�Ҕ�\�����d,�-�f�Ըf܉U��P趪+b�U#����T�U8��tP�n%�5u�Z&�$� �z���PZvA�j�6کWdȘ#d�M]+0〞[
�n�{EU!h�����C�Jۙ�S3^Qp�[R��plu��:s��\0����m�Y�[ej��U{`G^�l�sZ�[������V�6��[Gm6ؐ��:$�a��e�*phn�9��u�m�o'�V�w"���;z�f�@yxf�Ju�:���BM�m�=t+ݻ#�(�vݸ\��m�S`kRq�����;/X�w!��V����m'���i �'c��4�[�eN�����2@�KҰ
�� �T���6����L`$�ni��U٭�s�]��i�lnhS�/r���)�J���gf���χ|u��p޻;�e`lV�e@�F�/mt!*�8Z�ٺ����i<��.�r�6�+�g��3���0�ݔ����tkю�x�Eu:v�Ն;a�7��3�w�%�rGd���P�q]E"J���Y���'GG��O4�v�M����=��
�iz㰛^'m��_ ���^�>��t仡��N^�&�W��['9ûe��P��!��λ�'�]XBx�������ٺ�"�[Ack�.;^�{���yS��ኇ�O��iQ���$^��|�)��~�sy��f`  hh  ]mX���f��t��u�u*�Ȼ.�t�ڙ�'nGXjc�&��m*���*&ή�b%Bwm��U��ӗ��A�L�6؛5�eyen�< ��n�;<�����݋���|-����ʵ��
LͰq���mH�ȍ'cE�[�O���X8n��9�ڦn$�= ��n,�9nnʥgK��Iz]����|��<��:�
Mg�W��ƅm��[mT��l�c���g��h#La��5�c���2}l��up�W ��Ukbi���M�i��ِ����d�>����RF,F�\��R2R�T ����Y�����ِ������Sp� wY��� ���;��j���M4�@>� [f@���wu� �mib�<�l�l�;jݷiWAc��v�:�� �p�V���[��sؑgt�Tc����d ���wY����ޭ��IE� � ���~�r뜥͢hP��DX,F��A�:�	%)(����V�;V[v�T%2wص�q�Q5LN��X��V��L�}m� >����J=ׯSF��<����{�`nnڰ�:��3��v������CO�ě��� ������l��Z�m�٭���h�tn���.�.�[f��\v�d5�]��qԺ��m�6�4L�;�$�����y�Ձ�n֥�����rvNkJp�!�Ĝ�{�u{�r�I�۫}�u`��^�W7+ti�㌌q�W9J��ݵ`?7j�Q�I��I �BJ҈�����V��VK�x֤э,և�i��ِ���/u� ��� �բ����u�K5�7���VRY��X��Xmڰ=?>} .Ƃ�;+Un�l��[gp�)�i��mW:x�s1�5�Ye�!�ǭ�u� u� �̀����J=ׯSF���Sp�ِ[f@wW ;�p^�ZX�7���m�M��ِ����\�d��TT�Z�1=y =�\ ��ٹ';�lܛ<�!)��s��L�U�{��8I��NK ��>� �̀wW �libU���І�rnn�l�S۠d�j�g�	s��c����l殜�y�Ff�m�;���� ���;�� �j�S��t�8IVs2����q �f� ��� ��̀{ʭ�ki�Ɩkb�V��V��Y��"g��7vՁ��j�4�^�z���n wZ�wY�[f@���}�R�u���ki�57 ��̀z�2 }�\ �7$��(� 0^���y������� h	   u���y���z��Mm���d�^�4�&&y�XuH�=���0<̗e�k�87���	i�D�Jv_����ݢ�l9��un�u#����ֺ#; ��F�i9��WS\l��Hf6@6���fpne&r-��p3C���c�НSms�oh�K��v��mk�$k���9n��0�R^��,ٝ1�|��<��y���wv�� %dDה�f7k��jM�kp[NޏgrFJ�@E�{�i�3m�)ta�$��߾��C����f@>� ��Em�OE�*�Xs_�#omXomXm�^�s����qj61J		Q�$�-��@>� [f@���we�ճ�4�ji�����d�l��up6���U,�ߪ�Ÿ'�9�t�8[��ِ����f@>� w߾�v4f��BV�m�K:s���Y��gv�&+�O�ΈyO�I�ٵ53tnmԉ��wW ��2�u� ��2����q�Q4H1:�I`{�˫|�*����ؑ�vd�ِ���z�Ԧ=�3F\���.fn|ؖ'ݾ�Sq,K���ND��*�MD���eMı,K����ND�,K�^ִ{YsZ�����&f��bX�'=�p�r%�bX��ײ��X�%�{��6��bX����Mı,K�ힺ��[�fjd�Y��ӑ,KĽ7ı,?�׽��m>�bX�~ى��%�b}�{�ӑ,K����/-#�kqkc�}]�A��n��Dv���q\v3d֭·5���;Fm��T�Kı/{�fӑ,K���ى��%�b}�{�ӑ,KĽ�*�V�S9H�fV��_q�N8�s6��bX�~ى��%�b}�{�ӑ,KĽ7ı,K����������ow���2,�/76�Q���%�b}�{�ӑ,KĽ7Ǉ!T�$�E�A(���Q���]��K�����Kİ}�l��Kı?���'�)-�������7���x�w^ʛ�bX�%�}��r%�bX?w�17İ?!5��~��r%�c��~���������w��7��b^��ͧ"X�%��}�q,K�����"X�%�{�{*n%�c��?~}�꫑x9�t�,��HMQ6N�ٛrggz�7]�����D[��zfL�h�Y�ND�,K�{f&�X�%����ND�,K���P�9Q,K���ٴ�Kİ}5kG��sSW5sXd��q,K���NC�uQ,K�k�T�Kı/�~��ND�,K�{f&�X�%�����W٩sֲ��5�m9ı,K���Sq,K���ND�,K�{f&�X�%��w�6��bX�%���^��	ȹVr��F�r���r�s~6��bX�~ى��%�bw���"X�+��(�SH r'7�\ʛ�bX�'�~�����]]f�S5�ӑ,K���ى��%�bw���"X�%�{�{*n%�bX����iȖ%�bzw�������u�PnWv�gC�\p6Z�SF��\:��T����=^}.���$$��6��^���"X�'�~��iȖ%�b^�^ʛ�bX�'}�p�r%�bX?{�17�q���~�/��d�����|�~oqı/{�eMı,K���m9ı,�혛�bX�'}�p�r%��r�����Q���btI"�Y�Q,K���m9ı,�혛�bX�'���m9ı,K���Sq,�#��W�ŉ��(�!crU�9J%�`��l��Kı;�{�ӑ,KĽ7İ?�@I�������|r��G)���\IJj5�I�&�X�%��{�6��bX�%�u쩸�%�b^��ͧ"X�%����q,KĨDP;���33330 ��-�  �Ҥ�\��0�v�����vy���T�w[v�D�sg����!��9v�rrg��ח����;�k;�a�m��%�q�U���$4���T1b�>U��sR{V�pԫu��\ �Ą��	�ed�ʪ��laU����i�mWa��7V������ �k`H�����4���f�<�w���p6�{������|��������e�7�"�ʓΞ��.�ۧ�at�{O]���֣BS��c��w�w���oq�ǻ��Sq,K��}�m9ı,����MD�,N����ӑ,K�Z���Q�D�)�I*�R9H�#�����r%�bX?{�17ı,O��p�r%�bX��ײ��X�%�ޞ�����]\�eˬ�r%�bX?{�17ı,O��p�r%�bX��ײ��X�%�����r%�bX�׽.�WZ�C5�0�f�Mı,K�{�6��bX�%�u쩸�%�bw��6��bX����Mı,K�g�_bR[OC�k�{�7���{��?_��q,K����m9ı,�혛�bX�'��p�r%�bX�	�粮��MrP��-xn	ŀ(Î�V�]���vbSV�\A�삀���3��ՙD�I���7�Nw�`�! ���&�z%�b^�^ʛ�bX�'>��ָe�3D̙�-��r%�bX?{�17�@�A��Ԋ;���'}��6��bX�%�u쩸�%�bwٟU�9[\��L�"����-��75��f��bX�'~��iȖ%�b^�^ʛ�bX�'{�p�r%�bR��˩ʳ��R9H�y��H�p�µ�fa��Kı/{�eMı,K���m9ı,�혛�bX��r�����|r��G)��j620r�ja�.fT�Kı;�{�ӑ,K���ى��%�b}�{�ӑ,KĽ7ı,N���ffff[tj5�2Tn�mt�z'in�������j�K�D���ݺ�vvܮK�Y)����w�{��7�����17ı,O��p�r%�bX��ײ��X�%����6��bX�{��~�!'t��xk�w��7���'���m9ı,K���Sq,KĽ｛ND�,K�{f&�X�%���e5���(�q�W���#��R�{�{*n%�bX����iȖ4R�dhr'�mW&݉�!��x�"@b��* ��.�dMv��Sd!�_�ָv��`�&�CZ��568@�d̹�۩�a�	 BjkA�+���lN:	�j����؆�N;8�1��ʑ�2���`�mx��$" B��iF����,4�f;R5Z��SD���MU�d�X��D��Ӣ�D�v��+�
P�#�C�
%>@p"Wb; 6�i_ �CoT���+������y�l��Kı=�{�ӑ,K��v�[ֳZ.F��tL�ʛ�bX�%�}��r%�bX?{�17ı,O��p�r%�`*�MD׽��Sq,K��V����GD���NK�|r��G�{f&�X�%����ND�,K��{*n%�bX����iȖ%�ow�������p%�7@�-�v�����ء]�����y��r;.1v���݉rk5��f��bX�'��p�r%�bX����Sq,Kľ���ȫ>���%��~ى��%�bw]������k&�Y�fa��Kı/�ײ��X�%��{�6��bX����Mı,K���m9ı,K�}g�S55����3%�ʛ�bX�'��p�r%�bX?{�17ı,O{���Kı/{�eMı,K�=�M^:��W3XjffND�,K�{f&�X�%����6��bX�%�u쩸�%��A�L4*���"�$Aҁ�7��o�ӑ,K7����p���s�xk�w��7����{�6��bX�%�u쩸�%�b}�{�ӑ,K���ى��%�w���}�/-G*�
1�ׁ�T����:<YZy��U�����y))-���fk0�r%�bX��ײ��X�%����ND�,K�{f�g"j%�b{���iȖ%�bvz����֋�֦5�ffT�Kı9�{�Ӑ�*�GQ5����17ı,N�߸m9ı,K���Sq,K����M�Q@��	#������#��R+��ى��%�b}���ӑ,KĽ7ı,K߽��r%�bX=��}�"ٛ�W^��oq�����w{��ӑ,Kľ��eMı,K��{6��bX����Mı,K��߯ՠe�qp�|�~oq����w��T�Kı/;�fӑ,K���ى��%�b}���ӑ,K���;��w�>��   ����  �۴Օ�rj`�ìk�9��iSm�$/9u��4G���z��Q�Ӓ�c\.�(,�5`�ݢ�d��8^��]=�NݗiV�ܵ�q&pI������N�͕����� �*�]&!�EVһ�:7
��x��=��s�.��\�,��ж�u�/b������ǧ'��wniW�32�Yn�{����{��� ���/V��%�1m��ٸ:ۛ�ۗ�����R�n���<��s1fd̗3*}ı,K�߽�ND�,K�{f&�X�%����6��bX�%�u쩸�%�b{�����32ۙ�4fk3iȖ%�`��l��Kı;���ӑ,KĽ7ı,K�{ٴ�O��MD�?k��ur�桚�Fc�f��bX�'���6��bX�%�u쩸�%�b^{�ͧ"X�"+�̺��9H�#��W{<�F�jh�&��iȖ%�b^�^ʛ�bX�%���r%�bX?{�17ı,N����Kı>���kY�.Z�d։��Sq,Kļ｛ND�,K�{f&�X�%��{�ND�,Jr���.U��r��G+���$�$�n6�s��2d�ln�l�}n��f���u�p��u�s��:�[��v�S���w���d�~��bn%�bX�w���Kı/{�eMı,K��m9ı�w�S�<}�"ٛ�W^��oq�X�w���<��(Ez�q7ľ�o*n%�bX��wٴ�Kİ~��bn%�bX���v��5��]f�E�a��Kı/{�eMı,K��m9ı,�혛�bX�'��m9ı,K�}u�sY����fMj\̩��%�b^w�ͧ"X�%����q,K�����"X�%�{�{*n%�bX���?~��������&fg�%�`��혛�bX�'��m9ı,K���Sq,KĽ��ͧ"X�%���~�٭�e5<�[�b۫v�IX��N����asv��@���a�HK� �zk�w��X�%�����iȖ%�b^�^ʛ�bX�%���m9ı,�혛�NR9H�gg��ԍ@��)�*�_�ı/{�eMı,K��{6��bX����Mı,K�w�6���'���{�t}�-<\.��ڨ�|�bX�%���m9ı,�혛�c���iZ"��"�D�2'"{���ND�,K�{_�Sq,Dr���|�7�EH�䎛r_+㔎%����q,K�����"X�%�{�{*n%�bX����iȖ!���~��{��s7:���7��������"X�%�{�{*n%�bX���iȖ%�`��l��K�:�:����*�+c�K�N�n����f��wN������{#��u�B39�.B��6��bX�%�u쩸�%�b^w�ͧ"X�%����q,K��{�ND�,K��]z��f���̲�\̩��%�b^w�ͧ"X�%����q,K��{�ND�,K���T�Kı=��jj�˫���2�3iȖ%�`��l��Kı9���ӑ,KĽ7ı,Kϻ��r%�bX��}ur�550��M3Z�q,K�����"X�%�{�{*n%�bX��wٴ�K���, H`�"��!"+' WH.������Kı>�:�d���Ok����{��7�����^ʛ�bX�%���m9ı,�혛�bX�'>�m9ı,O�;Ϗ��v;��V��;���+�fխv�M6(����uv�O<֑������Z&feND�,K��~ͧ"X�%����q,K�����"X�%�{�{*n%�bX�}��s.j���5��5���r%�bX?{�17ı,N{���Kı/{�eMı,K���6���A]T�Kڿ�t~�\���5��S3Mı,K����iȖ%�b^�^ʛ�bX�%�{��r%�bX?{�17ı,O��;uu�f���d�.��"X�%�{�{*n%�bX���iȖ%�`�����Kı9�{�ӑ,Kľ�{^��fj�Z��.��ʛ�bX�%�{��r%�bX?{=17ı,N{���Kı/{�eMı,K��O!چ��������}�   -�:@  s��,��Z@�1��m�آÛ�
Í��h�1��0n�8�h�ݝ�P{R�fņ�S��Jq�b.Z�^S��g]rvvf..�7/G�령n��@�%@S����Xr��n���ʒ��^;c����G2	��3�'jW��1���7q�z��z����ʜ>nvZ���b�-#�Y������.N��<��y�Qk�T�|�٭�d��e�u�+�SFv�[#� ��ܖ�;g�+;dN�D���s������5ۖk	��4K��'�%�`�g���Kı9�{�ӑ,KĽ7ı,K��ٴ�Kı=�����j��Y)�5�17ı,N{���Kı/{�eMı,K���m9ı,�����bX�'����j�j�f��fa��Kı/{�eMı,K���m9ı,�����bX�'=�p�r%�bX�N�o5�f���d�kT���7ı,K߻��r%�bX?{=17ı,N{���Kı/{�eMı,K�}u�d�&ja����fm9ı,�����bX�'=�p�r%�bX��ײ��X�%�{�}�ND�,K�U��{�eUP:�r����:Ѷ����n�<����N���	���1sN��4��Kı>���6��bX�%�u쩸�%�b^��fӑ,K����{�oq��������G�1I�^�"X�%�{�{*n �?M�"��

�-w�,K���ͧ"X�%�������bX�'=�p�r{��7����}�][-&T{�d�,K���6��bX���LMı,K��m9ı,K���Sq,K��ǽ���-��5��fӑ,K���鉸�%�bs���"X�%�{�{*n%�bX���iȆ��ow��}t3��ls������%�bs���"X�%�{�{*n%�bX���iȖ%�`�����K<�<�<�>}� :��
�))��7L[<t�E3��[�m�6��[ss<�ͭf��5��ӑ,KĽ7ı,K��ٴ�Kİ~�zbn%�bX����iȖ%�b};}�ֵ�&Y�u�K��Sq,KĽ�}�ND�,K�g�&�X�%��{�6��bX�%�u쩸�%�b}�o��̗$�Lɬ�hֳ3iȖ%�`�����Kı9���ӑ,U� ����.{_���X�%�}�~ͧ"X�{���C�����]7Zm{�oq��K��m9ı,K���Sq,KĽ��ͧ"X�%����q,K��gn���d�j�5��0�r%�bX��ײ��X�%�{�}�ND�,K�g�&�X�%��w�6��bX������w����伴�J�[����X�*[���֎�j�l�����qjR�F�f�$�hLRE���#��R9K=�/�"X�%����q,K���ND�,K���T�Kı=�O{&��Ku�k.��ͧ"X�%����q,K���ND�,K���T�Kı/~�iȖ%�b{]��ˬ�3-��ML�d��Kı9���ӑ,KĽ7ı,K߻��r%�bX?{=17ı,Ow:j�5��h�5fh���6��bX�%�u쩸�%�b^��fӑ,K���鉸�%�@��趐dR0$@O�M �߷ύ�"X�{����O��Y�Y�pqT{�oq��%�{�}�ND�,K�{x��bX�'=�p�r%�bX��ײ��X�r���ʮws�J�IM7I2&�$ #;g��[D�6���6y��cmq���ځ�¢-bd���nI�+�)�r�\���U��ı9���ӑ,KĽ7ı,K߻��r%�bX=��=�55��a������%�bs���!�#���b_{_���X�%�}�~ͧ"X�%����Mı,K�흺����Y�d֋��iȖ%�b_��eMı,K���6��bX����7ı,N{���Kı/��׭�d�&��Lչ�Sq,K?5^�fӑ,K��oq,K���ND�,K��{*n%�bX��'��Xk%��5�K��ND�,K��x��bX����� �'ݾ��I�}�sbH$���
��ET�
/��(����PU�*���������
��ET�_��H�@�DP*T��E `	@�DPT��E `�@�P(�T��@E bDP 0T����P AP
DTX((
�PU�*���ં��UAV��
�AU_�T�PU�`UAW��U_�T�PU�PU���d�Md�n�L:Of�A@��̟\��� (�PWv T Zt   s�
 ҴGG@>�  z� � P �R)" BT%J��UP�����T(�QB�IB@)$*IB�UU**@)  
���   C  �   E��/������u��-�7]��� �R��7�o ;3�Pw}�E� ���Wy����   +��u��n�� =���ֆ�n�
{�@�:�T{��z�M*��s �w-҅  �x@   �� 4�
           9�       � U*��r�UX{�7-����z��:���C� P�J���_|�< �[�m彴���}�ʜ��W��v���gR���W� )�yS����uNN�W&�|��
 
  @lZ{�������[�|�����ʽ�� =��]��ݾ���rs���M�����S��� ���׭������ �Je�ھ�mvӖWy���ϏA�@������      + �Jn�^�_-��^m�[�)}� �)\�_O^m^������}� Oz}.����O'� w^-�i�*w�@ܯm��W��;�]�nz����y@*�����K�]���t�9_ ��  �   � ���f�}wKź����;��k}��=^ۓ����彼ۥ���6��@P�*X���y=x  �<��{���+�@y����t�Y�۟y����5+� �>����m�w:˓\������ ����T�(0� ���j<�J� 4hb'�UR��Ri�  ��U*M�J�  "~���IR�	� �$�R�" 3S�O������?��<��'��j��������{n;?�A@U�`nr��A@Uآ��� �*��@U�����( ����ڟIӎ�cI�#�'ӎ�4���c��5��bke�"�KO'f�;���|ه���¶m�N�?҇��(�`�N���-FX{�tj;�g��s���a��:	1$	4�e�����j�g��#��kuǐf��`{��޹�q���JI��X����!�= ^,U�.�����EQC20�1�3���h��מ����BL��l�f�FY�;���K4��>�v)uq]%˓���j��\���H`��F34�O���U��~�D���C�gaa�7(�)N���.�T�9
S�P�w�N�g��<,�Ґ�8����3K9��E��,Ѹ�F��b�����akNi-6ŧ���y��,.����p�#($��b ��Ԍ �~�����,��dR
(�&.c}����.g���Rp!!�X�0Č0c
'?p\���n��}������q��aȻ�ф�����7\DD���ƪ�ej6	i3(4p�~�e�ٟ�n2)�C �IĀ��`1"���!�*"	�"q�̮s������dm�
g	H���#2+�񃆢��J�ٳ?s�<-odE�4�l4j#ٯ9k\�ɢ����-	�Ijip��4da��,3Ph5�y�o����I8��`i!�H�eXh�Y9�F�������y�ՄˌL�����%���ߜ6^��yh�@��g�ƒ7���o��PT[3+R�N�f	�HcN�**bIr�Q		P���Վr���s#MQF19F:x�f���p�k��O�y���[.�K�0��d#[3�y�<���_��q�~&�a��I,�d�,�q�o^w�������'��7�S����x�8C3�@��8I���5,FVfk��v�����/�x�D�C+��<gD,�>�N�g�$pV ��՞��~kx��x٭���[�XE��s,��o�\�~�7�+�8Ic.��[y���Ǉ��f28N��p���f	�$"b��1�s=H�s��<�F�cD������8,A$���p�Ç�~<�f~��-6Q:I�p2LȒ�j+E�s8y���4��De��A@fh-l+{���k�ټ�T�ݾ�!RTR��§�Ev�
vo#�H<������se�A�w5���^=����8Qx�#Ș�121�v��	Z��@{�dz����1�)ɽO�md!��m���q����7�{�����Wg;�˻/������`0�g�b`���Z����3�~�Ќ�ۆ���"�WC���T���s�o�������9��^k�Y�a���a�����Ƣ#)�Uj��pߞg癣�4n0c�F1�!��8����U�SA3���Ɍ
MF�������xh.��ǉ'p��Aa�l�Ռg�Q�CLa��i{���ڜLI���FPh�8��6s�<F�xo���Иt���X�2�f���6��,0��$p����<4!������,tX���0��y�����`1IL�ӽ�f�g�����#��~C��B�I�,6�|�5��&Tk{x��x���l�q=�Q�3��%���I��$` ��&7$FI�o7���Ya��g<6��|=H�В�N,��q�o����h����1�`m9����l'(���z�C�u�~�=�������ٞ��#4`l'���6P�o����[x�80���Ȑ�<q@�8�M���oY����<��C�u*�v�W.J"R�%7;TU�|���|QT�P�JY���}���h�J��{гڧ7U		{��)�Mr;�E,�I�I�O�E~��^�ט��88CcNCkZ߼����a���"4:18�����+^sa��l�m8���	#C���D�aY��g�~֓�����b4��t�m)?����3�_5�"�Z��EqW
L�N�2YEp��2�r*�Ճ�;B��*�'߫��ITPA�di��y����9�X�����j�G��N`X��+[��1Ix��y�2ty�i5p՚�`U�5yA�z<�[4$NFd��f��E5G%���#�R'%Ԫ����|N�C���%��3�Q����a�1<�p��;�ׅ�[3���5�x�| ��Hc�%�GYF�oÞ�v{{a�JA��j�Xoy����pe	dqH�8<�1��=<8p�4l�Ã	)'�xJ�N�<��q�'����k|��pj3A��Á$��#&-k��g��^�7��&f�����ddg���Z`�d����ә�Zߞ�<_kar0�cF!���"*��p�<^\1�	�d=�o�v��&��#�"��B!R��u���4�㽡p��c1�$\��_I�ê����Tw]	˺���S�~�����m';,4���>�$���Y��3�fo�s�h	Ҕ�Y6���B�\+(N��uÊ����aޏ�9�vo�`[Q�����=c�p��B���JO_�� ����M\;�����'c,H��x:���Z��0�᧓�o�͛�����$��廹�M���1Ӱ�q�5��?yǇ�sds[�F:I-�<$��a����4o�k�8�#�v��]��*���J�W�WUA.� �����l�f�2�a�*���2�C�ֽ,{q��I`�k|���O=<8A��`6<"'�y�#5�xs{6x�gC`U�Ѹ�s0����3��bX�L�q������N(A�����m��6��}Q�zO���� �0�201�F6)�����Pn��P��'N�J���c�ے�UU�!f�޵;>f��w���2q&:m��kG|��l>k~�1����#X�Lj04�$a�1��a��GQ�q)��d���d�=��F��G{��g�4[�G[S*p� �	BJ�^��<x�:�a���u9�í�����[��Y���\���*1�$$_�!M^H�&��p,­i�SY�m�Df���Y�6i�!��4��$1a 	f&"L�1��	�ռ�[Y,cʜ��{��������1��$���g3��h���x�#)$,�mB3f����Nh�������K�Y}��Xd�cl`Op7���ob��o�p������u٭�G�߁f���6Nkl�3�������2�I1
�R� K$�HH���21� �03�C��5k~�s�,޶������~�������f����0�dt�`HC"AsΗ;��d�F�d�c4412RAPI2�d�)�A����ָ��vXoz��׻y&om���h�8`X0��q#֌
�^v���$Q\����p�#J20f��0#H�Q�F������yh�1�4r&�
�I���A:86k�'��~��#=H����F0b�Fg�Ћ��y�ى�G<���s�T�?{0�^���'���@��^YĎ�S�L�2�HJW??�o�~?=�f���M�p���:g���Q&^zsV�ݞK>�e�7�&?��{�o��I�����	���Xi�ׁC���h�K1$��3Df�Y��kda���[��НD�
��LN�.�U(\���2r1�0׾o���X�����[*G(s�:��ﯓ��N���1t�0L#I��{�[��k�{��=vaf��k�ڈf&��d�H�L��ܿg?F�е�M�Z�޺���0��`�	)�F3$�0L�8Ph��?U.���,*�o]�g|�K��0a��g�ᤜ��[�I��i,Ӥ�.�4�%�{����p`i�0�!R@b;�Б.ĂHe6����!!Qn��pR+!!I2�),��RB  t��?6:e��' �4%(l$0�&�JBD���B 0��<p����#&h���cf`���H	GH�:H0a���k=���{ -�          �     �� l �               P|                                        l  ��     @        �  hm�  ��  8m��s�v8+��6��]�OL�k]#��4m�)dѹ+	�N뱵�=v�E�\kԖ]��탆۰  i��h�l�6�v�m��-�� N�m�8�m�@ ��j�wa! m�   �b�t��Z6ٓ�[Np�퀐�`�4kd��l@ �cv	�]h �n�ۍ� �u�Xћl��q!��K_ͭ�'�	 �r6�+�WQo1��xd��95
�Ԟ�]*�����r�J���X���e\��N�Y-�{hpmHڹhrE���uK�:;"�l ph��ݳil[dt���g��U���f�gm��CiY� $5�',� ���W�DnL�]�iV�:��)��t� ����3l�� �   4��0��Oe�Y@2��5�eB�ul�J��	m���m�v -�6�&۲���@��<%�bW���@kj��m�کW�m���GW@[@Iz락��ޢA (-&�w:饗m��(��h��6�6��mUS�*�Gڌd:p �6����:r=�׀�v��]"2Y� m4Q���Fٶ��� l  �N  �ϟ�m�ͭ�i�[-�n  ��d[L�� q�kn   �� �`��m^�����r�A��!*�-TUJ�X�U^j���jZ��U������*˲�mP K�I�pl� I �+j,��Me\V���YvL�[lH���A6�l��l�  �U���q�V�Wi"k*sQG�*�����Y�~�P�W) sR��VΊU���S�+mW]bs�'B�i �	�ᮮ�z�	�i6�/I!��5 ���՜[q�Z���-��  �����G �PqUU.��=���ZzҬR�UUp���K,�դm��]�U��G"���ڪ�V�l   6�	�,�dڋhm�m�rNE^Tl�-�A�Mpv�-d�'M�M�f t�]�9�����ŴA6�5Z�@���*�M�Թb�� l� m&� k[j�6�I�l�v&�$�KN��Y� 7m�צ�A�W�;:Upq�p[,G�<��M�ڑJ[%&�6���T�@�ܸBg��)-����t�j��&e���eݵ�[)�+�m�-�8[`�m�t��U�Tj-�<h�L���p ��u��  hh6�� ���ެ� � ��6ۥ��A!;k� X[Vʠ� �*�pWAKW�  շ6�N��Izm%�\�U� lmu
몶�ې�2R����� m�,� m�  �j�u��B@$��/N`��� 6�  [@ �   ݻm�e�` [@�h
��>���Uz�pH �[p���5��&�%���IAz� 8m� zնN�J $��8 � H�H�6�n�[Gf��qضx��6����@��m      �� ��    �oU��Z��m��  � �i6-��x-��Ժm�i; E�ښ鎓�-0R��޲6���J�J���TpK��m sRީHr�N��rf�#<�U*��mP3mm���8 m� p��[@� 8� [B�#m��H��  �   H     ˭�  H	      �`�`6ض� 둚[���Z4�WT�R��KĀԥUV�T�Y�Kʹ� f�`�hh ���  H  l  [@m�r@ 8l�$i�Ŵ~�����0      �#]�`ZץCe��v�$� �J6� �  o�||��`[Am�8     �L��,6�[p m��ON�vlt�kS�}q�����&�㎕�]+��t�K��cqz�[:�-m�'G&� m��m@UJ�ڶ7Gh]���Pm����l rͶ�׬�l^�K� ѭIm��J�3M�D$��� �Ŵ h�/[\��"@pi���iR�t�$�n���+�夑+�6[@��� S����BK�@���黬�.�m�:��]4� H-ĢM��^$�"I�UV�+�i�^���@� ����o���k�"3I�ma�  ֻI�6ݶ� �ne�"������R^�{vi�IR��
� �/U�U//T��R��ln��qR�ʪ�ʰ�FAl�h�,kMv�4����|�|Xz�Y$D���Λm�� 	lf^ 6ٷlH�Ci�����À86ڦ��bC�6��8�H�CN�t�j�f�k��:A���H -�H[V�pm�	/Zm��!�]+e��H�ݲ(�K��ɣ�m M�[��UN��d6*㴝5�����7RT�m j�Vl  �����`� [\��     k�� 	k3$ �Б������8W�ڽt�  8 ��	��km&[@qD+u���G/OS�m���p���n�*+�T9� 8�h���&�ۄ� m���l���:�z�V�VV�u4��'m�4P�v   m�lrt��	[Ԑ6�6�J[$�ڃ�� 	m�U	��粈\���c�r����	ÈZ�V�H�I��֛i�	 	,]�L�Q��8��6� � �[r�ky�[Ikm#]<��6�E����.�d�bv���`8�2�(�� ���n庀�� rI�m��|��#��gUUr�:�<+ 5V������-b���չ�L`܋h$ٲ��`�U�(��o����
��5��U�hm��@Y��U�`��6�k|�o:�6��˴T�1@BC@Um�'g��,@�J���~��- �T �UJ�R�!��]Q@[u/1TT�iV��"K�:�,�	�&�� H�w[�AN���!�M�I6��`i��kN�l� h��J�Z�/PK)]�����_�@h��fv�YZy��/%ʻ-V�;�rFٷ6��u-���  �si,��I���ƀ�*ԉ��ݥZ�	�F�[]{M���`��-��&��n�   � �v�ͷkM��y��� .���h
UU�nZ�S��� �am� 6�ک���m��dب8�vUP�]5���m���R�U�R��@����PN�]�������A�-�m�b�W ��I5]U/(U@W�Ҵ�I�K(������
��
�]%����E��d� ���ֱ��倶�v����b���첶�5�۬	�8^t$さJ ��Z�l���25��ٺ	�*K�tm�ӜmtHpm���m�+,jj�8eh&�m[7 5���L [d.���8��\ s�@�]�n�v��n $H�m�@,�U��plV�[d 2�[���%o^�lr�U�SV�J�KUm������n�=�7c�=*�V;����E��,����Y@�ݩ^GkΌ��Q�)�Ͳ��
�A%6�茛��A�0ixt�'`���GJ5�9�u6Y�NL$�u۴�tu[o gJ
�K�3d��^:�����7>oI߯����B�T�D��פ��Ĭ��Ke%vZ%R��o���I�֔��&��qZ�X(�H��w�(+γ�~����l�\���Ua�@]t9ٺ���;Uv/H 4�b�ӡ���[aƶFl�N�]��`R[GF�C�uڥ��c$UR�l�UV�)(T��H-�ed��hM�{v��`m�q5��5�F�6�Zm�y�R]{��[@6݀�%�"ޠ7� �YV���fĜ+f��o��32q�� 7;> ����m�@ m� ;7���z�����;�͚��Է6�KP��N��   �v�vۚ���  -�����&�훶[@    o�^�b��` m��[ۭ�8 ��6�̀ ��u���vZ�[d�2kkYwa&�l  m�6�6� UUUV,e��Px ��ؕ���뱶9v|Eaqv�UVʵ*���ب(�m�b� �v���m��mn���Ns ����406�����֢�6` k�ZR�gm�F��ܠf��O4#J�؎���m{9P�4�.J0��VoӗVն�ݠ-�az� m�/ 6��b\  6��"�uUv� �shiv�{B�ʦ���T\�]�e;`v�@p��In�- �`ݠ*��؞nlS��E,��-.�5���_U�v�Ķ$ �۳7�of̲����"*J��Pd�	�'�%��
�����Q�U�R 6�!���N(���G��*���_�O ��� ��uCb��Tt��P��B^��:(���}N"'�=���_M/\��>��m_G���mD����C���=Č?�Q�	�?*��D�"U=WO="@�����P��@H!�࿀Gc�m�_�E���;��Ε���������C�� CJ���R4'�D<@��'�T��z>Q����UCjpEzc�A��Ht"��8b�΄�
��'�ۂ���C� ��=�QOC�B`� 	D`=�z=�:�0���~T|TE��:���[�))�Шxi�����|? :Ȉ�EOP�TD0�G���I0O��A҂�� ���]��	�IRJs`1�UA<"���7J J@J�  ����<}g�p
c���[D:;TCH�T��?ꀠ*�G�HU��P��b�.)*�*h�,T���A3���k_���  �  �       ��  8$��������[h�T*\�Wjv�IUmc�m��W>��m½��7PI����N���抣�u3�X7;B���b=J�g�&7
���J+�n`�4�z�s����b���XDX�&���7j�Wec�r D� U��lR�Xu�^��8[�����Uz�����_�P��b�7[n�k���k���U*�[Fm�1j1��n��S��Ɠa��כ�⴦�It2HVͬ]v�=n��8�8;c�gfZ�;o&3OijS����������H\zT�q�jU�en5!ujjU�a�L���@Wg�U|DL��m�KUP ��i"ȭ�3=�2��y�y�q�0���V��+�6u�b����P�n59^�-��o`��m@/)U�A�@WlY|�N퉵�p��Y飚��шs(V1��,�<���{��]��vyR�9q���Z�<Ս���yR|���[Xn�S=:V��mәz6��ϣ"���֊�����B��J�a�mP��n�$��OV���Ԍ�Tn�'�Z�3�N�J�g�����]�9����<�\���aR�1ہ᛺�6��'��(��2����ag�3cHy��arX.��7H���:����'ە�x��-ַ(�۷+�vL���@,:�'EU'R��N�C�v[�M�,��jıeS�]6��r6�m���i�F�;<�f�okv{hC��,D�Sj�7cx:E���ɘ���n8��`�*�,��+�0NnW]=l>�rmV�����h�Lkcp��9''gd<A�s�݈9��3҈d۬F��M�h�9f�N�n��l�3m�6�m4� �pLnJ���-mn�[6�0�n�)�W�]<���tn�`Q�۶��m{&��ѝ�ԭ��6Z��^G\������W3�]*���o����(l}O_� ��O�!�T6�� hz�3� ���
/� Ў	�t�~��dU�����n^�h�f&�j����<��Vų��8���:C�q�L�I�/%]ݎ	��<7&����͚v3f��Sr�p�3�LܨY�V
R��vs��k��I�g#�n����x힕�ld���ҝ��Ʈ�׳�N��HR8:"!ݹ�m�S���\�qn^�uAvg�5��:F�Y�I����סx�
�g��SK��6xkYh����Y�V�wc�<x;s��ϗvLvq����t�j�	�$�q�C�y���!���������6�0�Y��x��f��h�$�XZ���˪�;������
7�7}�`Yk��-L.с�ş�J�M�f�,��떦�h�$�X���jF���QM�Vu�q�0u���� �8Q	6[���j�7Y�eNR;8�
�>tۄ�� �]��U�Z��pi�`�!4'	�R/���x`[�-|`z婁Q�˙uf�R�pu7f n�y�=	�P�D,Y����s�-�|`vd��e�0:�NJ�T!�!q��,�۫��U���U�fn�:mrA7$A��U��M� ��� n�x����w4+�:r6�R�RN+q� �ݖ��X�78B�J骞�5*��Ѷŷ���gf!N3��u�2n����[�N�Ϟ���©I���DM��QH��~�,��Ձ�{���y��Ś&��� ��7u�}k��-L2T�$�_��r�Ď�T���J)�*��?yX��rP��UCe�1	P00D�X�C����*���Ձ���I�9%QQ�"�:���Ku��Z����S���2����g7�j���%����|`z婁��������		�V�C.h�y��cr<�����ӻ[dz�۬z�wcFnB�s��/ۆf�޵�떦���%��ޙFܐM�ܒ���W�R�2l�u`_u`��Xz�n�Wq�������w5��u���%��]X��+ ��KV��l, ��V��ŀy�s���P���Д|�Bĕl��`}���2ՖH���d��\�0:����[�m���ڮ4鹇0�Au��j���q�2Og�Ps�-Ӈ��.���⶯d8CLw�9����Z�R\`E-��u��Ձ���K���r���X.�����\�0*9y3.�Ks�6檮�u��>��XtBS;��8�o���++5:��s�\�nKs���_���>�0:�.0"���p�wDܑQM�*���`z������[�;���X���6�nԤ��I$�D�on��]"�2Nw�B-s��ӝ"�Y}=gtO-��9ծ������Źkc�����{�^ٸ �<&�0 �Xy2j�ْ��dnyU�����Ps��+f�T:���W���]�j�n2�nU���v�T���թ�!��h-q�����-�G3�<�(�G�3O�;url� Ѻ�l{[��w,_��{���~�������i{g3��6�wsO���v��o�L�
ܽ�:�u	H)'�b�y��u�w6����`uv�վ�l,�}�0;�_�j`uz\`E(�9��^i�ᛸ��|`z婁��q��7]��cJ���R�E9%X~�qg���_�������Wwxo��p���������[��W�u����*���)Bq��P�P���#�%rvzsu)̋��Q�0���q^�!붊�dm�EJ���V����sn�:nz!B��=;�X�M>�W$�q6;5�o\���{ß���B�,����e�@꘮�Y�o�ʼ���V,�w�i�z�i�QJ9*��?|�^�Kq��J���p��[�UpD�\�r������/��{^+��U�w�,���Dm��dq�������|`z婁��q�=˜�.WQ��7cl�E���<b��z���r0��\\Ptݹ\/;$�X�٧�Ҕ��{ݯ%)O��{�R������y)J{���┥'�����]��0�j�����?w]�qJR���{��)�{��R���{ݯ%)N��{����[u���y���)<�w�JR��8�1CP��{ݯ%)O{�{�R������Z��kz#anֵ�%)Os��\R������y)J~��┥'���C�JS̏O{�7�Zّ��k[��)?~��^JR����8�)I�����R��=�uŠ�(9XWV1�Pr�8��R��ɥ��M�L�qP��FƧ�5���0
�d��gf(QޫyVo[��R���w��)JO/�����{�)JR~��v���:�
�7sUpD�\�B��<�(��d2S�߾��)=��my)J~�79�D)��
7Q/���䪪����z%)O����qJR���{��)�M�D �A��Ҍ"D-�d�P���ݻ,����)JR~��v���?w]�qJR���{��Ǌ b�}@��k}��):קu�s[�kF�v���)���s�R�(��������s�}�)JR~��v�������(N4�mDR�(��bp�c�n˳=�WfTKg\J�h��z�9'oH[C��a��{�)JRy~�t<��=�{�qJR���{��)���s�R���kj��T͂��*��F"ηYR���{ݯ%)O��{�R������y)Jy���sF��[21٭kz┥'���k�JS�u���)<�w�Q�B����D �A	飛.�j跕f���%)O��{�R������y)J{���┥'��ݯ%)ON�f�h���i�ʌ��8�)I����R��{�~�\R�������)�����)JO�x@�V �{�7�Z� 跷B�M�n�:$�*Eƽ=!1�Y]�K�.�Wc���j^0�r�$�.{n-��lN�"f����D��O��ݯ�+c��ݒ�:ۋH�2{^�)���\&���]��
�wh��4.6�����Ǐ:���Wl�G^�͚;5�ٷnɨn+m��6��S�]���ms�lr���]��z������[J��yTU_*���_1�M � ��Q�#j����g?�*;7n�[�m��u\�KQ��b����J��
.��x�A���VD �T�{�v���?w^�8�)I����R��?v�h�Z�ڲ�-oz┥'��ݯ%)O�׽�)JRy{�t<��=��)I��Otew[�֍�o{^JR���{�R������y)J{���qJR��}�ג��F���w{-�������R��^��%)Os�{�)JRy���R���{�┠B`�mU9����"���Q�B����\R����{��)�����)J�|fk�Y�Ps��֩�9�9*8�hH�ɻe7:�dMdY\�j5��k��h��Ύ˜��;�h�YovF;5�o\R����{��)���s�R��^��'��JZվ�r����{M<�Pm8Ȓ���JS�u�� ��=?���6�~1ԥ'�=��s����)<���y)Jzw�7�-l޵�{g3{�)JRy{�t<��=��)I��k�JS�u�s�R�>����f%UUWJ>"D';�Y�!Ry���R���{�┥'���C�JS���5�Uk��j�0���R��{�v���?w]�qJR���{��"ηY�!/�#ɾ�h����jԠob6���K�	�{]�ځ֍��y.x����ܔr�GRd)I9ώr�������R��^��%)Os��\R������Y�Ps��)�I�N8p��_������y)J{���┥'��ݯ%)O��{�S�1JO���k_f���v���y)Jw;��┥'��ݯ$$:+��FaN"D��㉡�V`~"�6�1b1�~l6oHe�32�:�i��	�
z`�t�W��	<��=	FZ���.��3��h&[�zka���G���� �4�c�6����g�A�K6či#|3[ %L5,٣���St�i7f�mkҭ�:�Б�p�Km�@lv��F�c�l ��O1L0,4#��`�C7�4:}Sb�{��ozq(o߅�ʔc��D1l���	����B�qǑ�x�<�3 �������p�	n�{��@��J��|
l�,d��68p������:�l:�<��ҁ��"�LM���	��C�`d�����R����~��R��#���fe��e5�o\R��$�����)����┥'���C�J�@���{��|�9A�����"��q�$99�JR����8�)G���~��)Jv_udB���w�B���;)U�,["뇧�@�c�]��;.��wN�[���lp�(<��s�᝛�z�x�����<���JR��)I��c�����	��ߧ"D Q�'���0)UUPej޷��R��w��?�%)?w�my)J{���8�)I����R��=�Y!*���r���f�r�%)���s�S�@d����%)N�A��5N��R(�M��`�|������)JR~�ߴ<��=�{�qJC�/��)
�A���̓}���)��k�k?�f�ncz���)JRy{�t<��$?��O�~��s=�ӕ�}����t;������jev��Tgj���s�23\z�Wu=.�~{�*6�6���G$U��9A�V����);���R������\��]��*0�A��i�U�̗d�
�V��)JRw�{��|Hd��}�8�)I����<��=�{�qO�1JN�}W�!n2$�''9g9A�V{޻�(8�����$>X�N�~�\R�����k�JSӾ��굳3z7�淾)K�A�}�}�%)N�~�\R����k�J��߾��)JP�����������j�Y���|��;���qJR��_�L���k�R�����8�)I����{���O{����w��ߍf� i,LPSS�'gVm��q�:nŠ3[0� �Yx�ۉ'�H��=���K2�#f�����asZ�����q��讂��R�g���R��5���tjݻU�������d�,��z�f���77i�.�Я{`�kn^�e�{��`�,�=<�rvN������(<RӺ�t�)ݱ���Y�B<j�t��9R�;!Z+i۽�={�]�;������[��C�J�q-v������{=[�dv8xՄ���e����5�1�Y��VQ���┥'��my)J~��┥'g{��y)Jw;��┥'�3�+���V�7��%*!y�s�."H��g�Ta�!9}ՊR�����y)Jw�k��ֻ�6�s��{�)JRw�w�<��=�{�qJ��R}��ג�����qJR��X��ڎ��#�*��9X���JR���ݯ%)O�׽�)JRw��U�9�r�H��r!"A*Sn;�R�����y)@>����)JR}�}�%)Os��\R������y�э���Q��(������9���&��]����o;�Zܔt�:hk��R���w��)JN����$d�s�}�?�]�R}��ג�����_�EX]ʺDL��D �A	�[�,�@]@�|���}ϵ�)JO���^JR����8��"�kJP��/߿�ȅA`��W>9�r�/�����%);���C�2Sߵ���)JO���Q�B�i��R5MYD�����T�!I�~�k�JSߵ���)JN���%(>V^�}�)JR~=��>�����F���%)O��{�R���~�}����s�}�)JRw��o,�(9���s��MoҤ�ڐB#�pGe�cF��lV@�e����WD�e8�ק4��/�{���$��S�*8�]�(9�W�/ߕr�)Os��\R�������JU�O�"D ��!~R5�U�j��J�
���x>JR��~�\�rR����ג���k�g�)?w;�I��Ò��t�}��̷���٭kz┥'{��^JR���{�R� �b��P	HH N�B�,(��A<>\$���ʌ"D-�A�����U�UoV�2���ג��	����┥'�g�`�R��=�u�(O�$�~�k�JS��3j��7�xNf��R�����py)@|�=�~�\R���~�k�JS�u���)?�{Z�3_j�q�n�b�ۧ�<�`ID����pL�kcד�4�iJ������R��pLUt6�U�8����渥)I��ג������˒����}��JR�߬�+Y�|�Y�f��qJR��{ݯ#��LCR�����qJR�������JS�����P�R���fe���{�,5�����=�_}�R�����py!�)�}Ց"Bo��0�A��[35N��5���y����D�$����JR������)I��ג��_�J*��"C�;N/Ș��|�8�)I�];�}��f�[�7�����JS�����(�'������kﳊR�����%)O�������,$'���&�4Z^:�ō�[e���ݺ�c��=zǣN-�\ܟ�=���� +(٭kz��)I����^JR����8�)I����|7���s�}�)JS^½�M8� "�s�s��w^����}�ǒ��s�}�)J-��#\�D&���*ɺ��D���R������R��=�u�)��pI����^JR�����qJR���-���
.�V ���?!B��߫!)JN�ﶼ��?w]�qJ�P�!M����Ta�!w�fDT��e����\R�����k�J�P?��s��8�)I������)�{��R�� jE)�JO��n�Z� GCiQ�v�Y�Ψ�v2b��2h�v6‽:���sm֞��٫�5lQ���%�a����m�dL����X���.�s�6���[�����%W^:;؈�A��7 �F�a�'7 >�.��������p�X�g��z��[rp.�;r��.S�8�rz�=�m����Zp%t[�8��:E۲�1�ه$l�kY�5�DO�U:��럍kF��٪��a���Yu��%�Y::����q�u�y�Rt�z䭟�{}�,g�x�;������e?k���)JO��������{��K�����my)J}�k�����y������R��������d�s�}�)JRw߾��R���w��>K���z�+[�M(��*��������)I���k��c%/~��┥'�g~��)�����ffovYF�k[���@ �;��my)J^���┥'�������:}Ց"B�q�5*mUU�\�sw��)~�{�)JQ���߰|��;���qJR����ג��y���V��6g�[=�z��N�����<��n���Dsú�5������-�ś��k7���)I��߰y)J{���┥'��ݏ���){��o�R�>�'��찢�eb*��T|D �N_ud%ǿ��+��@�8�D+���lP8��4�R�~y�ג���߾��)?w=�$�"�Ē���e�2)��Ȅ!=��%)K�{��J~ 2O~����JS�߾��)<�Y�g�k;��a�޷��|�&{��o�R����������{�)B|�I�~�k�JS�9��W"�HV���"D ��:�<��>'���k�R���ﶼ��G�w�"B��sh�����.��5��V��)�3u,�"uĽA�i�6���9U�V��Ҏ�AD$qW>9�r�o���)I���k�JR���|�\�[��Ta�!yHӞ��37d�
�k[��)=���y2){�~��)=�;�%)Os�{�)�b��v>�)�DRNr�r���=���P)I���py!�"��?�@.� ڠpv�G����7���)JR{���ג���}3��Zݙ��DY��R��'�g~��)����)JOw�^JP|�w��JR���w��5F��a�ֵ���)Jw=��qJR��g�����JR����(!yιQ�B���:N��j�7vt�[f�gK�0d��-u��n�X趝���.+q;/��[ݖ�\7�#5���)JN����������|R��������y)Jw߷��)JOޖfe�ֳ���F����JR��{�����������}�\R����u�y'�C��{�f}��ٖ��[���)JO~����JS���n)O��� �>�����)w���|R"Bh<������-,���D �P��~���);��my)J_���P�O�Rz �fl}D4�𡬓�3��JR�2�?��f���첍����)JOw�^JP¨ ������)JN�g��<��=��K�(9�W�b�7��FF�PJU��k��a�0�N��z����� .�gDw���AR	�WM��R�)'9��Ps��~�p�)?w=�%)O}��p>D�%���!Bk��ʢ��V\�&n�R�������"Hd�{����)I�~�k�JS�u���D3��_R��EбUW*>"D.���┥'��ݯ$?�X�O~��g�)=�;�%)K���a��]uf̍o{��/�!����my)Jw�_���)JO��{��J�C�r#��ߌ�A��Lʞ*����*�u{^JR����8�)G��)����Ҕ��o�┥'��ݯ%(E4�:����d�"h݆��Z�/c�9sW���FwF��y�~I	$V��/�A��� ��$2�sl��W�Ú�&���Lm�S�ku$�pc/@޴�;C���J)���akI$o1v�F�+�s,ӈ�:3Z!3F��[,�3D���4l�sZ049��b٠��9����5f�0�	���BafXS�P���	���24������� �?HH�`HD�N��'�.f��"1!�����~�����zu��~��� u���            [@������6������-vHmG5��,
��p�9�çYI��wc�lx�<g��d����T�+kM����aɄl	�,��_lJ��}�~���c��9��s���oY�A�Y��5>�����ּ�����[q1|]�v1�on���m�u۱U*�D
�J*��"Ӷ��,*�rtpN�� g�v�w'IKXںn0qD��6I�px�i�B������Xʹ�����˒���僌¤gm�c]t�<;z��5ֻ��^9�,�Jt�E�v^ݱ���=����p*�6� )enpn�U*�T!��*�����
]�g�z���b���BZ�5dU���G(q<lq��r�p2�;/0 �]�v)θt��*�S���J�!5���%�@8�N��mR�j!�Uj���\�)����Օ��U�C?=�o����kuO�[!Ķ�K��U�F$K@�Jt��p�p�v48��qd���]�`�[+���hHf;G�6-��9a����e⍝����ۨ4������6ܳW/'g�=������c"�QƢ���oYFuO;T��[����V^�j N�U��C0���v{�Q��de&VUV�b<Vz0�sv�Wv�d^]9;���:K��k��l�M��=�*��B�S;-�e:�`��kM�ӃٴX�p�y�E�Y�H�����ˑMݍ�m�Y��� �4�hx�M<��;��z昰�Z�n-�;��Wm�d�<��K��b7D���V5��1[�Y�ѢƸR�u�r-�v$t�m����[d:���/�9�h8185�� kH��m�Rp�.�����n;&���1TYi�4�)��$��̠o)���9z1��ڪ�Lc�Z��hr���d�`$��b]S+Tr�����t�h�ʦ�)�Q�p5�۰L����[j�IM�%��ݤ=d��^U���t�h��'����w� z���,�|=����ʈ�������&��
�t�ݭf���{��6[ۡ/l�W��af�`2&�,�62z��*�-�M!u��i��4]p�zB���#h���-��2��=�l�����}�ޱ�畂�-צ�� �&���7]��UЛv�չ�Y�nw<�4^�c�mY퍷g:�y)C��{B�Px�'&��XM�0ٻ7)�i{@9W kf,�u�R�d]UCu�&j�5�l�� Qx�眷�35��ִWn'n�=�k�ۙ6�X:�����s1w%�6����0ќ]ds����f�5���y��R�����ǒ����}��)I���c�y({���A� ���n�hv�[JR������ ~B�;������^JR������)JO���I���.��Z�Y�ݖQ�3[��)I�~�k�JS�{�R����=�֣�	��2!BODӚ�6�Z͖�-����|�	��}��)JO~��B|4&f	BP�%	�%	BP������(J��"��(J3�(J��J��Z3�(J��}ǂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	��k�֭������<��(J!(J��30J��(H��(J���(J��=��p��%	BP�f	BP�%	�%	BP��%	BP�$BR P�%	��ϯ<��(J!(J��30J��(H��(J���(J��;��q��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B{��xy��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�>?��<8���K�S]�Ә4�Pq���t���7O�N��v>�w_[�F�e�lk[��(J��<���(J!(J��30J��(H��(J������(J��"��(J3�(J��J��(L���(J���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�}���	BP��9	�%	BP����(J!(J��30J��(N�}�ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�_Y��F��Y�#5����(J��J��(L���(J!(J��30J��(N���x%	BP�'��S�SO���6��� �&b	
`	����hJ��J��(Nf	BP�%	�%	BP�y��x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~��p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bw]��y��%	BP�	BP�% f`�%	BP�	BP�%	��P�%	B~��gm��q�0�o[��(J��<���(J!(J��30J��(H��(J������(J��"��(J3�(J��J��(L���(J߻�	BP�%	�`�%	BP�	BP%	Bf`�%	BP�	BP�%	�w��P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'}��<��(J��(J��"��(J3�(J��J��(O���3>��[w���{��<��(J!(J��30J��(H�hJ��30J��(O~��8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP��~�^x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	Bw߷�pJ��(O3�(J��J��(L���(�%!"��(J���ߏ<��(J!(J��30J��(H��(J���(J��?���k�y��6m�v�[8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP��~�^x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P*P�%	�~���(J��<���(J!(J��30J��(H��(J������(J��"��(J3�(J��J��(L���(J߻�	BP�%	�`�%	BP�	BP�%	��P�%	BD%	]�w����������ܑ�V��5�T�Վ��R�;ng^Mb׳v[�ɮ����|n�|�,���(ѭkz��(J��"��(J3�(J��J��(L���(J�����P�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	��}��P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'�w���(�F���%	BP�$BP�%	Bf`�%	BP�	BP�%	����מ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP��G���ќ5�f�yV�{��(J��<���(J!(J��30J��(H��(J������(J��"���(L���(J!(J��30J��(O~��8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP��~�^x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	Bw߾��(J��<���(JX��(J���(J��"��(J��>י�[��o���y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�����(J��0J��(H��(J���(J��"��(J���k��(J��J��(L����C���D6��qDT�(J��(JY�P�%	B}�p��%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�'�����(J��(J��30J��(J��(J3�(J���g~����kXn��o|��(J��(J��(J��(L�_��@L��(J��(J��k��(J��(J��30J��(J��(J3�(J�����8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	��}��P�%	BP�%	BP��%	BP�%	BP���������b T�Q�~��j+��7ё����A�A�����@�H*�BP�'�}���	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	������(J��(J��(J��(L���(J��(J������(J��(J��(L���(J��(J���(J��:{߹�Y��3Vk7�[�F��D�����ȾK�:�xxM�
v^�%����W39h�g7#F�����(J��(J��(J��(L���(J��(J������(J��(J��(L���(J��(J���(J��=��s�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP��~�^x%	BPBP�%	BP��%	BP�%	BP�%	��P�%	Bw߾��(J��<���(J��(J���(J��(J��(O���3>��o#[޷����(J��(J��(L���(J��(J���(J��=��s�P�%	By�4�B9}Պ(A	�u��BͼX�tB�����k��3f�7o5��%	�}Պ(A|鐰It!H�owb�	I���i�J̏O{��Y�ݖB�UWX���)!=��
([�ظ%	I���i�J��t���/�]��?��)JO����UYsTU�����D �^m�Ȅ���������>Ͽ���)J����F"���J�SwUJ�����=j�v�q�=/s�;/���7O�G�ݎ���湚5��v���x�)I���c�JS�����)=��vO��JS߾���(}�g~����֣u�k{JR�����'}�_C�JS߾���)?w��y'�9)�g��W��nբ����)JRw߾��R���������=��ly)Jw;��┥'����ѫ;��n7�nJR����┥'���JR��*[�(�!B~l�ӫ.EV@��{��)JO;�v<��?�'���g�);�w�JR����┥&���w����ϿSk�6[Ē�=K]m. ��h������#l�p�����;#�*i�"Dִ�fD����0�ϡ�TvZ5l76��1.�tD�8��T�gizݰ]n;�l/@�ᩝ�Wp�j�'u[kQ���ώ&�zu��i�n�-E�n�c��%[O=m��}n�d��D�^��N�u��y�g�lr�i�,�u��o���Y�դt#�YfC�����~w{�]~��C4��K+�� :�W��:t�zgO4\�I7&H�ދ�����h�����n|��>��8�)I�s���)���)JRw��c�JS̏O{��Y�ٖQ�5���);�w�<��RC%=��qJR����ǒ�����-9A��
�6IQ1�N "N*��B�oD �A	�v�K�RD&�qJR����`�R���w��n�ݼ"�{��)JN���y)J{���qJR���{��JS���8�)C絞�w����N���c�JS���u�)J?�������)����8�)Mnn���9YX�\JJM7J1�	;t*f��N6�&ԡt�'\�8v8M��t�m�]�?�{�Kl�ӎt���r����{W���)�}�)JRw��i�y)	ξ��A��fx�:�)V+�nJR�w�����S���R}߾��R��w�k�R�����<��C�TJF���kv̷���{��)JR}����)�~������I�~���R���~��)JN��-�-�Zݭly)_ 	�{ߵ�)JO����������R��l����ǒ���N���YkfYF�o{��);�u�y)Jy�{ÊR������R��?{�qJR�����{�.��V`F�B=:�AF1Z0�����]@ni�,���]/����d�]kZ�첷����R���~��)JN���y)J{���p>DB\����k�y)Jt��>�[��ȋ7��R����Ǒ��"����o�┥'����%)O;�xqO� �R�����I5$Z���D �O]�
����py4̕��� �<E)�?�_w���{�9 ��uB�wTRUY�Д(J^�q�{�b�<����!B��}�� �yD�E~m@��B'������+��Q���z�|��I=-�u��LA�Q�e�n-���^5�urIYۡˤ�S��t��Q��ܠ5uƮ��-�[o��� ����7���DB�_H{�b�:'P�QW�E5xϵ�r�P����{�b�<��~���B��ȹw�%Z�AR������`6�a�!B����5f����m�D�q�@���(ID��|��ـl��}�B��6/���Ͼ�U���>���\�QÂ��0/�l����%L��Ձ���p'�򒔤�n�h@�g�3�v�����v-��n��'�/n��6���������d$��S5w�:{�V ����o%��=���g���<��iI����s�(�=�ذ���6w]g�P�~�s�M���6��ځE:�R+?~�k z�a�"�r�Vϯ��ff��..������P���� m��l�>m��N�iܢ�@����ݶ`�"����{��`=y����ߝ���5�� )%�-�Ȗ��-6�Muhۇ��N-wQ崴Y�W������+rޖ��c���}m�7@(@�G[b�q5Kt��s:W2�v%cc��+0�B�2\�:nT����G3;��}z�,Y8b�N��6{
�c/M'�m;�v9���`r%�z���-���Ž�Kc�*�Ӥ,`�6zTY9��ͧIuƞ�<������=�N�q�']Gc�8]O8lcl5�ND������.�7A�4��7'����~��_�9�����������,�:!B��wŁ�<Q����� i�Xn����	D��}�����Հ=�Ӝ���S�鸚�DQB�U��o��ř����r�-��+����sA�q$uR�wx�B�M�`k�p�x�?DDB_��q��~�V���?!8Ā��vz�������/��}���C�_��/�*�Yt���u���nB��v:�%n�sE�s�Vu��[=�7LX��Z7S���l���>���/Ɂ�T�f��d
���`[��%��G�bJ1	$% 1,�$E!�,�C$�tCU��� x�D(E�}�`���0�x��(Jd薇�b*��*� r�V ��0��~�
�~�� �߿f�V��dʫRH*UWu�=v�� ����
��;�x��)��D��8���XD%���z�}Z� ��_���Z�֬�ؗ1�n1R'ingb7����s��o�w�닋��ݦ�׀���0ݶ`��<�D}!���`yg�yS��T��fM,��8ͼX�����
��O������MY�~uߧ ���W�a$DC�����T��ٵ��б,#LFHl�5�ﾘ�a��4�l	d�(xf!A�Aw����k�6~��t 6�`�<�!�l��a��$�!E�9�ZL���X.��!pѷ�,��HI!C�	ja�L�ŷ��xx�%�@�l8�!�9��hb���ȸ�(��/�q�b&�@���WHt������G���'@ xx&PvP���S3���uʾ����^w܉7H��H�=UUK�����7���y��޼�`n�$��S�*���`}�����}_�]Ӏ|ۺ�:�kT�84�$�$$H�����m�qԲv5�x��:<��ю�=v�w{�}�>���((r7�j��7�uXn��������Xȹt���eU�$s3w�j`v����K������$n�(��pCq ��X��u`9�u�����}��ο~�ɵ/*��jJ���=\K۾���+z�W*BBAXi��{Õw=�gu�mN SidU���7O� �����wuՀnf����Uk��1���9$��K�Z��6BnL*��q�ytt[N�an��-��(�E���4pN.��_����wn������ �9���=UwjP��j�L�_��I�`_e���ďx��&�*2��*8� �論��s�$��mwN�}� jO)�v!����rXz��[�|�c������X�l�:��Ů:J�� �M���np�	{�|� ����k����������6� M���-%�F�cq�F���B��A�Ut��<�A���z8s��Q3���?o���g�����]�v�ۍ��7=�ar�il�GV��6$��h�x8L\.8˕��79�n�<�&l�Q�v7De3`���.�G*�ZK5gAx���lU�n��X�.Mu���V��묉�2�!F��u�-C �gS٭���5�������E��~Կ��)���z��l81�
��M�s�nʻF�7��G��ѭ��tΎ:�ut	�?�ό�u����Z�����mB�(�9*�73e��ʤ��}XmwN�׋9D%2t�	���b6�E]]�K�Հ?Ss��B��"�{�Հ~��K ��V��[T�"8���~�� ��ŀu�B�J]k��=�Q&�$�
@J�N+�ͺ�=\�+�۾��7��������JRN	9Q�
tg�Ms����u�����^�R4�,l���v�H� �NIR�%QQ�%X�l�6}���l�$���>ŀr�T��U�hUuWxϵ�J�!$��L��ڨ���T3/����W���(73e��VV$�%��AN��X݌�>m�áD%'7׀=w��&jTI�J��p����s��?o������`�J!)~x�Sj{*����58,�� ��`OM�˴`}��V�k]k4�1J���V{��[o������Nѵ�ɉܷO��ӻ.?�����}����E)U|rI�~���X�4�>�x�DD$��9�^ /.����WS5$�0,�S���d���m߹��RG}�$�$��"!������|�8*h6b�C�G5�>ߕ��~�7
x�{%JD�EG�`u���u�?Ss�В�s��MK_������`b�k�=�W�{��;��Հnf��Q���G���j��et�i��5�ۖ�Ը��c�Ŧ�);;X��㤤HS��v���ͺ�������;t��J�4�P����>z�gB����������ݥ��#o�'%X�vX>�Xt)�n��=ϱ`}�2��N)$��&�����OS�Հsw��׋丸�e�Wի[᭪q�������������ݶ`{^Z�dft�x# ��%]�5y9��>�n��r�ĴI�=\�[�ꏁxW�u�k3o�ǻ�� ~n�ݶ������w
���ݫRU�+������rJ!D�۾0n��>m�΄�L���.�����f�n�-����m��0��:��Ų:"B
t������� �>ŀ���%�+����9��~�*&5#T�8XnmՁ���9\^���u�`�l�-(iB#�q
R��w_wwn���k�.�{v����˫h.?ٵ�/N!����]�ɋ6�.{0���k��;m7�[��b-tg��(/���ݩr�'[/hڨܗ�RY���+�s����1��n�y=�s��v�6�=9r�ۛ��'j�IB�Ԑ�M� �mr� 8����g�&�8YQ�7Jqs�u݃:-�cq���6�G$��4M�%'����������u�v�sk�#�!ė����\�#��ոJN����[������}��Gi���f�:>���^��h��ͺ�5w-�4���O����ܙ;]�v�ŀ��9)�^Nz���,*H&�p�|`����w�<y����7I���D�p��){=�, ���k�脡~����~0ߊ~I~�T�9TT��V�ݖ�M,̚X�۫��M�N8�M$��+YE�����z�0)&)�W<�nL�:iV	/=U)�w9�Pr9>������f ��/�$�z���~�ȿ.��6Mҹ�AR�����2�VB����!/DD$�GX�`z� ��tL���֥DƤj�F�,f���7����2v����0M�yJ���ʑ
f��G�U���x��������}��`~^����i
#��� {7���mҾ0�u�~���)sw3y�m0�f۶.C��ӡ�mh�:�s�Gk�sxK�k�{t�����n>�ɸ�_�����`_J��/��}.�;bԳ8�{P�IA�{�u~�$�zX�},̚_�=➤�$�Hs�I�`�׀u��JD���$���N��=u`f��p�G�áL�}x7|`����� �k��F��$��M,��Հowe��3]��rV�Sd�*�q&���gJrD��]�s���Ǜ�X��#����)Q6��q�m��7���7���ՙ�������n��l�&A��$��u�߸�W��}6��]q#������J��O����������ԑ����{7��>�T���mrSG���m� �������J!R^�W9Uu��9z���n(�t�{P�!B����w�r�������_V �f�txۦ��'4�B�T�B*A[W��p<]m�����uWZ����Fka7(]r9RI,{�,]�v�M?��پ������((�7%����9B�9�� ;_^ ?7y�(Q&Ⱥ�͒6�D �M��n��we���#��Ko���iFڕj9F�,?s�w=�`�zXY��̚X��[n��2QE�`��`uIq�d�0�u��߷�����d���ZG�=,w�Ǥt�*%���xe��)�	�ߋ������s�-.��3$v�D�\�#3s-F!��^�*u�𸩄Uz��M+��_G $|�"{�8�
J�y4�J�"D�� 4���kZ�{����{�m� 8m�           p -����� �(�5G��[�m���N�Pk�#F�L�v-�#m'	�S�ggrŮx�=������l^*�WV�/V��4�l\�L9Cvn�J6���`�j�ROn��hu��3f��]�6�
u�lo&a�r�A+e"��.U��n�[9KM��E��[Z؃���ug�۱�yۈ�l�m�z��FR�:�o7��iMvy��m͵��pl��R�,pZu�T����g%���9lm��j�OG�,�s�st>�.�oba��33�j��iUַ��,��]ғ(2�88@
VV��SgUU\��ٖV�uK�K��щw�R@�5�v����N3u��8ָ]�����
���g�`[�hYF���s=�ާ��j5��J��N�YYV�x�u�Uy[��Ntӫn���;kY�\��-�,\>��`%V�u��]b�!�1�a3h1PU�n��J���5Nx��d�-̊��L�Rڞʎ��(�<qkN]cF�ڵ�
X�u��d�.��ɇfV�l�,dZꔝ�a�XW��U�K,�p0��qͬL��y^j��SA�t�e�rnJ��=�l
��Tm���ɔ�8�(�e���m���]�pǮ�&)gi$)5\xw���A^�9ŧ�t�9	-�;qe�`�������t�nW�A���KNڞwL&КAl����^Np�2��x��9˄�GK�@n�lc7jo.�̚�Н�A˞����c��}�h6�Y:]dh��%��%�S�۫��ע�dD\m� <�gs�yM͗�ͳ���l��˰�*ؕ�u���a��ƒ�M<���r�pL�vJ:�t�Ng`�K�c�q�h���]T���n�^M�g`�]��[��We�n��/���WiN���]s��9�!�M�ݩ��͎`ɇ��9����,��kZ��PLQDw�H���:"�(��z�Ĉ��ip0��W`
�/@�N�^5�� M��YKk����m��j�n��3[0	��i�ϕs���O9ܑkv�.ͣ���.��!!�n���nR�;r�SW`������lk�ۢ���`5<(8t��x�b�����r�gD��<0�h<A�ہ�����r@H�$���t�:X�vڔ��&�8��4��$���t^K��U�b��njr�U�u�Dk7���f�~ʌ*ou�fxW'"m�m�g��6c�
�3��t�s��nǷ��w\��GI�
l����F�.�G'�j�u`vـ}:�~QH�׀]*]qmrSE!9,̚X,�v�͖�͗��q#=�$�l~�H���с�~�������m�x�OdI�#��l�:�5�ܚX,�vm1,{9�PQsu��%������<��}.�<~���͓������8|�.xEgt**zwn�8��cn�6-�[�g������3w�J�^�}.��s�<��,���*&9"e*I8���U�\��q}.�<����T������n����1f��K�/K��%L��U��VQ�������)$�Y����0;�0�u�w�qL��p�#���`Y6��-L��`yw5��Z\��dR��H�'D�M4�Mt]i�Nɮ�b�݇=�R����e��"B�9%��^���:���s�\����K�Sԓ~�'
#�����%2l���o� �|�`�cب��PP�nK�3]�nf�H�������|��W����Wr���TN�B
t��73e��<�`���S�o� zp�ɵr���p�����̕0�u��%�}.��N����Z櫠L[k�G0�v&u�l����1Z�VΝ��w��=�C����h^��p1n��}/���� ��X�*�7+(�g���.]R�O�����H;_^�O� ��tB�]*].*��#�8�پ���U�ose����`wqD�6-�H��Ia�UR�����׀};��6"�JcjaT&�`�`�ʳ�0w��$��s��9G*����`f��$��LRp�f,��/��W��}.�;�0߯�~���MnMi�����wgN�f�zpu�=�mc�/l��lZ��	��n�c�f��:���/��fJ���`b+���U�Ђ�9#���~�$w^�X�ޖ�3]��hj�)�Ou,8�nf��%L��`uIq�\͖kv��d��Ȩ�jEa佞��,��`K�ܕ0,��w�z�rF%7W ��N�)����O� 7���\��W;Y��1�$�I$�Hk�qٹk*YcMlݨ՞���*$�ukt��^fɲK4K���j��s�k��gN�[7+������\I�����̫�|�7$r���Ƨ.�r���k�lVq=C��l�����m],���^z�^��V�z�s�8-����6�l86�7�]����k(��[��p�9go6�ݒs��LX�# V���t��\��N�1��p�B�vqj�c���,�sv��{+p\ְ�7'e�w]��S �]`v䩀_K�	�0;��J��!R�$�>ך�{�,��V�͗�U$o�z�o�S�4�V�����y�Ϲč�p���LK(l��6������`���>ך�{�,�v�\�#��H�˻� ~�x(�u���;_^�y���X���%#N�" �$D%��0����+�X� ���Y�m��ݭ���VN.F�>ך�{�,��^�����2�Խm�7'"����ose����
��?� {Z� �ֹ��"�?z�D��q
#�T���?y��V��Lܕ0�u�{�r�o,Ú�I���
y���=��p���7�5Xn(�������$V��U�[.�'�T��%LH��ԳRY6��gN{fI����A7k������;.��H�狞�p��"$�	� �'�n��{%LrT���S_؉wN�5 �����7k\�DD(����N����`e#+5Ȉ�	!$V{�{�����_%*|*�1*i;ʴ?{��Xa����$)+����Z� n��k�J{��l��/[d�I��jE`���μ�`n��`}�5X��ֶ��7JU���d����-�h6�r�z��C��l�b�;j^g�6$�Q#��b�g.��'@��~V�0;rT�-�X�W*ʐ���7�j`[��nJ���{%L�TIpl{P�IR�+�y��7���μ�`n<�`gP��"�!�W8 �����8��8BJ	!)QBQj"}w�pqR7v"՗ P�nK:�U�������+ ����X���R:$L���j11/Fv�7�6�N�M^�8"g�vn�tk������#����*`v䩀_[�	욬�CUʌ�$m��4�>ך���`Od��fJ��U37R�\��ź������S̕0;s\�V���W�D�X�]]��y�~��>��M�$�{{� <�WUp�J�i�?!n��*`v婀_[�	��r�>������
�}���k�6[ۧ�Ֆ���bc6�
�Jڠ'������U�J�grK/-g��gH�b�)�Ll��^���^3����;��
䂕[]�������z����n%�ܗk�j�O�8�3'.z��=wOKMbwQ��g���k8K��	6N�tI��:md�b��{^�4���x�u�Ïm;:�!���ڛd�.�k2n��Y�Zխ���?'�VP8o�sf�eÍ������trXBq^�ς�����k�gM�`���[�h*>�~���}n�$�S̕0'��"]�B��pFu0�u�&J�d�����`f��D�D��3T��%Lܵ0�u�8��sIH�	!$V��V��U�owe���U��EmrB�q4R�ӊ��r��/���*`Y��d�^i��i�7N.GbC�/nn��e���<qػa���yu<⧢	HP�qJQR�4��q��owu�&J�d��ے���6�o5�͇[���]�]�9��0b����{�����L�%L��`�\U�N�d(|B�X�5Xk�V�ݖu���o���4�)"�;rT�/���J�d��?/!����N+ ����+��sro��{^�Xk�V�����N8�m'�͂+q)�[��8��`d Gokg�b���%8T��Q*Cq�>q�Z� �ֹ������xR4��B�7BEHI���U��r�;�V�����y��̢���!R8�)Tj�p�k� ~n��F$֤��DA�
�)f�3M~�A2~O�� ���ͅ�l��*�
N)�?�(�ج��@f��?*�Ҭ,�P�<�L�b�*��&BX�8�*BvlŐH��G|��DC5K�8IEQ��r�9����M[��U4+�i,�,��iPј�'(�f!�QNm��4 ���(&���>� OO�!�<W��T΂��� mQ����{���f��J�c���Ʈ����W�����N ����s�=Z�֯$���*�����p�D.v�~�O� �����V���D�Vqmٶ��`{l�wi�Z�V�ۛkiNsp�=��ECQP�t�B��)���U��s���D/����9����>� �T����^j���$�zX�|�ǚ��*�#x��I��4�l������S̕0:������{�IrXz�T��|�k�g*�=���~4V%��/灀��r�����i[�Ĕ��*T�&�*`uIq�_[�̕0;��,��7;5Xdk]���z�;��ލ��u����ls;����$|d�sI׷j�V����`vd��fJ�M�r�*諕uwX ���$���O� �O� �w]g��)��h���x�SibUuw��ߧ {Z��S>�����K �j��Sl��)��Z� �k\��w����J���N��$�(�P�IR�+�y��7�����{��]�^�9V�t��S��
hB��Yag{�}�{�����\ 	��$��L�®�����;1���XH۫��j^���v�ܰrͶ�ҍ�Z���d�������ͧ��cjW���w'D�,�n�YuVwn+���&�{;�G�%˃��/	�,�M������p�}��+u�#�n:�Z��	��t�gnCY�-��=gqv�ח��qQ�/n�N��5:|+vy�]��n	�� �v+5�W������&>W���6;Z�{s�k�[VP�ɘ� � ���z�8v#v������פ���7v�18� �{���j�7j�UU_ ��7�ѯ�P�"�"nK�y� {Z� �k\��w��~QG)���J5$��$��������j��)#��K����̣@ے�F���Q>v�p������ ����ݥ�!u5"���=\�vo��{^�X,�vt���R��\��������'��[hWt�n|z�gq'n�Íj:'�t�˪Q��׾V��VӺ��D/����](�ԩUQb4��r���{�С�U|bH!��" 4; ��y���U}���>ǚ�̉6�ȡ��$VӺ� ��:"gΟNΟN �|�k���*'��Ur�/g�,�}8��8���V �T���M\\���Y��̕0,�S�K���`uf�[���) �')8�x�1C�q�FrV�(]S�uҏF�E�Nu�S�3ؑ����`Y��T�����ɪ�̣@ے��M8��f� ��X�*`Y���o\Ot��WHU�`�w�}��p��B�D�U��5X,�v�����Ȑ�9uJf�@���`Y��T����9��,�M���U%"�7j�?��s�w��g�,��r���M�7�V�k��È�q7h�u(�l�붞��6@.c���鶓h��!T����fk����%LrT������tŻ����l����Sܕ0:���ͦ�oU)P�
$�9,��w%L�.0e��=Ȯ�L���ww8u�p�u��"{{��ԟވ.b�}��\(aF�1 c �pxy�k�3�}�{��s7���sy�50:���/���J��5X�W*�nyz4�Q!�N$�*����71��B����\������n{?l��g��eE@P�} ���K�y���y���f�5f�;"Bh��(��׾X��8ӭ� ?7y�G�@�}Q2�P�d�����w ϳ%��_�X�c��ED�)"�>Y����`zd��fJ���2���}n�=2T��%L�.9'����׽;�ߜ���f�\ $�%η��sW]#�-�&�ӀӮ�=�0�\���ے<-�X�5����g�񇮓��Sf�N���Ӣin���C�J�s�2��Q�XA�;��ރq���)۷����۶��Ţnq�Yv�t��A���N�݆�[z����<$:��9��8�Kc>�䋢ո�*�\k�.�'���],������^�:��,"�խ�I�la�;s�-��Su�k�.f��P�r��I���N�A���7X�J�d���%�D�ɤ��YL�f���lAR��}�IkɭZI/�f��I#ri-$��3W�z�k]��mZ�Jt�R�q�I%׻���$nM%���&j��דZ��]��[�d�B���|��9\�k�~%�������דZ��_<�|�[�����G.�G	�I.��/�I-y5�I%�����$nM%���\���1������K�I2ym�X��j�ˇ��ź-����TXn��rq�ӈ'H�Ԓ���$��s_�$��4��K;3W�$���1�z�J���I%������r�U��hܚKI%�7W�$���դ��>���ӕEA����7&��Igfj���ߞ�5i$���|�Ki�f���D�%�������%�&�i$�{���%�M,�KI%���k�Ӎ�*BH��$��֭$��s_�$��4��K;3W�$���{�|��-��@��4�hv ��F��vz�^h��E�11n,����#���RJmƾI%�����7&��Igfj��דZ��]��[�"R*��#��7&��Igfj��דZ��_=�|�[�����$×T���$���/�Y��{��9��D�3�� |oߊC���i�5�o�癙��o������jY�$D���_|��s��S���V�K�����7&��IfL���%�"L|{P�IRr5i$�ٺ��$�ɤ��Y�5}�IkɭZI-��Pt�8�3`Μ�ɮ�e�4�����<�whT_,!3[��n�1�(�۬���~~��|Y�5}�IkɭX�_l�_|�[Mгc	�R��"nEi$��5}����Smyl��$�}7��InM���Sm-�eo���#T��}�Iyl��$��3W�$�ܛ������K���)I)"�Jmƭ$��3W�$��4��K;3W�%�E���@��(B�D���`!�FQ���@!��֭$�V�-�ӑ)GÍH��$�ɤ��Yٚ��$��֭$��s_�$�[ߏ~r�]a��B�Ϯ���řy��tRpbd�Xѯl�B��ݯ��� �ﻉ�Ԓ^����K^Mj�I|�5��I�Ii$�kRY�E#$N�}�IkɭZI/�濾I#ri-$�vf��I-yc��ڄJ���I%�����$nM%��\�s��پ_|�^{<դ��>���ӕEA����7&��Igfj��דZ�����o��$��:�0��((r&�-$�vf��I-y4v�w]����r������\	ڝ|.�Wp�(j��D瘦�9���ں5��{�D�H���K�٬7^�r@<x^������8�9C0D1��K�ޟ6%L���(�""8�rs4N��RI8&� �������	�r���	$�w�BS����+�v��'�����0���M贁~��C�#T8J8��D;�?fgw��{����ְ��          `$ �,��Z�Ay��iҖ�$���q' �Jtt�l	�	P�-�֓w�s�u4���cD��Gtm9���]e�c���,��cu[�;�Q�-f�[�]�LaU�gg��n2LWI��v�)
Z�ɇ�wm�[\�� 'Xd^�V���ۧ��.�9yvy�Fg8Α3��m�
e6��m�5���u.�a/Y�\��t"I�q�M}s$�yh�9d�jq�2F�a�z�-F��h�mfu�G$���u�B��b�v�\\�3c�7����4"��dz�3��f�6��0���0m.�Y	cl2��UT��l�� 
��Y2�2dP���5<�q ܭU:eR�{@T�î�^x��rN�������%&79N�cd��*�����y"e
x��{�l�:V��&��k�!�7H5Q�jAN��;"�mbѵ��m��3�t�Y��=N�D��h�pr/W�zq�x�Pb�\�����=��
�r�>�\��qY��T����2�s�i�q�b��ݶݖ�%[S�d�� N�>�Zy�5�]����m9-�k�^�a����2-[J뫮y�(�W�JX$w�k�X5�M)I[�dm.����U������l=L훫^�X;���7l+�a���K*Q���v�rq$��l�8�����2y�籝��ݖ�%k^�S����'kOSڽOX��<����s�+'6��^��y�ny[�絺N�a}��an3ٷk���=���&v��t̤n\�\�#�I��u,6'.���%gm���Iқ��me6N ;m�l��A�%��mh�k�K�F��.�����I��1��*�ڻZ�d���{Z�p=���GMn�)�*�f���T�f�*qo�vD��-��Z[ԵO��,�չ&�-0-�����%ݱxK)������t�,Fg�xm��z�ۋ,]���ov��վ��� /�@�4�E*���ԃ:��Q�x�Q^�OP�OE{�����~w}����6� BGg�V��5�v�ՠ+<��tUT�<�㒵����q٦M6���1�Ϊ뇭�;x�w]i�s\�\�M�i�.�ͮ�	sK�;���N��v-�糃tkm��vw΃	qu�{=��v.���n���b"K�v�a��n��@=��K��1�����9�nl/C���[�b�8�#�VRm��ݶ�8�bB�߮����u��~�E;D���z�.J΍vG��ѹL:���ɩc���fѮ�g�n���ARE�j��`|�u�ܚ{� �{�`n�)jg�'%%�R�q�+n0=rT��%L�n0=�x��fĤU�`w^j�3j���Z��vW��`nn�/�:�I&�%"��~L�n0:�����S �*��H���R+w]����UW_����Vc�V���o�5��n񇛷c:1X�^���X��E�C�Q�'c�ӕ4�'#��{����`f<��������X�j~��*�����ʿw^�9�,��!&�^��� ՙ���n�6�яb	�R��"Y��$Ҧ^�V�`z䩁(ͭ�ʉ�h�X�������U����`f:)bf�NJK��UU���� �
����m�Ӏl�u�fJڍ�JR$ND98C�%Ɨm=��{�\��8�̑�fzl�m��<�QT|87��y����j�1wu���OwVϸD���♚ș���m�Ɂ��U��*`�D���n��!������`|�uټӜ��J�O^.�|��]����{��ʽ�����5��J���~�W9�.�{���=�32�=ʪZ��v�b��6������J�M*`E�q��n�0x�[�)I�!�(�����U�V�a����<����Z�-ح���h����n���M*`E-�U��uX�6�G*'M�PH8E`b��ΈP�)���ՀoWt��c�}H��b�)��$v�w]����`fd5X����m-�*(��.���ֹ�7v�8ϵ���y!B�Q�Ur7��7�Z���L*q|�O�/K��n0;rT��=����d8+pu�[vЛ`x��ӍԚ�굱nӻ<&�}�6v;[�����:>؋���یܕ0$�T��T�|ȡ"I	8����y����j�1w5��H�,B5?FەJ�ґ��/Ɂ$Ҧ^�V�`^{8k؂T	AC�)����`b�k�>[��=T��V�g��9Q'L%�4������یܕ0$�T�>���;���&� l���-��i� ��߾{������6�\)�ə[3�3+�n ݋C�-eu�7;�@�qL����6݆ⶲkZ�h"Q���z8�8���6jGv�rK�6�.9�����=-[�e�C������� َ�&1᝝7�N��Z�p9ל���t6^}���l�����$�{Ļm�t;�n�vY`�6��뻽���P��7�)r�ez.6�ǉ��.�]����sv�u�xuv���T:��_;�I�_}�0;rT��iS/K�"^+�*('Tpn;�y����j�1w5�-�w���ďfׁ~_Z��aV���>��?�/K��n0;rT�;�Fjd�u"J�������n�>ך�̆�jM��GR$��n0�u�ے��J�Iq�����a<�c�RRb�"tF�)�P�gno[9�������.�lk�\���1��[�T���?yX�V,�v�w]���F7��J
�H�̆��؋$��QN'�yy�}�\����>׺�ћZ�c	A!V\�;����X~���uwN ۳��κ)b�JJD��)�����`}�uX�V.��ͥ�H(7���3q�ے��J�z\`u[]�VwV��'RB*M�)L���ݨͧ��m9x��<��q�v�����c�>��w��f��m�������یܕXը�L��n�IR#"�1w5�m����SI�L�K3�2��rD�q�ۻ,��o9ʤW?}�	��k���Q��T8������>V/~�3��F7�6�R�n��%L	&�0"������]ުR�J
�$�32�]�v�w]����`|�kT��GZ݇��Z��f:ܶ�k�P5�Wkt�H����J�9QF0�X����n0;rT��iS��$T��Y����;廮�;�HfCU���P�ܥ�H(7�E�`}�5XM*`E�q��m����;��X`�f��m���$�XV�a�~�P'�0(�}���U~>˿7Q�n�IR#"���`|�u�k�VfCU���Xl���N��R�#H�ͣr�+�t�tR��v+m����TRE��U&����#I$����n�>׺�̆��W����7��o�7!�P��nJ��J������S�oU)P%D�Vw!��3���ν�`}�5X��Z�8�*�X{�no�����`}�5X܆��Ef-$���%2I,��Vε��9��w�yF�$���ԕp &�Y�J[[��I���T��rD;سl�a[<��ܾwf�8�[�s�A��h�y��[;[;1.�vm�38y�Ex�J��)��n{P��ֻ��h�l�cϜ��yƷ8;.�/��{gO�1h-�fR�UxC����ۧV�;�t��'ko5n�z5�7�����q��,Gb��Nv!�Z�v���N�2uے������Q���Pַ�٭kz��挶	�jݝ3��t˺���6xM�C�1������}��h���I%E㔨Bq`��~V��� 7u��} ��� ��?�i&`�N/��l<�s6X׺���W��\H;Z�y22$ӈT�����k�-L�0=&�0*�I�@�{�4�����7�5X̆� �͖qu��&�8�fj`_e���4��Y.�;2�������vXE�֋�v�5мt�t�f��nn��+�H�c�L[h3�=��K]mvݨ՚��J����-L�0;�6�� u�T��V��/꯸����) 3���7��k��9L��t��Μ�2l�s���M\!rS$����x�7�uX̆� �͖�6��TPN9J�M����U/e�N��Ӏu��v��r)��Դ�
�T)�g�V��,��,��V�y�yט؛N>6�#�#0����3g��8����H;q:��p܉��4�"2/�=��`gvi`o^�;�V��M�SM� �HnKz��*`z�*`��~^B1�rU	���y����5Yu�6A����k�k���kd,h3E���D��,/Sa�[ڨp�p�"�4����c�����px/�|2�~Y��6��BH�`X6D�#2��)a�C$�,H!�F>���s�l,&	�
 �d�����0���b`�6c+FeH��`��b���D6(��G~(!�4��T4z����eP?���}Ң�(I*��ܼ۶��R6�ʛV��j�LY�L�]`O]�z�U����H��"������F�J���Fg*�3*�5!*��mi�2������`d��zm�Zx�Hr$s�r⇲���꯶߿]��-LYͣ ��X�x]�QA��*,��Wꪤ����`�� �;f ����y3T�� M�����`��z��*`E�KMu)A4�"S���R^���7�p�np�	O�(��D]7fN �ړh����i$'%��{��޽�`wr�s6X�-����%f�&���^��cɯ<�[��{>X�.Y6ᣣ�B#��qT$n+z�U���j�9O7��k�p�Ht�Qj��"칫��ls����2�^ ��� }{��\�U$f��y� uT��V���m78t)���[�� ����:���$�>Ǻ���Vs!��73e�w�d��R���L�0=&�0%�T��ݻ�{��{����'i�  ����� m��^h՞��`X�yP(��O+�6���^l��i�U�Z�պSK�Y4�:�%��T�[�U=r��@mа��[r+r\�lX\n����L덶vuj���^�(����6GU�!��7��?9�rmӲ�ם��9R[zu�m�8�d��g����Z��OI��+�ݕ��c�� ��g����vH��ۻ�߾����yMt-��ɦ��]���u��]ې5m�U6H�m̦�v콘ۯ�믅x�v6���i�����'���J�v��\ӈT�N�͖�ݖ����4�5wRm4��$���z�`_e���9�`K����d��$rXUq{'��毌 {��|��z��ܢՅ��j�LYͣ �]`���7U��3[cz�#����ԡ��mf��{pg�3���ދ�ۋ4�&i�#�X�M�X�vR�0���w�?SsТU|�=��1Q^�z'Cs��$��n��ay(���j���ݎp{�,�m$���r�RKz�lҦ}.�	�u�e_��5���X
I����;���8���}�,��V��Zk���q$"2+ ��X�����S�iS��-�v���a����lb�nj�F"���%��;ˬ�5�����Y��-��e� �k�������D%����ňG����#�X׺���G{���o� 7u�t��i]r��V�e�\� �<��!$>�+��\\��������`}�2�� j��+��ف�g����׀?Ss�}ݩ���En%�:M�
\��K��q�}��}9�`���o/7�g�.up��u7#�.X͟���;3#d�'���i���,t7l�$�|�}�J���р_K��K�o_��K�m*�
��;�S���A��K�w���w5߹IW�W��&&�I�V`���>��XtL�[��<ݝ8��R����Đ���.��;�_V��pBQ
b|�^�>�GN�rB�5$v�3]��d5Xٛ,�f��7����q����":KӮz�g#YA3Zp1%7u���];g����I#�>̆� �����fk�>]�v�3k\�P!EH8E`���K��.0;&�0"��D�GI�AK��I`|�5�,�vz��Í��yXs},�m$���q�n�����iS ��~��췫 ��.�֯��K
����vt��!D�__�z[��>�k��B�)=���~7k�6[ۧR<Dtm�H�뛭l��ch{ ��Ǝ�7��S�h�m�G �����WMdY���v��e�A�'�8�`�̗@�*�`4�����#l`��ō1W�}c�i3����ɉ��M�M��+�[F�ۓlqm��#���T��r��#��hͳ�8������n�>:���u`���v�;$�ӧk�Y��\���N��{����gQ�ױm�i�.V�vi�qa�uН:؝O�!W[����z��-����� �w]`N���D}!�ڞ,��$�"M��Đ���3^t)���V���n��6'�H����DMI����`}�SK �3e����`muѯb�r@
$���Iͣ ��T�^���6@@�X�͖˹���w5�w!��śZ�M�!T�(�`,VQ�x���rnL��C���O7n��Y�y���n��N��rS�;噮��w5�fCU���k��l��t��TP�vӺ�>W���,�7ls�[�噮�I�QSߥK�I��8I�g���;�u��%�W���^*\��B�pFE`|����f����a�����<���$���s��RN;�K��K�ɥL�K���Ho�W?�vk�֡��LS�,�[;sz�tc]=��lAlGn�5�yf�n;B[��<���J�R\��+V�k��{� Q$���Y�k������K��/.n�� �*˜��u�};���HI"�Uv��[�����5X��bt�S��)�����`|�5�fCU��\����`��󒤔��TRR+�� �	y�:~ �}xӺ� ��&�z����S��m�.��:�]m���y��s�!��z�[��W���|+�vݚz����;%�T�R\`���l���q$"2+ �3e��<�`|�5�fCU���RGuDM�Ƅ��u��o�����iS �X��#vH)!�PjH��f����N����DBW�%��W��GD�I#�>̆� �3e��<�`|�5�[[�C�H�n� ��sM8cI�'�M:�f�Y{v�S��W%�%G$ ��}����j�>Y��U�s�݇����Խ�����$�>ǚ��[�vwa�`|�5�p�5�I)9 ����w5��J�^�R\`Yh���t�fg7�n�t[�Ɂ��q��%�W�]�v�����RJ2+���`uIq���q��4�����s��?D�sc~K�6a�s�I�J��45w32�OR�<!"�����((BBh��������b�~�FFόl� � �$���&�I�*@���#0"i+^1a���1��� jr8���Zqԡ��]������t�$.�S�q(jU6H��=c ����|��O���l?*Kd�s��*�~dC�~��
��G�?>�D~l�0s3 ��	�a"������~ �n  �          �� �$��miJ�<�<����V*�iWդ�6`5�MӶ:(g�tq��t�Q��`��gV����]�%�Z9���N�˒��*�Zya�vnIT�� �,�DE 	KcG^8��n+���E�7Sn2�-mۥ��"l'ӄ��UQ��Oh�u�(�î��z���+e�d���od�\u��<�7�֥��S3��T��J-��Vpa�EuJm�3k�8Ѣ6�v�� m�H4Eq��n������&�\�p������Jl��ZØs���2�nM��lm���[n`�8x-�UHR��]�6�*�,n���O�ݯ�n������c ���$��t�s����ٳ�[@u���[<��@ �6ۍU��m��ӳ�@(�e[jyJ��f�v��ۄ)y�;8�!d�f��0��5JZ�]�R���M������1�؄x�9M:��ƜJ�6�.Ǻc�d�X�g.àl6pZ�3\��n����[����8��0�AC�D���1˷X�&��Q�e(%[�SK�cU��'f�ll�m۝s�ಮ�R�g���h)!�=��$�	��,�E	�98ݞ��{K`5�����ϝ�َvq8�Y��C8�]��v��^��d$F�$�/�qq��F�4���>�y������"q� la�e�s��78����xMl=��pv���y��ٍ��~�]��0 8�-���Й�h6��������u}|�����q�L���ct&�W�&��l䛫��<=]N6N1n���ŝ�Ժ���N���m��|r�"�v ;8A��ӣ��������W׎v�UWoX��( #�vV����7]@@Uk�-mna�l�L�A�Sij�J�Qu۝*�UH�R�{�o^�<��훖74%U[-����V7h��8,k��=��m��x=T�Tx��"�*�O�C�~�`�z��M�iN��_T�EO�󻵬����]�:J���v���*����B�bw����p�c��1g���紉V�j�����q����&�ż#+pmJ��l����s��ze�͸�����fsR�����8�3��UВ:�-]`���<Wl��mW��Wd��f6z�k$v�6"�Z9��M�L)_�����x�z��e�V��I�m��k�`
����W���w�|��v�it׉׵hr\��S�Հ{1Wk���v��ݞ^�-q\t�	"��s�	RN;�w���w5�fCU���k�3��F�RC���������iS����K����V:<��$$����<��s]��q.��;�7���Fmk�Qp��4���������K��CU����[����NH��f�T��J�R\`ur��e���gJI�a�ŝ۞�5��mjѻ^C����w�>{)bM���I%)$��V��iS�K��.0,�\���>YU4�Wu�nΜ���)I)@i�0M*�)J��"$���

Û�e����u�UUUIW�yx�pQ2*������R\`uIq��4��ْ�#����BT����]{�vV�d5Xz�u���ňG��JHqT�;�K�ɥL�.0:������6E�׭.�;nF�e�'^˳6:�:@�C�.�# V�&Y�j�v�۶�f��vM*`uIq��%Ͽs�?s�Py[�0;ឯ7"�� �����~�s��OK}X������BS#�k��n�jp%9#�:�|��f�>�W(�e� �A�Pm���`b���p�5�rJrH #�:����T����K�-�.�Lut��wa�`mu��`|�5�,�v.ֺ�:i�4GĢ�95ٶ>nrP�W;zw���MW=��u2�ny5	QGRpJ2+噮��fk�>Y���!���wD.��r$�	ǀ};���N����Ӏ9�u�gP�[#N�PjH���Vِ�`j��`o^�7L�7�Q9' ������� s�� ~��!DjJIA��C��8̡�WV��؅�f��Iq�}���Z�M*{o��	���!(��qc��r&����N.�]ڴ�֞�뚆�v�%���y����0/����iS�.0�kt�ܐ�M'��{��\����Ӏt�Հ?Ss�=l�?��M7N�����=�+Vf�?W)/c����~��)f�r�#U'�"�*���-L�0,�T���K
t��r$�	�a�r��{���?yX�c����q	$�*Z�jMp �ŗ:�拮�m]=4�IH^����v9YNֱ���ӻP���b��X�Y��%��5=lęq�n\jx� (ܕ��]��� H�b8���nϞ�r�Mn���i�ҝp�nw��n/8�mk��{c���&^�)��q�9��:�RwcA��R\JFw=h؍v�ٸ��ms�V�i�s>���m�����&���i��w��{���>O��vI��ˬ)�h�YI�/N����{;b���uBk�	�b�OQ��"Ϸ[������?���M*`U%��Z����2�ῷyÙ��SɥL
�����S����r���g��9D��
$"�>V���0/����iS��1lPI��\���޽�`o^�76�8�B��o� 5���UwuSw'3��j`_e��dҦ^��i`}[[+i1�m�%D�*Rph���L}��p=&�vpc�m�)�k�I�%�\��^άq��G܋ή����~���X�����,��V��t�:�jN	6E`j�k�J!	D%����\�kY8�17L[D�����۫z�U��	%3Ο�t���6'dN��Uub��9����J�d�`U�q�e���L�7�Q9%QND�7h�BK�{��9�b�ֹ�6Mڢ��]�[l���O�u�LQ9ێz�9�Li��kc=e�}#A:�*4�e8Q!$�����=o ��� �����ɲ.�q$��.Jm�`{}�q�q�����`a�kt䍩��%X��r���{g,D�"V�	Pژ�@�7w=�uʻ�{ÕwsEB���M7J�����=�|+Wwk z�,�"y���0��J�+*������[�-|`Y���(����)��A*��LT���v���L�%��U�M��z���݉��F��i�I.��-|`Y���(���u�{���-Ey�A�%*%*���ܭs����]���u�� ���:'$�)ȜV���}����ɥ��y���A�Zӄjq	 �:(S>}׀w;� �ֹ��]� K��jzy���,�]���;oi&�r1�,ܚX�5X�tV�ݖs%mJhu��2(�$�e.����@������n�7\tq���Y�]v�紼�6�Cㅁ��U���E`��`6�,�d���}���KI�������������*`�)Vsp4�Y��h��������*�7h�]�6�[P��@�m��ֹ��d�~�IB�3��x�j)y�TnJQNIV��V����ou�[ŀ4,#aBM��w�M� ��ҥ:^��į%!AY�m6�Ψl����I�w9�n�4t�t�J&��隹���8��i	��t��1|�l�h9+��8x��Pf`�T�*K'NNہكʊlb�-tn������ny5W&��v��ܝ!�]�X�譊��wj�r�mq��ٶ�z2N�g4�J��H�3����e���rlHY�@:.�8�.4m��q�	���wwu��W��,ɜ��]��Bn�uv�g#՞�u��	%1��^�Y���:Bt'#	�*��'��?xL��`Yk�̕0%/.,�sp�i�t��0�u�e��2T��y��:��6H�np#����|`Y��lܩ�_[�м.g3dMH�C�`n<�`}�� ���{�u`n抅����S����;���0�u�}k�̕0=�mY�.�������>s\C�z�h��8v띛�g��c��&����[����nʬ~����4	�^�@sۑ0�\Æ,��e���|����M ?�u���\�{t� ����G�.�ש��	E7%X׾Vw#�`��`osn���(Oc	�*��'��Np����Ł�)�o� |�y��)��+ ����^�{��k�+���X.���%J� i���ip�݋Al!��kOn3!n��c�I$���L�GM��crX�۫q����z���ޖ�z�I*G�j�7x��%LٹS ��XҺ�7r�7�X�1���"����`��40�M��:+��"k)M%�a�5gCB���Q�� ��0t:��~����t��'ZCb~e��<H��4��P��Hz�G�PK���)���2b6D`�E�L��t�8HD.��P��t�SC�8ED���D���01�a���9���ħ��GI�Ѿ�3U���࿗}��A+�&��?&a�tġ< ��1�g�aU�d�w��a�0��hLt��`4�Y�kC�Hn�RƖ;:�!���I�|�~��ٶ"���TC��? �����QC����^���+�S������/D���LT7�}�U��{��p� �i�qX~�)/g�,�|`k\�t%�'y�t�;��2���@�rK{�Kq������w�����Jm"Eнq��a`LkgkS�{:�gf�tIv�;5�w4�mS���Sn��U����X�w�%�����9h�]t����Y���7*`���W�����fV��e8QQ�`������fJ�M*`y�.椛����7��V��V�"�a��vmPdt|B�*h�$�BP��u��g!�]����ͩ3w�2T����`�����m���~��WV�Ω����1ĳ���)c��^g�N�!�0�.6�/n����Ns�w?��zp������QHs���|�GDM�
mE`��|�J��݋ �O� ~ۗ8�2[e-�A��,��Ձ��U��ȵX�vXδ�Z68ꊔSrU�$���������� ~׋ k�J��rJ����`ndZ�{�.���xr���{���#�a@!_�u�~YF���}Y`�a�\�1[%���4��A�s��5�ý+�G2u�b��Ş�����	p1���ڟ.E�a�구��"Y*��i���e�E��X-����F��'6���]�z�&���+�V B�nM,pZ�n8�9��Ny]�Wj'q���q��|�GCd�pt��=P��\�x�؛�9#���'�H�m��`ݲ��c��~�������,2)�[9u��5n���M9��;����:�\��&�WG+��cg]3tN�ݩ"?Ͷ�x�x���/�;]�N�.��I��\�nK{�u`w^j�7�� ����)#4����D��`O����ULz�`_Z���p���r�T��T���=���gwe��ݺ�;�5X�B�R�m�&���'�����\�0,��`E���~\�r�ua�\&�ն{1]UR@����pDA��v�p��ֱ��n��W��J�MU0	�u��>�K�wWI
Ъ��ε�4��JY���D�k��s9U����&��L�'���EG����U0	�u�}6�\�0%'.nJ�2�@������7��Vu�s"�`u�f������/�|`z䩁d�S ��X���߽���/��Ą�V������[TN��:��?�����w�9��͢&����<�Ͽ��j��O[��_�{�9m�c�JE�͋��3������Xך��f�J6�
m\�����Ń���(���5
j�)D/�>��\��6|ɪ�2՚! ��`_Z����S�j��N��8��Z��QR��J�;�5X�'���׀?kŀ|�y7���9묮�s��n# �m�vg�k��l�S�#��dn&4u���fYs$x��_�O�����	-����\�0%'.no3s3���Z�0	-����\�07���VQ��58���`ow_�j`_MU0	-��xW�j�9ErU��{����Z�3v]x#�@�� �R�D4 %D%
�(K7� �l�~����U5s��� ��u�ov,Ξ����?W�y��h	S�%FƢڱ�l���r�v:�+�6͵�*.ݙ�t�ɮ�4�J6�
mE��,��Ձ�{����Z�Y�i�imBH��޷� �� ~ۗ8���$�D��b)y/)QR��J�3��V�"�g(S#}׀v�ŀ5�nI�Vi
���p:y��� o���x�:np�VV��8ۧR�A�+ �ݖ�^,Λ��ls�RJ�
��b=ݽ޻�;�}&� m?�e�~|4mA�VQ��tj^c��k��#�3J�V�&���w1C�i���؝O,k�$J��A�����(��:YSSͶ���ϣ��.����� �g����x����ݻkc1��+��^�i�h��\�-#ҝѱ׋+A�v�8��u�n��^5���a,C�8�ֈ�;r��cId��,N���d����;������w{��:>r����$��Rmڝ9-�x$.#WE��������u�f�۞̶�o��7Xz�����S�iS ��`zFۑ)#�DP�%X׺��CS ��`[+��E�������%���]>LKu�l��\�0����IDm�$��fn�w6����`n�5X�D���ڄJ�����0=r���iS ��`~�*��5{�:prRR
B�4G,M����{^@3:�7g˖��<��]�F���V�Wv�z�� ols��� ޻�k�D'��EG����j��� #Њ&�*���քv	��(�����_�(��������b�<��;���q�q�N���V���e|`z婁lҦQ��\�f�B��fn�-��떦�J�f�;�Ѷ��Ȣ(mIVu���� o���'��� �]k��B,�Ak�g�����}� ��O��+ӻ��ۛE��&�3�v��}[�ۂ��m���O��'����0=rT�;�
��@��p�&Ȭ;�,�۫��U����`b����$I`7��M��_!(Q�FD)�ι���,��)jZ�|A(������ULKu�m���P����?�պ�]U0	-���0;�uX��r���l^��rJT&�۴>��;��X�ڻ	�5�ࣳ�@s֐�kr�F�Q�)��:�5_ n����ݺ�;�uX���VQ��q��7X�����S˪�%���6��"RI$IP�r���V�ū 7[���`��W\�L��� �j���	%?��O���� m�XJ� ���?b��)
?�DD!D�_t�h��칚��3F%������Z�]��9\�+kf���F4�B��ҥ��7\L%գn�c<g����v��u��)J��9'�{}���U���K �ݖiu�-N:E�nJ�;�\�L������ z�,�rM:��٧㛚�S˴`[�-|`w^�>�Vָ�8ۧR�F�,=UJ�o��}ذ:np�ـ}"�Ů:���ܖ��Ձ;�u|{�۪���wʿ�W��W��@U��A@U�W�P_�(
�� (
������"�2�"�2* �"�2H��(	
�2� �$� �	"�2"B�((*� �#"�0��
�0�	"�2�	"�2��� Ȉ *B��( �@U��A@U���������
�����qW�D_��(
��P�A@U�h
��W���e5��6��#d�� �s2}p��    @  :��@     �     >     
RUPD��I   

I �B!U@��
P@	H�UH ��%0      UA@3 4��>��ܽ��=���oR����'x(��\���x�)o�{e�wJ}�� ;ʖ_}�K�� 6��<nn�پ| }<�S{}����\F��,� ��B�x�\�c�C����*�  UP  �x-�3�(�g  8� � *� soZ3��^ �� tq � ��    D  
@hi; `�  � �� � s	d@� � 	� i@ P��
J  l h�6`
@ {1@; 0L � Y� vo�4���_������Z{�g�j��O��ON�� �����y�����;�y��}� �O[��x��ν�wŻo'��� >�@
  6 )��݁�44S�� ���}�����&��&S� �ﯴ�|���7/ \�����=�-{��'Ӗ]N-��[��x�{G� ���8��r�����9��{�|  x   P �������{�W��>ν�>{z���Q�=nmڳ�v����y�^vS�}���Y�m}�Z�  �w��y�^^��Hg^�[�Ӌ^�5紼���� O�����+͗��d���g��� z����J�@ ����ʛʥR� �d ���R�*S�   ��U*)H  *�J=�R�@DD�iJSH��F�MOQ:��O�������������w����"����_��]UDQS��_�"*
����*�TE>���z���t��F���$h���D�&�
㎆�@�
����������)���xNs������y��ɘHS���|R^�(d�a�JJ*K*$�$a#1+F���`0`a�� ��&���H�R�J5��=a�*za�� L�$��!�#XGH-cA�A=X�����T 	FC-!D���x^i0�=�20����� �j�83\����g0�����58BD��!B,F�0�X�����k���H1Z@�HEa��0"A�
�hA�F�)�!��BB� @!J�����!B��H�V�f"BJ̉��'5���?I�1�e	B3�r)s	��n��
[#*d�b[CPTy��w{����H� �D�@b�k��
���!\ DC`#E�8ݟ�l��H�B$��,�#P �"�������8�J�"��~#�mas�5�n׀r�~���+����x�@���CË)�)$&p� э2>g��7�ә=�5��X3��wy﹣�
��1��8��7.sx2��np���Y�f���F��
al1��x@��p�0�F�K�)��\�sIL5%0�\֟�<��ؑbG��<|B5���S��!sy� ��׏ ��$�y�х3|����&�4�ѹ����~���7w�m�l�5����>�����|�}}���7������e2!X1cOW!BB\�\�猹� SR:*�P�/��M	!?RR�X�E�,9������+�HD��9���<x�
�7v����K�<�g8���P��!}�K�=b��\<�dg���V5|93���������A��)��^yIn��O��ʒ�I7��]����f>^�@�%�ea������(��0%2�P�%ap�A��j2$Zc,#.�.mcl�nܻ�Mv�ᶝ���$�/��C�&�t�Ǜ1��i�FF6�bY���	��i��=��w�~����.{�-�;��.C=I}?~��Y�JHIH�R{?{��B�Ò�"D"��)�̗�� q#s��?s�s��y��ig����%��wd?s2���%Q�[����C6����f�LÄi��R�BB�0���r�]��g���²�s��<�w�ܞ��ޟ���\���zK�k�\�fq��y��Iv�/����?���g������#+���y�=���Q1��ƕ�j`hRB��L��2RX�L���5%Md �X��S @�vS$V0%eraw�8<��3X��B��,�H�Iey0!+�#M=����B󑄓�f��g��۟�M`Sl�����0ْ�ws݇�nݶN�{편ί�{�����5�&�z��9%������B���>_�$�9��5 �	F%d`4`RR)4�H�B���R	D��"�����9������8`K��[3p%�5��C!LZ`�0e��۶����x��� �"Dc��9	�4�"m8ۜ�l��Ky-�ᴘ��HcXX�$aK��f�\�ww����N汮�汪D��'�᰸4�<�睘|�￳�u��zϮ{�ӗ��؟��U�0yə��bxCE����4����ƑjB�Y�{3��'�<;�����I� ���y9���?y����o����cn2�-s2{)��e�%�KB]3$fL���<e���-�L����y��.0��럿Y�?O`B�e V$�!�)�Ou����u�U��f���r5 �w�w��o|��h�,`�%p���\�%��?���}.�{�w�f?�������4�4!�V-%!u��ɥ�I1Ƙ��.�!7�:�K�r�
����I\�"ŀD��X	7	'��s|���Ç��fgw��?_L��$I�\�D��~g�h[��ic �		������w�FdJ0
@�$���?@����4%�o����\�?oc̬rX\�cxʘ���kBfe�I0 YP���-�
D�EP�rBe�\ae��@�m�C��dd2
r\�獄�V��\����y�q�4��S�����$�@`���@����7?��	KZ��s��,�,I(E���!R1@��R��h4`$X�1) ���\(F����LF`�
�*��"X�L�@b�B!"@p"��X	%2«BHV)U�X1XHR5��h@
A�A�@�c
�V�,Z2H�$`�C�3�Vۆ�Tb���)���1 F%(����%�T�)a$)�B�R�4�Z�H�M�h���f��Rs���jq�,є���0�q��b҄)x�L9��RbS�&fa\
�J��D�A��)�nY$$�	BH��k�d�l)C'��ӓ�y��/:l�^�����|���	F@�,�!Cd	a1���v9˛K$�C[�q���$i�a��3��fgA�n�}���"H��,����!N2����9̞g.�<45��������e�&��.y��\ԗ7���IA�,��*B�!����u �J��3�0�JI)�
���f����$gi��y9�W�R5�"I�~��k�?m�&m� O<�=�36~݌[�5�7��?Ƀs|fx��y��.�2-�^�4��}<ba<$�,
�!H�aX�%P�`Tb�
)Q�$��!��HB�	r��#
�Bd�!
yfl��<L'�H�H�8 E�1bH*0k�����]	D#�@�W��B��Q���J�l
I0hTɞF�@� ��䐦<
x�eaP��7���Nra��x��)��D�@#��)b�
B2BA�KXX�(@��l�\�`l�,�`��5�qCaRHQ�T @�H��X�X�#@��bQ�� U�<G�!�y���~��%=���ď?Mx��'�Jc.�N0!.>&�������
J/1��]6~	'�Y��>���$"P�'�
����o�s��Ƅ��Ж� ±bd-=&9��C}S#L,�h���X�@��
%c3���޻�Y��6�j�����@�H�IM;f�f__ߡ�d�y0�H�Ri�	�W����))q&xrg��pOXd`���!4�"Xa��K�S5�����r~$���9	!O��L�ؒw��R~V- &�S���U(��
�²��8p�����y�/�P�X�H1�)@D���"��C���oH�|�I$�ie;����)�*D(~�g��3�o=)��ǥ�������F$�{���}e'��'�2$���WB2E�1 Д�����6�'��s7?K��z�<HG�sy��i�A�D��jH�#F c��	X�����yF2G�8K�W)�szK��$�A��AH�Y-D�L"�"1�� 5�Ղ�D�#��4�x~#%��2��$��1�H�H�@�8A��0�V�ο�vߎ�_��                                     ���                               �     >�                m��   [@ 	��                                                                  ��     ��@l�rWU��W�Ns@WUK-V�ʪ�T�ik�k���7bC��D�!���� �8�km�	 I�� ��ll*�|m�l�� $  ��-� m�H��@ �I��`�u��� �lm-6[m��pZ�    -6����ܦ,k{m��$`m�m�[u��ۭ[q"��`��-�l �6�[B�� �`6�B����6�h��[Kh 8���� �U���.�����^e������� M�m�m�	���L�`Zt�@V�J���n�ڪ�� p�J ֊ �nٶ�	��j�7bR^�J.m���*��U��6C϶�v�Ͱ�ɥ�v'I7V����<�K]UUҼP �`����|ڳkA$����-U*�Yj�]�B�5P,�*t�&��Hg�5ɱR������t����u��h&�̘��ʭ@Uࢹ����!�+̻��U�jj������g$t�W]�(&���9�/)sڱ�W���ܹ!��  p$�GS�]m�۵�$	  mm� ���j�'L�m�{l�l�m�f�e���%^�$Zj�I��ù  :M���Cmͷ���j�Xv� +j �')��մ�n�2�Kp*�
�m[UJ�6��H����'D�m�  �q��iۉKm �e���d.pf]����mm��`H�j��m��ڔUu�B��u]@J��d�m�%+�����l��2� m�6�M��@m  [@-�   �`�폆� h m� �R�$6�m�  hm��m  ��@��.�X�k���*����WeiUU	
Z��j����rM���7:�`8-�m�]�m  m��l1A�h�U�++X�ll�@mZ����펶yp   �Kͭ��   � [I  @   im�B@�z�� [@-� ������ �     m� p�� m�mm    � 6إl �l�8���h��	%�ml����͵��g�jC�hH  �h$m�h0�	�m��I  $H���mw�`u�������eb�3��A��JʁUP  km�n� 6ض��� m� �8  m    6�m� 8  6�� �� ��Ā��I��  h	8 �� ���lH $�&H��irm�r��a�C�m��u�cv�  ��[@ $�	   $�� ���m1���(��@�UT��#�8��m��� �   ;m�h	�G@5�   @p  � �ʹ��m�mm�Ĉ�/4˲��U*��4��U�        <[V�{ku�5��q/�X%����4��-Vӡ{n@�k��� �u�Nץ�V�-�����^�mmp I��&;gF��\�q�Y��F�<�[���C�qw];��+���+�^9�gCJKUm8v�M��%�T��p�9_��o�N�a�Swl�ʼ�]�]I��\&ա��/<Ҡ&�Խ��UcK�e�g�H]e��Xډ�#�,!�m�9v�+�f��m�m��9m�J9i�6�/iBI��lڵ�8Xi�5U-�� �[@m��S���I�gQ&��z��l���R��3��m���m���Ӛ^����k��� �M�3����f��]�:�(4U�����;h�z��m��R���Vx�}ʅ����(mT�cu˵��Q�Gj��.�e��j�
���Heʅ@v��6iZ��&�yY	T4ĭ6�m�z�vTl�a&@��{6��ڢM�����W��u;GK*�qU]TvR:m*R�2�JB��Kl�ڶ��6�� �:��ۣԱң�iYn�Ҷ�`   %����M���W;8c
g#�9�y�@v�������u������⾇�scey�ִ�d�ݖ�"�TyYHq��5˹򔵲��[Tjz��?J�,S۲�s��mU�wlM/3׎A�$�j������6��0�r���/\F<p�y�a�,`(�k��$H�ͮ ���K���6F"EX8/[�յ�d6m��6�K9�U�C���U2�5v2�jjW����3B�m��^Z����cM�۱� DM`*7M���Tݼ2۰�M�UmWN�#�V`'e�G�sUu� �l�S����] 9m�]6  [@   m�4��v�G�G-J�Ւ�����[x�&� ֚M��KӪ@ �g]� ��  �`   [@۶�8qUct�]����]/�}��UQ H f� lm� [M�m� p��m��ŶK��     8ݶ   [`�   �`-���[@   ������� _Y5�m�h�&e�j��U^[Ý���  J �q:z� 	  �ض��lm�I�hmp  �c�����   ���� �KMl��ݷ=�27Y)�^��i�h��� m2[Xi0-���� �����m��@ ��	h pI]U@R������=@� ���m�-�h �]$���4�t�l�8,�Z��E����f`�[gMuB9�^�:2M�	cQ�x{6�1m)^��@V�D�k�[mUJ��ó����I��`   $�,���Ԓԫu��&���-� %�������x�5lm�m[���5�G�E�6�m�v��6�դ [@^�H�vհ  ZNٺYx	��c`�M� [IpqS��oR��M�R(�EPUTg��ڝ"��0�+�T�	6ʷ�*�� �kH���4\r��0%��ak�DX8{}������M-���6E�p�mz�E��k�M#l[hl�c� 6�^n�p �gkM�\s�6K��t]Q�m��p $a��Uu��ާK(�i6�I�5�N���(n�	��ۜ6��,Nٳd�T����H�I� snۭ�7��ge��)VU�����@�b��M�6���G*������#�m�LO(�N�nm��*��­�U��վ���e���fHK.�F�I/M%�r�D� ��-���^��ӥf�����)L�U�25T9eZ3��s��bR�'d�V��gL�ț�VsP5� ��]5�	  �6���v�$��k3�ª�PR�Q�sH۲��mv^h�l�l�H�Q��nGg½5�j�5�F��`F.�W.:鎚����#.[��ܒ�F�t�� ���Hf�51�F춭�Y�����;��^�h4���t[Gt�/�j�n٫i�ѝ�0N�mٺ:�I�l��Vq6ԥ��Yg`�������6j��^�M�-����M� �� m��l ���f�||����h ��   	�m���� /�f��j�2f� ��	�Z��l�   �m���p �"۶�^�^&�:� �j�8p[Km��m������X [Au�CI.Զ��t4�Kt�Ic��h�Dnt4P!'M�[@�c��kݔ�p	"����;R�Vd���v�,�[\$V�UyZ�mzLM��ִ���ͪU����e�@j�A!í�) e�V�l� 8Hm�Tdm�  �p�KD��T��f�� ۴�m�o��N���+��s;3���1R����ɞ�6ҏ[R�<�f��U���ȶ�J���J�ܤ�U��6�6ۛV�8[���ѹ& �cl��n�
����;Uͪ�;cW�I�Uq�*��Kp6ٻi0a΋u�m&�4IE�{cm�n���*�^Ɇ%YWղ�K	�K�Zn����� 7E6� ����i $؍jۛV�9�'�MͶT�猁�`݌�!i�M�m� H   6��m ���#�m�   '�w�[v�ީ%i�&�wf���*����AO�^"�^*��H������UqB H��0�0BE��$ 	������F��)��T|P��(.�LU��  s��x�AX�����Ȟ�']H@<�O�'}��4����_:�J��t聩� �"$��Q��(���P�OU�C���u�����a0P�W�����~ ��� O�D�x(�(�� �&�� �'���<_�~`!�S��#�����qS�/:8������*⊾0�Σ �*{�D����G�11~^�-}F��Ȋ$��N�@H�D`�";�=@����>�x ��^�!� �J��/�P�� �#�+��*U�0u5�@Ƚ}�A��X���#(J�JBEb�)���#��?>����2�(8E$�� ~ ��h�D?�$
��@��WP
�V"���?���TEAW��b��ꊥS��
�
�lJ�	xDJ�T�'{���       �`     ��  ��             �`H�itɚ^ok��J�R-�\n1e{E�/#�dɨYZ���bl.�����u+>|�֪�v�v�PA���p�G�Et��1�E�N�i�+�]8��IƋ���ϐx��R�q�T�6��
'�*l����ۚDKD(6:��v�Ԇ֬����'�9�����s���,xr,]lTq:��^窶�uD��l�S�ΐ�q*ۢ�E
�]�j��WURM�q��ummX�I j���۔���:��5�ŗ�ϐI��*�2���iUI�%Z�j�b�W��N����-�6�]MѺ�L-�h-�W�ʵ�յ+��r�Se��x��ܜx���=��I����B�����Biz	��n���#���vH4�=�:�><md��Ǝ����1�����y�,����<���GZ]�2�8w7�铍�\�����iT��za��������|=N��$mZ�k6Ss�b�华1c�#d;U�j�-�j��kg[m;���$A�(
��^�H�nI&�@W[UWOm[YɄT
�����y�fٷn���4J�9���)�-K�I95��&]Mn�t�2:���@�K=� *�ݵ[��nOe^�˻I΁{nڀ�֪{ 0�[g[�]�f6j Ǝ9c�q[ֹ���*V��&������&]v���أ��ƥ�y���D6�sg��v^�M��"c�B�DY�$ҖZ*����`u�0���+=��4/:����ۛ=������-z؂���yw�`�ᫎ���cPW��&x���B;��M�y���5'c���r�v:]̓�sc��6�Z��n2Hƪ�+����+ve��=�L���T�y�hہ�Q�r�[u��@=8�/*���1Խu���]���w'��q�CS�A0(x�8�(��%�A��@�q�"?��{��޽��{��o�m�d��  mM^��[u��l;ٰlqp�r�4f�k#[3�����fg��jË�hq.z: ېX1�fm�t9����.�Q�P9r�����i��.[�z
1V9ݰ��vٲ>Ek2n3�� Z�[Y�u]�
7-�n�7�6h1�{'U�\��'�z��u���4��{���<;7�m����ۛ��(��fKrKf;/=�_;l;q���=�w#���Gm�O|r�㍻<탟s�K������O(�3�>П�����q	90X�D��/e��Q�=+�,��閆�j9%�����	b�zW�YS���[�k'��I1�8h�w4YS�/0%��M��R������c �T��m��	b�y�\J��W<�ڽ��y����70�n�. ͎'��l��;u\�����]���&��d�Y�$�&Lx��"�I���>z^��$�� �T��gCK��Fa�8���I=����߂�V�@s�B�S���Y�o�9$����$��zT����gr�V�\��׌��x������;�g ��֭��@�O�5� ��h�h�W�^�s@��Xɉ90X�D���=�=o�8��p����U_�ÿ�e��on��������5���;��b��a�ӥ����8��%J��d�/�������`ʘuˬL���O͹�91$�z�w4�Y�^w*�9u�~���A�W�Ex(�	e� ��x�|%ꤒ@�$/�V!F!"U]ݾ��䓿��������IE$�@�ܫ@�׌mx�=mL���˻Q�0���ؓK^0-�� ��0nY�wuԱI��M9�$a�,I5�Ӓ-c���,�=�ܖn����nn���u���r��ܖ0-�� ��0nT�����g,W�d�G#���fʪ���H���ˀm�\���o'&!����^���̫�$��9��ɰ��v�n��Ŷ]���<���<���~{��Ҫ�Z�e���)r���-d�ۙ&$7��`ʘ�*`K޴8�.��vЧ
'��ه��S�1]3�?���O��h�u�����ۣV�e��� �i���gʕ/�$��:��A)��A�RI4��4	b�[^0	eL���˻Q��Y��x?k86�q*����E7����Lj��Wy�y�Jܓ�p�o y��������Xzյ��@�g��YS ��L	b�K^0/��o�$�I$�I I&�P  %��KtڇW
ׂ�&a����c]m��k�����-�y{}�/K��N�([Ã� &��!xbSpnzLn
�B��Wh�����1�4$�������D��\�t.;hdr��d1���ώv��ڹwm���.ޮv��t!qtkmv�����nji!�<�"�;[��x��; �:#�����w<'��Ն�ڝ��-�F�ʹ��(�ŭ�)N����\�,ܱe��ۛ���q[�@�\���F��`��{���B(�y��4�)�UR��� 8���������'���I0Cp�:۹�z� ��^����Q9����	I+�� �)����m��?y<�!Ll�&8)�m�4�)�6�. ���RJ�_��n�yz�̷Ls����k��m�[�2�8�q۷�;�Wk!!1<��چE�s�o$����|���eU%�`I���5hf����m�撪��RV�Fbh��@x>��7�sy$�~��x?k:*��E��qem���nnf� ����-�SX���׌	2�^����-i��n�D���"��8����׌YS��G�j��r�Z�&�Q�m���mʾ�~���Y*�Ք[�w;\�h�K6���������y2q:���iו�Xi܆��`ʘ�*`K%4/.�TNG�q�D'3@:��mʘ�F��`zgd�5gp��y�$�%�SX���˙�b�n�u�hwD�mC"�9���h�F��`ʘ�ʘd4��� w#yn�Z�K*`ۖhzS@��TH8F9�I%&mI8]t�'����e:��M�I����6��r�~S����s4�Y�ۖh�F��`I�s�gf�Xn!{w�?6��Uv8��r�?=���Ʀ(E��#�&�~��@�k�,��Kr��/��w,G%��r��K*`ܩ�ffg�~?~����yM �֌m̏�h����~{�EnE7�À�o���Ϳ*q7f�@72�m��[7Z7cղlq��1k
�7WFGN���rLە0%��mx�%�h{���#2~���4�)�^�� �T�,�SlɻC5b0��o-�C�^0	eL˕0%�����?��5?8�s4�Y��T��*0,��L�۝�;7��q[�0.T��*0,�� �]��} �b`�
{ӻ�=�����  H��  l��[/HmʹU�u�bt�+B��nxƳ\d�ح;FF㳴���r,��]w>8��U4�(��M2+u� k�M$m\�]ۄl��b�=v��ץ��Vݞ�ED���ڐ��A쐛���jX���D�����4��Ó�T�� U�9���v�K��2ŧ�Gh�����=����xk-�7%�V������Wa�ц��Ҙ�Fێ�V���L�9Y��n`�F��MáŢKS��K�_�~��K*`̩��e��ܟ�s �Ć�[�s@:��oe�^���U�܄xG�iܱ�K*`̩�,T`[+��ǜ�Ƙ�ӂ�ɠ�Y�OUF��`�������9ov$����ex�=eLٖhWhI'$�~JbP��`/<�b�ۘ��m;)v�=!�NiQ�q[�]�[�7��4z�h���{,�����À�����6��Xnm� ��w������BGvN�� �*0-��L�۝˃y �B;y&lʘ�F��`ʘ{����J%D
d�^��-��K*`̩���n�_ݼ��n��`[+�,��[2��Q������C�"c�&E #k$�cMb)^{/l�mv�l��C�<���t�'i/-i�m���~�oe�^��-빠{�󕘓pR94��ފ��Àq�\�����j%�p�����w�q�8?>\~J�Ї���Ģ��ǃ��	�j�A$B0�	!)����X)���)R(C��s=}���"�����i� �-C����ڗ���s�A`� ���������L�a��w��mX����"L�䣄���s 45�	G�p��L&O6��͂I7G|  ���bo��'� e�D��	��XQ�<�xt'9���B>�F�z��ё���<X$R+e��T�S1�jpC��08"z��O}8��DEP"�ġx�� 9 G�T�N�Dh�+W���@�U+�j
����y$�{ӻ�'����X�0���I�@��s@:������U*�C�r����6��\.X�%�0Y�0%��	j����JH�x�"��	�o!
Hu��4�ボf�Ѧ����m��������,�wB�e����M�<���<޳��X}�4s����"DPQ�BS$�<���v96 ��m=�*��������me�/u]��p��<����]�E7�q�8�v�3t�F��^^�y�J��q��"��y�Y���� $HT�U䊪�����NI?{�}s�̙76�͗w7y$�R��'�����?���������k�{��II���F�-��5�CNʽ>�[�ͷ7I�F��n&Q{u�Ϊ�Ç4�,ܚL��s0��I����y�g y��T��"��;i��,XcpN$�u�����~�dSx?k:U��cŔmz�����&-ʘ�F�Q�&TV7��294ۖhzS@��h^�@�ܴ��"@�id��n�~�p*�$� 8��m=�I�}'ow�����  �L�� nj�ƛ�k�vMkôض�]f�\Pi�k1(vJ�����]t�۶�8K kq�v7*7E�NӹfP��o	�Eu��ع^��9�r)��M�օ�q��O=:wS�x�rͬ-����e�I�ă�5���{m.��Ӯ�ۚ��
E؞�͹#��';t����v�Yf��Y�q?��?=����.�W7f�K1�N(�@���̐�wM���n]ɓ7�l:�v���-��C��mˇ�#,m;ֿo۷m�������?4�AI���>�ƀu�4��4�)�ܪb�o�i���`ʘ�*`K�F�<9�mc#��
G&�u�f���M���oY�y���\Dd�����&�T`KU���Kr�.�I�cp��87���oY�nY�w�S@��T�ԉ&19�]v�Ν��S�@8'=��g6^sEL]�z#����O�f)��?LdrHh����,�=��>���`��pji0��.�5ɳ.n�I=�N�=~��>�P��a�O�a�������=� v�q��@S$�=����-����h�,�=��&!��rbƜZ�I���� m���\��|"��L�nne��fi��{�K�)��Od��6���I$��r�^����`d2b�Ƴe涽��,۱˘J���6W;\Fӣu����?*��lS_�������?�7|oY)XK�g�yc.+7FZ3j�� �7}*�J�l8	rL��{ҕU���y,W�hY�w��v�	&Àv��2�-BT�
��H���@���V�E��b�"�U�O��(�'�g�@����:�|"��O�&2I&�$�d�8H���w���&�h��1�ě�,d�8�ۖp*�d��$��o8�_�0��ˡ�-]��E�r��ܙ�����ӛ0u��8bv�&��{���|��Wձu���g�_ ��p��D�XE7����+���Xf굗�|��w�K�0���g }����<��*��
A�#�����W�|�ۖi�b��s$�I��<�/^;���xf���pJI+�"��9�_ ��p*�:���V�X�:�|�/�>���t靗��e�Ze�3� �7|�$�.I� �Vhٙ��|�'��$әX1zv[��$Z��f���.��i�Pm��7����qa�Ě��?����r�� ��ؿ��/����E�m��wwt�=m�諭Y���/���g�_ ��tJ�M&����E�7oss��o��*���̟}����8ߓa�n���m��iw�w�*�5�������ʖd����j|
�j�sV����|��pRU�)�O������{���$�{��=����  �]  $�u]�6�L�&�[/�\�Vc�;)D�f�N��=�4밻�4D�U6��)��i^@i���X'�Ƿx<�M�9��ncH=�l�6�j�;�������t�uy*��ۮ�g5*�Sۮ{/o����8l"���Cq��7iP�qs�[�K[���g�J7l3�v�ZVGN�G�U�N����c��3$i����Q�L^��ڞnݘݻpWK[/�>~�����v�Z�o��_1�9���Zcp�����zm�4�������a�8�L�.$n�����m=�UWc���M��~y�RT�����}�6����I�_��hl��~��Wn��E7���톆�f혮�o��䪒��}���}O��i��UUUW&�|���,�h7V��� ������[�M�Lr�;)�{l*$#�G#m	H��IR3�QB��X8R����J/@IrGK;���{���v:��71����H�������-}V����U$�����p���e�m���t�䓽�{y�H�E
�H�b���@�@Ѐ�q8`�Ju~EY���rI.9� �OzURWg�2+/��75a����o��l8o�8�UvI�K��^��$�0�6��4>�_?�� �)�~|�%R�$�\��čݽ3B�w8���UU|�����������*�^��Cd���E��ʍ�΍t�m��zUv]��n��.��Oh"+m�
n���˳+�\�n�$���Òm���<��XE7����-[����b��\��w�R�Y����8}��x��tT�]�V1\YF�f�7wsW.9����6�ﮕQTR*�(pH!PP�Q���O�����/nhr±��4�"����T�]��G9pm�����\��p���e�iwY�ޭ��>\J����.9�������%t%՜\�v�H	��3�]^-*��Υrh�uf���w{�|���q����a���$��;~y�m=�I%���nh�/��D�GC�rf����JI%vE7���\�|�%J��"�0�q#woLн�� r)�~|��$����,���r�>����/��-����+/k/�J���s�pI�$�����<N����	H����-R�`t@��<��y$��;~A�vгv�W����o��|���~�?@>����[�s@��TH89�4����d�6�\q�B�M���@�tP=+W-�lJ�u�:���6�5a������� m�x��D�K��G9p'��3V^^j1a�{�� �f���R�$s�#��o�:%J������4�33L���7���\~|��J�]ˏ�}���<���[��#��$��IU,�����}O��l��*K䪪��ߗ |���[�w������^���<�>��U�RI,��7�}�ܸ�{ÒM0=����s�p�n�8�F,��:B�<���I$!�"V����0 B�8����F3���	�Y�{O �( �����o�R1O4XX��0Z#�|"�/��Ī��?{�� ?�|               l              9��K�p�I��R�e0,v]:
�H��a�Ugm[�6�����fgy�C�8mk���pYƔ�r����N�S��n*Ǔ<�F��݆YM���Wk#sk�1Oc�v��������6䮳�^��ڳ�LK:K�n8BJ}cp�;�gs��f�
�zؓ�d�A���l��v^����|�� <p�+��kj��jM���&�@�8ˬg�끺@U�yUT�;@pmum[X�a6 j�MM���7+�.�Ty�`��zT&A8����� �5YY@�YsՎ�@�s�܇O1���gVMMq��F�a٥ӓ��y։B�^�7��5[@�ۡ�39{Y'�4t�E��MZK���в�[�s�g�uU'd���p��C�U�;م�r���mc&�������pq�vz7��<�*���]�p�"�ۮ�UyĪRve�T�k��s�w<뛐���d�k��g�L��籬8�[Y]�'6�ms�b��mO�eA��7����E�8�H��-p�v�Y}"�qB��0��Њ���'b���6�ݶ�t����3e�5�ԭҢ��\�.��Y��&�b� ��)Cu��� �wQ���Վ�rKӠv�v�T�l�%�V�ڷ<a�u�u&��)�Vⱡ�Dh�q��u���s]g��U�T�V �m��1����P1m�����6[�� fi˳�1K�:�)V4�q��i�/mb���	ǲ��6+�*[�% ��=`赚��:��n6�Pћ1z���@j�������Gi��@s̮��
qF����DV��$f$;�z���Ѥ�5Q�@�uR�Sq��+�*GE۪����^+ms��n��'M���7mmlk������; F���<u/v!V�����G���#��ZES�U���"��S�'��{������������   �  ].����ͦ���5��k�ӡ����nr��)^�N�rktO!��Y�"�N��5[vґ���5jT�j�7c^Ke��D��6�=+�t컮�On�����WS���{<�DW��;3ۉ̠YŶ��Ӝ�n�ٴ9熺YJ��O%�mmƍ9�\�L�Μ��$n�4t��}���r�y��#\�~���w����xo��U�.�+�R�[R�+mb�;V��v;a��l�99-�X+���wsX�q�70�,��?�/}�M�up��W���&p��r���B����7�m�]�	UW�UY��O�p_�}� �f������%�5i��v�W�����\��q�%�Y��}��}�.���meA�����\+�$� �Cx���W#�ˀqM&��2�Q������7���s�#��W��=�*PjLǒrA�e���v:�=]���d�Z�wI�6..�����q��p��'�}��s@�������W�� ��7���+���Y��[7t䓽�{9��?!E�F��� ���0 .�@��\�� �p��>])]���������̼���N\s8���$��s�#�p�Mf!�n��������r����\���R����}�O�@���PK�S�S@���������������Z��5�2H.A.2Zv�,�v:ӳnt�Ӳ�뎺C�ҫ�Ɯ�>�ٚ�4���@�"'&x��8o�8��������}>��}Z��Q�j�wwt��<�T��#r����\���$���a��bna2(����M޻�{�30��T��UR��&��.9��ɾ�˼��6�hn���I|�$�g�O�.�7�v���R��U�$3@��K��Ds�cC�4�� ��~���]��m�M�w4k�d��HbmG�q����9��MqѷnZ{q3��ڞ��vffg�Ku-yM�m5�<���g ?y����%U_���"���D�ݽ�2��� ~��J�+%V6?}��|������>�|�������g �X � � ��M�Y�,���\ۼ|�����}�� �`�`�`����ӂ�A�@,l~Ͼ�8 ��~�� �`�`�`��{'��i�Hn�]�8 ��X*d����pA�666?�����|������}w��A�A�P� ?���#�j���@#�A������� � � � �zl���1�Hf�7wwg �`�`�`��}���� � � ء����￿��A�����>A����ϧ �`�`�`���~�f]�nL�����-�
)[��q�7�ۘ��ь�#��v6��ھ�nl}�9�u��������w6667����>A�����Â�A�A�A�A�����G� � � � ��}�pA�666>�}��fn[�3f�6Mͻ�� � � � ���xpA�#�0� �l�������lll����8 ��~��"�`�`�`���Ϭ/��ni���Y�� �`�`�`����ӂ�A�A�A�A�>�����lllo���|�����}�� �`�`�`�~����nL��ۗ3r\��� � �� ��}�pA�6667����>A�����Â�A�A��A������ � � � ��Ja�M7n�ɛ��|������}w��A�A�A�C�B ���ߎ?��`�`�`����?� �`�`�`��}���� � � �����{���=��?��  ��mp  /��o�}��&[.]��V7A���j�����W\
���!�i����p k���l�llm�2dkRu9D��v3c�i��-�-����wOnd۳��ƕ�Dj�� �k��@z
�g���fG
Y��x�L�1�@�����U�]�46�ӗOn��pH�G���a�}���f0t=�B�.Z8�{�����[F�j��ɐ�qC�v�E����0n�s��I�z��^s�ߞ��7�Ϲ��ˬ��x �����>A����ϧ �`�`�`��}���G� � � � ߻��x �s�>�3M�Cwl����� � � � ��y����G���A �`�������� � � � �￿��A�666?}��|������>���i&M2nn��>A�����ﳂ�A�A�A�A�w��A�6
66?}��|�����w�N>A����r_��ɗ3I����� �`�`#`�~��]���lll~��8 ���>�|���`��}���� � � � �����2�34۬����J�XI'.�T�*���|~��ﳀ���ߘ'�t��Dn���O9f���d�O=�ۗ	�d��s�=k�Ǐ-���B^NX^Xniv�f���M������bIW���"���x�ưR4��NV׳)Uy*���U�O��{$�����'��������v�f�� I�� �7|D�U]���&p߃<<��/n���ݽ�����6K�#{�o8"�Uw����	F�$CĤZ��*�� ��M�j�*�R�R$���5&@1��wb�(���'`�u���I�-�Y���Ć����qn?��d�G$��|������W�ܤ�����8����2�46�s778����I}J�a�����}&�p[^���f$wg�h7�n~p$�hd��?{Yڕ��%Ki!	PR] d �b055 �O��"}�}�q<�bX�%��mڜ�bX�'��{!|5�sK����'�,K>UH��}19ı,O���'�,KĽ�v�ND�,����׉�Kı/����.�IwrܺK�u9ı,N����yı,>Q9��mڞD�,K��Ȗ%�`��{u9ı,O�s�~���<T�p�LM���v�M���ݰ�2����Ύ�#,�#������nv���w�%�b_~�n��Kı;��oȖ%�`��{t?�A�DȖ%���}���%�bX��M�}�l�mr�.�ڜ�bX�'{�vq<�� �"dK���br%�bX�}��O"X�%�{��ڜ��ʈn&ı;�'��f����ۅ����%�bX�������bX�'{��q<�c�ș���v�"X�%���s���%�bX��N���e��,��ݘ��bY�"}��~8�D�,K���v�"X�%�����O"X� ��,�?�R╔��e'�a��e��6�sni��%�bX���ݩȖ%�bw��gȖ%�bv{���bX�'{��q<�bX�'��d�w772�\��)!��&qe���<�Fy��չbv�&��ww����,���յD{�{ŉbX������O"X�%���xbr%�bX��{����&D�,K��mڜ�bX�'�N�!|5�sK��3gȖ%�bv{����ș�����yı,K��mڜ�bX�'{�vq<��
��n&ı/����t�K���ܗt��Kı?����8�D�,K��۵9��Dȟ}�>�O"X�%����19ı,N��e.d�&�ff�O"X�|�ș��mڜ�bX�'�}ϧȖ%�bv{���bX�'{��q<�bX�'�M�w&�v��݅�۵9ı,N����yı,>c����D�,K��É�Kı/{ݻS�,KĜ��~~~�?@ h$ְ  m.Y��4M�:%�4�͂GMYٴhl�kK�ٳ���d��gZ�1j�r���z���ZU��yz6㞲wJ���x��iyAq����1�<f+��v(���w���r;�P��=@�P�&�.eH�v֪�\ؙ�KQ�2� ڠ����nz��MՆ���l�[;t�ƺnu�a�#���v�/)�(o����Ϧ��B�V,�p���7e�tZ�TR���؂�N�-��vw�=٤O�^��wVl�?D�,K�p��Kı;��É�Kı/{ݻC��L�bX�N�R�)YJ�VR��Z��h�������,K��{�'��#�2%�~��S�,K�����yı,N�{��?�ʙ���ܟd�ܙs6M6nm�8�D�,K���v�"X�%�����O"X�ș�߸br%�bX�}��O"X�%��p�e�m�wn�7v�ND�,�`dO��ϧȖ%�b};�ND�,K��|8�D�,�_�.�����S�,K������[.�6�fl�yı,N�{��,K��#��}��~�bX�%���ND�,K��;8�D��oq�����%e��^,���۱�{tp�1m�ݧ����/���T�iv�Z�f �K�K�l˹.��Kı>��8�D�,K��۵9ı,N�����"X�'ӿp��Kı>�gm.}!&�70�34�yı,K��n��?�~^�hϒ�`��Y	 �Q�B$�"��0� ��F B*��F0�"� A`����x�	�Fd"F DBE�c�Y$���:�2��5�<��,M����O"X�%�����'"X�%����O"|�TȖ'�7!~�m�k�v3n��Kı>��}8�D�,K�����K�?���؟����O"X�%�����ND�,K�~����v���p��8�D�,K�����Kı;��É�Kı/{���Ȗ%��$ȟ}��N'�,K��>���mfif��i�Ȗ%�bw��Ȗ%�a�s�븞D�,K��Ӊ�Kı;=��ND�,K����n��-�Ը:��]JN�Ք\k[b�+N��ץ�z	�I���������I¶�:b�����%�b_�Ϯ�r%�bX��y���%�bX���f�șı>��8�D�,K�>Æf�%ݻ�l�۸��bX�'{�vq<�bX�'g�ىȖ%�bw��Ȗ%�b^�;w�?��M�ؖ'�>����wI��3gȖ%�bO��br%�bX��{���%�D( w� Q}�h.E8���s�ؐ���!��
���zg<�ںa�E@fRbt��'�p 'f���������¯����$���� �d�ڳ�a�Q,���"Jl؊D�	 ) �H�b�)2�����`@ ��Y��8��\�8XA@�A �Ѕ�a�Y#��q�8�$G��K�j�<8��辪� u�ht�V'��pS��:��E
������Q/M�B"_y����Kı?w�}8�oq����~?�n��FI�g�Ȗ%�,���}��yı,K����ND�,K��;8�D�,K�����Kı;ݞ�rβi��\�8�D�,K��۸��bX�~��>�O�,K��w~���bX�'{��q<�bX�'�od��̗ܻn�u�":	�JC6�]7�ˌ��;Hv���k��� @s��TO������D����yı,N�{��,K��{����2%�b_�Ϯ�r%�bX��}>f����˄����%�bX����'"X�%����O"X�%�{���ND�,K��;8�D�,K���^�����M����,K��{�'�,KĽ�v�'"X�aK
RN�R�)YJ�VR�����%�b{Ӽ�K�乙�a�sn���%�bX���ݩȖ%�bw��gȖ%�bv{���bX���2#��/{�'�,K���ߏ�,��|ڢ=�oq��������O"X�%���xbr%�bX��{���%�bX���ݩȖ%�c��w����B�]�cV�Q����$g/����ێ�-�*�6��Y�Y-�Ω:��)�ne��<O�,K��w���bX�'{��q<�bX�%�{�jr%�bX��y���%�bX���fe��R]�f]�wLND�,K��|8�D�,K��۵9ı,N����yı,N�{��,K��'�zgr4ܹ�is4�yı,K��n��Kı;���Kı;=�ND�,K��|8�D�,K��k;�۶�%݅�۵9ĳ䁑>��>�O"X�%����19ı,N����yı,K��n��Kı?g�;:�7i�.sgȖ%�bv{���bX�$~��O�,KĿ}�ݩȖ%�bw��gȖ%�bw�{��?�|H6�  N<�[�� Tlp����Įn�X��P{s=�p��1�ѕ#��Z�4���wlҠ=$�Vs$�W���EH��t[k��+I�ƕY�]���
�����egeܤ�u��]]��ph��U�p�&�F�G@k�`��Ny��r����;�<2NwU �\��i�qm�79�'�	�	˒�)��{ޞ��/Ȱ�&��g��bz�cc6C1�tq�/b��:�zV;bq9��K$��3����,K��É�Kı/{ݻS�,K��{��'�,K����19ı,Ozw��p�.\�0ɹ�t�yı,K��n��Kı;���Kı;=�ND�,K��|8�D�*dK�>�I��m.�wn��Kı>��}8�D�,K�����K����؟����O"X�%�����ND�,K�ǽ���wI�2�͜O"X�%����br%�bX��{���%�bX���ݩȖ%��L���y��yı,K�~ٙni��nٗr\ىȖ%�bw��Ȗ%�a�Ͼ�n��%�bX�}�>�O"X�%����br%�bX���N���D�H�]�[n���ڳ�8�mì/lq�]�@WW���:�F��n����bX�%�{�jr%�bX��y���%�bX���f�șı>��8�D�,K�٬�e�m�K���jr%�bX��y��� =X`0"!��P&�ʤr'�,O�����Kı?}��O"X�%�{��ڜ�bX�'��'gY�6�ۄ��'�,K���{19ı,N����y��V"_��n��Kı>���yı,N�'izn��3L�����,K "�C"}��jr	 ��۴I�=��u9�:
��'Ӽ�br%�bX����d�i�.�0ɹ�t�yı,K��n��Kı;���'�,K���{19ı,N����yı,O��}ņK�"ˎnݯ*�A��5=cxÁ�r�l;��	���E��{���o�/Vƛc�7v�O�,K�������Kı;=��ND�,K��|8 ��L�bX��۵9ı,Oޝ�K<5�wM�-����%�bX���f'"X�%����O"X�%�{��ڜ�bX�'{����'�9S"X���nf\�).ݳ.乳�,K�����yı,K��n��K�"1��@�Ʀ���&�߾�Ӊ�Kı=�ߦ'"X�%�韧s�s�̹�is4�yı,K��n��Kı;���Kı;=��ND�,�������%�bX��͓�-�i���76�ND�,K��;8�D�,K��Ӽ�byı,O���'�,KĽ�v�ND�,K�����v���Z��V�t�T�M��s���,�v��k��s�tW�rt�f빳��Kı;=��ND�,K��|8�D�,K��۴?�	�L�e+)I:K��e+)YJ	j�ݢ��2n���ND�,K��|8�C��DȖ%���ND�,K��Ӊ�Kı;=��ND�,Kޝ��in]�a�sn���%�bX���ݩȖ%�bw��gȖ%�bv{����bX�'{��q<�bX�'���I�nIeݲ��wn��Kı;���Kı;=��ND�,K��|8�D�,}��y��v�"X�%��ӽ%����r�3gȖ%�bv{����bX�G�����ı,K��mڜ�bX�'{�vq<�bX�_Ϳ*8X8s6��Alb+!�e쑎��qTS
/+��h�������U�{.乳Ȗ%�b}��xq<�bX�%�{�jr%�bX��y���Qg�ı>�ߦ'"X�%�ܞ����vR�]�K��Ȗ%�b^��v�!��؛�������yı,O���LND�,K��|8�D�O��ؖ{�?�F�XV�V�b=�oq���?����8�D�,K�����Kı;��É�Kı/{ݻS�,K������]vCwl��l�yĳ䁑>����,K�����yı,K��n��K���������yı,O�d���7Yd˦M��ىȖ%�bw��Ȗ%�a��1Ͼ�n��%�bX�}�>�O"X�%����br%�bX���t��⓽ݽޝۧ������:??~  H��  m��[��QM�;���t4�ɢ5ͱ�٣m�� g.��qm(�p�j2�^T�cr��8����psX�m�O4�M7/Mܩ���-�I�^�W/�l\-�1��1��v�]�'%;�*�WX[��J`�bg{<�����~���;���ϖ��u�D���W�l���9�v��V����s���b(��ny�-ٗvۓ.���m�� �I�渘����Ƅ�i���b#n�V��9��Y��s7d�&�����ı,K���S�,K��{��'�,K����19ı,N����yı,O};��p�%��%wf�ݩȖ%�bw��g�|1ș��w���bX�'�}��Ȗ%�b^��v�"|�TȖ'�N�I|5�sK�2�͜O"X�%����19ı,N����yı,Os��ڜ�bX�'{�vq<�bY�7���~q�;'ϻ��7��+"}��~8�D�,K��ۻS�,K��{��'�,K� �E��}����Kı>��O��ɲ�2�]�8�D�,K��wv�"X�%�����O"X�%���xbr%�bX��{���%�bX=�{m�ܶe�-�r�]Y���c9�
�o0.���6��6���]Z���������*�s��Z�w�{��2X�}�>�O"X�%���xbr%�bX��{���?��bX�'�����9ı,N�O��u��.sgȖ%�bv{���SLCbX�&w���yı,Os��ڜ�bX�'{�vq<���L�b}�R�n��.�77sLND�,K��É�Kı=��wjr%��(C"dO���N'�,K��w���bX�'�{��0�33t�&��Ӊ�K��@ dN��n�ND�,K��Ӊ�Kı;=�ND�,��P�����Ӊ�Kı>���L�m$�v��m�ݩȖ%�bw��gȖ%�a���~���%�bX�}��O"X�%��w��S�,KĿ�vC���ws6�gY��q�űv�82Q�0o(u�z㧵�=zn�� Js��5�3K�2�͞'�%�b};�ND�,K��|8�D�,K��wv�"X�%�����O"X�<oq������"2N+�w��oq���{�'��9"X�Ͼ�ڜ�bX�'�}ϧȖ%�bv{�����2%�ܞ�ٟd�)s.��Ӊ�Kı;�}��9ı,N����y���"�hb	i`���b)ȟO>�Ȗ%�by��8�D�,K����fff�L�vl��ڜ�bY��"}��}8�D�,K�߸br%�bX��{���%�bX��{��9ı,O���-��f˅����%�bX����'"X�%�ʑ���q?D�,K��ۻS�,K��{��'�,K��w�N*�+%u�ܵ�\�7`u�l���q��p��j�Ή��ۉ���g"���[�Wh���O"X�%���}���%�bX���wjr%�bX��y���%�bX��{§"X�%��^���v̻�7v�O"X�%���wv�!����]��,O���N'�,K�����S�,K��{�'�?�r�D�>��re�i&]ۘ�m�ݩȖ%�b}���q<�bX�'���Ȗ? "�؛����É�Kı?���wjr%�bX�~=�/��fiv�Y����Kϕ`dO~�xT�Kı>��8�D�,K����ND�,pJ��T��=E�Ļ�vq<�bX�<~?8��=�p�J�����oq���|8�D�,K�������ڟ�X�%��������%�bX��{§7���{��?���⤩�y�����^"9����s��y��F����Z�LՁi�&�\˸iw4�yı,N�{��9ı,N����yı,Oݽ�C�I�L�bX�}��O"X�%������`9�k-G���7���{����>c�2%����9ı,O���'�,K��w��S�?�C*dK���_�.�!se��l�yı,O~�p�Ȗ%�bw��Ȗ?��2&D�>�wjr%�bX�}�>�O"X�%���aܛ��˦M���ND�,K�{�'�,K��w��S�,K�����K���߯�9ı,N������w2n��8�D�,K����'"X�%�����O"X�%����*r%�bX��{���%�bX�_ <A�� X����T�� �:	D�$!�8$'���]�	������'��w��,`p'>�q)�,XX�	a8v�DT��!(A"R��RBD#	�B-"�@�@��}���             �   ��              9ųY]iN�s�K.aXr�E�+H#�
���r�Y���6��8���֝�kC�M���.���qH+<�6�m������˵ӎ��s��*�7�&VS���[��:<�ax�`VV��u��1�kYŞ0.!��Kc'A#���
�T��\�46�������ԫ��<��D��Ge���V�@66U�Zꮀ�՜���b%i�y66�5�m�XG* �`�6������(iS�f����۰v0M�ոҏ#��h�)� �z�R���
v� ��\��@��=���x6�i��:"N�l� �k�
�8A�	ꀖ��̨�W@'i�;E�� l������7�ǵ�fr�[�qz��:�u���.���M&KF�*���\�-m�^{mvMu<��cv�ݵ mp˫�K�2��hi_b�r��Nۜ(>#�v6�z:�j��7a6�N��:�]�d�.+4VqW[h�	�m�;�U:���e9�;�=N�^�f��Q	 Ϋ;zf��͎��+�j��kF�VL�V���MYPvݹ�q#m�K͵�$�ke����J��B�	��ɘ�4��uJJ���,�pui�s����N���5ol]��������Ѫ^L��c��le�‧����q<<*����+ė�`�) i�\�!^Lm�8�\lZ�n8��Am#g�͵QBJ��X�%ۻV�����v���e���,����4o)��L ��.�QJtY{\X��ݵq��'g�V�����R4������g��.�R�]6��2�8�q[���7�d@�{QfѨ(s�!S�L�c�͈h%�:t�n�6Y`lv��]��OEs��l
��m����{iNV�F���ѫgX^.v@��h���̲\$�ʡ�D�����@�4#�z�>�#�� ��CAJE=;ǀ��G�A�v{�� �J� 
����Y�uۇJ��(^���x�qq����$�����\p�S�9�[�E��=��n'�Guv�X��S�|Ak�VI���-�M�0$�6�����y�uu���D\��=��Yyu����ƠanC�.��^���ݎ�R��e�.����r��7���*��C%u�m)���nf]3vm77r��W��̟�S7-��um�a�su��Sf�Sݎz�<D���n���������u����(_fm����ı,O�}ϧȖ%�b~��
��bX�'{��p?�_�/�6%�bg�n�r%�bX������\��]�e�6�<�bX�'���Ȗ%�bw��Ȗ%�bw;����Kı;��oȟ�����,K���e�vnI���ܷt�Ȗ%�bxq<�bX�'����'"X�%���{x�D�,K���Ȗ%�b{���tۓm�&n\�8�D�,�`dN��n�ND�,K��Ȗ%�bw��9İ>������%�b]��~q�ai^���Q��{��7���w��O"X�%��oxT�Kı;��É�Kı=��wjr%�c�{�����;�-J��k�R^�1L�Z�k!�!�Sv�<�7h3k����v�K�����Kı;��
��bX�'{��q<�bX�'�����E�DȖ%����׉�Kı>���f딙�2nf�9ı,N����y"5| �8�y"X�Ͼ�ڜ�bX�'�w�Ȗ%�bvw{19ı,Oz���c�e�0ɻ�t�yı,O����ND�,K����<�c�C"dO�����Kı>��8�oq������w��WGd(�,U�D�,K����<�bX�'gw��,K��{�'�,K�=߾�ڜ�bX�'�N���L�.�2˛x�D�,K��ىȖ%�a������Kı=Ͼ�ڜ�bX�'{���yı,K��K���͙�������e����4���O#u�a�	�D��#�f.1u��N)J���{��7������O"X�%��;�ݩȖ%�bw����"-�&ı,O�����,K��'o�۹r����K��Ȗ%�b~��wq9��DȖ'�o�^'�,K��}�LND�,K��|8�D�r�D�;��������e͛3ww�,K�������%�bX����ND���Ǫq���ș��É�Kı;����r%�bX����zYu�K�.YwoȖ%�2'��}19ı,N���O"X�%��;����K�� ��s�Ȗ%�b}��&�i3rd�ۛ19ı,O{��q<�bX�ʱ�~Ϸq<�bX�'~߾�O"X�%�����4��������uҢB8�$��Y&��X���x:�n8�Y��[u=������[�����w2n��8�D�,K�w;��Ȗ%�b{��oȖ%�bvw{0>E�DȖ%�߾�É�Kı���_��;!D�a��}����d����'�����ؖ'����Ȗ%�b}����Ȗ%�b~��wq9ı,O==�|ɮe�3neͼO"X�%������Kı;�{���%����؛���۸��bX�'�����yı,K�zۦ��%ܗw2����K�䁑>��O"X�%��}�n�r%�bX��}��yİ:r?'Dŀ�B ?�������G�wbvyىȖ%�bd����f�fnff�O"X�%��;����Kı?w}��yı,N��f'"X�%����É�Kı=��Nn��fK�̵�!�A]:4u�v�q[t�ҙq��{���'hI�����1�r\��{��,K����׉�Kı;;����bX�'���'�,K������r%�bX�����뤗6ܒ��'�,K����br$r&D�;�~��yı,Os��w�,K����oȖ%�bv;N���&i�w6��ND�,K���'�,K������r%��C"dN����<�bX�'���br%�bX���/nXm�w2n��8�D�,K�w;��Ȗ%�b{�����Kı;;����bXȝ��~8�D�,Kޟg%̻I����3nn�'"X�%��}�gȖ%�a�*����byı,N�߼8�D�,K�w;��Ȗ%�bAz=~_�  ,�  ��&ٹSIRY�ҧM{-�i*�.��n������S�јD��6�SX;is�N�U��w�Q6����gs��\W�ZU}D�+ʶs�qL�rQ��p��Wk=�gsC�r*�&��=������v6rv!#0�fے�xs�tݫY��`��I�yƽ5u\�z`qm�񵎜�@�'v�1�<�hjo�q��{�~�Ad:2�s���轖�*ۦ�h׷a��܋U#&�&����ڛ���ʷ1s������%�b}>����bX�'w�O"X�%��;����_��&ı,O����yı,K���e�Mܒ�K��w7�,K����É�Kı?gs����bX�'}���O"X�%�����>EL��,O��}���7l�&��˚q<�bX�'��}��Ȗ%�bw�����K,[����I�����I���L.fJd���D�$�(�}�w���%�bX�}~�ND�,K���'�,K�������Kı=�ǲ��뤙�\���'�,K��oyS�,K�����~8��X�%��}����Kı;��V��؏؏؏�ܮ�BB6���҉�6��d���ˮ�!�ۡu�j�w.�h��)3L˹7v�"X�%����Ȗ%�b~��wjr%�bX��}��}?DȖ%����T�Kı>��/�2�a��2nM�8�D�,K�w;���j?)��B�&D�;��oȖ%�bw۽�9ı,N��|8�D�U�q6%�ߏ�乗i2�۸�m����Kı?������%�bX���ʜ�bX�'}�|8�D�,K�w;��Ȗ%�by���<ݺffi�t�����K��AG���?���ҧ"X�%������Ȗ%�b~��wq9ı,N����yı,K޸�ɒ0��#q�/٧�G�G�G���q<�bX�'��ww�,K����'�,K��n�T�Kı=���aȢRc@�9	��1�m�'&���v1��{96;l�s����Eqt�]�'jl˚q<�bX�'��w"r%�bX��{���%�bX��w��"X�%����Ȗ%�b{�v�ܙ��p�sf��Ȝ�bX�'��{x�C��L�bw�~�9ı,O~��'�,K�����ND�,K���^��vB�$����Kı=��eND�,K�{�'�,z�yE�(~H�"aA�p4�%���ۑ9ı,O߷�Ȗ%�b{�Ӧn�I�f]ɹ��"X�%����Ȗ%�b~��r'"X�%����'�,K� ����T�Kı>����M0�4��8�D�,K�w��9ı,O}���<�bX�'���Ȗ%�bw��É�Kĳ�����SS�4�����V�,��ɞ����vE[��B�.�p�R;)E���܉Ȗ%�bw��oȖ%�e���^0&�y���xƖ���X�����	mx��׌	��`Y֭ ���ɒ0$l�f�z�������@�n�}h��F8�s4Vנ{]�@�n�~��H���P � os��~��)�G�'9��v������~�<߾��9^�@��BH�	�DE�=q�q,���ĝ[^���t5����z�*=\��!2
bJ~��D<JE�u빠w[��r�^��v���+$��cz��,`Ik��/0=z�`OZ��������ǋ$��z������Z�閳{�nږ��ͼ��?<n�~o��7˂%IR�_���Ͼfl�cnBE1!8���\��.��<�?<n��J�*�{�����ݯ��  $�P  %��Ye��bFݰ�$zFu�(I{us�z�i��6�=�ϗ�Ms�0l��p��m�m��UW(bm�Hv������8�Ɩ��[�E�jm[�WXm�`��Y���>z�Ҡf;9W�%�;N�n5�^.7��%��[d8gD�.id�r"�nE۵s8\�]�����iÌ�����H��w{w{�����}����/9���E�^{�pqv�qT���Z��WOF��Y�٨K�o,�ex���y����z���uq6((�7nf�궽����d��7'.����{��m^��Ž��B;�0>�n�$��I^0=Vנr��\IO�?)ґh��hJ�������q7/	n��;�q�c�^0=��`_u��������$ƔɊHdJ �9y�ic��v�[b����۴��sյ�.N��]��.X���y�g[�	-x���s@���y���G�w;W?�c	$_��y'��9$�w4U��.Z���܄�bĜL	�^0=mx���y�'[��Q�@�`��MI�����z��ڴ?���4�x_�O'�����o�8�$�����~�� ��.6�������*Ny�mu�ʤ�Q��V8�n:^��i٫�{uί��}qsL=�#�����;�w4��g�r���
�(�Ĕ��R-��s����\s8�n�ya�OڻFj̽�7W ��.��<������P����#	$R��b���A$$B$ �Z� ��,�����"D�)p9������'�77T-�Ye%�Y HXVK�� F B��+n/���OX`��H��cBbS�4�0� A�@�$F��f�l� F�+(�t+�f�$�	(�ZǗH���	I��) �M����"U�j�M�$H@1D���Wp����b�'�AA���N�:����(jt�@<�� ]����^I?{��䑺{v�ZՋ/KXn��>_,{��8���@�m��/[��{�n�<�I&�m��� �����_�G'.��7��Y#$�����$ciĶ�p%6��ru�^v���;���o��קu"�BԎ�Է�,����^0>�[�:ՠ�Q�B(`ډ�ԙ�^�s�J�����K�?~���?�#�5��l��s4=v��h��s@�n����Q<�8(�Z���I?~��9$����$�H��~RQ� q(��=��y$��{/Ku �Դ�Ե��J�%�{���ڴW�R�$Ci�A�23�<��9��E���l�6�j�5c����뮡�'\����mF93@�s@��j�=�ՠ{�]�����F4��L�<�������ϗ�7˥R�����4�!�I'�N-�|�}빠w[��y�hvZ�[��r8�Z���x��׌����ٳ���X��cs"���MI�u��������?~���uRuHI~^�G�Io{i�~���o�@&�  ��fۦ�nƉ4屶�d�y�/%�qsq�V�\��y�+ٕh8���޻���m��km���*�r�����i����V��u�f9E�����e�wBG!6㣇z��ePh������ìe��e�Gכ��5ƻa{]�v��&�Git���+	�1��l并�,�Iooлnc�L��rѲ�����{�����U<p����ݲ�op�����SF�B[I��� �e5F�1/k�di��<��h�j�=������g�-����@�F�ypQH�k�h��Z����`M�Cnn��A��CJE�{�]����>���/y���;���@��9ed��cj1ɚu�����׭��+���n����n����K{���[�zW��w4�����O�3N(=!t�k�Uun��y�����䎈�����sY��8���iŠ{]�@�޻�u��~���y���=���Ű�9#�1H�'����B�Ġ��B	��
� (���ȃ[��?��5��^0>�n�=z�`�70���n'3@�s@��j�=�ՠ{�]��\T��&ț��3BRIU���|�I|��|�y�\w,�D�$࢑h�j�>�π������zPƒp���]y;�c�e����^�nC�nݹ���mf�ms15�)�S��D4�Z����;���<�ڴk�h�g,�����mN9,`Ik���u�����W���J�Y҃�FI3@�@��o ���H����g��8rI���f�ݖ�I�FH����v��W�	-x��u���e�hзW,����/v�����D�r/�?<��k�h�jX���&E9'�C��g�[8�����<�\��陸s��h��:�u�9n!1�����~�s@�@��V��s@����H��dM������[�[^0$���ۧ���j'�N)��?�Z�������ڴ^�%pJd0��CJE�z���{���=�n�?��I%\RQ,[���(�E�N�y~��y$��'V'����D�Hh�w4�j�<x����p��Id�V�n��,��A�p����`^�2Il��t��������y�Lk#P�$����Z�ڴm��;��h���I�F7!'�n&׭��T`I+��n�~����F<M��2�}>4}�}}�@�|���1��&6�q��J�'[��X�Q�sݗ,�1'LJL�;��@��V��%x�y�����fff__�I$�@�I�`  ��k��ę���t����t�]���4�P��O\��v	k=x�E9��A���yM�-(�c���瘅;��ᳵrf� ����;���b��իD`�J��w�m��t(������bxź���EY�W��s���kFSu�8�1�[n�92s�=��f�3u��.umysv�r�����Ψ�`�www���V���n��+���v�Fb�mu�n��NF���4Ʉ�Q��A88�^��ՠ{l��^0$�u�6dݸn�Fږ�jZ����%x�����[��f���U���� s��h[����Z�ڴm��-�`�7��(<f᛫�U*Um��Od��~oY�?u��=�-֓ȌnBO�&�Z�ڴZ���W�	:�`{�]�v���Bq7ݲ��T�3]Q���Ɔ�<�U����	3:��El�eiK������I^0$�u���u�HJqܰ٦Lٛ�nl��}�j
�E:�o���h�ڴ+�m��;=yr���dm1�3@�v���Z}��.���[~��<����Q��A88�Z׭��T`I+��n�&̛��C�LLR-�v�����;V��v��߿~��߾�����F�"8gfv'&�l��p��t"M�ezH�X�6ö�!jb��b�9�[~��=�j�<�ՠ{�ՠu�`�7��G����[��[�N�XJ�=��I�F7!'�n-��Z��Zz��`BR�?���!�u)-�J�bBFl�ˀ�y%���˵�m�f��ͽ��o�UU+��/�m�\��Z�ڴ��1��&1����XJ�������ӭ�����Z��� ��0ss���A3�vg�]���l����v��6�����<[�ҎIcӭ�׭��[�	%x��d���D�	�qȴ+�o߳:����9p���J�v;i�Ŧfh��Y�jZ���~���`zu��������9&�)�A&)�h�w4y���O;��䜨�#E���X��*+'E��|�o$��=�ܙ�15<dc�4yڴ�h�h��h�T�Ԙ&�)�I�P��m\7m@L��m<L�ts�H\�Zm�A��I��ۋ@��V��t��{���;V��e�,�E�$q<jE�{�Q�d�N�X�n�		L��&1���!�^빠y�է߳�����@�gƁsוX�ĦF��8%�{%��%���gUq���<��J5�'��"�/�ՠ{�)��{����m��{��m�2��?=w�}�j0�"�pP����)!O�����|0���D�Nwx�7�Iׁ����&��&��6�b�Hċ44O�p<�Z��<��a�&i8L1�I�p�VI$Q��OY ��}$��������p'O@����=�ā2'���$-�C�?ozL�? �B���wt             �    2��              r'^I��ۨ��v��('b-q�	�BҤ G!�kz���T�H&-��@��EUZ)�U�]9�k<�p��L�� 0v��];Qe�X�=���d5t MUT����x.ynїV ����m�]��Մ׸l$:�̶��*��챭g�6���#3!��WmۺNٕ��
m5WUP q��Q���g-����n�`�l\���9M��-��k� j��YK��H�l�l�LZ6� ���Z�X�4/U�$� �t1A���'(3��R�AN��A��VP�7mEd�RP��nZ�U�tG\�]�R�m�
��] p�뒶e����Wt��=ll�l�I�*/g�\�i7]#�ac�̅�`l���ݴx�kvۯ[�1��Nٍk�t�������p���plݳ�Ei��q�9{f؉O�D�{R3�x��1��[9��g�� ��fhݵ<�X���S5�1�:�����,�U1{s�K�V��� T��a���j�vw:��:��fۂ@[����xj�B�U �p����5�J*vq=�Svi˓���U��e�8(�ٲ��ݪ�(��v���v'EV�鬠Vs�D���(v���+�]�J���8]����Bj�l㤺@��������n�����<�����J����mu�ݶCu��kq��=�%@
��K���k@]�����\�^yΎ6#�&�
ڃ��z�n�wnÉ�Lv5�n���V�ì�T=�تU�����Q��q1$����`����ѐ����q�O.-[Fv�X6�M&捓���gH�N�,��v���<�K\�.ʥ�u����D��׀�{5�0N� �m��$��
E}��h���:��=T��� �uT* T��	��È��=�����  �m@  �r��CR��6"vy��3�+�.:���ƙ�f�,����ɦ-���Wg�t�ujz^�[,�1�țX�ܩ�:\sd@�s�\@'F����n�Ub�\t56i���X�F�	�.ײ�{Yw��tG������u�8�[hפ|�L(����2�ۮ����X#�Hssٖ�.o{����:��H5�42�-����������\�z�Ӈ�7#���\�p��2$Oѐ��s5"�I+l�5[o}��ym���w>T_3-�{�}|��{��_b��b�'0ԒW���x�K���I+�y�Iu�pԒV��*�MǏ��<I%���$��Z��}����pԒ_[���%�u��$�O�&܏RI_e��K���������Ē\�RI{�kK<�Q��Gb�y�Iu�pԒ_~���o�群���Ԓ^Yj�~�?��{��_�j��1�[�xF�/=�d�ű��ȍ�{=RW�rtj�6x�$��I+o�f��K���J���w*��컷&�:�����yr��x^��[�y��s���D����f�NKW�$�[7I%����Ē��LV	F�y�8�RIye��K��������o�$s�MI%ϳ�/��a����E�%�����y�I�SRIye��K�9!�'��)�5$�w_3�K�ٙ�ϾSĒ^�>�y�Iu�����?��d��m5����( �"�v����M�l�vgGF��V�>\�#�L�Ē9ڦ����W�$�[�~�������y�x�V��ZO"$����ۊjI/,�y�Iu���$����x�G;TԒ^�Z��!nd���ȷĒ��xN[m��{��u��J <W���ٍ��ǩ$��Z��$�K�i� �6I0ԗ߳?g�n����$����$��Z��$�ٸjI.�f��&)�!)3�Is�=I%喯<I.�n�K����$��) ���MȈD9�˕���s#n=F������e�N:uƭq�pG�"(�RIye��K��������y�I.vǩ$��rE�?71d���-���xN|�9�o{߼<��os��I/,�y�Isg$;�� �"Ra�$����x�K���I/,�y�Iu�pԒ]]c�6�ǌ�rg�$��l|���w��ym����r��tZ�߳?K|�3�K�.�I�D�9?8�r=I%}��<I.�n�J�_3�Is�?������;�hLs&筐�m��ތ8d �����c��<]������}�7n�:�KuL��{�I_���������Ē\�RI_e��H��6��Q8�$�RI^��y�I.vǩ$����%����i}��_���X�����$����$��Z��$�ٸjI.�g�$���
ĵ��Q@��#Ԓ^Yj�Ē�f�$����x���~nϾ�RIWr�}��?'11H��$�ٸjI.�g�$��lz�K�-^x�K�~V�$�I$�H��  m��[�Xլ�&r/�pJ[p���M���\s�F$p�8��؍Ŵ��5�砢{�JK��s1Wf��k�X�i�rc[=t��a�m�Rn���na�<A��%�	X;`Ԃ�B��,s�p��%evL��d9{>�Q��5'"`�F�K�﮾�'\��^|�	ӛt��<��Y�g] �Y����r�ݵ�M�/����ٯ���]�]g7��c�lG'k��;`㍳8�`�<]<Y�۞��!���L�I��$����y�I.vǩ$����%���RIu�T�$�Y1��L�Ē\�RIye��K��������y��~����V�ۭ'�����ۑ�I/~�|��$�ٸjI.�g�$��lz�K��ZY�"�̒269�$�[7I%����ă��@�V�֗Fӟ�;;�j�9,`}%x�'�L�K�o]��ٟ�w�%�H�$�l���8:�,=p�h�ݍ�UVB�Q-��u2���"��,jb�&x{女�>�@����+��L/���j�{��$�{�����"$#*1��
�AA�g}�I?w���!��4U�H�����&)��빠{ϗ�Wc���?c��~��1�`n�a�n�������=����s@�V�	d�Dԙ�֦�K�Y^0>��`}苢\=s�9.���n��aqM��f�8`�z���ٷGU�iY�I2��1�폤���u��+��W�z���-��hZ��$�]��k�W�����@�_U�u��m��'���%��y�{ÒI���y8}�8J��p
x�����%K�U[�r�H�p~��,�Y�ڴF�0KS{��������篑`�pLQL��&�=���׌������(cU�Ѣ��v�v�ʹ�D�moF7{C�n��\=m�X�]XNB7����}���^0>��`���K�l&�բ���R]�Y^?f�Ky=ҭ���g,9�	d�Dԙ�Z��.�=-x�����[s{D�\��[��0'�]`{ּ`}ey�� ����_}��'};ܴ�ͫ�bK��ܖ�=�^0>��`���޾�@�l�A�1�24�ܟ�Q'������S8�ѐ�s]Mr�������:zJ*�ε�:~��&$ԙ��~��}�h�꿼A��ۚ�:/�I��5�����=���W�����J�����Z�orI�OJ���`}ey��@�\�1O�?71�h|����0=��x�'�LzT���n�Z,�,5-Ա���� ��0	�W�O���������{����@ h&�� �5䱺E���&ݙ�o$r�;�]zvn�u;��V�N� /p�-�̊��+X���	Λ��ᤑ�کR�����ڔ'vn�@J
.S�k���7;���;��X�VΨ�dYK�c��mG,��1���[�Qm���ro��~45���j���9ɉ8f�����k;Z5y�`5�i��v-��R�:i� |Q���ݜ�vn�՛��/]w6x$��L�i9���e�e�K�v'9�J��y�.�}$���o {�����/��/���\a6���5#nO�&ܚ�u�����y��~ozU$��ԙv�M��՛���jI�?_�J�OZ�����K�k'�1�bC�4�ژ������x�mKNՆv�n��z��>����J���?�~U��°�[��m��Na7c�\/F�l��<���6�1]*:��O��w$�m����`I+�=j`{}=��e�r��3w9$��{ÊQ �!BDR��b��}ˀ������tI+�֛.^�7D�ԷR����=j`[f��빠u�U�����Ldc�4%R�v�&��&���.����{��q9�H܄�"mɠ[f��빠{�|�ߛ�R�^��w�^�75j�bo�96H��^j��u��hZń�䓮�Ƭ8�(҄QF�9"jI���s@�+�=j`[SZ\�|/彜rn��0$�� ��0����+��
�&L1��	I���4������� 0 �|=%H��%EL\�X�c"F�V0�d�� Ў�1���9�FVT#X�IIB$R�"6�1��������n@��(lC�*x��#!f<H��P�G����P�����IU'��񏇘 n�<A� �u=��'�D�0Q���� ��E�C�|Ey�|��$���xrI�ܞ��L�Է���.� ��0=ex��W���h�9+�)�D�'?'$�=�w4%x�%�0�S�֋D���)r���{\Y6pv�����"��pHT:V;l�8�V%�iҒ�����������x�ob�_��r�$XKE��Z����%��T�/�L	ey�^빠we�s"��	�Dۓ@/�LY^0,�� ��0=2��bջ��.�ԓ�W�	%x�'�w�ja֢�'��TX���������ņn���\��ˀ�V�&� ~�o�����	��xV�H3lc�Pv�r��;f;[����,��S.'�լ�)�PJD�0Ƣ %&h{l�����+���`zq.�7��{�X�s7w�?�{ҕ*����\nr�~oz%J��vӹ�/kv�v�7w��s��y��U��&����~���h�wKKu,`Y+�=j`����s@�P+�"�c#��֦}j`z��d�nfh5
�b� �>{����������쀒@  6�̻\�O-��d.�4im5�]h�f���ci�������-�h۠�v�S�ew�P\�r9��m�]����.��s��o�wʛ�!^#f���kt�$LWG=�gsgtdz�Yo[�y8�;D���6�t)mj-��� p�;CuAh��Yd���eu�Y�;%֬�<�:�G�:3�����5;T]O�������Y+��f�n����]�ۨ	�:7`��!8�gN$]�fᱧ2)���M�= �ﾚ����W�z���J]˴�ŉp������`I+�=j`[S[�ĵ��O��L�;��h{l��@����/��+s5"M8�>I]�I�=&���.�ϗ���F'�G�7$�/�ՠ{z�h��h{l�<�Ԕ��2%��ܝ���S]�8����FM�ue��ymv<�զE���K�R-��s@��s@=���UT�/�	��ZlW4V��ݻ�\��.�]*I,H���}�hz�h�*q�@�Ldg%�YS ��0%���^0$�.4�E#s$�"�ɠ�f�׮�d����e��]�����rI�,�J�K*`֦��6���Y�!ծy��8k��vDθ��m��;-�vxd�1�Sttv���9�4䱁d����_Z���`_G�N��X�QA4�h{l߳?~�v�o��.�ϗEWg��3Q�����w3wxzM�??>\4�L�R�U%�UIZE�ˀ�����x�i�F�^n��J�����F�. ��h�٠r�����'0R%&0,�� �T�/�L	ex�����J0�V����Ϡ2l78��N6��%�٦q�j�&���ڇ��n���t����L����W�%x��*���##��294�l߳/���79p�������ٷyy{{i�����0,�� �T�/���hj�2���a���7WUq����M���ऒ��$�I!WUU	hB!@��{��'}��ov�i�v齼��OZ�����+���a�����T�Y݁����V�K�]m�u̽cΆs����C��tb�u�:��WiP�仒L�������^0	�S�g*�S��I�9&��빠^��'�L�����9v �XjW{��~���m���Wd���9&�n:�+�"Ɍ�rf�u�h���;\%V۟ˀmM"�՛��Vm���m��%U'$�_�6�. �oxʕS���T��� $�P  Xٳ i=U�9E<��3 ,V��9.��&5��n;���ٗ��kB�/Pm���n�jj�۪�1ـ���{.�ݓI�����,�;3��h깺�/l�\�!Q<�6�����tr�{8�ؖxv�S��=�n�Ɉ���˪��z9�Ν�gk��M�(�;o���v��G"�V�:땝�9���F���ݽ��߮�~��{V���yt�-f�/`���;��\BgS�\:=�}����շL��J[���{�|����RT����g����m��7Qy{�����t���M���=��s@�G�V&��Q�{yc ��0>�n�'�x��W��}\��
4�G#�M��Z{k���`��ٓo��%�r\����	%x�=eL��������qP��K7@of����ч\:���g��8�mYۉ�k��6ݹ뮡��g��a�	�`I+��*`}z]`OUF\|�VH�&21ɚ��6����3 ����)�w�w7��s�}���8B�I�{����Q�=+� �����L�iƣ�&ɠ{��p��. ����RI]�9��Gص5?E1�LN���{z� ���{e4�~��_��$h�(��ll1T�؛C�U�q�t�Ӊ��F�6H�����E��1ƣ�i����M ��0'��ϴ=*����ù���ܒI&�� =�P`_J�_Z��9W�f@fE?ɠ^�M�ׇ'@S?	Q q�7��@/�f�VZQǄ��)�_z�`֦}*`Y�Mмl6֬7�\ �7�U=�_����/�w4;�Q �d�'�H�����v����.�{Ѱ=Rt9R99.u
�]��˘�#���B�h��h�S@�����@����q'd�D��dT`_J�_Z�^�_���,��ص8̊c�&�4��� ��4+��)�w<�T��5D�j����������JR�j������r�$Y&j34.��n��fn�>�.�,��	�^0�SIC��+��-�8�q�,E�Ͷ���;cC�a��Z�ՉâTW�ڴ��&�W�������>\ �7�$���'��,��� N`���}빠�c���^0%Λ�x1h-Ŝ.9,`֦��0,��zW�{,.71����B�h+����0'�x�/�LL�1��K��$���Z��W�	�^0�S��	ӈ���"i,@��kEHI $Y��� `� )��=���Wy��/��Q�$�IK�>��s��4<<}�="}A�a��B�&h8��!���qA�������Z�I�o��?W�~Ma�����3���!���_����0�!iSw��o�#~�b�4���;Ŝ����D����Z�g� �(R0������~�M�B8�"���(�` A��=e�X,�b��B	1�	b
�bl	��4�H��	�������<1c������fI*��*�NcEXE D���B���\P2��<S�{@tR	� �;�Ͽ��             $                   �V���+�WRUF�-����%٢���A�:.���)��l �-�@����Wfu��.�'n�]#�BX������%��q�����&�Vv;E�"�۬�C�6�iN�.���P�x%.�:V�7z�r����o�&>D��˭�^5;,h��U!��Slم$p4��*�u���h��@@��f�Jz������M�M�-������I�8�#n���A"�j��A�5��d���3Ns��Ѫ]���m�Uh� �� ����͆����X���=��ȿjU�n��Ԃ���Ľ;T��,�mJ���O9M���8�둸�;�͝9�ut��u�u�N��<S�!����.�ʡ9�;7[�
�����%=w�u�XN����7�l�v�퓳snnwn�	�=bn4�m�)İ�n�].gv�m���p;���W>H4���:S&ۋKXفyK�1@�έO�ˈ�}�Ձv���PK˸����`�m��F�&zy6	��W{N^�]�g��5��U������� �җ sUUv�E����F�kei%jyrђ�.�+q����dqd���u m��[����iUNۭv$�9�t�[nj��y�E[5i�k��xrY>лDu���bP�d^�ѧ���t�MU⨸�W����h[��Pg]F�.É��V��9`YX�x��v��]�[���yz�l3�]���u5�5g��u2iKuc�x�<k����!��$�O��v=��n�Ɵ����l�ѝ�軀u@�UT,�&���M�d҉nM5�p0��Bs���64뇬"2��2z� �&���.�媔�f�n;;KR��qӲ5�$�d�K��l�ё�r���E��7i��m�"�m���w3$�0T���}Q�~D x��"|
$Q��}Dz)]A��`j)������M�  ܭ�]�᭺�����5���pm��~w�ٙѻ:���H�^c��[\���r�uE;m�N�$��Ut�
9�R�˨u^���yqғ�.z�,ۅ��K�j��).;4�p3(�a�{v:�=��]�Uk9H'��`U
�(�<��z�v�m	�t�$;7I�B"�%�7�=(������#t<�Yzw\�r�o﻽Ǹ���Wi�#���[6��M�#�8��6溋K�~��;����V�Ʉ��Ȧ1ɂjL����� �ژm��J�'e�ԃ9v��ܱ�_Z�m��J�=+��?���qߜ�8��y#��&�{��hJ�=+�}j`I���.1��W�o$��W�	�^0�S���ZS� �冥�czW���������W�Z��BX�R6T�u�ϧ.Y:\��Vw4�Q4f���%�9�n���$�Dd�F93@/������^0'�x��ʋ��9%���6˻��w�{��O��S�X(���R�]t��쏧.F�p����T���}���ٻ������G<`_J�_Z����=p��y#��԰�Ա�}+�}j`Ү�����#�3%^�,ܽ����\}j`Ҧ��`_J�'P�Y
�A07�[2��coM%��lc�<�����L=�X+�Nb�1���ҵ���y� ��ˀ��D�T��	�7�osniu��fn��|�R��y�\=&���)UU�-HC-j�Ay����\��ox�IrR+�YKI���zr�Xz�k��LY���e��w���^0/���<참��NB~q
I�޳@�׌�^0-Lz���԰��b�z��p)2��z��ݎI�	�M���X2m�Y�fuIԌ�Rl}$�����Ҽ`Z����=p��yq�VwjXw.X���� ���/�L���
��0��"m���T�/�L�XҼ`zgM�M塘�n��fn�JUT���{���xrC�� �(b���;�o$����S ő�x��@���@�z�h���<���=����D�lo�lP���d��.8����mtb9�ҭ8o6Ąv���F��	�^0�S�������3�.<������\ �y�ET�]��9|�9|�y�h�aq9�8���@RM�����*�~s� F����}���D�Z��Z���u�=+�d�@�@�qjq���L�Z����ץ��[���a�_� �J� q��8]�d6�ױi䎗��V\�n�Is0�D�"�Vw9,F�s�6��,��yLe�z-�͑  ���_i�-�uӹr��×e756�a6��ν/V�2�����,m�̪��$�/jĝ�t�8|T���D���:ڝ�O8ឳն��gl8��u���ѐu�z����k����b�'.M7��{�ݻ�����j�����ę��D7+����%;�����3��!�2h췱nd��[����&ץ��[�	�^0>��X��bxdnFܚ��[���>���@�~���f��-eK�J2X����Z��;��`OJ�Y*`}z]`]�J,A����o-`OJ�Y��<�$�%W=�_ ��ݑb�sQ�8\rX�,�0>�.�/��`w�w4VԠԘ7&cRb��b���m۠��׎@آ��N�H� ѫjp�ܷ�p�RL�K��XҼ`����C�8�$�(���/���T�H���. ~�����y.k�\b䄵,8Ե�=+�d��J����/���/�=�C�E�r�ow,`J�^�X�n�'�x��f6���܍�4+��}n�x���_m��ڒ�4�}#�mU�1�(ݞbH����t�g\����xx�!�DD�
c����{�4~����{R���1��%�n ��Xj[�`OJ�_Z�^�X�S@�䋏�XC&21ɚw��'��{y2�B, HUkh�33{�4m��=참��NAg5$������*0'�x���fj���hs��8�$���Š^�F�������u�[B��r֙G7\$��/-:Y���v|e\�rѮ��ْx��3��WW��:]r}$���>\ �7���;�RK��7����%q�0��3@/���1#ߝ�h[>4���݌�LnS7m&ץ��Q�=+�}j`IǮڻ՛vZ�Ջ/6�%*T��}��\ �7���DШ��T�u$gl�Z���ՠ��Q{��p����=eL�K�	����wQږ������g��f��������b)�իŞ�c�D�"c����&h��`}z]`OUF���Qsyg.$vp��I���u�=UҼ`޳~���>�l#�!�"lN-������� ��0>�.�=2��|/��$���CzW��T�����R��Uoӡ��.J��f�ޣo35p���K��/���=�ϗ�6b������n����� 4�� It�����nJ���u��iئy��ڻ62��(�q���eed&୶Ld3���W�ZV�fPO��V8N`ˠx����i�c.ᦋL=�g|���x��;��m�����	7+�ַc��2��l�������=�����녺ݓ�ڞ9��\`�n����܋[��N-p�94v�k�q���.n��ȧ�D���-.��s.�J$��kb�
��^��$�۝�y�����gk���\�2dI�diL �rI<ϝ�h�T`OJ�zʘgCnj��������'��zW��T�����<{n�`o,5-�0'�x�=e���Z{e4��H��D&1q�c ��0>�.�'��zW�{,.'1�G2<d"rhW�h�T`OJ�zʘ6HRK�r5E�=�Pb����s]�s�<�Be'�D�'�����&&��8�$#cqz|� ���{Ӑw��=�-�z/�ܱ	,.\��'���z�b�,���M����������ߒ�8Ҙ-��~�����z�0'�x���vY�diL �rI4+���8~���]�9�kq^�vZ�Y���X�Q�=+��*`}zS������8�y]dV�;�PnS�N
,qs��l�ͨ�MۉuӴ�m��P�.�u�l+Ky	�^0YS��������A�l8�+l5a�f����0>�.�'��zW�L����I2Ld"rhW�h��ǟ���W�,*�b�R�UH$X�BE= %`�FT�5%��s2�H0�!�9���+�=��jE
���4�����⟘����� j<'�Z�E?a����2�$��^|�P���~Ay��1?�-?>�`�/� �A?	ס�8������{�%��DV�((J1�h]�9������1Mh��B���.�y_��mx�(B/�YB�`�k#�_�6SE����ADE�@ �Q=�P���O�t@�$Q<��
E��_Z��8��R^�T����� ~ox�M��[���ln-�^�~4��� ���URU��|��Y�mnf���Fe�	�^0YS���z�0�hqRVk8+�Xv������b�KiI'6Ǝӣ:ul�-�H�h\������<��笊��W������Lo#J�$�hW�h�Q�=+��*`I����ۇj÷��'��zW��T������	�� ��Xj[�`OJ�?w��$�w=���O��H�jD>	
 `��/7�����NھbȀ��F93@:����Z^��;޻���]>D�ɒF��Ԇ㎭t��h2�)�,u�捁ꓣ��8s9�+uv�"�nI��!��=�ߖ�ץ4~��R���7��R�[�����na���y�Y�RIR����9���Z���5��nd�L�4���,����u�=U���3�o��F�fj���]�9��_��Q�=+���6�4]��]ؒI&ץ��T`OJ�zʘ��?��w����  
P  .�Ifפ��..�Kα�Y4�7\���s�aLь��������?<�B�m����tQ�S���f�����S���v�n�������[��QK�;jtv���9�WNԬ�L��Fͷh�n�Gn�H�6�r�-��+�h�뚸�x��<��hMɎ��9�zS^��FD:Nc�f�n�;,Eu鏳����F�������׻��w�e3E�n�ŌV��Vjn�o@x���m��Ӎ�v�"���Ж��a�g��`OJ�zʘ^�Xa6�r��B�0'�x�%�0>y�|����*���q`���mM\.9,`���^�X�F���aP�crL�����ZX����� �T���C5�]�#�Xnn��	b��W�YS��>�~���Y+�*G-l�7Fl-��*�F��s]E��?W=��n���9��7u�o),8\���/�YS���X���w�q0Q�s4�Y�?/��a �,⧠�.�z��*0'�x��:e团�Է;�rI&ץ��T`OJ�zʘ�����I���ץ4���,����u�6nB �冡rҼ`ʘ^�X�Q��w�������jͮ[�@R�F�R�<���j���&�Y�t��鲕r�fۭ&��_ܸԳ�	��L�X�F���vXTӈrI	��NM���X����� �T���C5�Gv雺�W{��{��p��.%%]
�<U"{�#�)�w�}��}�>�䇽��5��n~rLN���{z�������yb� �LD�o35p��J{\���À��h΅�1G1A�r&$�i$s1����n���k���2L=�[ħ7M��)��Z�I�}��X����� �Y�wq0��Y�LM8��)�_ex�%�0/�]`M����3�a�\������.�%��q���Y���G3@:������O{��rJ�����H20`(��;�w�$��XVӈM�����Z^��/�w4�Y�}����(5&	�DӮ��l���v�T���`�i�)Oj�@�V�9�&HF��,JE��>4�. ���_����jJ��k36�ua��0/�x�%�0,�u�,Tr�*Uvڹ�����5yy����ΗX�F����/-�ݻ��ŋowwx%%UT�{\�ǰ�/�x�%�0$ȳo�Ӗ�����	b��W�YS������{���}��ޞ���w�  ��mp  -�o!n�3���am���S�]s���k4'SsU�
�^�0�y�2!�k��/}r���%���2쭻U.�DzQye��9zֆ���"ԠO�A�6�f�X)�n(�5�&6x��y��-d�r�+�<�	��V�Ӑd�-�',&�;g��f0�0:��km�i�p�5���)+�kGm�n��C�#�>s��ͳvY��[���=�.����.s6�5��]��'*RZU���@���#��}��s@:����Z^��-�rI\Y����0	eL�X�F���`�Bn@x�4��<���:�F�����[��ąڎIa�jZ��*0'�x�%�0>�.��[�k'����4���u�����~�pUUI�&��{���f�iV8m�da���ݭۜ1i�j�헳n'����d�,�T�F�B�~������0>�.�%��	�^0=8�ui���ۓ����'��{y� z:�� ���$��IU/�I~�k8������9vr�DC`�6�Z{e4�������u�6hbB��Xj!�=+�,����u�,T�:�9$�,�d����z����X�����m�u�p�5�]�����l�������6(�:��:IQ���'��1�$���NM���X����� �T���C^����tԵ�,T`OJ�K*`}zU�{�o嬟���I��@�z�h������Aa h*�ο*�:�M �\�p�����Dۘ�%�0>�.�%��	�^0=8�5a��KQص$� ��0%���]� ��h~����)#H��F��'\V[c�Ȳn�&�ss:��\\��dL���G�L�(`�����/�|h޻�,��_J�rB�$,0�冡rҼ`ʘ���,T`[�rq�@�O�1I�׬��Y�u�M��s@��X�r`����`Ҧ�Q�}+�������`-9�� ���DM����L�|$.�rKI0%���ϗ y�� ?'��T��
n��i'9��Ep/��4�`29����]xY5�x{2��r��գڒA�?�O��9p������O�À�7/s1�Q������zU$���q���ύ�빠{��	��EI�}fT��*0'�x�%�0'�x���0Fmfb���T�[���Y<`ʘ�eL	�!C9b���^��p��ˀ�X���,�?{�}��"*
��"*
��A_�"*
�PU��EAW�@EAW�节�������,@"( b( �� Ȋ ���* ���b("�0 �"�1��"(* ��"(
�0��
DT�"*
��DT�*���*�EAW�PU��EAW�Q_�DT�*��"����_Ȋ����(+$�k ��o����0
 ?��d��.o�d    (        ��     
  ( 8ԊR� �J QR*� Q T J*�J�)*�H
U$� @E$R� P
P ��    ��  D�
PF���=���j�=z����g���@ܣ��w�����yL��p ��J͹���j� �&�' ���OzB�uʸ�͟_}�W�9�Uo@��y�9��X��p=�  ��
 ���Q3:t���\Z������6���  	   ـa�}�m����o�i�-׀ ]^g�os��`�;�r޵^�M{�<�q�(�}P>�|ۛ��8�8���ܚ�� >��((P �
���}��x��l�ԫ��V���Y�>�A�/���V\�����:�������S���0M6YJ  )� 4b T:R���14 1 �`hQ�@J4������R� =� @ 
PSA� @Q��i�v@Jh �Ph�B�шh��Iˡ\�M�m������׀ ��wM��4=�>�������7v����]��ڼ�Ҩ�_K�}�O'�{O:��K� w�    P( @ =�-�ew��Q�w+������ ǯ�;R��>^�0��w�K�x}h���qs�r��  ���o]�=Ѹ zwz���{��.��ݼ����zu���{����/K�;��.�y<w�l� =!Sx�*��db41�P��T�@  O��CL LMD�*�"�1 ��BT�ԩJ� h ���IP���)�O����֗����V{��{ì=��B����y�UEt"����
����UE�UU�*�*|�?����$.�3�/��7��lY)�
aB�BH��L��3E��fi�8@���De*���U7���	�6����_OU���_�����u{K�f�T^/�$u	|{���n�z�q���\7sR��0�@�ޛ5��K�2�}y��}
���s�-3�
Z�#O�:7��^�̔�Zp�֤̚�F�
�(D�� \	X�hIaBE�	B � ġX�4�FT!U6��(�:A��4�4�C�I55� �.�&�X�]k���V�,k�iv@�U[����C��I.kF�Op��5��P"ge���B��B�k, �IKI��4e�B5$	m,�[=��߭]�伔B��;HHHbL?`}sSHJ��2HE�!
BJa$�<}��<��{�4B>��m%!$���Q����\H��H!rW#�"C�(�
,B�7n�	p�0!ak-��!P$�Q# b@# !YO�a���$"U+�P>�U�SD��7��I�.�ĉ���\5
&2繜7��(�$hQ�� q(cp1N$)��5 Q�0�F�K �I��FΏ!\ D���@dC! $�4#$b@%qRVFa'm��H�c/F+R�!N��(L��]���B�B�J��)!�K��k����υ>�r}>=!�Bނ7I`FaX{�����pԃ
��n!��-�4�$Դ��!�p�&WA � FF$	�Fa�d�$��������*ơ

��2%H�B$���_�!=*�� ��A`�H`	�@�LB5�Y��f�p��~f��a�l�|��HI�w�g:<�l9��'5���
*q"pɲ��m�d*�d_g��R_"{�P�d0$R!6�-����R�J��@�"�0I
eC��0��8JI&I����4�J����)���}�fwG�ٶK���o3|��5�	��Z��B��#ޓ�CG�!L%d!%�@ K�e�.�}�B�F��BA�X�A�$8�,B�"E��H$I���Ab��Dd�B-:��' �-������C��.��ԙs>zw�q�BO��A�1X�"H�a ��$`@*��@(0$#�,.�S	VҐ
0�{�Y��$&�ފB�ӱ6�)Hc\>v`B)�T�B�F!����6a��U�*\f0��%C0�R[���]	�~�;�HB�7����u�h M�ּ>aSJ�@� �Hţ�(F���n@��4`^H,)<�u���F�u�Y�Fڑ�rB41k!$iA#0����Y�dvpaL6yփrnpጦ&!� BEܡ�d��I#a�ip�D�+&i��;�vo��[w��\�p6B� h!H�!T�P��a����%�p`T¿+ �$0�K�Ea!�����!�$��_#a���5�D�@�F)%�HU�``�`@"�"G�Ԕ�`R48��)p�a)0%at��"MJ�B��r&k��M�n�f�jW��wE���)���%bč!B0�,���d�K�%2wr�@������;� Irr������ A�6�`��)�3&�ѳΎ)�hx�a�}aI�J�"E)�2F�)SP2ġr�p���L'3���	������\�Ʃ��������}M�� ��
Ą*B�L���y[���p��o_|\�2j����!0�R+ HJ�Bl@޷M:3��4`P��H� �[���0�Cdh�)� Kp�o�=�hB1D"%�0љ��]�百g��s���B�$l0�L��&l��Mk~���!s�9��a��&�Ōt �����`�d�`!3����a��*B!$i@(A"��I	$9�,�H;��GM=~
Zu`1�_BH$J�@
ģ $�B0��a
V��B��Ɖ#���!7�4�j\$�0�?.D��BbSJƄ
��`�@8�$hD�ޒH
�bdP��>%>Ѿ~��9��L�f��H[H�J���#�I�"Ec;e!$�P��3X�
h�DWU)T��NG4俧��'b��~�BƑ"Ĉƌ`�#)JD�u�T�������sw0�76I�k\�'���פ6}�%l��+_���\�8����p���2����M:��.q�k���sF�Ob�m�'v:��߱�C+�%J���
�9"A�!#��wc�!�$��BH�h�h��%��1�P�!�� 5�D
8��I���62	� ����X�bG0�y��˄�U��C ��daR��@��ť�>�G�$X�H��q4��K���čM@i��eHv"M&=z�l2�!�jH��E�>۠��Ex����$	0�a�z�0�u�p�� ��:HpѢ�Y�c�'�5K'�\��������7��߀��@�jD�$$�X%:�I�'�D�B4#S$t0��B$��޻y�gܒh��7͚�NCp2��K�b@�@�I.����0=��ed*F! �3�$.f}������E��3Z&�2\	Љ��753��bF�@��?lnʬLX�>�rI"C<�=�&��H�i({	�&�C`1(ȆSt��F�ċD�F4���i�F%(��#Bh�#1)(���Z�HИ��ih�����H�0�,%6��R��j�C[3sR��-���6�7��0jbS4��
¸�t��tCH��y�l�?��^�
!1�"�+
H�e�����Z� 0h��M�J�(�����`D(kD4	�
��l֬����a.XВ
ƕ�-BB	)�)�G�×
A�$i0�a���@�RI�`��
`3;����	��ن�\�bB�*@*1�Ja.������~ P�T T#RP!J|��C&�i	 A�	���aUaR5"�5�nBJ�P%�-˒���d5����a�Dc���R((�!I!*f���,K��5������M�����_4:��.���sP'iaF1�D� ���b�I\m&j�|6�JH�d�04�H�-�V���$�+Ss'�Ĝ�Z��ӡ���5RB5 ��h�"��"T��09
b���sЋ1����z�a˻�R�!�2a%e&&������5�����	������J&�M��au�L�8�!v�K�����lKkd�fN�N^?t����*D.��v��4}ee�CI `0��by�D�>z$H$j�\�q	�-�
m�C���s~�	����m�d��)��\a����z#&�A���r�i ���0�!LcR�!p��o)2{Gq&k����/3a���H��H�O��_���t=�gL��ǮN��a�$�T
LSn�K
��Ȅ<ߧ)[�K��Y�q��bF\5.k��n\0��0ԛ���B���� KB�� tG8�@�*`F���߾�Ό n0�H�!XV�i.hdc�5��u����[����F��3SF�$0�q��!���#:ȓ
e��a�H�M_�o1�P�Zd)��aH0�A"E�$*�
�(� KliZ+$�dc6�@��9�!2e�
���L%275��e�kp�orl!H�P�
nS5�$�Ͳ��
�����      �  �@    @ m� ��K(   �� [@H�  m�~���t��[y'iagm��=a�� m�m�H������5�@����յT�=!P�R��Ԓn�s%��yu���:6�����`k��ra�쯶�c���@V�*ҭT�R�8�m��H�k,�֎�e^�m��6�-`E�9�v�ճY��c�r;�LRKJ��t��ݸ�,��Ѷ� ��ڶ  �}��m�  q�N��    l A�	)V���y�6��U��a��P-�l�I��kYd�.���wc�T�T���ݲ��k�J�[6��MͩUV��k������E@�v����hlH ���n�l�`8�M�����l���J�I�h	 m�_nZUѠ�DEPTTձ6� 6�  ��}��   �����kmm[sm 뭹��@��� �ܣ<�,��J�J�*�R춀m��j�m���	6� ��@ :۶m��6����$ �I�m� ���F�m��m����iXl�l� � 8qn�v  ��	���T8�j�k5�`p�� )B�d����mz� �`  k���`�96�� lZm�Wfؐ  z����m�i �ʹܒ�k ����*I&��蔛\�۶��8  mk3��F�yZ�WfA�f���L��z�5s���r� 8��������lȑ�������6Z�$L�kt�m�M����T�m��
9`:���ʧn6�U [Bu�:[BA���m����_\wֻ@-4����U��_�W� *����v�m��� m��s$ &���N�m��	/UY$�H-�U���#cb���:ķa�T�������j����5J�Ljv3�=S��2@�+�Փd�vj��V��U��jV�H�� 5*�[k���r+�Pg�[l�F�98a������
��(��� �\<���;m&��cYۣ&6� �ʃ맛�ڙL�+�������` ����n�n��kUJ�*�t�9�:*v� 5���%�vֻ riu����� U�!�T�(�տ[�k��jMjô�n�Vl�,tv��2:x�����u9͵��Wr�+s��E+��<���M�[@ -&�E-5�� �@   $ n��0[@$ mH$� ղnò��TQ�[�� ݤ�%��m�`Hm�8��`��m��n֍*�	D��UT  � v�9��9 8-�f�`h�[I� Kh6� m��`8$2]�[&�[`H�WYv�&�p�f��2Y@�ݰӬ1��ܶ�   ��	��8  h[R�W ۶I�lWX�3�@  �>��Em�R@ � [d�m�&�m�۶��m� 	   @ -��`8��5p@��U*����� $�6���lM��RȦ�V��0 Em�$-���6��U-1��S�J��ʻU*�WUTw�0<�P  � �m�iU�$���� H���li0 @ i2j�`�U�E7i���4�mk[E�l�Sl�[[m�@�j�V������̪��}����yY#Z�#k7mKT n�[(+�PUT�p��@�5)mU���	@�f�ރ]���uvL�xV���OյP9��q�mps��E�t��ۤ묡�Ѷ�u�2����ӗ -�$<	  m��J�]�mN�)$�!�`��}�Ƶ��V�:��6��/,J���<mU*�q��]��m*UU[C�U���i6�U�m������)VڪX-���O���)y�d�U��*�YW��T�>V�2��-�ph�&�
�*Cv�u����*� ��-` Tڕj��e]�H!�Vܓ�ڐ6�mW��[YEV��T؃bW;�-� $>>��-�6�[@ �`m��R�.!�@�W=l�l����Vr�T98
Z��j(�m��+�m��-�j�ɱ�Aj��X��8������   l�m� m&�%MNp��ekVݲ� �iV��
�*�٠'���{ETB졻B۱L��Z�6��&��Bn6R��slm������۷l說�`DUmh`��m�  �@�c���^�����q�l�1e�.�B�v��
�p ��   5���� �����UFt7+���j�p����  [T(��v<v�xwM#�� v�    ����-UWU+$�]�YUI�Q6�� m� ��m�l�   �t��l�r�m��ob�z�l gt��mkk5Ĝ � m�l ����nd�  l:�e����  � �6����W�n���ΐlۖ�פ�� ��[wnر�:$ �����]����m��6n��:�
�j���X��VV�*4vP����P�p2a�4n��Cض�F�(� �@Pv�јb���J@U[�8iT6 :ꔝ'��T�o � $H�jNp   �m� $i�%��uu��4]�]�L� -��i��M/3m�  BAɵ����[nղ�]�6�ܶ�D�!��-UR�ʪX��2ǎ` 8 [M���n�6^��l%��J� R���[;�Q��i�,�l��c����[$h�U*�Ű��1��r�V ܒ��ͷ��  m�u]� U�����Ak=M��U���>��V�U*ƦU�V��i6�+	�9��M��79�JiA����κ/�l�l��/TU2��m.�lm� ����t �`[wE��Y����۶�l-6   ����,�m�-�Ӵ��ݳ��$��Z�`vٻ`mz'i���4��m���	�Fٶ ���5��Mv�U�M�uA[-m���h��iֲ��q#��U�a�Ӫ]�����T�o]�6���  t�Md�@8巒��$ pnt۵�Z�8  � �`'A��;.K9��yz8��:��K$�`K��%���q,�7�b�+I� ph� H    mq��[vݻh�o�� $�@ �m,�-�Hí�h  ��sm�  -*U��{)<�*T���T�h��Pr��m�A jtZ���8ڐ���UU.v��۔��� �֖��bڝ�N�[[d݀   �ɹ��.� j��[�\m �u�u� 6ؐKh�Ӻ��9,��h�����6ٲ�hp!���� @�l���I#i4�&&������8B@[A�ks`m�m 	   m��[���6�m�P�W�b�	��P�T�dyU�%V�ڠ��UP
��Q�,uK�� �p�!mm�h���T���۶�ݶ�m$�H a�tA�HMJKPW�kj��@q�`6�mHmm�U���$���6�h�٤���v�\��jsK��/3.�>V�e@�UU����h�0�kHm��-�u�g-�7��V��k���� ��Y��l�K��J�]!*�p
�[U6턴Ć������I����,		 �9�l��*Ѧ��Z��T��@  m��[u�pqU*�U�*ʷ��Za�d.��lβK�F�k6��ƴf� �]���,�{-`��m�� ���m��-�`m�Km��I[-�-��m�p �a��lh    q�r:�L��m�j�jڬd��,�ZP �l���n��  �4]��H8H $.�T�np m�F�*��g�
�i)Kh ږ�� �D;�*D�m�$8�6�d� -6��p6�9v�̴[@�E�5������m$k�����l �M�I-��	 �mr��*���U�v��-$�;|���.��V�t-��ŷv���h	�m����N� ���E�ku�Nn��6ݵ��#�� p[m� ֻ-��nm��[WI���tUU��,�<�]�m�tS���Ki"C���� �#m��J���[W�񱏻'�[��Xi�m��-�Jl2���l$p[V��`-�D�m�H v�h  ��hH�6�M��m� s{V�崑�m��h [AJݶ	���bK��Yd��� 6� 	å���ֱ��0I��:�l 8mf���ݶ��� Im-��bN %���m A&٪��T�\K:Bx�q�U餠�l ]�kA"F� f�m�lm��6ȧh6����i   ۴�F���[�ɯ� �5h����V�t�9z�sm�H�e�������{��
�ت�"xE(���@���	�_��i�DRDB �"i"/A6���#�9@ڦ#�� Ғ.�'�>B�@0B��O�J���'Q:���?i8 =���`'�Ђ���ŀA�H��S��@���0� ��P/��F CHt
!����iNy6���A$ ^ ��Ry L]�Da�$E�t:+����GH���D9D�^��� �"yШ/E��h
��N��8+�u O��!��P D1N'6ȌY�z�mT=A4��M��j)��DC > uX�ȏS�B�+�Ê����t*|�	ȉ��Xz*�
�2��P��`�U�6��j>�>���O�w��Z�࠰ *G��J�������q���pG�'��:u1U�a ������@�刔pA4qT���:ۡH��������z���@z��:"V!	@"��P�Q�aV�KȊ� ��t���D@��@D�(@"� !��>@H"�Z�����Yt @�V��Pt���]\O������_�W�E����*@R!D� 9jA1PZ0F����i��)�� �L�Ò �m�i��9!M����1�Iݶ��R�=f�����r%v�ۦA�����{���*�骨
��*��[;C��nv�6�m6��*��w�m���9�VBn��!��mA�*blݷh����1ecR�t���n6�kDͪvzY\l��W��@m�Ƌg[�.�\�q�m�O"�K9�f��W1����)P�;g:]��+D]���c�
��ۚ���e�	��8�F#e��c����jm�q��l��M���Ҫ�w2���y�=\�P< E	�E;�g%��:0K��iٜ����:(ƻ(�ٵ�m���X��g��^1�n(��H\Y&Kp6�����(�)fvٓ�B�;j�ˠ -�nl[prsuiLܸ5s�v��7i�h�t���r���J�)
��n�"6hC=L���l�M�u�S�r��ۥW��t�0������<��@1:�G7�<k��7WRA��K.��$Z6+k.�u�v� ��M��nc��"t�$��6����J����f�U�K�#+M�<��eD�fÝ��r�3�6늻JF�wT[�Y;��ӳy�n�M�#��Bli��s]� ݇SY؞q:�	yU�X4�;cP��T�΋��S���7��+$��*�%����u�Ī��a�k�ܖu�5F�b�m�uJ�S���Ҭv���:��f������ݗ��������䖶xzKHuSHr�t�:t=mN�t�SW>�Z-��u,N�]��7>)Q���g���MY0��� ѵűe6��n���/C�	��4�s6��A�V·%m\�ERr�S���8��3J���ђI��&�{i��i��"VE�d��R˶�X��/=Rj�βu ���ń©��$��,u�:ֶƨ%tfڑZcBV��v�3"��k�0�<8�M;m6-v@��D{T�*=�r�S�Zxy@6���hC�P�x�b�~?*��)�C�:��CJ<���t<}��Ң0"�`�_jR�nм�	�s���۰�I��7�4I�c`.��u�89]����͵wj�fRz�6Һ����ЛV#���[fଖ.{Uۆ�"���z��Ԫ����n��s���Eo9�]�^.���֌Ӻ[��>�gX:ٶ�0ۡ�� �N�k&Y�u�|Ơ��b�Dȩu�7i�^W��:��35&fMY5�p�-!�W�*��󜌤��-ɓ332坝���\���;p��n|�ؘ��<f��,���h�� �>u�? ���@����Bsq�Cqh�V���8�j�*���_j�-���{"q�'�qȴ�}�@����}�@�ڴs��I-�(Fز5"�*���_j�-v��|�eՠ�\�&�0"JDӏ@���v���Nk�5����"!.���n������C[�rh��*�tC�9���k��'��Yk�1ؒR�u
�3o�~���Z���& <��@y���E1H�2U9�v��,�S�@V�@�j�"<�����o<��j�-v����L_bq'"�*���_j�-v��_j��ϒE�`E�D����V�!D&���v�;�Ô'���`|��1�$���p�Z�e4�}�@��l��s]��D(}ϐL�)�=-�����:�NwZ�8׻:$�顮Ӹ�O1=sfI�H�bI����r��uw����V���M��l�4�b��v�ۘ���-�6<r�ﾪ� ～�6(�D��iǠr��~����=�(�U @b.������~]�z��Ҭ�1Fԉ�����`���- �<r��S��bȇ�9�_j�:���<r��`�}R�6����.�:cL�g������1��u�HxFۮ�\e��7:���<���)r-���@��ڴ��h��V�g�I)�2'�`~��w�	&���v�;��׻�`~��j��
GŠv�V����i������W|��3�ȜbW�^�n����& <��A���C����x�MsZ��rN}�fI��iB$?�R-����}�@�v��_j�;�r�xcI�bY>#y�g7mB�W�Ӏk�ܛ^4*�Q�-3�O]���D��iǠ~��Zk�h��W����*���Q�/2d�FF�hn-̒�x��1�Z����=��'�ő�Z��M����]��h��Z��i�b�	�28	�C�*��=��-�ڴݲ���$w)�_�G�s��h�V���S@�]�@��H�m}#I�C�l'jW�dWq ���74�2�r�-�ktJ���|�{N�cNwn޳��ibg�xJ8��MS��+�n��zٴl�%اf�B�f�B*�L��B��͒H�^�DY:�;{�3!�I%�`w��]���VNɘ9eX�ۂ��#tr{tS����Ŏ���-�.UY��dy�˂��t`�X�M���Y���{����'�����e��m���um�K�:�&�uz�{O1)M���r��b�k36�L���6L����@\�fȡǊ'���S���cg<��_?U�w��h孃��R�Ϸ34@zc���ZG�@y͆�rܸ&�YR�����/���Y�@��)�Z�V�yؒ��Ldi����-즁��S@������`t%	,���*��r��GBmVgq:�����s��f%��ggvK&Q��<�t��)�Y��!�_O��h��^���wmq`v��ݔ�S5-��a=����� 3��HÈI턗�P�Fa9?[�;�,ٵ��(�Ìr�P�d�S�3gy�${�� $�-�mf]]��Nj��9�v�>�,���vsV�޾ՠ\���q쉑�x�p�=&�&9h��@H��W{Wg���&�ш�gf�=��%q\Dt�|*�ʷ���.NYH�>���ߟ��Z�9h	2K@zc��=%J/2�fZ��QSUN�ϧ5�B������o��k�h��W��⍩oqi'���ܓ����!~$Ra�R9�����Zz�V�{���DcD<r8��ڴ]�@�}�@�ڴ��0MbZL_cs"�-v�����j�/j�/mCǚ�6�cwk�.��GK�H��v6VW�6[j��d�K�r�H@�$��$Z��Z��/j�/]�@�lƖ%ALRGqh�S}�bG����^>ՠ\��ǲ&F1�M�@�}�@�v������h�kcX޶����@�v������h�:��Ch�n����I>�O�[��j�!�h��h��������^�V����4�R ���Q�Kh�(,:�s�;������֗�z
j�-�ݴ�x��*�6�7�=}<h�ՠ^�V�z�V�{�����"2Hh�ՠG�Z<r�͂Τ��ʻF���n-�ڴ�ڴ�)�^;V�R�.S"B�$Z��Z��/�@�v���%�1I1��Z��?���/�z�yh��]� �"d,P���S����~wk���W]�mکT�+�V:��g]`��`�Zx��v1�a��Nw+�v���XU_h���P2/n�&���#��v=�f�HpY��
.�����s�/O/<җ����×�v=��75��]u]����L�����FRnՎ�8$�	�iu�(^�m�l��vmb�q�LJ�I����>��k[ \��h�j�d��浙�|��*�l;�b�=��s��p�v�U1�wb�#�m����r�*���z��o5��m ���y%�#�-� ;�����H(�Z�h��h�S@�v� �{��#k"Jd�8���@G6	�%�:䘀|���'�#mțx��@�l��x�Z�z�ϱT�V��v��&A,bȇ�n耝�Z�9���@y͂��&���5L�$��7	�[g�OgD��&4��B��띈���k�w���������sa�������g� �yA��X�'�@����GJ����A��b�����"DF"�F"1 �������!��������bPs��Ǡ~��-즁��נU{^�ܷǲ&F1���#� :ۘ����� Hؖ7�p�19&���נ_�W���kK �ͫ�/��p/�MKj����(Y��FM�ь��:Ij�"]��9�n{O&	4F�D�Ȝ�����@��)������@�{2��cR'2��M��6��Q�v�X�zl:??_=���$^��&A,�<i�ㆀwoU��Nk���/? ���P�!"�#	� ?��W��ϴ�8�vij��x9�=H�����B�T�+��	���'�H@ �E9@M��aU
�>5(l����!B�����TJT"M]�8����')tU#c���$�>�f���$b�1v�z'<HR!���(�ui\+
�D��1_��[��)��G!C�R$$bA��%z��`��lCɈ��:��TƄ|*�T�E<ֶ,j�D_@H�Px#�����p�!O �@袯Ȯ%P�!!B�J?�!%��rl�,�f���b�}#nI4=��b��@���?f֖I/B����`�i�^ ����*��@�ܾ��=��qw���v�`�1 ��cLĜM\L`�Y�m�N:�ӀN��Ms����;�\�x��8�홊I�D��/�� ��h]���~A���\��1{șǃn��W�ُw�����`~ͭ/ޙ;}�,o[QD��ܓ@���zU�z{>�._O}}4�{��4F�D�Ȝ�6	D=�ޛ����3sj��E("�Ѐ, ���A�P]�&�0QW��[���ܓ�}���-ˑ�\�sS`~ͭ,^��P����z~_w�������X&�\�%��׭cs�9��f�s�����籬GF��k��B卡)�����*UNT�����������l�=͞ID~a��q`f�	VRj��t����l�%	���`}�\X�f��%�2�M����
����M��k��ޝ�g�&���*���9��LoG��1^��`��`c�ٰ�	����]��uU2T�J�sN�>�6�%����������9���XkҨ�؄�On�Y�1u\�Z[�$�l�����h���b�^���m��렠��u*�\�9��k� ���Ŷ��<'7u��ڋ/�;3��;^�����k�����;�K�G:�9\�&oU�۶��5t���t�������c^��e-���8b��e����&i��lA�i�a��[e�M�G=t�N�T,���&�`�4��ӷ .�-Ϙ�� ����3,×Zº��*��d�[��q�d�^�"h��\/m[��f�����Q!�9$�q_�~��6s_B���ޫ ��92YS-SJdNH��v��}���h{}4�����E��y��ҐM47�|���}�mY���(��������;���j)��d�*ULӰ�P��ޫ<�7���>��vP�$��y��r�*�MIN��X�6lJ�+����- �;f�߻rQ�& ��P�%����pb��;9����vúџL����+c��5V�M�� T�j�Os�3g5��fהDz"!/�9��6���#ĺD�r��`f�k��IdBP&DR �W�`��D9�3�~���`~�w]�K�BIL���'�F��<m8��M���}�}����o�~��/���9ΪЇ���Қ��P�=�ޛ��`f�k��K�o��s��؆��Ȓ��=��`tF�o?���`c�ٰ<��[��n���ͥ�on��q h��+�tK��۞�X7&��mv�:�,$?�w����^M �"ɚޞ��ͫ��/�>��v�Q
7|�s�b�r�ʕS4� foU�&��,�{���9����wA"i1c2E�94�<h��Z\�ϳ q���"�9�HJ��d��A��=��%hK�n���`wuX�Si��@ FĤ4=�����/���s�h{�}wƁ޺bK<���x؈���- w9����-����^���4zq���m�n
c��4�-�֥��D�6�=�4��5�;\[n+U:s�Zq~ �o����M�����/���;ڼЇ��Hy�I4��o�#�}��ޝ�`}�W�!&�3�%2YS-Sn�34�ͮ,��vr�	&ϻzh��h��VO�%�&�jCC�"ޭ�`v�X�ZX~PD8��H��`�
"Q�<�N!���7߽�-DO� �H��Ǒ����Ձ�%����76��3g5�P��3��SND1ȝl�DҔ�j[ѭ���\�u��HxA��ۓK#�u[������wg�q���I�=���h�e4�ڽ�~@s��@3�%�g� D�7��vR��Ӽ��ޫ �ͫ�	zd͕ĵ��50oR�Z���?��H�}�^��@�h��H��<m:v�sj�7�ڰ3�,9DB������{����$<�$�yl�?���o~��{ޛ ���`b�"�HBQ�333�kr��
"Ǆ�����nQ�r��6��z��nL.��t��A��z���]q{]mr�n�s�X��A�;��՛OOizus���F�ʆ�	J�6�SKn����6�4�\<���j�.�К��+vvz��R��=/dd�w!��t�8e[6F�S�i��;��n�K�3v����C�����L�̐t�;�C���H���B�n�׽��w�zy� �����n��ɖ7P���S�.��krlz�.���lמ2iN��i��=})�U�נ�l��3�ݾ���y��F9��F�hs��䃻z��z���W�6fk)�R��U2K�)������ڳ�J���<��=����&,�#�I���脔9�w����֬n͇%
P�v�X�M�.S)�K��w6Ձ�B���;��v�X�mY�����~v�p���<�����׍>S�n:�m2����i�%3]�����wq%�0o���yw�zol��������V-�C�*���$�#��	=��[<�6��O� ��D4h(�(T\7T`�T�z'h~T/C�禁�_nhr׾�>� ��lC���I�$���M���=�yv���}4���h���)��&���ݽ�X�zlw6�:!7ٽV��<��ģ��#s4
���/z�~ ������]-����,4�8<W�m�������c��H�V��͍���-�����P�US$�R����z����~ �ޫw6ס/�5�����A,�QI��qI4�پ��=����{�@-ͫ�M��M�.S)�UMU�ݿ�nI��{7*��1F�b�EX 
���ʟ}3����$�����嵬%�&T�2�P�:������l��f|�n��.\���I##�Ǡ�l�=�}�����������׸�����9۱�񝞉�MA����d��GA�R�8u�K�n}��gل��$�6�i!�9$�}�M>͵`c���IG�ݽV���,����I�UU��fڿB�
d����{�V������H�*%7RM'.j]Q`k���6��Q�:��M����`g۬�5QLUS2J�uNÒ���ޫ�oM��eia��LlB$�+�Tӂh1
W�����w�7�Z��_��hx���RI4
�l�J=�߼|�=�`�mX���c��[��5ַ���y�^WB�#�t�n-,O,�����wa�k�۴hh�?�{�x�-v� ������<��=�yZig�50X�ڐ�-v���|�6��`s��7�/��I�Vj!{I$dc8�ݾ���4��g�|��g��~���׉'#mƒҪ���JD�w�V��Ł����(Iz$�Ϸ�V���S%�2�6�9���7�,(IG�Q}~���ޫ �}�nI�Z]��q_��Ĕ�B,X����a���iNҮ�`D������Fv(E(o��y �� l����%0B��Mf=9�!�tR4�|��H|`rIN�|�1U���O�f��� p�6�޳k�muԺ�]�g�М�c��m� ���-�7#aJ���zs�S[�m���� ѳ�
����#s�8��zoA.���d������O,�Ŕe5)��m�����mR�5WS�u�,�Hn�(UR�)���wc�˷n���jj��%fў�*��n֝�.�(��j�8�8�	�S9Ô��c��g���巶��ݜb����-�k�����G�i���\02a�z�i��68�l�A���q+ɓ��g*��5J��*���^���m L���B�R ���km�6��uhmr�e�Z:%�n�t[�L��C�Ҭ��m=�cC-��Nݥ(�87N��X�zI�㝎�nw���3����#i-[�۫6���Ƴ����\�Yjd��gk[#���R���1��+6��=c��o,��F��(���VuyUiQ�(��]���{
w���`��1pd�K1�\��u݄'Z�ہN��.M���  �5�S��s*���@r��(��Sv�ԼD�����ݚPA��}�}78�������8�JL9��:���JEv
�ꓢmq�8�&PP-�Y䝕(*��h��Ѷ�f�T��=�;s/	��4c<*֬$�Ѧ��	%��n62I�`]���vj̸%�uU![;*����
t��gMgh�p�Fӣ[mfC*4�*��n��s�]:��(z+���0�1��'f��J��i�p)��6&�����t,2�nn��y����L��kY���n�4�^��Ƭ�5����
tX�q;v��=Ip�����gj G��ԩ���F�f��T��QZt�Mq,��imD��JP���`U�f�I[4�Y����:�^�Mɴ�q���n�Ү�u�5�9�jx���~���=�G7g����aD�iek.h��k�>����gӛiB���(V��;v�f�͆���p<sD�M��=[ �� TU,��<A5�|}N;������'D�><;A��������~�:x�o������J.�5'��X[A��v[�*Sk��/%B�3].=��,�_�H��k�ٶ�b���hDӵ�l6W���N�M;�v�<���۶0j�<���r8y�Y'c��>���d5m��iePY��p��i{kp�B���b{I�h�Q�r+/����Ε�@�dR�V�8�y�v<r�T�V���v�j�&�۰��g�����J���̺À�"�Z�5u�ֵ���.B8�������8yq�9�_-Z˒�655A����f$��|�FӘ�q�
�����^fՀfn�(�ók��y��)��fIR����W��!��U����`}]�}��Q�{��&,ɒ2I4��7��Vt7�=��;7��Ƶ�a�A�uD����I>����������V�!7��V<4���66���v�ٟ}��o��o��y۹�w�Œ�����i��Ĥ0��9�]��B�s�δ;��QޔoU[��wu����j�J�ID����z�36��6הG�P���O���ޔۙ��5-�b���$��}��~�V� ���M3�+JRQ	.�K�����zw��oٵ~K��{}�9��e�n��j�oW��v�=�bG�}4�zh���'�S��'.j]QaС�Ws����ڰ�
<�O���=��[���*��')�~��@��b�ޟ�����9]�@��Lx�q�i(�́��Đֹذ.3�Ү8e�Oh�`!�v�ayt��}�=��l��&,ɍ`ܟ�-���y۹�r�W��Dz} {{�`s^byxL��r��߳m_$�ft�; ����37j�	/(�2v�Kk�%�l�sJ��O�w$�����������D����nI��j������UT��J%�;D/$�S=��Xw�Vۛj�DD(�;�� [|�I��q���M �z�
P��������>ݫ�c�p#욣˗PڐӸYz:�8�c�m�ĝ-U˹.���%	�������y�9#:��~;zՁ����v�(���ޫ�~�O����M5��~�վ�3�s��wz��6��$�ۼ�̫dH�0R- ����w��Of%�}��}�����A)ʺBR�5.��=
#�3�ޫ��Z�?l�н�'�P�,D ��)
�D �X��F �U�A�U���?�����ܓ����M^S*�����77mX����y�����33j�Ź���)��-Ԓ�v��t�7�y��;uq)�:�}5�c(;Ҍ�k��ݗF�3P50X�&�~�~��[f�ff�G��֬�@β��J�[�74�sv��Jd;��`{��V盳~ă���I��q��1�&�v�M���=�q_y���4��"1)�nM/_{�hW�z{l�w�h�W'�D� �b�f��vנz���_�3w���ݵ`\$BP	&�
D-b�(ѡ�{����V���f]�u�U�n�9���]�(�P1�.y�9ஈw��[�iܻ[;����[���VqLo/X箉ֱ*���Z�u��ԩ�����6��;e`��߬�|��S9�fՍf����'C$v;\�$�f�\[�Wh�oN"�ݦP��S��Nv�����Yg\�g�jl��6�Egz��;Y��L2�k#�]�!��Ki�5$v䜉קm�rnUv���Z��k`�b:���6�,$�V��j>��<b�:���@>�ڰ37n#�~a�=��պ�1�*������7u 7&��R�Ih�پ�*�#y"$�7$�-�`}����	�;��w����rص��CM���a�'�]��3���37jáD=������	��UJjFܒ���<������ߵ��A�A�A�C���L����[~��������6 �666=��߮�A����7{���;v?�[���p"Msp�X:ΜnM�ɉ4�\D�컺�[�{7����W��e��˙�m�k5��<������~��A��������A��������"�������ߵ��A�A�A�A�~��8S,ՙ4[�sZ��A��������Dvc'_"1t*ApA�A��s�؃� � � � ����lA�lllo���� ��ʑ�A������9ur]j\�.�F�A��������y�߿kb �`��67���[y{��y���%�yc�fd�$��؃� � ؿ���ds���[y�~���<��������<���`������A�lll|�߉3&S� a���kb �`�`�`�}�ߵ��A�A�A�A��~��A�A�A�A��~�v �6667��~��A�����~?a�nI&e�U�*F�]��b�Lqۘ hxә�QzR��ڃ�7a.���Y�35�lA�lll}�߸lA�lll{�_�]�<������ߵ��lllo���� �666?��L���2�%��.f��<����k����b dr67����؃� � � � �߿����A�A�A�A��~��D,ll~�!rkZњ�m�[��y�߿kb �`�`�`�}�ߵ��A�Bt��G�~A�tAA� ��p؃� � � � ���~�y�{�.kY�5�nXkY�lA�ll�~���<��������<����k���A�A�,o~���<�������5fM���f���A�A�A�A��~��A�A�A�Q;�_�]�<������ߵ��A�A�A�A����؃� � � �"�D$��?4x�t��ɨK�Rt�`�*�tK���v&ݬ�+[u�I��]�����9֥˭\���� � � � ��_��b �`�`�`�{���lA�lllo������ �`�`�`��~��b �`�`�`����$��%������Wb �`�`�`�{���lA�B����߿kb �`�`�`��~��b �`�`�������0��
!L�ނdm]!)R�5U`��X����P�y���;��h���*m˚R�ÒP�{�+:{��}��`RP�����"*�������e.`�bx�&�h�ՠ�� �m�f��wH�s"�)�T���=����\u���r�s�Ƒ�+tX[���[��c�I<qp�M �m�f�Q�gOs���D���f��,USU`��|�Bl��`gOs��v�С$��DL�.��jYL��uNjj��zՁ��볢"!�;��w���Ű�\�T9sN\Ұ�J!�Ws����@ɨ�T���/2�w��6<`�Z�l�=��ޟ�����>��vV�H�Q�xm��	J�Jn��T��hQ'Sm�kU���7mJJ�v�����2���2�:�#���5kn3�lW!+U�Y^�ⶶ-r�:n�����=���ۊ�=�U�9.x�f�˽�@W�3i�3<Wm�*�;Y�f�����c�I�.��:s�T�	�"N3��/�p}����Fڻ)r��e�d�ʘ�<��=U�.�S!�mЗ<�u���{��~w}�~����������i��d���^����nLe,�^��ޝ�_{.��J�L�p��V}�j��gu�K����L�0^�aӍI4����M�����(K�}ޫ ��~�m�VF'�nf���Z��4��H�ޚｹ�w��G##�<Ni�t$�v�XouX��D$��'�~���sUD�9nX����77j��[�ߗ�3���ۛV�$�J���{d3��['���S	�/�B�J]�z�rlz�.�qZ�]�GW��pP5~����H<r�G7������:�oWD�r:�˚r敁�'5ި����A �X�A�G�T�F1�$��@b$ R%�L�@I(���E���H(@�� D�H��#�0"L�f��(����߂��V���>ݵ}�f�pf�1UL�*A�; �ޫ ���g�<�����X��v33`���ݢ�+7/wu y���*@y�k��M�oU��+��#|
�fi5V}�j��D}��� goU�~�f���pz�@İqa��SE�O��ێ�M�-2�#=��v�bQ+i��������|�Q��@����|�����m�м�I}!���X�=eMT�!.T��m �Ɉ�M@t�R�9k���Ty(�2��	&�I�rܰ*�l;���{�ٹ��!"�,�R/�(	��'��#�� u 	�!�v���њ�	:��p4�$�����Ez=b��LP8���W"A D���z���$(��%P̀X�h�� �	�DG�P��|�I<��Ќ4!��xth�$CxcX�H(�*2�P��1�����^�C 5ڇ�����?�"�i�{���� xJ���O
���|��É���ziا O_�V������ ��Q�(s�}��ܓ���f䓝���n�%&擙��P�y�ߕ��=�@��@;m���\�ģJ`�SJ�͝�`rI%����w���Ib]����w��Q���2bH�Ҁ(���<�����=���	�]dK��ڊ���k��w�o�az��S-H:��=	>����3����wmt%��C�}�`s;��ڪBNU)��@$�I �- �Ɉn�`���ۘ��@�s@�]�O(P޽� ��6rT�[$�#��/3i&IhnL@ɨ6�������"�=�pܓ�v{sY�2<�8�����f��n�k�h�����3� `1��5�����V-�)�ؑ5vq�c��]e����i�I�$����M����j�:�k���PLJ!�srM��H	2K@;rb rM@I�˛�](Ҙ(�73@�v���� �m�-���j�h��(��
E��w�zo�4[w4Wj�;��bo͘f'�#��٠�@��)�qvנ<���a��PFF�_8,cl�8-ȷW��{P �n�n�5�b֦,xNKJ��W�i��q�:��o[�O��|k?�����+CJnj���st�h�s	<����AiV(��6�8�G)�b��yp��=Y��y�N�ǻ<�,ғk��3��sۆ�E�nw�`�yhw;Y#q��})��U��������:�l�J\�����qЩB�;f\���N<~���w���.HfjM8�MK �מ�)筎F��[pi�����ܡ�͓�ɠd$lrN�������S@��@9�٠v��o2��x�&�h�dܘ�=�j�� 'Q.�77d�D����<ݛ ��mY�Cy�<h��@9��r184��$z��4+k�;�j��3w�z�\�&%Y1'2F�hVנ{3-���W�z-��:뱡2,Ra��49f����q��6y����}��e�{���Ł�Nh5�b�)������-����ݵ��{�6��2��u2�%֮�^�ٽC�E�%
�%	
!lz(��~�����}6�e4�{~B6a��(9�w��绳g%���,{�6<5��e�䍸���{���1��(o����6�	��v���S)t�R�+,77q �9hnL@��\���$��S#��䓄�)�!�s�znT��m�hvX�Q��z���ww�����M:x1�MȿU���w������}�g��Z�|Ɯ�N!�I�>�PrL@t�- �ɋ�U}�]�s�	�D�LȊ��W��r�բu4���!!��E$B�J.P�>�ί���{�X���O�#j`��z+�ZWmz}�já(y=�6��2����ԕ5N�Ǜ�`rQ���~wM���k�%%	~I	F�/T�:n�R�J��c�ɮ{��;��r�×�{F��ˋn���m")�1�"r?�w��hVנ}�������ޛ��hjY�TN0�f��m{�=]��*���ϳ? �}��˾��<�Li�CR8��ڴ}��y����4+k�/2�Y�G�x!��"�:�k�/-��8��C���}��BNՠ��c�������	�*@u�1��bۓ����O|q˫[�)seHF䧣���獹/MT��MwWg1T��-{��p7U3K���l�۳`c���$�0�{���O�#j`�rM�����dB�Jd������� �wj��yDL���LŦ*n���M�Ͻ�?}�j�9m�;^���&�5L_c���BI/�Iz!Ef�ج�ޫ��l�z�%=]�M���45,�*	�t4��ݫ�%����{�6��7$� ||�"�! �����v�r]d�v0h�^�E4]�Ru�-����]"�h+��M��݊ݜ�-����Z��N�8�����6M��'����*�u�(qjS.��9��g��\RS��kb�ZI��3�A�$t%�ӳB���M���=i�ѾM�6���t�����6������e��A��8!v]4��R榳�^w��rH�9$z���绻�����?w��L���-t�Q�4o5�x�^�<J`N�(����D���wv��{�sL���%�'�ܘ��H� t�P�Y�G�x�<iI���^�>Ďw����ޚ;^��H;o�1��pi;wq���H�����1����b�9��e�M�)��V����1���=ݛ�Dz!B��{�`o��_�|�SԒh\�z���*@;rb�IEwJ�+@��������	�|���;���Ƃ���u��GD���7��ݙ��Q􍱱9 ������m� �ݯ�<�$����7��&If�ELѣ5�f��}�zq��D�9&{{V<͛���D$�1�K8���敀owU���ٳВP����{�ۚ\��ec���!�I4=�
O�{�`s��6��j��%�
&w��X���.i�T�ԩn���Ǜ�`zvo~_�3�����l���P���ʃ߄@�b}v),gHy3�$jz���e�t��v���7�;9dXC=���� �j_9�nL@���Q��s� �m��v�hW�z�n�����y��
6���UU`��`|�vl�P�
����QTG���� ��uX�uJjf-�U*d�uUa��{;�6ݽj�9m��v����7�����*@>��~� G?j�I����þ���2کn$�����vnL�m��p�Lȉe�)AC���}����$y������v����ٟ�s�֬y�e.�i�r�&����3�ڿB��ή,�zՀ}��~Q٘�]%�:
�ڕ#�����?nm�:<�)e����_M ���r1��MIUaВv��`��`�mXLRI(G`u�� V+@ @Ť"U�
{﹭}��';��\���4[�1�Ұ�6�%�
'��_ v��`o;w4�AS�cLC�X��1���yΉv�[c��k 
�z�$�DT��p��bmL�9$��٠�@����}�ߐ���9}�x����<l`���n��$�l�޵`��`�m_��_$^�`���s�2B1�4v�s@9��g�M���`��`nJx!�ކA��RL�^٠��@;�f�����~� 罍y�&�ć�h�f��js��G5��U}�VǠ�$c	'M�G��8�"���<�G"b)��4��2#b�
�����60�@pČ1V, C���7�Q~ �4|]8#w	09��`�%%�X�GK@	���"YvE4&ֲ���0��c BS��BC��9����"4!�hL �@����$�i!�0�o �Ck���iBC���ܜZ\�����)A��Ҹ�my>a����;��w��Üm��&�UF��;'m���;��:1�F����6�,NS��y�s����HHEU[A%�,���8(��ܜn:���)� �� p��V��L�dk`(��3G�6X��f�:�rڤ
ڍm1�wV�s�)c��*�]�vYs.���r���t+Gj��W�n;IѺ`�b(6�UiV�ɮ�ܧ\�l6�c�����@t�N��N�Y{��t�[]4m�v#�M�39�VSU;�)`����n��vpZ��4�Nɖ�U�V���mj�iT��5Q�@F�i]���ui�k�	.YzR�-��KηI���P��[1N��mӸ�S�ڋ��zĎe^S���Qͷb��c�Rw����M$L��Syu�a�lꞐ��ш������KQ�"v�hg9�W#iYd��Gf�q�9x:���S��uW�,�82f6[&2V��<��,���qV6�涱%��ki���u�j�B@*�.�8���y��˶�+���K`���8��v��9B�g�(5�!J�Q�\�=<�iot�s��A;T���z����e��8w�d�W�vU�6�*C�f%�["���V{3jL����F���el�������rlO+q�H��yx�� ⢹����1g��O3a[��Kզ�ܬ��@N.0�u7��Dխ�Y��ۤY ��z-C��s�I�FK�5�U�`n����o]��=�v��tݍܙ8mKn�C(ӗV�s��y��j4@q�����9��irW;�u�9X%y���9m���Ɏ��K�4�t���/�,�4�k+�3�u�8��)���-5����0]iT�&�nZ9:slʯ�st���*:��ˇ���TXj�pq]�ԝ�:Pνjj7%�]��=,^�Z�\���UVIʻc�s�փ0DNה�U�,��͉���\�1��6��45���97vvV�c���q� ���ƶk������9����h����(�_�H��x��A�|UP>� i(PGA��D諠>O�7�ݽHi��9#Sʹ�R��lQ�v��)>��]P��0�W<��ݴ�n�*qe�HG'k�[`յ�g�����	�T�R9NSk��Ӯ�n+�d�;�����q���X��nƸ�Ms��"��ˋt���ꃮ��Uո���p�D��&X�1#�"F �v��dl�pQ�]PX��+����aҗT�T�aJU
�f(Q��r�JnSJ�j����.{O��m�֖�nc�X���ջ+I�"D^ĳL�k�x�<b�J��K~͵`���P�����V�ސcq��i4`��v�hol�����7�3����0P1'1����?j �9��5�{�A6V`�j`���&��\�����{�� 8�:9YWY�+>���0/wP㘀�W���x~�� {�������}��G5���g��0.{�ٻ<=��}r�<����R�Ak�1v/��Z�l�fڰ�ڰ�f�(��}��u�0LK��m$�4�ٳ1�Q^�U_U�Iݚ���1�qR��L����x��M ��٠��=��֬{���k[%�:*Q$�/wu 9&�=�*@I�?]�m�<zґ�<��4����=�b����v�hm�@��lѦ���ݸCm]pkY��$�n�����g�Qt�n�,����
&$�8�� �h�j�37k�yB�C7�j��Od�JQ�0JH�@?s�o�g���_y���V����BM�����LT�L�UX�uX�͵c�+��BP+�+,�r٠w���dx��!�dc���O����;���ٵa���uX�6`�K��Q	9��l�������H	ҋ�b���2�KXqq���m>��C�l�i���[�ibQ+h���&}���!�����@�rb �9����n�u0Y���eʑ�UX�vo�<�L���V����=�j�,0�[���ٟn� �9���V{�&oz�~���?fF���"dmA8����>J�ޚ��M��f��#�ҐVU3:��G�٠s��6\��j`���&�~㚀w$���H�5��翿^����\m�`�6zy	�[��@�w�˯NK���S�u�n�t��tt�A����?��؀�8� 9&�s���ŚeP*5Jj�l�fھ�I&�{����gؑ��M�{�@�}1�M%C %*�6��j �9�rL@{�T����ϫ�$8�C�%��M�{����m�(������G5�njh�	r�uUV=ݛ�"��7�/��չ$����$��>Ab�E�w��fkXw-��]&�t�kH`0���zy�W��#�����9�l�U:o#���=a#������c9RwJ��;ö�lU4�1-��Ʈp�.R������t
��k�"�T쇙�kj�k�[��][4�d;nt�
\h�eGj�-��v�b�Һ�⋇k;	rin0����`d[��uD��v�q�[m<�2=�8S������V�w���6㗗>�a�l���4���&9K*����U���Ɣ�&�#��ۚ�l��f�$�~a�����ʂe�c)7I�T�{�7��}��`k��?}������M�E�m��R)z��M rMC��sk@w$���w���X�I6�y.�f���x�:��@?s� sY[�y��m�������& s���P�>&U�y���)�0{W��k�a�/D�#�-���byu��K���i( ���v�4�;f�f�ח������y9#�IR9M�Y���=�jﾯWʪ����x&)���`��~��%�N�y�M����%�a{����������j �9���J���Kr�&��<�(Jٽ�4�ޚ���@;m�W� &�B&F�&�� �h�v� �h�͵`rP��rd�g���Bj])�e�ո��i�n^;���'��Yr]ֻjj�y��u �#m�r9$�o��u[^������~`owU�����U�)����sSE��wf��%	6}�֬{����:_B�D��ޒnUJsH
5SUS`f��nI;�{[��1<���Ȣ�b ~E��刺s>��v���rOs��T2 ��4?�į����=ݛBf��`s͙L\�5$�Hq�&�~�]4��Y|���nh����s�� C� l�m�j��u����r�o\{%��4�Tu�)[��[;��nT��h�?d���6�²!X�%�{�m9ı,K�s=*n%�bX��}dɇ5��YnX[u���Kı>���M��客j%�{�~�ӑ,K�����"n%�bX����O�*dK���5%�t[tk2�.�bn%�bX��{����bX�'���7ı,Ng{��r%�bX�������G؏�e��7r4�m�r=kZ�r%�g�D��~�7ı,O��~�ND�,KӾى��%�b� ��T`5Y��[ND�,K�u��ݎ�MkR�nk��bX�';���9ı,?�?��O���D�,K����m9ı,Og}�"n%�bX�>�=��ѓ-��I�^�v��s��|��y���tw]�:�Ob'�RMJt9�
�:������L��Zg�bn%�bX��ﵴ�Kı=��������,K�{��"X�%��t�A�o�P5M�)�d&Bd&Ay��[ND�,K��k��bX�';�p�r%�bX����M��O��%��ޙL^LSRL������~!2�b~���aq,K��{�ND�,K��ى��%�b^w��ӑ,S!1G��ٷ5*�A�R�U(�d&Bg��4�����p��	��	���a\Kı/;�kiȖ%�������uJ!Y	��	����D���˪�p��kFӑ,KĽ���7Ĳ%�Vwz��	���ީD+ı,Nw���Kı:`��h)�%FE"�����"�3��f��	��
�eC&܆X{�A6�*�����׶I̒t�!4[oN&t��9�:���jA!\=d(Y�v���Kp݌;#�+]�o9����*�J�U-Ѷ��+],�^���ͦތ�x�՚�v�2�ҲPb�ܽ\�6i�^�%ˇh��^XX�+f�[���d^ݜ�kv4��Aιj��`�M[z� �\���n]S4Y�k):9 :��OE��8y�n:[H�.㋺���f��)]mîB�N�S��oq���������"X�%�����Mı,K��l?��L�bX���ک��%����߀��8�n��U������,K�fzT�Kı/;�kiȖ%�bw=�ʛ�bX�%�{�m9�T�!h��Vȧ%U[��+!2�b_����r%�bX��g���X�%�y��[ND�,K�ٞ�7��#���O�PN`dx�NM�?bı/�}�Mı,K�����bX�%�s=*n%�`~	�>��|m8Bd&Bd.%=K8��53U0�%�bX��ﵴ�Kı/���Sq,K��}�ND�,K���Ĳ!2!|�e�i(mH�G2���Y�4oT=�Xv��8wRN����s���ݾn�v̆k&aLֵ���%�b{?~�7ı,Nw���Kı;=혛�bX�%������bX��vޮkZ�ɖ�Iu�"n%�bX���i�tN$Y	t� i@�M?��蜉br~��Mı,K��~�ӑ,K��{��&�X�%��{�&\��˭e�YnkFӑ,K����bn%�bX�����r%��DȞ�ߵ�Mı,K�~��iȖ%�bw;�	�J[�S-UTҘVBd&Bd'�f�ӑ,K��{��&�X�%���~�ND�,��������&�X�%������/��J��j>�~����{���{XD�Kİ�B?{�?M��,K����f&�X�%��u�]�"X�Bd.H��m��U*�I#R�"��d��#��־��۱�����6ݪ��s�z�2��r����a	��	�����\/�,K���bn%�bX�w]��r%�bX�������%�b}���2��IR�*��_�L��L��m��q,K����ӑ,Kľ�g����DȖ%���o��r%�bX�Jz%p*��7T���	���뾻ND�,K����7Ƌ�B�+VR$�F&�Z�Tw 6��41:(G�A�hVడ&'&p�����
�G mفM���vD�@5m<��8x��'z��|�!X���#FBH��D�bԍ@
i� �0D��gD�4sr1kD1��B"�XS����~�a�08���T�a�Z/9vB��a��-b�0b�@�P�Ika�I���"����S�i@z��@����@���);<�����_���$�5����Kı;;혛�bX�%��L2k%����r%�g�?{3����%�b{���m9ı,ON�f&�X�%����]�"X�%�|�sT��m�c��+!2!2��z�9ı,?,O~�Ȗ%�bw����9ı,N罬"n%�g�������۟��� �E���I`�:�p�/jz���e����.g���=�t� �KsWiȖ%�bv{�17ı,O����9ı,K��zT�Kı;����Kı/��8ܚ2�̦�u�q,K����Ӑ��r&D�/�ٟ�Mı,K����iȖ%�bz{�17ı,N�^�3�2[n�KsW5�]�"X�%�}��J��bX�';�z�9ı,OOk�q,K����ӑ,K��<�I��u��j\�5��7ı,Nw^��r%�bX��צ&�X�%��u�]�"X�
`uP�@�(E� ���@B�@ hD����aY	��	����?���IR�&��9ı,OO{f&�X�%��u�]�"X�%�}��J��bX�';���9ı,O�?{��ܙd�2���UI!!X�5�ɠ�xΔ��죗�&[\;=m�i&������{��7���{��r%�bX�������%�bs��ӑ,K����17ı,K�z`xɓY-�����r%�bX�������%�bs��ӑ,K����bn%�bX����OȆTȖ/�����hֲ[p���7ı,O����ND�,K��ى��%�bs��ӑ,K��=�a�G�2%�b}�~��2s2�Yn�Z�r%�bX��_�*n%�bX����Kı=������%�b^w��ӑ,K��w�tܚ2�̦�u�q,K��u�]�"X�%��{��&�X�%�y��[ND�,K�����Kı=��Pъmd�4��h\���v�9���u�Z�F�O;q"��39MhF�A�9����oi���(�\��dvځʼ�]��;8�x�=v�8��m�-"�Y*�hзG��xS�;�d"�ָq�T�x�.f5D�t��$�V��e`n2��D��qgJN�բ�P����+u��q��9G��[C�X�4�êx���ɴ�l���5�Wؤ����{��=�6��ڮ��v�����S�.�-�n�LӺ� �2�U���v]����w�{��7�����Mı,K���6��bX�%�����'"dK������K!2!p��dT�U[��+!1,K��}v��bX�%�﵉��%�bs��ӑ,Kľ�g�MĤ&Bd/�5�⩓H
$�R4���bX�׾�&�X�%��뾻ND����ș1 g�f~�9ı,O�����Bd&Bd-%<�L��k5�Mı,�2'�߿]�"X�%�{3����%�bs��ӑ,Kľ���7ı,O���<jd�Kp��k5v��bX�%�s=*n%�bX~��߿]��,KĿ��kq,K��u�]�"X�%�{o�,�eֵ��:���06�]�����v�Ѥ�z��=��������n���<v)���{��,Nw]��r%�bX����&�X�%��뾻�&D�,Og���%��	��3�Snd�2ꥹLm�;�Ȗ%�b^�{X���>I� ,D{G@��$6z�_�r%����v��bX�'���7ı,Nw]��r%�bX���N��F[�Y��ֵ�Mı,K��}v��bX�%�s=*n%�bX����Kı/�}�Mı,K��e���[f�KsW5�]�"X�~AD����*n%�bX�{^�v��bX�%�﵉��%�bs��ӑ,K��d=	Vȩ���548VBd&Bd.w]��r%�bX�׾�&�X�%��뾻ND�,K����7ı,{�����~������yꦍpxݛ����e��=<�[$�'%ɭ�m���L�]�"X�%�}{�bn%�bX����Kı/���Sq,K��9�7�	��	�����Z
���Z�kq,K��u�]�"X�%�����Mı,K���6��bX�%������%�b}����S5rۆ3Y���Kı;������%�bs;�fӑ,pЈH�@Q5�����Kı>���Kİ~��Ƶ�Md�p�]k��bX�'3��m9ı,N�{f&�X�%��뾻ND�,�Ȟ����&�X�%�������˭e�YeֳiȖ%�bv{^���bX��?{~�v�D�,K�������%�bs;�fӑ,K7��������ۋt7P�[X�wqi|�qv�ɰϜ���k���.B�i�f�q7ı,Nw]��r%�bX��{XD�Kı9��iȖ%�bvg�q7ı,O{�.g�R�5�[���j�9ı,N罬"n%�bX����Kı;3����bX�';���9ı,OC���n�Y�֥���7ı,Nw]��r%�bX���\Mı,K��}v��bX�'s��7ı,Ot�r�E�I52k�3WiȖ%�bvg�q7ı,Nw]��r%�bX��{XD�K���P>S��� TSA���"Q`�[�������9�L��\JxD�@�US�s
�LK��{�m9ı,N罬"n%�bX����Kı;3޸��d&Bd.�K{��ǴSRT��T�P8���џ	\Z�-2�<��7\��$m�a�Y���̹�'�,K��~��"n%�bX����Kı;3޸�'"dK����ͧ"X�%�����kSXe0�]k��bX�';���9ı,N���&�X�%�����r%�bX��{XD�H/��D�~�K ��l	��b�
��ʄ
B���pI�N罬"n%�bX����Kı;�oN���2�̦�����Kı9���ND�,K��k��bX�';���9ı,N���*�L��L��Y�������ә��\�bX�'s��7ı,Nw]��r%�bX���\Mı,K�ﹴ�Kı7�|G�p�*X���q��v�ʷl�[��[�Z+5��˅{l�����t��1)*����גk���v��;�7Q�H�.�m75g�4�m1�LvB+Km�͓����r��=��s���;iC��B닫6p;�-��2<�nP-lすi��ܙ^��*���l�y�Z���+\)g-�q��t�+�����,ɫ:Sn���.�TT������e�RS ���>�w��iM���HX��bt"V�n9�9�͵��M^�J3uȓ�R4h�:��j�[��'bX�%�ϵ�]�"X�%�ٞ���Kı9�w�iȖ%�bw=�aq,K��ݾ�]h���.�I����Kı;3޸��bX�'3��6��bX�'s��7ı,N}���9�TȖB�S�a)� ɧU48VBd&Bq>���m9ı,O���7����>���9ı,N������%�b}�zX��ɬ���]k6��bY�E���aq,K������Kı>�ץMı,K��}�ND�,K��g�kZ��)��XD�Kı9����Kı>�ץMı,K���[ND�,K�﵄Mı,K�"�~�a�>��)�&vnʸ��7c4R�s��=;u�K�c�yTu�K��������׻�����ow}u�T�Kı/>ﵴ�Kı>��XD�Kı9����Kı�����Ӣ�.�|͏w��oq������Ӑ��F	RF""�
��"r%�����Mı,K�뾻ND�,K��²!2!fVk�52���7USu�m9ı,O���7ı,N}���9��2&D﮿J��bX�%�����"X�%��y����3Y�ank��bX�'>�}v��bX�'f{�q,Kļ���ӑ,K��̉s��7ı,O�w�9sE�0��u���r%�bX�L��&�X�%�y�}��"X�%���6��Kı9����Kı? =�~��n��mi׭`��f���/'X��Y�tt�<�	�Eqll�����19ı,K�}�[ND�,K��m���%�bs�w�a�}"X�'�uÅd&Bd&Bͮ����T�T굴�Kı>��lMı,K�k��ND�,K������%�b^}�kiȖ%�b�;��ѭh��f���Kı9����Kı;ۯJ��c�� �EJk�SF�!��_"0\���P]�r��ؗ5���r%�bX���6��Kı;�����[�e�Ym֮ӑ,K?"02'�w�T�Kı/���m9ı,O���q,K����ӑ,K=��~�����rU>fǻ��7�����}�ND�,K����a�,K������Kı;ۯJ��c���r��Q~q�ȲLCțB��8{4rx������,3JwQ���O}he6:�[�]]k6��bX�'��k��bX�'>�}v��bX�'{u�Sq,K��}�fӑ,K��<�xՖ���j�\�aq,K����Ӑ�"�"dK޺�*n%�bX�g}�6��bX�'��k���\��,N��윹��jd�9����Kı=�Ҧ�X�%����ͧ"X�%��{��&�X�%�ϵ�]�"X�%���L+	OX�M:��²!2!~��fӑ,K��=�aq,K����ӑ,KB�	�.�J0�V��&-�@2IM 鷑3��J��bX�'s���4e�����ͧ"X�%��{��&�X�%�ϵ�]�"X�%���zT�Kı9�wٴ�Kı:Oj�	 �eӕ����f�c�`�[g�ZPf�(:ݔ��\w:�ngL��}�X�%�ϵ�]�"X�%���z�n%�bX�ϻ��$�&D�,Og�k	
�L��L���(%O�l�m�cn��r%�bX³�_�\ND�,K��fӑ,K��w��&�X�%����w���I	�����өn�Uk�kWq,K��;�ٴ�Kı;������?�ș��~�ӑ,K!2����	��3/Jr薆�D���Zͧ"X�~���aq,KĿwߵ��Kı>��\Mı,�&D�����9ı,O���~5d��f�T��k��bX�%������bX�'�;뉸�%�bs��ӑ,K��;�aq,KĈ| v >���G��L	�`O>i�N s틂ƈL��bxx(�L���0��C�!R6"D;�c�K�Ǒy��)I�����N�&��||�I��k��>"���pO�#��n`��	�(O����@�P0t��v����H�R����@�pA���)�M�D6	f�#�t�U�~�������: l�h�������d�۠�Y^���V9d��n��N��s[5 ��VF%ٖq��Q��V�{B�q�v�;X�	ݚ�H�q
v�3Hv53��b-�nr�us�ZL;�ml9�����a˶�X��ݫ�V�*�2��Tjj�Ѷ��ur�g�a'��Ҽ�yN�Wb�����*�:6�6Wn������!�db�u���J��U������n�����gg�d�M��r��0۷a�ηg)h��gm����Sq�1UJ��+1E��ҭ��j���� R�q���i����m&���ctH�	ic�5UKj���ѓ+�"Ý��b)bL��Uqq�Q��s�ru�B�S.,&��#��cp�C�'j�T�]U�vvVtDs��8��,�:�BM�@ճ�Y9�`KRa3��c��	�������m�MU�
�p[I��q�]�1�U�em\�����s��y��^�9�n*�.��k�@b��U[*۲�2� ��)�����Z�;�K��Ue��"�<[,���񋎥R�������q�ַԝ�z%������+�*��)�l����r)���65л
D�u�]Th�:�e�����@�ƶ�lJ�]/�k��M������3�N-��[��[[i������&��.�k�.7'n��3��vXNcI٥��Cj�<㶞�۪�%��  ��.!mXq��9˪��6��pw<$[<p����)5O.�o\J��Eg>��.wK⧌��15��ƺEM΋���*���=��;f���,�r�fy���L�͖a�ͳ�Vٳ 5�Q&�#lܮ�ef�M.(�$���N�����K%nR�] e����vk)(����;N���{up\ 
�I��A���ژC&-��ݻae3D��Q��gtk�v���h�#98�Id��M!�lrn5��R�Ú�U�asv���������iA�xT�	��N�� �(tt�#�E��AT�DJ*?z(��A�U���1#������풣��_U��ǂI,p�lbc�F�FtRg\ݞY�3�8Wۦ �k��;m�\dI��%wn��`6{:12��s9�K����ݍAY�h�e�=�^�v�y�S:��P�]<2�)7&x�&՚��,���7>��kV��7C�a�_:q�6T�3�&�Mf�2d���7.LV��OD��=Ϥ�n�v��'N7{��w=���6m&���ַg%�c�G��_/j]�t%�ӡv[$\N�ὺΞ2������oq��;뉸�%�bs>�iȖ%�b}������ȍ�&�X�%�kj�Bd&Bd-%���!�T*����n%�bX�ϻ��r%�bX�g}�"n%�bX��w��r%�bX�L��&�~E2�D�=��r?�C4\3	sW5�ND�,K����&�X�%�y�}��"X�ș���17ı,O����ND�,K�u�Y�j���nI�Y�"n%�bX��w��r%�bX�N��q,K��}�fӑ,KH��u���aq,K���~�L3�K�e�X[�kiȖ%�b};�LMı,K�?k���O�X�%����aq,Kļ���ӑ,K���w�;��~���μ��\m\ld����*p�@��d�:]�u��r-rv���W��AZmѭkXf�jb}ı,N�fӑ,K��;�aq,Kļ������DȖ%���~���bX�'�����u2���f�]k6��bX�'��k���>N&Ў�n%��kܻND�,K�����Kı9�wٴ�O�*dK��~4[kZ��as5�Mı,K��~�ӑ,K��w^���bX�'3��6��bX�'��k�Bd&Bd/�f������ʔɚ��Ȗ%�b};�LMı,K��}�ND�,K�﵄Mı,�"gٽW�	��	���%6�1P��kZ���bX�'3��6��bX�������XD�%�bX�������bX�'Ӻ���Kı?+�����/g��I�Ք��z����=�5�3��n����FwWO��p}��ssہ�~;ı,Og��aq,Kļ���ӑ,K��w^��9"X�'���_�L��L��Z�>�t��nBJ�aq,Kļ���ӑ,K��w^���bX�'3��6��bX�'��k���S"X�{��I�s-�շ-ִm9ı,N�k���Kı9�wٴ�K��+�'G`�D�'3�k��bX�'��p�r%�w������si��a���{��'�2'��fӑ,K��{�����%�bs���ӑ,K��w^��!2!2ٗ�K�Zn��ӗU6��bX�%�}�7ı,N}�p�r%�bX�Ok�q,K��}�fӑ,K������S2n��2e+��64<�y�H�5�,5�NY-�΍4Z�{RzIÝ/��j橗.kDMı,K�w�6��bX�'�����Kı9�wٴ�Kı/{�h���%�b}Ӿ��Ѭ��f�˭ND�,K��zbn�c�2%��w߳iȖ%�b_{��D�Kı9�}�iȖ%�b}0��	OX�UUUQ0���L��_����r%�bX����D�K�2&D�wߵ��Kı;?k���Kı;����e2�[����r%�bX����D�Kı9�}�iȖ%�b}=�LMı,���8V�m�K�sٴ�Kı;�B�Y�L2�nHkY�7ı,N}�p�r%�bX�Ok�q,K��}�fӑ,KĽﵢ&�X�%�y�d�̄/�CD�V�v���/';���^"d���hy����v�2�x5]�������D�{^���bX�'3��6��bX�%�}�7ı,N}�p�r%�b�~���0V����>ﷸ��{�Ng��m9�r&D�/��Z"n%�bX�w߸m9ı,O��鉸������Y�}$�%�RڤN]T�/�'ı/��Z"n%�bX�����Kı>�ץMı,K��}�ND�,K���D���\�2��h���%�bs���ӑ,K���^�7ı,Ng��m9İ?+2&{ߵ�&�X�%�㿿NhֳL.[5�Iu�iȖ%�b}�J��bX�'3��6��bX�%�}�7ı,N}�p�r%�bX� �AX�I=&Me�n�x��J��GP��lt<�e��1�7Wg\9�J�pqv�F��g�����9��i�O:�`�	��p�,q�����vy�:�ka���Γ�s��s�j4ZR..�\������V�gu�3��Z��Zn�S�!���n��{Td�8���S��ܚkc���v����e���ҝsSt�{m�r\C�!H�Z{j��w{�y�r�r@#Kf�u�X�5�.���e:^���c/JU�bh[l%:b�USUC��	��	��No��r%�bX����D�Kı/>ﵴ�Kı>�ץMı,K��쾖S!��!nj�iȖ%�b^���q,Kļ���ӑ,K���^�7ı,Ng��m9�2�E2k����.P努j�
�L�ı/���m9ı,O�u�Sq,K��}�fӑ,KĽﵢ&�X�%�y���2kYf�m�٭h�r%�bX�z�Ҧ�X�%����ͧ"X��2&g}�����2&eO��6�}Q��=��/��Xmmr�ƛ/�왕2&eNk�{6�}S"fTș���j��fTș�>����}�L��S"vf�.&�fTș�?
����|ܴ������Q8v�ל���ݨ��-�Ɂ��t�(|�lP��iKm�?^����;��L����Ѫ���S"fT������dLʙ�5�p?�5��2��߿{����r��{ǿ���Ǫ�9��M�̩�3*}�}���g� m�(A@�T+b+���P�Nr�D��}.&�fTș�9�����2�D����U72�D̩�N�ߺ�{q�%w�����;ܧ����ޗq3*dLʜ�}��}�L���MD���Z5Sq3*dLʟw߾6�}S#�{�����`ɏ��ئ����{�*dLʜ�}��}�L��S"f{�Ѫ���S"fT������dLʙ�+G0��2�I
eݖhƤSRo&�Wi��2&eL���kF�n&eL��S�w�O���3*dOLץ��Lʙ2�>�}v�}S"fTș�}	f�k�f�v����ݸ��[��:��|��y�I�n5��nZ�#���<���̩�3*s���i��2&eL�������S"fT��i��2&eL���a�M�̩�.T�w���5�f�m�٭h�}�L��S"{W�ɉ���2&eN}���9�L��S �{�f�q3*dLʜ����}�L��S"fwڒj��k��"�}�or��{��~�������Tș�2g}�i72��<�B�N	C�t+�UC����D�bwu=��|m>��D̩�8�����\)!L�_a���(c��A&�s5��}�L��S ��fi72�D̩ϻ�Tș�2'r�fbn&eL��S���ͧ�Tș�2-s�4Lu�j�.e���Lʙ2�>�6�}S"fTȝ��q3*dLʜ���m>��D̩�o}�4���S"fT�{���Ӯ��5����kWHF=�s��v�͖�95��m��N�v[��i�lA��]���2�D��l����S"fT��i��2&eL�{홤�Lʙ2�>�6�}S"fTȝ�f{-�,��Ԓ浚֋����2&eNk��6�}J�r&D�o}q5ı,N}�p�r�bX�L쩨��O���Lʙ����jI*@R���/�p��2�H��l�&�fP��}�p�-���l�������~I..���4ěr9�R_��7��p�-����˻m�ϻ��-�l@c"	S�D5���ݶ�����3Z��$�"I��$�+��RI~|��$�[�x�$��v��ߒK��1-4<Ǆ��4>t78��8���9��	��zɲό��-�+�k!䈘܏RbԒ_�;_��%��Z�m��ٿ����m�OZv�o8ޑ�$_��"nG��Iu�W�RIs�����\�ũ$�>Z�~I.��ۓ��'8ԏ���;g��$�e�D���k��$��+F���s���#������|�������t�l���}�j���P���Ndr��^���^nI�����9���$��bEP��,�_K��!�����fj�uڳQ��cv�����pm��WU44=]-��=[V�M��H��˹�Ḱ�*����`�$����X�F�'V|@���6<]m��;Q��x�3����s����F�dy��|�u���	.�N�q���7��>��aɠ.�C�n����L�^� 6yڷn�ˋ��#<��ɬ�d�tNɒGg�`���{��wpu��Z%07n��L�M�MMAp�l�>���h�-W)<��7\��+;$ykcӉ��?y�7�s���+��%�|�lz�ų�J� �J�Uz��qR�Ih_I���UU$���x�H�$�)&h�����svl�Qٹ����޵`~y��*��Y��W��h_I��� 9]�@�;q��Z�@	r= �;��噽�~:{�����6����7n����4C1یs ���S���{��f�o=f�ꡎZb�m���?>�\����/P��鹵$��k�Z7$���]���F(�`���	��`��w����ٹ$�o��9��������J#&��$v����ۚ��D$�f������36CF5$Ӗ
\Ӛ��KЦw��	? =�`������`U�2i�LdjE4s�s@��)�~\��ۚ���DwwD��2��*t�D˞6�>nx!^q��=s댗Y��UnU.���{}���x�H�$�)&p���h�-z�ڦ�s��@���D�䈘܏4_I������=�`�}���}���d �7#���M �;f͙ȝ-:v҉s\ݟ
kBI>7�>��`�B#��>��;a�㤳O�1 B0Hb|^n �Ũ�p4�b$�^;ںM�A��,�p�T�M$�["V؍RC��V,T�}G�!%
T�����4b��LхM=�`d�R(�Z-Ӻ�+�/���Vץp�BBk�$ɤ~�P��,��HPe	�*`�|:E� �~ڣ��ڏDz4��CCO| |&��D>O*'��lh |�P\T8���5�M�9}�f���t���� ��H�X܎)�w�ۚ�����C��ﯔ�;o����И�ݤ�P��G/P� ?������t��ְ�/ >S�t:-e�� qgz��byt�#2F2b7]�g5U`~f̀f溰?}�k�/B��{������Lyō8�z�ڦ��qR���syAeL�eb`�#R)�s�����V��������M��ϱ �_'�D�M�e��
I�ռ�{�6���âPh:�~��@�\���'}��5l�UL�5U(�T��ń����y����X�s]��a�A\ҢJ�P�z�Sc�-��h��=i�e�w�?�	��;SU۞�S�SP�Q�� __)��@�_j�8�k�;�)nH%��'7*iՀ}���!$��ɞ��5��6�ڦ�f}�bGm�6B9�Ȅƣ��s��h]���/���9�����tТ2a��NE����|���M�;w4�����h���ƞ�n �@{�T���-��1�ڥX(@"�� �ڞ/&sI�j��4��K�	�+�n8n0�Nx��Gr��s�5��T��eY����v���)Z��0�[��Bhvq�W���V�Hk&���7l6���27i5��}E~��%j1�M �v�i�Iu�N��<�W�r��ѝ��n�c@mZ���:�ڇ
�j����j�2\.�l\���R��S�ʕ�X�K��\�K�.ݻ���ܿc� 7.���<���fI1�wW^{&��lyf�f�(:ݔ��m�܃Ƙ&�Ԋt�]��}�@������M ����x�H�$Ѕ7��=|� �@z��@{��$$D�$xE"�?.v� ��S@��������;pm�q� JE�C��>�J��M���@�_j�?.v��)nH%��'7#�h�;^��Z��b q��n�Z�3L+KA���[�3��z�r��_/j]�tk��B�r�2HG0�����������6l75�(����ٽj��ڧ��e��$.h��]�9~�~P��X"}�V������ =1�@�	�� �x���@;{T�?s�s@�_j�?.v��^	ev������=�*@zc����r����oĉM��4�����k���V�mtB��Y�e�P�K*&\�Lv�.6]��j�@�����kK��޵��Ex���4��(�����E�qv��oj��� =1�@yӔfak4��ܪ� ��u}��������y�<͛�ؑPx��A/��8��S@����w�s�G�*% 
R�����\��Ѝr���ܒs��9�5�ds Q"?����s����?b q���� :㬁f	B,Rbr-���@;{T�?v�h��Z�����k���H��W6�P�>�{;���;;�&�6r��(�`�)B�'�q8� __)�s�����V��rנ^Y�X݃�8�܊h}�j�&Ϻw�������W�6}�����H�$т�f��;�~\���"��M�~��9���5LQ%1I�C�f*�����4�ڴ��������s]���Q3#�-����� �@zd����- ��1�~I2��d���G��NQ�n}��c��M��`:�k#�r�pLu�����9wso|~�߭�Z�s�^�9��Ml�&LQ#27���ՠuu�@9z���-�d0��n�:����6l75՞I��{���;�s��U4�2<1��@;{T�>�kK��k��I��t�wR%����pq��9�)�{>Ͼ秼���߳rI���$��B=
-B �"�.{T��kR��a��]��G�Z�!%�H�V��8Ҁd%�z�L�^�׷V�Zf��k�cFT&�-�\c\Ac�7�@nu��lQ��:Xq;*�v62Ss*��<<j�ݨփp��Q�a��	��j��:Ѯ���C�say���͌Q��[���w�r.֊�7e�\ش�nJٮ�r��R������c���q��R��������7|k�@8F.���E��[�;�t)�f��.�<���<�Q��P�h��{���Q';����P����~��9o��1D���d���پIBl7�uX���ݭ/�JE�K�l[�(R(�zۖ���1 �� �1 � �mm�n��E�ɎM�v���h\��n[4w�[&I�H�9��e4���&�;�K@twy�f`c��I6���-��br8mA�)/U*v���8���#!)1'��� r��vIh&�鐲��u�f�������'}�k[��H?9�|��{V��YM����bG}�X�"�n(��;��-��h\���l���_'�D��$��/6��>ǹnfՇBP�+��wt���A)�ɑ�h\���l�9�j�/,������3~X4��4�|F�8מ�ۜ��D�ն8������%t�5�za��Q��%"�G���h�h�R��]��YNܐK�$N,m�&��n��@u���#sP�\��$Ɋ$dx�"�/,����^�ϾX	��X���T�R$D ��.�F�mX����ڝcD"��&$�qrנ��@���v	�u�`s�.I\ԡ74��73j�興̮��ή,�ۯ�o�����7���p[=iw�@q�c�4�Dq�|�]���^��Y{'5f�n(��9�j�/,����^�^�� ����y$"I�IŠ^YM��� ��8�[� ����"	LNL�E�uw�z{�4qڴ�j�/3�طP�Q����hN_{ٹ'��z�H9�E6�<���|�سǮH%���<m�&���1;$�_I�75�.�V�S�&��Y�����n�����aj�'&u���[7��p�j�7O)O�o����X�ͫ �ͮQ
?0>��1�)�f4B,Rbn- �;f�^�� ��f�x�Z�DV��Q�H������1;$��&�#�S�) �6�M����ڴ��h�l���_'�E�F�@'�;$��&���_I�Y�}[U�.��ޔ���Y�1��"0��$�k�pZ�Ї���O���T�!J�}���IFb� �", ��Ԍ ��ʎ.��ژ1�8��S�� @��������j&&����g����s�x���K(�L4����Ch��l�ɯߓ����y<�D�D(�  ���!�$#��V�Dp��"lF#!��H1�h%��¹~���P��h��W!�����?!�F�n~?�U���	����DB� 	')Z��B��*��@D�M� �$��E�u��n�m��h�9��0�NT���!�Oj�!�jUBR=5Ul��r ��QIq�5��bY��d�E����S<���3;5,�mA���wk�ⴏHC;"�Ȱ'D�=�����īe61���-�3���n��y,�..㍃��{R-g�0����;|����=��ts����ͮ@�p�R��ԕK�q!:Mr��d��bA��]�:��;��Y5A�[Nԝ���$z۱��#���8�e�hԪ��2�]q�T��\�-]���S���݈m� ��s�+�nɖ�8�C�)�~�Ɇ3@�,�J�f�7*�3��Y�m�^��)��3T�2��r�Nvt:��rT�gum�����/n�ڳ��r�5�m�mu�a�5�ۙ7S��˛r)VMH�,l�]BA�<Z783K�:*��8��.vڪ�@�K,�;��8��ۊq���M�N׮]%\y���ז�ۮ\Ug��Z���K!�+T��mW����+5y��6�K�:�t�:��.XS�F�m��:�RΓq*t��c6�n�llm��rM��fc���*]��G��TD�A��ݣi�
�C�ez0$�p�UKt�>�x0r�슪��ú�����F��繭����b��[p%^K,iX��J�$�������p9v�	ܝ�m	��t&�kVݧJ�]mE�&�pJ�����n��~��}�~��op�$i�:۷U
�өRƭR���eh�1����s[!�Y�!NjL��u�N֬�db����u�sv֍ͩ��������_��}r�F���*iz!-uz;rk���P�z�a6-�u6PlF=2�B.8"m)�3�x©S����MӴ��J�P*�Ies[G5��1�B�&AWS;q�0������iJ¡��J1�f��V䍅x#nي\���L��5j�{`D�rp@5ܤ��U�:r�IȽ�6sH���� �Ȉ�@��Q�
?l >Q*��_+�)���� |>K���~���w�%�n��M ���	�V19�*i��Z�]���^�&0��8mn(�^Sv��΀Ҩ���q���q�\�WN�z�rm�k�	{ƦM;�����d9��ַg�
���c��:-I2��Oa'\ٺ�Q0�g�Ӿ�n;���Q6�<�ԡ u�N"��Ա��^Ax+s�G��������mc�n�%U�=���=�u�����	�m����m�<Vvgs��o.1F;%�Y6Y��ns^
{I�j�Ͷ�?��@�����%�'S�feڬj ���&�w��@��@�v� �-�����$\Y��&D}$#�iɠ;�bvIh	2K@��	�U�$ɑ�ɏR=�ڴ]�@/{f�U��\��#!)17�&Ih75.I�	�%�$eߝ���j�ӭc*�;g��u�6&8�K-��M�A�zX��獱�c=d�8��G����& 'd���$�[�ʶD�Nl�rh[^���}~��,�%hC���"L�������A7?��Ӛ�36��BQ��r�<���i<X'��?yh�V�w��@;�٠���Dj2	79#��	Buw; �ޫ �ͫO���������ɂR2H���hnjvIhL�������̲��7�:8����{q�l9�oi�`챥�q�P�h��̙�B8񶜚�����v���	/���;;�˷UJ�h2c�G&�x�[���Ďy��@=oU���l�$��3��b�YMt�K�v�;��73jΈ���!	$�%
�__�`w���>`�b�]Ji�Y{�h75�nbvIh<r����Dؘ6�G&��w����B�	q]����ls6�͇�Nplg���<n�{f�ү8�]�<�ny��u��Y�Q��[�7��U��!�����ܘ�:9��& 
�&Yu��8�n<rE�uvנ��@ⶽ�v� �s��(�L�#q�뚀�bvIh���up+kQ�B8񶜚U��z�����rLE|cI]�D7�]ﵹ'{��&O�J!���@�v� ��{�4�Z�[Cbf�$J}>�1û^zț����0��i'��޺:X�]s��<[!"F܏@9{f�~�l�:�k�?.�� ����D�ŋ�94�f��Qٯ;������ۛV���`ؘ6�G&���^��w��ВI�;z��ޫ��4L�5-:�w�{y��[sG5 y���s49�ZD�8�n7$�@?r٠�}��>�wٹ'/{�ܒ����������"K	��/�&�b��j�\ې���)����7H�'�$֦I��N���].+[�Xy�n+bۂ�"lްb��j�Nw=xϮ�p�ܚ�]�v^BL=n��E۵f}�u�:�a7=q+��I�d9����_o���ںѶ0�e�Slmuv���K!�Ì�"�Ì��j�f�7b���]av5CK�;Z���.��ԣ�&������{�w�����i��p��ˎ�Ӝ4v��le�x�w����JwW���Ǳ�݁�sK�x��禁��נ^;V�~�@�*I�$#�iɠqs�����yh;�M ���#��[$�>�Vnn�?<���nj ��@�j�n_���`b$��Z��� ��V�7jâ�	�Ws��OW	G�5"rh�l�ݶh�ՠ�l�?e���Ē1��5�� �h�Ls���g'n�u���&�9�J�k�A��h�/377P�����1 ssP�����jD�⑤�
I4ˮbt���O�� �sPrj�I���ő)�$��A����h���=��%W}�q[��n	�F2Qw�����<������ �����"2HG6ӓ@��@脗ӻ��;z��fՁ��S�r�%��^���P��W)봯<u<�qt�Iv�tNî^���U]x�3�)�m�?��`nmX�ͮJ?0ם��BJ>��|�Ĵ��#nG������W-z��נ�b�Q(�bƔ�k7$��}��>���s�E���� ����GIA�Q����>5���:�����3��<���su�$�����5类�O�@����5�D�����{^��Ɉ��@u�1 w]X�&ay[Z,��(Oi�,Z�>�eC�lt��D��.�]��W�� ㉋"SI9���]������������z��6Ҍd�)27�w��}����y�^�zWmzŜ÷&Dd��<lnM�Ɉ\sܘ�9�t�ykwuT:n�(n�l:J���`k����kr'�� ���2��$!�G���7����9���,�n�.��� �1 y���& =m�@{ﻖ���1'�4��8����-K�����۴u�δ��N;9Aޔg0f6����e��nx����& =m�@;rb �S:���H�rhVנ~M�@;rb �sP�!f��^V���^�n�����& 75�$����%1ē��9���^�~�ڰ>{�6	(�O����x	�H��U3S`�6�P�'���<��ܓ���nI�w��p�`���f,�u����=g�A�i��tҸ1Y��u�A[YD-֘F�P�9�lj�.6����Ƨ,n2t���H�Cn^�st M�,���C0(�G,�j���L��D�/.��R]����˪̘a�7G[����8n�v�!��M�^؄�4�u�n�΄�ò�.,�e�ܛ=r�l=���6���Z������9.���(c�MsE�d%��A�?�y�}o����W�9:�{	c+�G������:]�۱�6%�]�������f���\����^���?.v���������;|6�92|�Q�z��נuvנ��4+k�֗䘔&,��nG�;rb �sPrL@zۘ�Xi��
���������1�t��ez��U�y�����l�`H�r :䘀��1 tsP���ڹ�x����B��[[P���x��t)�%3my$��V9'b��:s@<CO�[��y�;@�_��T���m�TҢj���g5��D$�>P��K!$�(��7�*���t��f��a�_ �id�)"�[�urנ~]�z+�Z�qhL��1��k7P�L@zۘ�nl����
��&O�J!�M��˽�@�e���9o���mzy�h�Li��ح�����Z7=�k��g[;)�	y1��wC	FO��LY��܏@�l��~�mX=ݞP�%���w��7���4���/t@nj�I�[s3�h�K��I�#�rh\��N^�ٹ�
�h�$�.Ԅ%B�@A�FD��x>N�|����nF;Z�Ւ�֔�@G	4<s�P0��	 � �)����� RtŁ�$I��4?#�R(l�Ӽ�%ڦ��f$��;��]�p,D!) j`6�P��"H��+e�+H������I��MR"G�8�c��x�L���Q�T��xČO�a$VLpD0�$�@:+�D�ay�H0�(G^;���Z��H�!��ia$�s	�b�X<��8���(A:<�N���@�4�C��hm���A9 |��G�%|ip4#�0?���L\SJ{��w��Qyd����4+�$"21Ȓx�r=��k�>��v�3jÒ���wM��{�e˘��L�����h�v������k�9�ܳ�h�,��n|�ܢ�ޢDۂ�}��^tJÑub�gV�\Kj�ꛪ�`�6�ń��l�B����:w����o_2�1U)s32��w�b���Lr����U����5�2#�C�)��o����V�~�l�:�k���b@�	�2I�J���`�6�G��l?DB��	5`�Tk�& ���4#���?�w��=�i��
��SN�?75 �������<��+.��43��X�a�.�z��wWlt���f`�Zכ�����O��
y��g��m�>ݛ��ٰ>��~Q�n�X=�leIRMSnS�5S`~y�7�(��fs�Z�}4�Z�R�mjSQ93+��Lr����w�b���s��&�Y�JH�=��\��@����?.��������]DȌ�m���W-z��נr�ՠ�6��*�D$$ҞӃ�M�j�/�vZ�xSh�ӳ�.^J�-<ۭ�qsqS���])���㵣N�]t�����͕����V�	��y��,Y����=xmm�p��P�c�u��:h�6%�w���N1�hK�a�b��m-[C�T�x����'ڛjuΉK�9gA�N뫞lE��v<9#Q���ke�V٩�������,��zƥz���b����*�B(���gښ֮LɆ�p[��WbK�z��ve*XG���M�%�&&��"2$D<��/�����9��?fm%���� ����	N�+������Lr����w�b����Q���6�\AB9*i�I�P�L@zۘ��Z�(���d�G�4��:�k�?.����� ��٠~���H�'�����s1�@nj�I��W{Ww�8G�n݉7;��]Yٹ��.�+�1�-�@�>]Ҍj.ӥ΂�!��4����c��<������ 	\��:���7UN�?fm]��!@�  ��.�� �@�7s�ܓ����Wڴ��]u"2Li��rh�L@zۘ��Z �sP�[�"2$D<i���w����h�ͫ۳`y$��:	N�&��s;��쟭 y��}& =m�@~�����~N�=ߠQ����[��s��=]������m\��qibV�6�6���ra�����������1��x����L#��&���^��w�1�@nj���PC+�wW)�N���f́�9��CJW��(ʚ�@������ܓ��]��UƖ�1���c���ՠ������9h�J�^a{�u������ͫВ����{����V����,p11cb�l��#4Ocq���s�iI�t���ۊ*�6oc�BF�#��m���-}�@��j�-}�@9�٠v�R�ّ�"8�@��j�$�- ssPc��=*J�*�����n�6�c��9��	1�@y�V��p@�.S�dL�- �{f�{��]�9�����P�JAp���E>]����rN��I-��d��mɠZ�V���}�ܳ�_��N��6�����k�S�6��Bs��1�u�E����g�Ӳ����<�;ҍ曕���MD��8�_��w�@��� �����=�|����Ūb�'#x�ݴ��75&9h<��ꯪ���xB�,�R%$Z�}4_j�٘�+����?yh8vTL��*\�̹���
!(}����{���ڴ��9�����#�!��H<��d��9��	2K@t�����;��Aۖ�f�v�q�e]Ha�v�ū��l**{<UUZz�yi�aucrޣ��2sNyXֶ-�n�[�]�x��[*���{q�j�V黩����g8ٓ��u�!x�W�;�K��m��#\��q�H��QΡc2��Ɇ�:�H���F#syѐ�rO@lX�P�8�s��x��٨F3�S�=�����i�.�	�a�R���l_��அG|��e��4MI�R�Ԇ��������7)�[g���tOF%�:O],O.��(�ݍ�"��Q��s���h;�4]�@����?�7�M��P�NJ�v��h�V���ՠZ�Zz�	X���pm�4]�@��j�-v� �{f��p�lq�O��h���%�njL����Ye���M����k�h;�4]�@����P�-��Q���D�2)��(Z#���0�ű�)������(-�\s�Ļ��=a4(��%"Q���M�j�?uڴ]�@�ñ�Y2(��6�NM�{��]�PNE���N��+�S��P6 �^g��ܓ����s��@�:�59>�Ƒ�n-�$��& njL���p� �I�1
E�Umz����j�?uڴ��bH�O�a�8�z��@I�Z�$��& ?�O��<�eܮ�K�4��s�zq˻Y��vJɹ��EzR��sۂ�5�͕k�������y%�%�1 ssP�x���I?��E�~�h[^�s��@�ڴs��!j��M���������O��ksáb�ሀ(�V�(I"槹����gƭD̊1(�z����j�?uڴ
��@�ñ�Y2"i��rh䖀��-.I�����}U�ߜ���;`�n=z�;*�מ�\�u!�3�֓���:K��B�:��LƆ��tg�c���~�h	rL@���%�'�C	e��' ꝁ�wf�% fmX�V���ՠ�E�|C��& njL���W�|�+@K�b�.�S�q�m94]�@��jܓ���nL<<��
�Q	
EbR���)���O-DC�h��c��I?��E�~�h[^�s��@�ڴ�z���85�@X2�[=�I`�=�Qc���▎�{��p�ӽ�!&1HZW#������ ��$�-�Z �ĩFf�)�N���ٛW�BI��{����r�*���ƫjd�m����%�;��.I��&�<ܱ^UE1H�2U9�v�(O3o��wM�~�@�ڴ�;L4i1}��qh[^���r����� �>uh�UU��UU��UE�*���UTW�EUQ_���UU��UU��@C�H"1Q��@
�1@� �"(��
�1b(X"�1A��@"(b( b(������"� �U����DD I��UTW��UTW�UQ_�UTV����EUQ_�UE�UU�qUTW�UQ_�UE�UU�UU���d�Mf��rl1f�A@��̟\��| � D   �(     U   @    Cp��AH�R� �P�
��I P��P��%P���D*�U)D ABIB@	H@�     L  P �� a`�����ϫ���u��k����� 9Ҭ[͔���;��}������D
<��ܷ��^-��  �ɞ��>�筷� �v�]��r/N!��q�]� �|��ů<v^ڸ��<�}�_1� ��@ �	   @wЯ�o'�o>������zq��. V;�-͸��͝@ �� : �8@��Z�x�  ��M@1������׶^}����r������)����;���ͪ�ۼ{� =�(  �@ ,0 �}_aͽj����;��oo3W��@oW�����v�t�۷����:}^���篭����o�� ���7��ܻg�|*�<�qϼCO\��[�w#�� }|��W���z^=�^�k� |�     @@ ���[ź;s}3ɧ��ܓ�@���m����׶\Y�H<l�� QѦ�J�LE4  DR�>�:R� `�M.�Ac4�A��1�3�� щ�@��  �   �
T Oe)�" � h�M4A�P�تh" D�������w 
��Jr}�NC� ��.���=� 
p	2=�/g�'��+� t�so0��;5Ϸ+�wżkx ��J�b�T @����T�A�F�"x�T�P�F0���R��EP�#@���*���R�� !2���F&�#��'����������➞��>�=�T _O�� 
�� "��� 
�� *��� �@T�'���)�L@�L0!W!T�cV@�����7�h����SO�	��ƲN��D`8,��hK��y��ɾ!�ϷYo�o����2�M0&a�4X�aV�MB�
@��5���\�I˯7]�@����ɴ�f�283�|4�,J(�4�G8�K���|i���5������6>�a�2����B\��d��Rċ��%����.��U�*����.oG9��7�C2�H�Re�P�)m/
�=��<���7w������"D��������J&S����dJ����bAB����F�Ē�8K~�
i�
2��
�hۡ�5���Mʱ$a�iB�9$,�LI�����5����p&ad�-i����?C�B���1���B$HD�����!Ja3��B&!H��Ą����7��C��\�F�����V[���M��!FFB�J�hd.R�Y�aW&3�_$/~�D�c ��@����-9=E)S6�B��_{c*s�����������&�^��9Zb&eR%TJ&j���U�Q�!i���� ��K��`W"t1",�X��Lt��G �q5�vA�0!/\E��7��� �w�������P��D�Й���ow�HK�1��
�H�F���c	m2
�Е%����#d�:M��:jGOdw�k��0��8��4S�H7Q	k��t��Jb�+Fm�!�2$M��� @(&H
�H� űjD� d��nH��3t�@���p�������D�"�j0�KInd3"������7�vhԦ��:@D	�zT�Üe�u$��m��)�4�� ������H�daԋX��V�iF2H@�	D�F%` �FH�H� 1$6�u!����-:(e�cd!�!�PbbX�1>L\��ưB�
�XC)�� �4�)�W�䦈����� �n�JBKa,&�@�H�H���cJ��	5@�˛��I�.�r淽�>8��˾$a�8K���
�a�ayL�$�nD�&���|r�E���d���z)�����L�U�@��ݶ{Y��$왪ph�œF��oL8Ӧ�O��='FO��,F,�BF$BK����0`�2c,�@�$�dHD� �Yl�!`��1	J��"�+0`Ă��	0��Y"�D�@+>Y�Rv{�D���u���I;�ٯ�w��á
l;�t�|C��6�<'54�C���nkyd��� �� �%*���{��%]���9��s]�a&Z�,�$�R5�q��͓*|FH\\��e3�GbI��$	n�g�����~==ҟ�"Q"@��$&ay�o�@�GKi5H����4�y�Ŋ�
@�5��kf,��k�O(F��!#BE�K!
[��=ݩع��M0!8B�@~��0�1�&��1�} a=`@�:��!c�섅vB�iz?RCI !�P�a���������SXԴ#H%.7���~"@���M1�䲐�VF����߇�;őjd�66BR�pE�)��F��b�a0
�ԑ
����\�����Ū@�� ��@
 ���i�3ۯ�|a�b�a��	��k
}�sWqNiٰX�ZJ@"X@�E�ȽL���@0v�.Ż��2�BB�e]M�hB�����#��G�5�_t�r��B��̆Ɇ>L!XXd
LH�Ӓk��;����MJS��@Ł�Ir��_�}'�y�7�����:�u���5�}5�F�	���Q �'0�5��v�dIR2E�H�%p��6sG�i�2�~�jyG��Hrc#IYS����Ɖ�I��(�>'i��0�G�̥	8f���tW������XUbP��A�б�@X�H�a"L*H� �1
u��>C��C�
�!��@��0J��(@��kN�-۽lٲk\e�f��N���$f&�b�FY V�	"h`BH�N��0�"F#JiIB`U��H҅F2!#���!L��A(T�C�cr�P� P�+
�jK	����wc0�y��6ki���(E"@dH~�d3[�٣\��[�����r�s���zN0�r6��0��F�2�|���]��G��$��b%0#D�����'pk�B�F�`P��f�a.�C4L����T�w�}��z&�U�Ww�f�\�\���FS�jK�0�kJ�>�2`�xRg�DdyޣU$)�+$hȎ,(c�)�c.�������ٮ�!%��	��$JxS=����>ic���vl�\A)�$b�F�jD
&+��B!b#��`�0"1!#4�$D*F�Ď1Ӂ9g�oA��adJ�$X0$ H�`��EbB1tB� Ą#!
F0"�(�(�w�E*bI�`T�B:iߥ։$i�		~��Y��	&�a�jB4ą��01���b��)�%Ll`Dё.�&d+�C�zf������xq�q�D�ޔ��)��6w��&Ka�g�I�X�22��!	�JNk��g��t.?bѿN�	HZ������z��ceeaHVVP��n: �:�ҙ���
zBnd��o�k��f������
¾��
c�6J�I4)�<���e��� E�C���\3�ޮ�r0�@��$�D�4^jdXHu|�HH�$ �1H$ Ё@�	�27\�+F�#B��,�K
@�Nl�R!B��Ԥ� �s�f�q;���(B�HԂ�0!Lp�����i�|o�&Þ��##J�Jm��2M�$,Q���FU�!
���ҝ�>�Of�����Fw�$��X�)[��]kh�Б)0�!)J�	�?D�(�����0��9����P�|���/Y\fl���ɻ'L�����U�H����7���`�f����IM��!I�� >5~a�	4�I
ᥐ�
KɆ��gtn����B,X ��,�k�g�l�>�&�L4$��&�HC���[� ��i�Za")������;�m��K�Ƒ��!#���|+p����B7�#�"�>\H�#^���	r8a�4"0�G"�`PĤ�0�:`�$�P�"UƘH�"إ	$p���LH��C�qc&�M��
���$�	�,I��u���YˣT�(K&��
��F���R�v@"�b^�%:��ݚׅ)}�>�B��fq�4FJc.B�4B�`Ё0�! ��4B��v|�~H�D�F0�?0dG�*�N)�*��$hc��)K܁�R@�F$�Ȱ��JaS	bk�$$#��� ����5~LF �I4q8�GHF�r���sDޚ;�5��g���n��P1����Yɴ�CI$zd�i*@�F(Вҝ�e�	y5,���$XV�#Ө|��P�P[�L���_�Ӂ
�$���c#`@��D � #�V��7�z�"HC!U�lHP�/�
��ƤP��$���#u#c�#F�$���$X���#!5aHBl*2�d�!6��'�E�;)��m5�7z��ĩ�5�t�-�ㄘa�Ȏ�z @(��k���D(�D4Z��}Mqڻ��^\��Ʉ!5������+���>����H^�HWBF`�Q1��d3iH:��,�ؒ�EaJKy����!�ߒ}�%L%Ͱ�oR��}��jD��lc'.`F�S��H�
H�`�D$���"@�^�UU~m��m�m�  m��  �  �`    @0���  �  @�  ր k      l   p    ��� p�2���ȡT�W*�!���Z�8�8튕��b�5�i0�Ut��r��p�C���0�*�j�G�B���� s�K�VͣV�ӡ���-��nʶ��I�V���-Tp۶��L����f��h�f]���*궪�-T���^ �K��p�m�����#��l�o	�T�˵UJ��	I�mnԫ��g
��@x
(������q��@4D�0
ۣt��x��c���&�!n1t�s���z=wJv �  К�g*�:A����V�jt���n��t��7l���Iі�:�����  m�E阻Y���`��   ۶ � �ZU��35����R��
l�� 2��[[l6�m�t�p�cE�5�e� �6�v��  �gG*2�u�-W�*�&��  qmK�h�-�W,#���lF��i�¡|��+{kiTȽ�:M}XkX�-��JN���b�jw��n�԰(�4�ì��$�] �  y��Pm���M��Ÿ6�m� 8� ��wa�ø|���UJ��cSR嚪�R8�i���ҭuJ�̙*���W>wʵU�I��p�V�n�^J.7��iU`ԃ���fu����~��^l@U��ڃb�k[&��P�\a�	��lJ�F����]qKOFm�F݄��ۀ ں�i��Hl ӗ�@WT](�y^e]�
��rk�ᢵ�;H�V5uT����B��9�d�l6��k �W�R�mr�mFT_%�����tR��mR�x���J�U!> r�UUUuVU�W�]�V�� ��Hv�$زCl��+.�q1ږ��oh[`v�x�@����ma��J����#��[�F����8��<�̻5��j��Ywʾ��u�.���^^n�^S\�ak�T�UJN�`-�u/[� [�֖}M��v����L�j��\ia[[�I%��f�l��i��)�ߏ�^��m��ѴZ ��l �+T�]m/�74����'�;*�UTg�x&���y�6*���k`  �"d`&� B�Q%.  �F���m�\�� �`-�e�Q�knׯ۴�   �Ͷ[vۖ�-�H H p � ��4�E�6�H�V�޸V�� ��հH[v�i�l m�w��@86�m�� �ֳ�m���"�h�kX䁶� �- %� l[��!� *���YWT�*ʷ*��[@mH����qm��m�8 �T�U[@�5tk��@f��m�8�ڪP�eVIm��d� � �e�[e��`-��&M� l 4�f�E��.�l m�ӵ�۬�@*C��m����  8 -� m� ۰6�At� m����`	���t�4�u-��V��U�*��^�6� lf�u��$���ŵ"��l ��m�� m&�$$ � ������ 6@l�l6��+d��WTҭT$(����Un�RX.K��s��Mv��ϛ�[	Ų+sۥ�v�cu�w�8���}O�=me3�k=6���Hd l$ꮺ��٪U�XL��&Q���  	�Y���]��Q�EJ�n��8�ݪەn �`$  m�Im�h�Ylm��am
�
T��Q�m�i��ePK�PM��g�� 3k6���bZ�4P���I��eM$���f�s�B�#G]��ҙnV���Yy��S�.�C-�[��@^�m۶�������$�'&0 -�t�msom�m]���8l�#Ke��!�hji�v�\��WI�����o-H[��l՛`Ie���v�Н�d={��Z��{ 5T���nx�*����&�j���]vxO���/)����m�6�$#7�l�/Z�T�� [@i4��\n�a�����Z�1�l�۶�v��l��z�I֊Q{% 	6�ݮۮԺ�^�2�C'I����HC]n���'� ۶ ���[m��v��	 I�bK�k�6�t� ���#� �-�m ��$GXl����+��Ͷ���  l�ͶH-��i��I� -�~/�]~�m���`�a:v���l-6�l�Ͷ@��t�[lv��l�u��"@ ��M�yu��J n�H�KV��l   H��m��)<��J]�Uڹ@Z�eej�Z�^�[l m��m��mm� �7m�ۻlP
�@R��[����g ��m���kz�66���s2��x���|` �l u�z� pm�j������� kX-�Ͷ6�@   ٶUU@T���Ue eP$�����f	�d�UU@�T���32�u�8�� m��l�{l�2�U*��VZҭ)*��b�J�UTW�k�۵��H	 )[fͱ7K�A���� �������[m*�J�K�<g�6l��� �@M�m�-���**յ6�z�KU �٨�i���n�@� �� ��f�V�G�� l *U�#UJ�U��3ƍ����c�ڥZ7`V��.@PN��y�^^�:IdI ��I(״��uN����EHku�f�#]�`i,F�� p�m�I�m�[�p��).�d7m�8:�US�&�m�u���@;I�uRlI�Ul�U�d��ewI�4��7n�������%d���v[Ye���6���n*�
U�u�E�T�֩�z��Ӣ���vY6Y�%����h�A�3k��7�X���e�I(��V�tΆ�n���oQm��d�[Q�UU*��������[�+��n����Hv�l��l�G�Pvj8*���� ��� ��Ԁm�m��-��M���N2;e^7�n�J��F��f���2;G]����ֱ�=-���m
 K�����-�-��C�6؅�n���)V^��UVүU�ttѝ:���R^�S6���X �h�+EUUP '�iS��V0��CAڞ�ڮ9V1�n��`  p-� ���^�Scm� $�����
�Pp 5�	��� 	e[x a��dH�@t]����H]%ݥ[@: ���x8 ր�$�Z�Xv�6� �c� H$�� ڻl�8H  �  Z�psv�m��$li�u�m� -���m&� m�$ ���j�n�:��f�c�6�6�  � -��   �[r�m[ ��5t�,W*Ғ�t�E3f����l�6�E-� ��M,���5( :M�[@�$ku� m��5h�m٭b�j�[*�T��l.�l h $�-� 8m�m�8�$�ݮ ׫�j[Gl��\6��m[�dR^C@T�l����j�3iU���V�U��/:���lm�Num��x���E���S+��L�sg�u���K��EV���UT�� &�J΃��m�7NM���!n'&uT�d�� m��I6��l�XJ�6jN���J��d;x�u�*�y���[x%�!� �r�5Uu��bl	�͇�1m �8ͮ    HY�K�j�J� ��c�ѭ� k-���+OM��������t�*�j�I`�����5uGU��.�O:G�/�SڣH����*�]���P���ڐl�`��[�%��	�%$t�$$   ��  �>��l������m�  �M�����`��@ ��6$ �`@	�m@�ko�@�2���ͬ�aoV�&��x6�t�!�哚,�e��;-Զ�ԽT���z��r�@�Y���U[l(z����6�k�gj m"��	�}���l���9!&�$�m������� TӦ�i�!%���[�t���  ����  m�  nͳ��$  hn���o �8�j�2�����?W}W]<�K�)��Y�]S�+�v�Bj�Bn����`��҆�ڹ@�,�\\�L7bV�jAR�MUU�]R�gz�$ n�u�H  �<�Mnm��n۰ �|����{�w�M�����m� �*m�Z�H�J|�ml�n�lE I��C���	V��9�U[F���kFmpb�,vz�
]t� @�h�`7b��Y;moW3�&��  A�@ �6�  8 �I�  p	 �m �c�8��+NWU�Imq!�e�4i�����]�4�W����ǥ��b��������r�ۻa��鵬���((��ADUT��?�����)��p_��ʫ�*�½t� @ �(���7 ڲ/�|  ��DB���@g���^U��BA\؎�N���(�t�t�F/E>D�A�I��	��j� ��E�VA�Gc��\ ���$�MT+�8�m�@� S�AD� D^�]���qD)؏ ��iH�t�ȧ �DO;R (? `�<$q:k�a�ФdC�8�#�9�R�b ��R�qS���}�W X �T֐a~T����B�OuЯ�X�@�J5�������
xE
�Ah�����4��S�O�~
)�ォ��LD*�b4@����(�O�&�Џ_E�O(��M ��	�R�� �M�D҇����I��8��(���y�8�D]E� z �^��D�R!�p��PHDF��v�����ʆ��]E�pA>T�X�P����~@!O�`��_������@���B ���h {1QC��/:C�V�A��+���BA>~���!�t��� M��DH(iE�1Eh���uv��[F��� :xlA�Uz��8h@��|����@ U�G���q�8#k�"�#*ʀH�E ��Qb1$� E��@0�D
�P�Y���$[v�m�$�p�5�6�	��i$�r�sc5��]h���F�jT�ӂ�ڪNw1��[�o�'(.�s5�j7\���ڰc�;n�X��N4s0�UR6��[,P��C�z����� ���ۉ��Daˣ�5Þ��л�����Өp��&1���'t���^�����2���B���7�7P���zv�݉���\�5�
-,O%��Ǟ1�/h�;W^�:%6c[u��zu���v�k�\l��c�]u͊�آ�*�cD�AJ#��B��f��K��F'�Q��lt纇2��m��ғJ/J=K%�s���em���䪪��A��eg7l�}M,gk@Q�p�gZ���˫{a����yeQ�Ō/K� ��Z<��;s��P�bd+Fܜ/X6�'F+�����sls6�0�qAٙᤇ�' =ۮ���q��4z��H�(�]�8�q�8{w%<K����	�H|��V��հc�9&[�gtv�����Ca���n�a��aWY��!�N�!�ZW5�-/�pZ�[��f�u�&�I�ZII��t&�iT�$
��ک�#�D�� ��+a:1�g�p��m<�.qœ����v/[T[v���U�v�n}c>rZ��h�K�Z��̲���f�F�e�^x耰fτ��k��oPKZ��mn^ɧs˱��ɸa�%�(6�p7�^fȵmVw:W�;.��;X��m��d�`����j\ĭR�UU�B��T�ИuI�֋4Iv�u�4O�fUQ���v�ۣ=���̩ټH��].�A���>�狄6���eTs[��Q�q'�j��'�6N��:���m�u�q�A<B�Up���-��+�偶�P�g�[�՗unlݻ[s�;�g��{c�H�B�c���O+O����]y�������hW�����lm�J`b��=I' Kq�a��ψ��%��fˬr�`ؒ3��A��6h�w�������4	���5�Q	��ȋ�!��8��:��P����W��� ��Q^�L��]�,Ʉ�.���њ5h��m�m|\�Ӧ�:��7�M�˶]�s"��N�]ka�T�M�������̦��#�к.4�����1�z�3Wv�\���r�Si��9�ڢ����a����k�4Ra�6��Ŕ��㱣�v�+��e�b,t�f�l�c��=�FK��15lG^T9�9c�|`�$�֐v'TCH�B7|䕘d1�v�.��ݶy^L�������8S���r)�xIR�������s�l�́�m��p�}!m����K���I���$Z��9�&I�l��ŀzX���ښ�9�H�"��@�s@��s@�Rՠ_��@�c��0�<&I3@{��M�����7[ŀy�ndp�	��3@��Vh�j�;���/u��=�3�~H�I�qD�$N�]ZE�Z�ݹ�x��n'�՛��C�+g�n�q��񸜃F9��?��?yh��h��hWj� ����$q�2L&ff��{�پ�k���H��@���D
)����#�g�x��k��?Ss�{htU
ۍ$7��]��ڳO~�����@�{ۚ�[��0pO&
L�;�d�ٓ}[�`{wmXl�n�V��gUI�I�cNH�@��Z������z�%X�D-Y��~��NjhuL�=�Qz]U�ۮ�Z��-�I��3�z4xs��n.�U<sHs�E����{s@�n���Y�^v��-O�l�`�J���=o�M���s�y��9%�M[Fkc�Ӧ:CR�mX��+rO}�������B���$�d�x����&�S��(��U�Wr��np6�`u��7]�4�9K�G�&<#mŠ}m���ŀn�r��np��NPW�`���S�k�`zK�Wδ������'G��6$�N�yҚ2�������� ݦ�`���m��=���*�5J�h�Ձ�Vd��2o�vl����^빠}�]i�D�&�6䒰�np6�a�"g��Xu�+ /e��?	�rE�}m��/uٹ'{��7'�T�@IC@6�t@"���w˹'�=�ǋf��9&h�U�w;Vh�j�>��h�LHF�1��E'1]���c���|�<��5��e�g\l�/6d�Y28G����;��4�hfe���Cg3j�<�T֔�U,6��Y�_��@�۹�Uֽ��Y���G�)q��rdɃm����s@s��J"e�}+ ���='��h���G%S��6""'k3j�̭�V|�Z�������(��ɍ8��nV�m�O�owb����2T)VB�0^�NjY@锚bl��Y6�8�ˈz@c\��R�[*uТ&H�)��nܶ�����@�Yy�d��D�A�Tr�6�nt��2k u�'^v��2;�i���<q�����Y$����W>�.:.����o��g��{�kK9�asUۇ�q�{33���A�B'��ح-�P���tP���4YuQ-���Z �+��v9/	�{������oy�7�$0����Z3���ŕ�g����=������[���H�v�����&�6�>�~�@�۹�U�^���Y���CI��DxC�h6�g舅2t�Հ7]Ұ��8�u<cF̈&䙠_��@�v��/;V��v��gY�dp�	�w8�"[��X:��m��mh�nGV98�r19h��@��f ���}M��9(����Z�1#df%1��"�㩺��#:7 ��;/"]>��d��i�����m����0����nWD(_Hs���=&�K�yq���o��b�����:��@���MDʑ$@Ȣ&��Oȫ��}W��:�8�m��2n�e��(�&L�@��h��@��)�Uֽ���bPj4��ێ,��)�}Ӏ{��=�s�o�\� ������"1���zS@����/�������Z���b��H��V�
4Ͷ����0����WD�$9[r3�m��&��j)���ap�/>�@4�h^��.Vu��&F�HjYT���ՙ*�BIL�;�V�'��j�?�܎�nc$K�NE���`{l¢�F�(��&�2f���ڳ@�;��#�G&L�6��@��f �X����9m������ohM�F�4
��@4
��@�����gԛ���c���jG<�@���k��t�ƚr�[�#���-a��D�D�2cN=�v��*���ҚVנ_�]iA��jcnH�@r۬䒙7��t�u`�nVr�ă�=�4�� �C#q��<h[^��;Vh[^��J<cOZ�-���X��`tܬ�n�6 8!�+*� ৃ��C?��~��gY�A�L&(ӏ@���`�$������X��`)��;~t�i���oY�k��c�ʜ��C�\�A�0&Sv��v��ݎX��ӆ����`����� ��`Z�e�t�m4�%7V��j�D)�gwj��?yf�WZ��r��Ӎ��8�wV�:�`tܬηX�x��ݍ��(�&LiǠ}]�4
�נw[��^v��:4���i8�4]ܬηX$�}�/��]Ӏy׽M�:��)
���	-і:�'��X׳Y{֗ڣZ������݈�0���"�Ǌr�&�nWV�%K;ml�����gY�uI�[�t��툞kQ8E@拖���)���H�Xr�`��y���y��&�:�5{��C�w@'.��fZݙ�]��ϱ�2n����3\���1���D7c�F����S/GgB["i.Y{v�I)���w��wx��7�\9c��L����wY������P�r��첐�6:��{���=���yڴ��f�WZ��exĞ�L&I3@���Λ��9�� �o דu���dR1F�z�ڳ@��zu���j�.[�Ս�d�c��ȳ@��s�n�� s�u�
�� ��R�:j���M2��fe����f��-����ZiɵX�m7�&��V����.�;a�d�x��v��N&/n���8�Ӎ��8�$��W�^��e��W�uD%�=���>���3J�irh˚��'{�h����B�
����B��y(�ǝ}��6�,ϵց���5��A�ә�_�U�}m��*���;����jN~ �ت�� �o ��� �o �Z�@��+�$���I3@��@�o �Z� �oТLV������77�qg�h܊���g��d�ל������Wd{v�n�Ί�\H��m���ذ��8�x�>�XM���W�(,r8���_�U������4s�V9�����1b+T�T�M8&e��7��`ծp�Q�y4��	�Z�s���>����À�����<��jc
�T�-'���5q|��l��H���L4�H��N�LdEX0�H @ 2�	+)HKaD�U��ڂƆ	�}�6��X&����`H�`�B+0�Jӌ���@��bsb�7>��
�, �ٛD�<Sa�)�U4e@��A��"$`B\�)���JB��egu�c�vp$ `�H���K�HcZ�"E����k.�tѦi�meM� �!�|��ā@��*�H�Q�:!6@����q�}�|�;�xl��F0�ƈU7�b@H`�o�v�F*a�bC8+p"�1bM0�B�P)n������ �CHD�F�
��E�
|��"��p��
 2 ��`,��(�*�X�`�$ z*���X��
������w�	�'�@=���훒w�|��|�di��Oc����fg��y�`fnڰ2~�U�B��gw|�gu���3T2T��M:�=��V�B��n��=����{*��~^�-�eP<i�@6�^�۰���z.\Ѻ�.��<�rNn�o�#��4YR��S54��t��Xfe�'ٕ�t/�7{�Xrޒ�\�$A�I#�>�w4
�����hwW��ٟ�:��<bOZ�&� <�� �o��u�y�� i��H��E NI���V��٠r��rO��lܘN,�ƱP��AD�yD~J#�~���v/btqT��%St:����ʰ<��������{�0ۿ����*eݨ�ӎ��-��֛�۳���gk@�k=%�M��6�3�C�ه9�$�����`���7[��Hl�Հ|�U{#N6bx��f�u�@�s@�wW�}��o�;���ȓ���T��Df�~_���mY�>��V�����tK(�F9�Nf���@��� >���_w� 7��*f��)KmՁ�fZ�::+���w�Ձ��@������6��F�	�s1p���1i�9�Q=��Cf]�����Н�����@H#Xр��}��퍸��-�ۘ�q.k��BZwf�Ȝ�sd�u��Q�!˒9��]c �Ψw �R�k.�Mֺy��ldƻ#���un^�V��>��}�cQ�@��{J[�����H�JWkl��Q�k���+2� ������cR�yu;أ�߽��=�ۯ���W1��˷m�q>[)�����d���\�x��yx�n�����?n�pj�L&� }���u��˺� �zx�=�zdX�8��I�4��gL�-�`�|`���kWE���##s4�uz��i���f�3wmX�"���m�I�$�X�l����5�� ���>�g��Ӎ��8�䆀u�@������r���:�M��U�t���������wm��_lZ��9;9;"r�
b� z#�g��7�<�x�X��O�/����ֽُ��(K�7�����4qR��L�34nI�｛��.Q��߇�ޖ��ٙj�B���3���3M�)Kt����ŀ}��c��e��9}k�;���hz�a0�746gٺ���V��ʰ�9�zX�u�c�(��'$�:۹�|�נ{1�`{1��t�wI4:.tp�!uV�wgj�F��7V�+��nݺ,��MU+�]SM�%6�M|N�U��ǅ�}�ǰ�Hf�ڰ:�!�j���'�N���K舅2��`f�ڰ>�fUꈈS'�d���ӪҧESl�f�=���iBD(Q�)%!%��4ESR�Q��5hUH�X�#(�5",P|��~@6�>�/w�nI����?}�ni4�iS�SC�t݆S����6_u`ݳ�%:�� �ԩ�J��ʚ*��>�fU��
9$��~����`{3-X�B��6f�P�Y-��n9C���x�vr�v����q��GV���G��_�z��� ݱ��-�����ϋ �َ��fZ؄��NnՁ��ڊ��]B��K�X��w�#�*�{�Ձ���`{1�{	)�wCj��U6�!Jfi�`f�ڰ>�fU�����O�ޚΰk+s!�qXj���ڰ3u�`{1�~�!$��,�D�`|~�)��o����zbRI�N=���=��7_�3wmXO�*��[�d��,ĳq��ѻDs�B��k{m���})��E���I�vɿ���F����n.Ij�ݱ���;ٙj��}�Z��n�,��ni4�f�%M��v�2��:*���{�����"d��:�4aR��SEU�ӭ���0��M}׀>�ŀ\�'0A�H��:�M ��x��`tB��}Հ7�ꊚ�n�!Jf��,�f;TFn���NnՁ��0��! JR��]��IE!�1����-a��M�m�dgW[�5Y���T�D��=�����	�j��lggF/n5 �9�q�|���vy�����5b[��8H���Sڱ�Wk��@��e��:]O��$�9��'bu6)z��g�sb�g�Z���83���[��Oi��r�h��њ컃�C�.qS
sn�E��,���+se�\N�+��K��If��6�&�l���\�1��=]��e�c8fX��grl��crH�$�����s@�u�@�e4�h:���H��B48�h�n�m��kw�ko�O.C��1�$�'�o���u�O(Q3�ݵ`zsv��}�174�b��]7MX"#�EVos�3��XO�*�bDNn��`}��sI�34�*U:�M��ŀrIB[O���v, ��xߟ�Ǐ���Z��c��q�W���{]�(��^�[���H�v�����v�Rp�q*�*J���/��n�X�n�/�>�����c��a��8���ٱW�� J������
${DرMU���"��8�*����N�M~��ܓ�����>�k�~H�y��6�5$� ���o�(��}Հk}� m��2,nHDNI�u��˭z��jæ}���՚ʕ�-�Nhu(�Ձ��2���7{��os�?{2Ձ����m�tp�+1<��ƕ0�m�Q�Ѯ��c�ʽ�y�؍q��:����%W6݌7_��, ��x��.��6_u`'��M�6ة��T� �َ�!.QT{{�X;�V��Z�P����m�&�%+%J�����<��`�n�ĈD%	�,�- �#YT��h����J׽�X>��:�4aR���*h���I)�}Հ7݋ �ֹ�؈����`l���U5,9$UT���oД{����_ϵ� {���r~r���W��%�t�OX�T�v����n�^V³�������z��<��f��i�k�mf́�c��?{���_�-��4���I�!<Y�@�v��%2o� o��ֹ�P�bG��{G1̆D��� ��M��jΈ�QU��3��`b�+SUM���4݆�D%9�����Vl�{��ܟ����D�8�A2
�G��"%��_�?�9�}�;(Ρ�橶)hr�5`~�{&��
!B����|��v�2Ձ�=�_�켊Y��y��зV�i	�F.�K's�:۶�"z;1_��Ͼ|���h��d�W? ��� �u���]�>�ۓ�R��R����m�X�{�DB��ŀy���<ݳ9BIL�릺F�0H�6������Ϫ�߳�~Ļޞ4�}4�ex��&�a1*tڰ�^�ޛ;����a�B\�I*���X�V�MM7.B��T���1�`rP�DD(�n����V����I�b���P�HKA�F3E�Rh�s��:	��C�>Wfh�n��`X�0�"�����Ě⑰ɳI����W�H��)�'�~�� V	���Y�� @�������6A��	�kО	���tI���!B(�c(�a.icpbMK��D��H�"ϴ/�m����x�|&��B0�b�~���<]�����&���� ���h� �X@�J�N��C�E�H��X rM�ۀֶ� �mq��0Zjp5�����k&��T�y�'�ή׭
�^70���mh�������;ut�=��nh.'G^)�VA&sl�km��V
�w&�KW.�ö�v%X�`!�k���v�����GF.eR�ok3�F8&ۍ�݌WR�%�$@�n��;����Gv�P��&��u��t�f6j헞`�.f��.u��]�M�N��丛N��"\^[�E�j��5e8��=�5�Z�A0�OKUlfk�%����d�1��L�ђgY7U�;+z(��.���W.*���M5�]K�aYU8��Jڲ�Z�p��uv��77$q]�< ;��Z:� �v�`�l�U�"j��C��pss<��Z6ͥݝ���FQ�6�8���l,���;.�Z�B�6c�Rp����Md�nNwdiG�"�zp���cS:+U��g�W�7lZQw1�m��AԽ*�������u��鴙��,��䏛�K$�$.�,�2����I�wcv-ͳ@i��x�.8-SUP��۫��j���ϖ$���g�*�ݲ�hln�m�J��RʤX�%8��n�lO=���a�Ƴ����-�p\8W�2�#�m�-o+Bm	&��NK`-�JHi6)�j�v��l��˨�z��xN�;v�s���$@�z�V�W1ɶ�3��:쎕�᭕h����v���:4k��� áX�J	�s��tpܲ�-� g�.��'��n֒ym�WZ),�A;���[[V�%\iv 9ی�jy���7 
$v7H�sє�I���z���f�������6b���
·6�2��n��;!#Ud��;R�H4]�u�ڐ��Լݝ���V�]�s;X��ڷs��sAn�v�jyZQ���=�-?7�S:˶nMi�Z���gc�G���8G�3��Ν��pSzv��}��Kv68{+�$�2�b�:��j�y����h_���?
u; �Ƒ"�_�>� �<���:
(�y W����dX�L�V�Km�����m�I����o^�ԉI�V�γqq����V���$�-��1�w���
�/[������RLu����'^�Gs�N�6���v+#
ݮ�ȭ`r��{��3�8�ꧦ���e��M�6�7,GX��Et!ֲ�=����<&5Pu�r��v�S�6����t���T�gG3ѱ?���V�L˚8��+����&�au��)�<cKjݎ�.3�)GlQ���=�T݇�lݺ�
.lv��E4�*�j�����`ko�ֹ�/�u�rh���m�L���fe��%��T{kzl�|X�{�P�O��Q���m�KC���ٰ=��(�=�����`~��ni4�j�J�NJ�6�Nu�N y��u�X�|����VU*�T�j��ۦ��?{��P�37g�W|���h�S^brbcq!�C�u�ܼ^nJ�ޜ�sod1k�vYd����wk�z��0H�6���[�nhwc�>�̞P�B���=�����uP�V��h�-�f�nI;��[�xn	T�ì�T�AaVE�P�"��{��~ɰ��`{ٖ��9(��{��М�Sn�JS.��:���>m�	)���`o� ��ڛ�C�"X�ۋCٟ�����-��4���rQ�U�}�`b�Ws�3M���5w�6�,��m��uwN |۾�o�����Q{Z�ד����H�rh�7nm͸D�9$��ף+ӌg������qq�47N������̛ ����G(��;��X��sI�3T2T�tM7`fVd���`n�ڰ�1�DGD(UFn�]R��J���m�nl�ޫ=�l����bA AHr 
�P��fu���p���U%����B��XrK�(��]��+ ��vefM��a$�"�si���ڡM\��5-L�wk 7�VIDDCv��O>��w4��TV�FD��1#b���nE]�]\Y����&q�=gn��Sw�w{��;Oа����D���~���f�m�[�H��`}�f�mQM72��UT��3��{	L����}���̛�J&LX���d�ڤ�R�wvՀ_��{3�^����z�M ���rD�B����V��J������6���ܟ���a d>C�@UyE�����η4�s4�̩T�n�̬ɰ:"rUۼ���Հgَ�?w��~n�[(<i�F+����tk��%�9��q��:���{c�����rqr�U�������� ����uwN��V�U# ܒQ4݁��j�GB���`wWt�{��fL��
h�A�䙠�zh�V�H������@�A]���CĢrh{1{��Z�}4l���1/w�4�.��4SM̪t�U9�����(��߸������6����~�IB�س��Q�0�'0�#X�@Q�NZΎ��8��Q-�(B���J��6����b��4�;/Pm�v�+l� Һ�Mm`�q����%���x����;����Nvv�G�\m*�m��)ԁ�sk��^;v�v���w�v���춞|֖���`���b٭ȴj��n��l��c�#�lt�4�A�m�A�Zgl��cl���] �/g�b�q�����w�y��jp�]ڀme9�v��9gc.���6�;A2
V7v�נ�q���;}󾕚�۷7�}����1���?ȅ)(Q�0�޵`ͮ���M�)hn�e�gَ�%&�ń��j��ǅ�L�f��dI�b�ܚ���^빧���<h�ޚ��R�&5�̒d�6��b"w3+w^��f;IN��Z^��D��
!)3@��h�t$������U���Z�>^̫�+����{g���v���K���l���]�YĞxx�n������ۥ�;�Pi˚������n���rJ#��0_�Ɓ�$��ɠr�^��TBK"2"!lB�U�o~�`{u�`�c�P��D(�=�o*nh��ȩӪ�u`v�Z�>�xY�(S&�u�9�V��X��:mSK�Ն�I%>����7ۮ�=�c���"�w�V���H�9&�8�h�٠���X�x��'0S.T�MAweH�������S�-g]�Nܻ�^Ñ�@���6���w�����dI�b�ܟ�U}�^� �oBP��ou��dʻ�R��m��i��3��Wˡ%F�u� ��vә�{�)�'v�J�RK�DKj��ݵ`�c��J J��A�v�q ������ܓ�����;�JʡM�2]N[j�TDD��u��ݫ=�aВ]�����=m��ܒ$<J'&��ٙ�=o�����V�f;�"|i��#T��lrp�s����G���b�����Wt��v�=+i�Lr&)�#q�����s@�j�3����=;�V,EmV�K��2eL�mX�e�ԡ)��n�ӻ�r~,{߸lA�?��A�BQ"��}�]#d�ےT�tꚵy����lA�lll{��~͈<���`�`�����b �`�`�`��~��b �`�`�`���~�&�[�5)L�L�kb �`�b�X �?~��y���y{��y~Ch@"��W��"��~�����A�A�A�A��~妵�)sF����5�؃� � � � ���p؃� � � � �߿p؃� � � � ����[y��߳b �`�`�`����?[���ԋ�]�{;<�:��� �㫉�=���6�ݓŞ�6�u�~w�7�mc�k*�:S��w?A�������y���kb �`�`�`�����l9���y~�Oِ̓���̗5u�y���kb"�X � � �?~��y���y{��yO�  .A �`������k,���kV�-��kb �`�`�`�����͈<�����{��<���X � �߿p؃� � � � ����[y"E	G�f�:�j���sUN�BQ�P���Ql{߸lA�lll}�߸lA�lllo�����<����s��ٱ�A�A�A�A��k���.�Z3R��kZ6 �666>���6 �666��~��[y��߳b �`�`�`��߿p؃� � � � �m�x�l���S&9��ܐ�u��׎�VU��2I���Vb�nL7�+�B�
�ԁ	r<�����s]ka�$��t�[r]��	���7�ķ��Mũ<6�f����z��d��ݍ��H�6Y�������l˻7]��z�����q��t�f���<�+�ڈP���0MQ�WBTOS���<psάꮳ�MlG\�T�x0�cm�a������-J�_J
��*�tԡ��M�k�zG�R-�������C���3��&m.�߾����b��u��5�YK����؃� � � � �~���A�����߳b �`�`�`��߿p�"� � � � ����lA�lll{��j�j��)rk%�kb �`�`�`����ٱ�R���߿~�S��9�߷�6 �6667����� �664P�n���M�R��n�u4�Z���(�A�A�A��߸lA�lll}���6 �6"�X � �~��[yg�~͈<��������fe�$�Yue��4lA�llER�߽��b �`�`�`�}���lA�lll}���6 �66
 �A2?����v �666?������㚳Y.kZ�M�<������ߵ��A�A�A�g�~̀��ݭٰ3q�`rP�ԶM'T�l$p�`/Jv��+j�`�p�ǵ��nӤ��aXF�۳������7$�"bQI?����@��M���â"#􁻚�e���%�v�j�f�rO{;뾉� �iGB.B�Q��&W�?�Ń�ڀlW�W��Ю�TV!�i�RW�}���wk�=9��J"d��V���rc�X�R-��oY��3�%�D%U���`wV���eV*uU-�)�����+����C���g�}wƁo��<�LME�21I4O]`����o��;� �x�?��\�d:��J��N���L�j60I�������zHv�uN}������U��st�������6�� ��>���BQ��oU���]%T��%�"n�p{l������ �k��	/�BQTot��R-1��m�,�y�I���70�vI��
�"A����!p%�O#� h1�2�	��D~`� �H,aYCB0ɒ������NEZ�`A �!$*E�&F�f����.�wxC@�f������ �J���b,b�}��A�I��ht�ώ�H��@�M���+1@�T:���b�gh�lf�(� D'�|�����M�)w:�"@�|3�ؐ ��X&s�D"�$�L%B$e�����aG��Lt�u�z�t"x�^(8�hG��O�zAT���!F������à*�7�'ʝF|�p?D(J��W�M��������rӥ5M��F�\��6(��ͫv�f��y�`����q��SMdqF��>�R��
n^��37]�3���`l���n�	i�n�����ˡ蔌�Fx�.A#�G��b5ǲ�����]���\�8�L�n=,��v�=��
]
>���ŀ{z��:��ܒ��S4� �����z��hzS}�����ȉjJd�u2۰2w6��t%U��� ��vfe̦کSM7I��n�5O�oK7��f;T�@�D
%P����V�f5R4�ˢDI�JhV���
�|����o������Ʊ0�������Ƀ�[�ݺ'b��c<Ƚ��O#�c����.�����I��> ����r�^�������x�=���ܒD��E$�9^�@��M��hu�@��[���1�c�&�z��h]�@;��+k�;>����rc�X��4?ٙ�_Oyh���9[^�����յr4ԑ�ӑhu�@��j�>�S@��U�i������5Lp �99���ms]��ҪF+9f�gr;a�'��=��-�%ܶ�3>:pwg�ڶ���Rf�-�7����R^Ǘ^��sl	׍4祎1�=P��K��f9cr�����k��X�ʗK�v�k�.zݮ2�n�d;u��.Q�Q�]v�1ҙF�ۆs��9��j�SC֞�S��kt��m:g�۷e��N�jݓ���w���2r�eC���bt����|��\$�'[�6�,,[�a�z���j��Ғ|��=�e4�ՠ����,vcX��H�9����Wj��f�����h�h���R�$m���&�=��g%
?��g�������Z��cz%�"4��E������[)����{�@���rI&%�@�mz�~�{||�����ʒ.G�D�6���g��]���"��Ӻ�5�aʛv��mm�ֳbpmLq�n=�e4�ՠ��~����4���~�LpK�jnI�g�w� xF*���T�.IDn�|�� ���7l���: �!)��"��f�u�i����b]�O�����}�by�2LM�&݇�R��U�vX�zXz�0�I/ىw[4މc�Ʊ9�<��r=���npu��m������5Ŗɡ�NM�vQ�\�v�F�����]q)�e��/����{��������c6πޮ�g���̭��D~����@���<m=�m9�@:���n�{l�5�s��$�d�rOb�r9LJI&�W��u�M~?f���RV:}�� ��D(߾��N >}x�Cjn�Tګ�\����:����ڴ�Y�����W�y�v��j9��&�r�^�ДOs������`(uL�T^ָjx��W)۞��Q��7=��n}
�K����H���9[4M���7�}�vә�`fy���/�6w������ģ2LM��@�[^��G��K'7k�?H����k�U�T���y#��z�)�uv�?ؑ�_M�{�@�wR&�#B�,D���~W��8��e�X�F�L%0�'9���Y^1��NE"��l�?ي�ޟ�[g���h�*i�7$N���i�)�s���f=x�r�|q��m���M߸@����ݵ�56������7vـk���(�@�w^�Gr���j���r�������B�z���=���=���%�U�V�tԺi�dʒj��;�~�8�n�[w�n� 3��wO�Ǒ'"�����47u����'5�́���sI��BnJ���v��vB�
f^��ͯ߮䓞���"#�OHs(OT4�uAVh�����`�5�5ckde�[�:s�q=L��o���]����k���#=pV�mONe�ҺJNŮ[�U�'L�yD�EU��+m$�6띸2\���ù6{=]�
;ͬ6b����Yq�,�K�q؜��q]�����s�W���E�u�q�Z�n��+{N+X��\.���e���7���o5��ˉ�g�㤛��X��Lٳs6�ɫ�L����"_��5	�o5�2��6�a��H��n�ɰ�c�"��C�ua�v���Q]̪�*T�T�6�ށ��M��h��h��@���6���L��R6��Y��䒪ws�6{��zwJo��E��y��,q��R- ����9[^��ҚWj�-��pMȜ�!$����{�@����&ÒQ�U{����Kr4�2I���;�S@��Z�m��٠{����i��"8�p�	��rcs;��8�	�!X��G+^�nq���|�	9��&������[f�u��B��%��,{z���T�S*����ܒs����`kML�<�@��%��� �v�]79��MZ�"s��$Q�&�__M��4�ff%|}�zh�c���8�H���7�$�wq`oV����v�F%}}4+|Dڈ�(��I�{&�舉�w_���`{�xX��3���K��/l�r�]�Њ����l[��j��<�m�<5������/�9�"r)�������zwJh_U�[�+����s���h�W����)��|`���ͻΈJ&O:;�ՃM�Jt�UMՁ��K�^ɲ"8�	ѢPV'��� �������/����p|�C�c��	�h�?b���p��x��X�(J[y� {6�F�mT�'3M̀~��`tDB����l�u}V����_�2,CI�M�:�#,WJ�b����e܀�(<��� z �+RJ6��9�t&�m˧M� �͚wJh_U��٠_�%��iԺM�*��=�</���""�ޭ����@:��]ԉ�1a%X��`{+�6�3�Т���v�,���cz%�"4��E��٘������V���	�50�T	R!�
�6�©�W��.䝼�{�
8GJI4W��?ٙ�	-����oV����v��#����'	���V.mW)>��r����-��t����v��Tm]7k�N�ʳ�����ߛ ��,���%����Jt�*dʒj�`{3-_t%Tf���=�V�c��%!�ml��SmL�'2��Y�`zs2��Q3�k���ݼ�>��I�Fd&IG������0m���)�o� �w2��T��H�G���[w4��Z���nI�ڭ!���@�oǂ<u��:u
A$ 	�c�k����Sh����6�]��t��"[-��a� \�ČT�=�|��Ɣ�xa,�@�M�%Cwk�H0��	y���0>O�,���E�+LX�c)l��L�.y��X}ĉM,���TK���������H��9����.H���{׽������� �ʵWHM�k[m��$k�gC[��C�u�4��&[�j�+�e��f�oN֑ �N���˪�a2�>�ۗˢ��$tQ�S�Wn�ڐ��wU2]�HX5fӝ�[UP�r�ʵr�n]Y��<qf�,�Ǝv��uͦ�.��6��̷�Nۓ�ֺ���	@��a�ݞ�x��*��Ki�]�-�6�Y�Z組-tv��M��0�-��VxA�; ��#���ܲ�Z�-��WU'���o�en)SUY�`FT�Թ���K�8p�m�&�.e�,���4�t�	ͺ��^�k����.v�9�Ul�LF��I��j�ڜ=�u�ݬ�Y�vbK�[/F��y�e��ڷ=� ����1=��S۩Z'��y��l�9�&$c4q���z�/�����l(K&s̸ٮۊ��q�L89B�9!	\g�:$�e:]����,lcI�c����<K�g�Ÿq��]R�\��*Õ�]t���:N}��pdx�H,���KɪtJ�KV�ؕ'nN�B]�8)��/�ܛr�j���`���-��Z2G�Ӥ��zz�,���������lm��T)�VmV3�˲�*s�'Gl��A���!�̆���{K�,jw]:��	4�6D36�\��yW�$�i��c;�-.�&P�v�w7���rmCOn���.��1�}v�"  1p5�Ueתk�,�k_*w:,b�@j7Eͨ)T�H�MSR� m��@A\��j�6Y�U��C�bi��$ k[A�ʕ[*�왶�9ݦGP�;n7k��Y�0[��*o[s�;n܉a��7Nm,UN9sOڤ�l�X��1q�,!ʉgbh�Ąq�m��-\�A)������me��tk���C�"����ö�ڒ�,���Z�AU�ZU��3�oBtv��[s�:��]�ѻE���Y�`d2Fz,ݮ`n�Bi�ccn8��g��c�a�+j�m�(sU��<Iڿۗjb�A�
�+� ���$6/����h��~4"�/8�!TWh��uW��ϳ.�Z��Y%�2���w38v�=��z�K<��7�V�aힹ��Ƨ��ն�̀t��)�� ���ų���ݣ/����8ix�����/l��prv:X�ՌuZ�1�T�/��&ݖֲ��W.�f�Lv��=Z](�.N9UѶ�.ld��Lꌋ���<����rp�u�ڥ��X"�K=�t	��;2�'*	�*�"��S��������99�sYnY�\��Ք��sk1��k��c�\��5]�x��n��Wﻼ;4��1a%X�!�>�ۚ���ә�ДrK�o>,�Ԫ���N"4��L�>��h��@��)�vfZ���P��UGv��Z�MSha*��p�߿V��f��X�����܎a2H�F�6�z�����_{ۚ���g�_��z��ߐ���,Bn[w4��Z+k�?��hW��,Jq��@���%+ۦ�V^:ۈ����$9DU3��&m.�������j�B���Z���N�۬�v��B�B����;-��&
#$D�qh���+��-'�E8�P	ϧ���w����}V�~�7F�9�R��5wX����a�(��o� �����Tژ��@�!��W����V�۬ДO�g�ԛOF��(�$�4��^�����������<hm��*ˊ�q<�?L�qsք�y�X�/.�J��C�Zx��*�76ݜ�6�((���8�Vנ^��=���������=�w)m:u)�5UT����x_DDB�3wmX>�=������{���ǎ	bpܓ߿~ٹ'o��nP�J@ XU	�4�5(P(�k5n�7l��щ�Fۢd��]5a�:!V�ޫg�������Q
sw+fۦ�ˑ7#�2�X�̫�/�oO�f�ڰ9wW�vR�l��i&H�cc�1��ru�';�s!���ۥ��iY��NzP湦9�̑�n=����׮��������*����<�&,#ģH$4z�gDL�:��ϱ`y�3�(S%�X�!h�8�I&h���{-Y��U{��`ooZ�3ޜ��,�J꬚	S5u��(�ϾX���x�&��%@ґc �@�$1�'�bZUP� ����I  2!��R
��a�B	�SPL
�D`IF	IH�p�? A������ΪL��5��cQ��?�Jh���6}��z�`���N�d��a����0���)���5�v�\�����7�k�e���S�q�x��!��/��4_uz^����M ��.L�9"�\�լg��?(S#�ذ�g����s@��Ȉ�pQěq�z�`=�a�e��X�}X��ʧj�U4�MҩmXt��6nm����V�����4�O6ɋ�(�9��^,��u�k׋ ����;	yG�w�{{��l_ē9��]�R�,d�3r���v���o]��6mY�
��c��m�z�T��-��y�g�:�6vF2�\�Tlr�3���z"瞣mhԂ�E��In�.68�͙;ee��}rf�g�Eu�gf�^���Q����q[��{3�+zN���U�����u��ΛH6I
z+��<\�Vۧnː�.s��p��S��\cV絝�w����w�}�{��o����`#]���>���;�oU��<ݸ&�]we�$p���8��'1�QWwv��}X�x��M���	(�����fz�S�)�:�S*f�X�<Xަ� ׯ����ߡ$�U�wKi��Н4ʗMX����g�~K�U ��s@�����ƀ��Q	N�,g{� ׯ�������M��nBU'2����V�DC��/���t����<�sEeMT�T�<t�R�ZMulp����=�F:m��#oi�'�9�Dc"�y�@��s@��ڬg��DG%Pd��X�u*���Tֵ�Z�.�nIϳ޻������j�Q	T(_|Kǋ s�� ׯ~ID~�T�uUP�)�S!%76�����u�k׋ �����T�I¥U�.QM�Շ$�%��7���޵`~�ڴ�w4y+���ۍ<Kq����:����>ŀz}������7�O=t���0�=�p'��xS�k��q�lay8�|l�[r���\���u�n�>�78�x�O��G��b�;�[5�Ni�ӢI��6��j�(��2zu�`�b�>�79�
"d5>����]ܓ%+����l���5�ŀ�B��$
@��� HE h����+�qW��}�ٮ��;��v&DDc"�y�@��s ��������Jv��`�u*���T�m7J��`~��&�四�~���u빠^��XLPn$82	�K���o����ݑ^�ե;��0�{bҺXdx�k!ȴ�w4��^�׮翐}��Z�X�!h�8�I&h�k��Dɭ�,�Ss�k�s�2v���M(���i��8������j�:��@�wW�s-RLk$�I!�J��}����\��7Xh��$�
*I�X�M���{��{��ܣPq#�qh]�@�g��}�?�/���@;��V&�M�	�B�T�i��dX��,�M�:ɬ�#�N��鳞��ìq$�Hyr-���@�n���ՠuv����DF2'�r� ��,ަ� �M� |ۼ��;1�nd�$x㙠w>�@��Z�m�[w4︭�,24(�,Cnl5uo_t������V	)�y�@��y���8��R- ���Woo|�v����W�l�(I	(!�D�eh�X$�N�&f��<Z�=#03N����eyz5�Z�,�k�V�[�AI�d�v�ە�$�l狵���o�檻."�WF;N�N�s�L;�����1�[��1�ln�˝�=�3��شKh��, >/Y˵��n�뉹P[��iM�ʻ�
��7#d�]F���k��sVu��r�hYe$���-�#g�ccu��S�%��:]k�ܙ��4��A�C|�}r��X2\]��Lsp9E옢)�o>2\�C>8���Sa��	܉���p�w4��h]�߳����}Y�G&%�C#lU2ڰ=��M�Jdٰͭ�u���o�?bG����521	'�}]Ӏ6� ��,v�� |�Ӓ�NF���'"��l�:۹�w>�CTNkݛ�5���rE2�S�۰5�ŀnֹ�5ֹ��w�x%����۝�⦹yú�8N���z���]��2p�\Dk��}���r����u<����Ӏk�s�6� ׯ {��F��.eJ����^ɼ�8�LQ�z�G�Ϥ�7�nI�훒w>������މc��'"�h��^�^,?D�t�p��p���'$�nDĉ$�:���;�U�u}U�GDU{����v�K���M���.��7k\��BP��O����5�Ł�{������.9DN��m%n�l.�c��1��Z�ť�Ӌ�GU7��q����;}����D��$�_����h��hz�hϪ�����NF���'"��k��&nm�2�g�~�ٰͬ<�]N�%�j�*��� ׯ���%�cM�}��"|�(��"��cQIIB�%��"H���#R �@�
چC6G�7sVh�cH@R%&��}>b<i 28������5��«�!g�Y	߅�F� "	���X��
/Nø��"�(0^m������]r��!� ��� �L��x�4r��H����<:�3nh�}�P��
.�����:�5M=	��� ��#�r�'�x��X��&�6� bqUM|����O�b. � QB���S��pQׄpUt�v��}���]�'>ﵹ'=�e3�*h����U-�J#�B�y�V�oN y�^�X�hꨵ(���ʕuws�k�s�rJ'[��ϱ`m6���Zm�op��Ȣy4 �EƸq:�Hz�ƫ8��m�<5�S�`�4����� {u��^,��B�A�Zu�ښFGnDĉ$�:۹}	)��ٰ3kvl�{�Q2d��5&<X�1�E����u}V�}�f�׮��p|��@��ԋC��}o� 5��^�XI1!D/J�� X|��uLM
�}����g՗$��!�Iȴ��4��`m78��8�N`�W*B���Bc�I.�Ҽb��t���@v�y{D@�A�W(B�u69�ڦ��{zՁ��ՠu}V�}�f��z5��i�b�$�ԙ�s�o�ff$_;�o����Z�P�L����T�(e)s*S�������]��(�|��]Ӏo�Z���KDi9�C���}4붬ެɰ��+z����j겦FS��nh�n�=��`rQcݟ�f�mܒ}��[�q�=�q��2�aA*�E֔j&�2l����V\�VNe�]�\ε�4t7U�n�]����G.����6�,�SD���c<'WE�j�	�Ӥ�e��r3�[���y�͋���X��/\�"���=X�f�y��i:^�G�\�7;�cۤ�Ꞷ��[^��^ȉ;�-��CM���\d�'*;i�F�f��r:dtbT�6�{Ybm�q��cg�y�[�P���sA�(�w����t���p/�#&v����=��sf�Iwٹ���$�cp�³��$��_k�W&�CiG$�;��h_U�wY����@__M�c��MA�L�B$�@�Z� 5� ׮�����O�� ��	"NE���@:���1%��������-���\��&89$��W��@���u}V�}z���k��71ɒD7&���^���΍�ޟ�3���{=����ɑ�H��sm�n���p���@��4�F������6��6ƻMZ�t&��O�o����0�]��w�!B_H9������*��Ur]L���� y��%�Đ(Hx��L�ୠU��S���n��9^�@��� ��W��&�L�h[f���^��ڴ��h��jF$�b�ɡ�߳��U�����- ���䯽�}�u�ɨ8���C��]�@�g�]���}�M�����X�J&�d�lЎ�}�\�t�[ml����!�"�g��̋��ݹ� ��Ǒ'"� ����٠r�^��ڴ���
3���8�@:�4W��:�V�u�7�?$}���cs�$C�hz��]�gSAȀX��+�K��[�O}�kp�����&�,X���{�+��- ����٠r�^��g\f7�X�L�r����������d�mh]�@�>G
�y (��$����S�l���i2�����{\e��%���`/���ș�0RI�}�M��h]�@-�4E�5 69Q�7&��^ɽ���3kvlw5��1�DL�{���D��F�Z����[���&L��`n�l��YCs4ۑ!�Iȴ޳@:�4_U�������Dw*�+���U��W��4�l6*��on���?H����)$�����J7^l�6�f�3=���J#������vxAc�%r���.��y��`m�����ۥ�㴑&�͕9�NV��ث����N��� o]���������M)�dMX�NE�u}V�[�h�1�����9DDCf�H����I��v���`{������� ��*"d�i��M �l�-}V��ڴ=�3�b^���*=|5&4ҐQ�7&�k��ՠ��w���$l!����}e��]e�vy���:ky9�,���m��[u�f����t��z�RhkN{6�:+��ync˭���k�����ӥ-�W�s)mg��67`*��=���۳�`�ଂc�+���XYێ!L$.���q���������l�q��X�F�Eۅ$�Zm����^k �v3�4�D�۞g�g�F�:�SJb,��WKۖ\ɍ�^=����&���uv�K�yzZ���<8��(�5�"���y��#\v���ww�����2db#R/�>��- ����f�k�쵫�$�Hyr- �7x�]�u�pu�s�S&����Md�I$�@/����}V��S9��6��v��U�T���Ӫ������(��ޛz���=�d��f�w֤ҟ�D<�łr-]k� �7x�]�u�p�/Q���n�k�v6k<��э���tnP�װ$�����.�����M�}�/|g[H57s��^ k�x�k�]k� �����q�I4�Y�����ت%lt%FuwӀ>�Ӏl���6G��̎%!�1G$�>���:��O��ؕ]�= �������A�L�D�nl6B䢷�zl�� �{�W�h�kW$M�LH�r-��Ձ��"oo?�έ�=���(��~����T�Ӝ�j���c��|Q�ݯn-��^�ݷm�pD�:���'Yn�$����hW�h_U�r�נ^�c���$���@������$_;�U����f�w֤ҟ�D<��D����\�>n�!b�$�D%� �bA��*b �� ? �E��g��ܓ����rN�/dQUd�M�9��D�{v���hW�h_U��1̂�mԷ3-��g���\�g^���o-�ֽ�+�J�<N'<p�E�5ldO+����ޝ���{q����Mm���t)Hb�nH�����Z/�~�������@����%��L�MH�Z���~Q
ds�Հz_u`u�s�$�C��5�7!1"dIȴ
��z��^��߳�;�uw�@�>��Q5���]]����u�|�\���8��ؖ�Db�
F0P�(%,Q101H��F�!�T�D B�@�$�������:�Z�J�lm:�f�X:�8�����u�}:�`�	Z8ߕŖ����M��M���u7q
��PI�r�&lmP!x�Mc��G�omk�g�� �u��P���S��7L��1�d�1��@�e}|���_y�:�8���~Q
&M�}2��EYUN���t���sv��^ɳ�DB��Vl�u��9�JL��!�1�#�����Ӏk�Ӏk�s��%>��X�~��&F&�N-�}V�u�4����nI�g}w$�Jp�"�S <D��K��t��J@�U��0�;G̼�$�&�41u�fpMT�'�h�� H	#>��kPI! �?
�ba�M�#��ҳ���F@�ޝ��IM��D��B0�шC�{h�z
K�8�G���a$Ϟ�1!M	]<��6lM�'��:�Dڃ�iz�&
�kbf��e�i�RB,`$nq �ʮ��@�L�F!'~S�RO� .MX����z�P���~@�G�^��AᡈY�48w}ߵmֵ&�m����@��ְ$i�gK8��N-��m�'Y^��5B��^�zNu��X6�2d�A� �*�;Z1��q-䳡6�u�gP���UXr&�&�u*�����r�/����m	@��MәZ60��f�vƸ�Ge��ŵB�g��k$��r�u8Q9Ӊ���+��p`	E�&�6Ch�lZ������g%��z��룳�ۃ�d��>����2��k�W���R{GT�n�a�MW=8ҷUV�¯I�A2sh��šg��˖0�A�_%��jf�r�tg�=8CQ1F��A�������U���+ղ�D�;Y�^x�we�C�)�M�m��N���.�{tof��ɖ1�I�s��1;7$WY0ܓäݦ�\bu���Ą�,账��nMv��ͪ$�;��1��į)�{;�hӮ����ݺ�ۂ�QMź������]�[s�k��4�)ԫ[�35�a����]�ݐC�=O�^V�un�r��F���+�L%�!�/f[�m�b�cŪj�8�c�
��y�8��6{nƆ�b��H
À'�vw���ʀer�OF9����\3C�Z���Ax�V���um�<�@j%�C�(q��(d}�t�<��˳` �t۴kvwEZ��s�*�ɖ�6�㫝0n,ƹ)��3�՝=�ͽ��;T� �2lrݪ1WUgv�ds���(�x��wd"�������v�IL�6Z�j_.�KН��a	���lP�ũą#VW4�f���Z"�M�d�c^�Y�A�[�v�m�.��yt�7@*<���Fu�է`��i�3ngGl+Hkay��Iu������̜iZ��5t��&W�N����k�\�GF�����n6�0mgxFYм����|�z�$���W��ı���e�X	඙�\����q��m����[�;vg�
�0qʷ�ٔ�]� kR[u��.��4�(����4y��5�^����(xwA����#@�P�A0�/���p��j�52L��&h�h��\-%�m�Ț2�+'Qm�������c*8I�Q��݄/��]�q�ې�,K��b�*�H�ۭ)�n��c���'����`:�N4���Z�0t��n���Y�Ju��x�a�ݱ�66����d\�]=��@)��._�ݳ�7��.�b�JK֟f�8]i�UZqOkm�Mi��lq[�p��w{��{ϻ�̪�*��Twr�۳� u�+M�@S�$��Ξ��鳞��×W5�"&D���w�f���נu}W���˔$����6,�]L�uR�T�۫��m������� ׮�P�>�F��cX��&H���ZWj���}}4�ޚ�։�~YD%J&�� �M� k�x����a�K�ZSߘ��2a܉Š���BJsw_�=���=��6�D{�oϟ�WQ�����p݁E[:�%�ks�'.��nx}<n����{���}�q�sf�I4��{��f<,efOBQ�@�ޚG��Q�M�Q�7&�����$R��$�M� o�� ����2\~�#S#��/����٠m���h��#M��2$�Z�l����e4=���}=�}��~q%Y�G$����ݜ|�� �n�� h�a��ra�i�<`u�v�����s�=b��p8��͓]��UmT���i�������k�� �w]~J����wq4)�dm(,_�p�:�V����@:�4���$Ze��=�2a�ȜZӻ�`��g�>��.�%IRT�)B b8f��znI�g}w$���2�����t�R�N�9$�BS9����ǥ��ɰԣ�W�wU��v�L���S��(��wJh]�@�Vנm��xn�cck"��"N�j�s	�4j�OKe�������E��ﯞ���1�����$?��~��?���[g���x����di�"�"NE�NfU�DDL�n�31�`{+2o�O��~q%Y�#����4��:�V����@���f4��H������]78�۬���j���([����ۺM�S�%̩��e��v� ��x�n�ݶ`[��ba��<�|��[R�Y���]7C�o	�>\�n��-��4�N�����n�����l�5��{{�T��R8F�#�@>�f��g�H���{5�`g�ޥT�D�i�8)�������c��P�d�� �o��_�U�&�Jdbdn-~]}�4�}4�h{?+��Z���m�	M7T�`fc�6D�7_�3+vl��ay(�R/"e�I��+q�]��3Өˆ)�����n��y1��\�N̥��6�!r-F�!,��J7Ab6ݑ1s��l�T��Ϊ}3=�]��6l�pܾj�<�E�=oJ�#���hppZ��&��=�.C���ɮk����J�۶엌�5ٸgXj��S1�<h�-�v�3����c��$���J���:�ۃ1�VP!���ߝ���kѷ}tpb�jІ;L��j��B�ڶ��<�#�˲�<E&lY���`4�s	����4�j�>�)����4��X�1�I�C�h���=�ـm� {[��!B�Ϧjf~YK�ȴ��4��i�H��M�����e�1�I��l��@<�� {[�}M�N��0}�+Lj)#FI�u�@�v��ǅ�}������d�l��IU2��Τ��z禺Iw�d�;@R�]�XVu�p@r4��ӟ�D����-�f>���u��'kd��i�rk3WrO��zoA���`T"�b">�J!�%|�� �x�78��\���ǒ7!�[f�}ֻ9D.�ݮ�3y�`|�β�̍P��ɠu�@�v���h�cX�d�9��9&���Z�e4�l��٠Z�ʑ&<JI-�luvp���s����& k�v��n6�k�����D�s"K�ȴ��h�٠u�@�v���Lcؓ".�T]՘������7[ŀ{l����R��BG�I&�}���;�{f�: ��q`�`�%�!B����ݳ >z� <����I�pNM�����h�l��*�H�#"�4k�`�w��� �o�^hͬ`�'Tvr7��s�yF������I<�r�~�,4N���Mӆ�c�����m�׀�� �7� ��f���]����s���l������}2��ƀw���fg�H���cX�L��)�`g�mX�$/c̛���$)!IｭD�Kı/}�kiȖ%�b�ٌ�� StML�C�����&�I���wM��B����;��
�RB�,K�{��r%�`|x�ČdF�B�TS�=y�o�&�X�%���ޙ�ɢk!��\��r%�bX����q,KĽ����"X�%���l��Kı;�{�iȖ%��{�ǿ߅��b7L4���A1�[��m=�]/K��E�֞rW�`����?_|nvY%��H:l���$)!I
sw]��AbX�'g��q,K���]��	>��,K���j&�X�%�}'��SN[��K�n�~!I
HRB�kq,K���]�"X�%�{�kQ7ı,K�{��r'�.TȖ%[(��S4�Թ��j�Y
HRB�~���iȖ%�b^���Mı,K������bX�'g��q,Kľ���ə�[%0չ�]�"X�ʙ罬�M�̩�3*g}�ki��2&eL��n�M�̩�?"�Z������>�s��{��~J�ˬ���0���S"fT������dLʙ�^ݘ���S"fT��]��Tș�2%�{Y����S"fT�� !�o��):�F�\��vC�p莟�Lﰚ�C����ݝ�:�N����j�nX'�t�(�d"@ql��,O1��wn�c�%�ѡws	 U�[����g:c�3U�h�Ѵ4X�l�\c�Ws+�\�\d�x�u�v�����tng�w	5װ��d�+e�Zmi9,g�/ظx^:x�$�4��g�V;0�J�=�[��B�fd�eeְF
&�?8��}��s��ʳ͒�N�}�ɲ��b�-��v5=a2���<m+!�=-YS�wU5ve��k�ߪdLʙ���ى���2&eN�~��}�L��S"\�����O�~���ș�3������}S"fT�����k�P��v�ϻ��S��veN�~��}�L��S"\�������2&eL��m>��D̩�=5�ى����7P�
�af6�GΦ��B�nsWi��2&eL�s��f�n&eL��S;�{[O��������n'������Lʙ2����]��Tș�2&e�vEͩ��Lǻ��S��r�����ki��2&eL��n�M�̩�3*w�����dLʙ罬�M�̩�T��3�CR��)�����L*!VTȞ�����Lʙ2��?�������i�Tș�2%���f�n&eL��S;�{[O���3*dK��!�R�R��v)��zy��8&��Jw`�2c�</]���#�7N.�������=��-N�~��}�L��S"\�������2&eL��m>��D̩�=5�ى����{��?����NZ�z�����&D̩�.{��T�* �A^� #�T�h��p�u92�s����}S"fTȞ�����Lʙ2�}�z�>��� j����s��|Ve�i�w�ܢdLʙ�߿ki��2&eL��n�M�̩�3*w�����dLʙ罬���{��;ܧ������r�;��]&mki��2&e��Q?M�嘛��S"fT����v�}S"fTȗ=�f�n&eL��S;�{[O���3*dK�{V屠��
���P��U0��U0���6�}S"fTȗ=�f�n&eL��S;�{[O���3*dOM{vbn&eL��{�{�߿��������q�I��ۣ����9�װd���g�8�6�w:��k!��\��w�2&eL�s��f�n&eL��S���6�}S"fTȞ�����Lʙ2�}�z�>��D̩�3/}fr.���@3ﷹOs��{�����O���3*dOeצbn&eL��S�߽v�}S"fTȗ=�f�n&eL���^f{�R��)�%�p��aQ
��D�]zf&�fTș�;���i��21�A�p��a>��ؼ��hVP"ЌP�YIm�*T�!	H�#VI$B$XcC_nP�# �	q�+A�|��O�ͤ�Ө�H;	_���6$�@ۡ�M�%j�)�����"�@��.�w�a"1#!���A��78~]B @����p�Nf�,����e&m!�JP�u8��	W�#�ґH�BWIH�A�!;��B�n
�G�!��hE6�D:���\ C�}��}~Tb"�4DA��*pO �@�jn%�}��M�̩�3*w���ӟTș�2&�.{4[���F��Y�����S"fT��]��Tș�2&g��j��fTș�;�{�i��2&eL��]{.&�fTș�=�g�թ��=G����=��)�w�?*<n&eL��S���6�}S"fTȞ�ײ�n&eL��S�߽v�}S"fT����w��TD�ӝ��C�\�8���F�ۉ�0t�:n۶츳/���(�e֥���kU92�D̩�߿|m>��D̩�=5�[����2&eN�~��~ g{SQ3*dL�ߵ�T�Lʙ2�����//빬�5������s��{���׭��Lʙ2�}�z�>��D̩�3=�kU72�D̩�{�O���ܧ������{=V6�@���3*dLʝ�����2�D����T�Lʙ2�}�|m>��D̩�=4�f�YR��Bd*���-�I�jU6U�fkW5v�}S"f^�5Z��Yq,K���߸m9ı,N��Ҧ�X�P�R�V��)�ʜ�&~��]�"X�%�^����5���\���&�X�%��{�6��bX����]��9ı,O~���iȖ%�bw=�dMı,K��=-�MaXz�����A��3�Θ��oN�{ ���[ul����-憩�$Jw�����bX��ץMı,K�׽v��bX�'s��D�Kı;�{�ӑ,K���~s�x�H]cc����D�;�{�i�~9"X��ߵ�7ı,O~���ӑ,K�﮽*YT$�L*!I|�֪ln��R�UZ��r%�bX��ߵ�7ı,N����K�2&D��Ҧ�X�%���f�~!I
HRB��T�uS5BuN��Lֲ&�X�%��{�6��bX�'g�鉸�%�bw���ӑ,K��f:!Y
HRB�}麥U�*l��M���iȖ%�bw�^�7ı,? �߷���}ı,O~��"n%�bX����iȖ%�`�����$x�b�*��M#@�Ԟ��L���ݝ]Q��>��nA�w70nMT�[�L�� ���bt�
���ݫ��5\a������j�z�l�+d�u.�L�˻�+dy����7������^��;U��;q�����{#�¶N�A��ݙò��,�n��nF���r��-��Oc��sՓ0���HS�\Ͱ�y9��7"�Y�"U��7lc��m7{�{���mYu���5�mWo&����:�2x�'mfєT�vlm73S#��l�T�l�XB������~�ND�,K��l���%�bw���"X�%���zbn%�bX��<Yf���jfc��\��r%�bX���dMı,K���m9ı,N�k�q,K���]�"X�%�{��yT��GFk����7���{�����"X�%���zbn%�bX�����Kı;�fț�bX�'p�cs)��KL-����$):����LMı,Kߵ���r%�bX���dMı,K���m9ı�{�9��?�a$.�����{��7���}v��bX�'}��q,K���ND�,K������%��w����p��V�Rw�%�K"-˧G,W9�f*E��u����{tȏKsZ�������r%�bX���dMı,K��m9ı,N��҇����,Kߵ��iȖ%�b_޿��4\�k3Y-�kZ"n%�bX��}�i�j�h(D1 ��j%��]zT�Kı;�{�iȖ%�bw�͑7ı,Ow�y�e�Z�0�h��ND�,K������%�bw��ӑ, 0ș߿fț�bX�&no�p���$)!f<s528)6�F]jT�Kı;�w�iȖ%�bw�͑7ı,N����Kı;�J��bX�'{6�s!����2kY���Kı;�fț�bX�'���m9ı,N�Y�Sq,K���x\/�)!I
EzqӪ�n)���Ocra��ce<6�Ev��h����s�ƃu�M��<��e#5�����oq�������Kı;�g�Mı,K��~��ϢdK���ٲ&�X�%!z��ne5M����ڸ_�RB���kڱ7�	��,N�׿]�"X�%��߳dMı,K�{�6���ܞ�{�������c	!u�ow�,K���{��r%�bX���dMı����#�:A�b����D�'��6��bX�'�kڻ����oq�ߟ�_��T��V>ND�,�@Ȟ��8D�Kı=�߸m9ı,N�^Չ��%�b}�w�iȖ%�b_w�lѢ�CY��n�Z�q,K�����"X�%��kڱ7ı,O����9ı,OfU����$)!jJ��5 Q���k�mɆ�.nv3vKz�ٷK�\v5���R#��X{V=����n��n�{���7���x��~Չ��%�b}�w�iȖ%�bw�͑7ı,N��p�r%�bX�ǎf�G&� �SnHVB�����k��NC���,O~��"n%�bX����6��bX�'}�j��O��L�b{���p�5���d˚�ND�,K߿fț�bX�'~��m9��2&D��~Չ��%�bw����97���{���ߏ(�t�K��ow�,K?@Ȟ���ND�,Kߵ�V&�X�%����]�"X��B�> ���p�8(hR��'=�h�d)!I
HYG��r'Ce9E0r�Fӑ,K���X��bX�'��}v��bX�'}��q,K�����"X�%�};.zY�,�.�bz[�:�n(rz�j�b����l�]<k(�}�E��/�\H]c����oq����]�"X�%��{6D�Kı;���iȖ%�bw���Mı,K��_ֳ2����ff�ӑ,K�｛"n%�bX�����Kı;�{V&�X�%����]�"X�%�}��CV��pM]��oq������=�ND�,K�׵bn%��!�2'k߮ӑ,K���ٲ&�X�%�Ͻw�f_d3E�3Z5sFӑ,K���X��bX�'��}v��bX�'}��q,K�Ȟ���NG��7������5���ny��﷋ı>����Kİ�
1����'"X�%�����iȖ%�bw���Mı,K������aD���{_1I����y�6c���أ��k]W���K��q��Ugf3=�Z:�Kd�rY��&7f��M�h��dI�U�M2:4�ۖL�vs�]�ݹ�^scl:۳�)�<�d�Z^7����F�"�������.�J�:����b�	��ج�K�<솽!.MR���,����}2�ӡ�gT�lF�H�� �ir�t�5��',o{���{�ݸ���ba��<�=�G7j\Y��=7UvD�]��i����A���jq��k+�������bX�'����q,K���������%�b{��j���NDȖ%���6n����$)��j�*\��R�Lֈ��bX�'~��m9Ȅr&D�=�_�bn%�bX���~�ND�,K��l���%�bw'��j�Fh��5&�֍�"X�%�{�kQ7ı,O����9ı,N�ٲ&�X�%�߽�ND�,K��.{5e��-ѩIsZ���%�b}�w�iȖ%�bw�͑7ı,N��p�r%�bX����q,K��ƽ�ɭk3)�h��fj�9ı,N��Ҧ�X�%�߽�ND�,K��kQ7ı,O����9ı,��I����=�Bm�7[PO=F�`θ�t�"8ܻ.ys�RfŞݞ1�����ǻ��7����{�6��bX�'�׵bn%�bX�{]��r%�bX��ץMı,K�z�0̾�f�a��j捧"X�%��z{V&���SQ5����m9ı,Oz�Ҧ�X�%���ND��S"X���ڷ-�r��հ�Z�Չ��%�b~����r%�bX��ץMı,K���m9ı,O��ڱ7ı,O{Э��,�ѕ�5��r%�bX��ץMı,K���m9ı,O��ڱ7İ?*�7~�_�RB���'�U5.Zt;�F�Zԩ��%�b{���"X�%��z{V&�X�%�����r%�bX��ץMı,K�~=g�f����^YԖ��Uz`�e/���b3����
μu�	�V���'-�������x�,N���V&�X�%�����r%�bX��ץ��$Ow��n	 �U�u�'�4�AF~�������n'�X�'{u�Sq,K��}�ND�,K����Mı,K����%z:�)��7���{����K�	��%�b{���"X��V@倄j4A�R�ȧȦ����Ng�ڱ7ı,Ow]��r%�bX���SY�2ᩙ�Ku��J��bX�'��p�r%�bX�g��bn%�bX����K���Ȟ���Sq,K��}w�f_���0֍\Ѵ�Kı>�Oj��Kİ� �����v�D�,K޺�*n%�bX���iȖ%�b}�fY��d�Z��c�ղny���-Y�v��v���i�0g�ЍP!�6�=Z���Kı=�{�iȖ%�bw�^�7ı,Ow���Kı>�Oj��Kı=�B�_p�3FVܷZ�ND�,K������%�b{���"X�%���{V&�X�%��{�ͧ"~T��,K���2d˫�Y5rh�kZ�7ı,O{��ND�,K�h��Mı,K����ND�,K������%�bw'{�MSE�˨[�5.�m9ı,O��ڱ7ı,O���m9ı,N��Ҧ�X���8,`�D���؟��ߍ����oq�����������b&�X�%��{�ͧ"X�%���zT�Kı;�{�ӑ,K���=�q,K���I��շYr��ֵB�#s���u�N�ٮ89AO"xH��b7��8R�%z:↟����7���{����Ǎı,K��{6��bX�'���X�șı;��~ͧ"X�%�~�~�T�Y�Kc����oq���｛ND�,K�h��Mı,K����ND�,K������%�b}�����j�kVkZ�ND�,K����Mı,K���6��bX�'{u�Sq,K��{�M�"X�%��?��Fp��=Z���{��7��ߵ�]�"X�%���zT�Kı9���iȖ%�b}��Չ��%�bw��m��3FVܷZ�ND�,K������%�bs��ӑ,K��==�q,K����ӑ,K��TN���}��1<|G����%s_���TB M�	kd$(�3�Pǜ�ޤ!�,�h�}�/��A1��8��4�&�WHh�*ȠBOUd	���yC灨��w�@��G�A�>R�c�~��+*�'@xl�aхO���t^�!�"���w9�4�A]�X�$�8�͉�
0!򤳫�A���7�"��R��Ô�%�a�,�+���H�����mֵ#m�� H8p�*�]U*�K�;�Q�f��-��.d([8�[x�E�8�;����>{b-�q<r��Gn:�:ܛ����R���4�Cdݕ��K+��@2m.�켭Gm��m�ʮ�b"%�P�[�[ٮ���۠��וpZk�N}�t
��F{z�v�.5Z�y�!��:+��ݞ�f�4�2l���p�<�J�h�^��1D�=4�c�=-Ɲr��S��a�瞗����:�`54���AE�£�'2��4]kdy�Y�=�,��ԫ6�j�4�]
<��Kf�[��z����[��b�Ѱv�t;��*h-���c�X�h�j���Tp}b'���on���0W5�xt�L=�]�u�k�c�7EQ���kv�u0Nх�U.�⃇mqHq�mmm:s����ڻ�/c;h;]�)�H;�d�G�l��e6	���$�x��ѵ�vMs�۰5�1n9��ʙ�^��C�O<���i:6D��k���[v���/*�U_9�_��U����l�*V���{/�����u���;1�ke%]�٠�vh�ri����{��m��Y[���R��3�� �8ki8������R��	�#3�u���s�"5�Z�F��͈;��{���=2';���,"ݛXnn\rq��V���kj�N�K�0���ا��d>D\q�snU��]�^����v�1f�X5ѻv��U��1��٭�6Ȭ:�-R�v,u
K64�J��+�U-��`��Ђ��˗cX�)~K�}1ɎUCC�u]��m��|UZ��$�n7e�v�ȯ0�>ѹ�u�����X���WUT��\��L ��ٺ���ZIz+e��l�E�QS���H!^��gf����}>6����k���Yϋo!d���^n�O�����j���c�����Wgtp�#�l��
K�W���V�(E����+[cM�X���X�]-fN!�=�ū;P5p�.��c��љ4����(AD��Q��(&A��퀴A�ȥ`ᇅ���,>h��΋��۞/��&I�'Ltp��D�9ڡPK�tZ]v�����z���]+ϴ����;;7:6���i'gh�?~��~+qA�`:���6\V�ni^L��V�{c�˻��ϑ3����&"!9��2����>�;M��j�Ma����랕�D-�݅�q�:���Ͷ׶ᡠb�Ǜ]��յeF��k���v���v뵥�Iج/c�h6�{�b��@3�'�3j�e��V�f�����8�݂CN�F�#�Oa�'XY��JeΧN��52�m�ai
HRB����p�ı,O��ڱ7ı,N����9ı,N��Ҧ�X�%���pԺ�b�aN[.����$/�r&�X�%���}�ND�,K������%�bs�ߦӑ?���,K��[NIi��$$�$+!I
HRB��?fӑ,K��n�*n%��Dȟ{��6��bX�'s���q,Kǿ�����uW�?{���oq�����zT�Kı9���iȖ%�b}��Չ��%�bs;�fӑ,K�q���N�����ǻ��7���x�{�M�"X�%��=���V'"X�%��{߳iȖ%�bw�^�7Ǎ�7��������Y�<(��l��,sn���%�B=�y�I����EyeL��d�jm9ı,K��k"n%�bX���ٴ�Kı=�J��bX�';��m9ı,w^չ.��sZ�d��5�ț�bX�'3��m98?5��X	I�1 ��S��(/q@�W�5���ʛ�bX�'w~�ND�,K�{�ț�� L��,O{Ь��Mf���f��ND�,K��Ҧ�X�%���~�ND�,K�{�ț�bX�'3��m9ı,K�g�&L�]���tkZ֥Mı,�2'��?M�"X�%��ߵ�7ı,Ng{��r%��KJ!n��0��$)!I(��N)ԙ����5u���Kı=������%�bs;�fӑ,K����*n%�bX��w��Kı=��!����l�7%s�燰eS�����e�'�G�5�ܼ�a1t����g{���ı9��iȖ%�b{�^�7ı,Nw���~V}"X�'�?k����$)!{6K��M̶ښC��k6��bX�'�u�Sp�
ș������Kı?a���&�X�%���}�ND��eL�b^��]L�2��d�Z�ԩ��%�b}�o��r%�bX����D�K_��G᪃��`�� 4�D��^"�X�D�{�iȖ%�bw���Sq,K����S3ٗ&�a��Y.�6��bX�'����7ı,Ng{��r%�bX��ץMı,K���7��oq�������!x�p�=��17ı,Ng{��r%�bX�����S�,K������Kı/������%�bs>�񙑚�F\�əq�qy��]��g�c��í��p�1\���-����B�]���h��&kY��%�bX��]~�7ı,Nw���r%�bX����D�Kı9��iȖ%�b_���s�.��UX�}����ow;��m9�c�2%�Oߵ�7ı,O����ND�,K޺����%����=�T�S�
r�p���"X����D�Kı9��iȖ?�C"dO߮�J��bX�'���M�"�oq���~<��e�X�,�w�ŉg� 02'���fӑ,K����l���%�bs�ߦӑ,K�+�P��*�P%"�U(;A�Nn'�=�dMı,K�훹|kR�Z��5�5��r%�bX���dMı,K�#����i�Kı?a���&�X�%���}�ND�,K����좙����:3œ�gE��h��`��t�m�v��_kI()ӮG��
�����,K���6��bX�'����7ı,Ng{��r%�bX���ʛ�bX�'>��̹53.��5���Kı=����� r&D�>�{�m9ı,O߯�7ı,Nw����B�aQ
E�e��9��d�h�k"n%�bX�g��6��bX�'�}���X� �ș�{�ӑ,K�����ț�bX�'{�VK���[d�k6��bX�'�}���X�%���~�ND�,K�{�ț�bX�'3��m9ı,K�g�&L�]Ԛ�tkZ�7ı,Nw���r%�bXh��Y�,K��=�ٴ�Kı=�fț�bX�'@B�o{������aC=�	L��8���s<�n�m
�&�V����v��k.pl�+�`�`�+�b7u�;��N	�9ڜP������,�����Mשx��ʖ^d���\[��<q����"�C�ʷ��blD�ڱ���+\��%�f�������krl�x*�҇Uқ�q�@ݬ&a4ʘ�s�'k�kSY��Xfuq�Z�DJ������L��%Ԧ]M�4[$�,�n�q�ʽ�7��k�e@���][r���7��Tɖ��/�)!I
H[Ku�
�R%�bs;�fӑ,K����"n%�bX��w��Kı/�as٫5��]��3Yq,K��w�ͧ!��S��RB��B����$/n�"X�%��=�dM��Qʙ�_{6O�R�%�Ji������$)!H��~͑7ı,Nw���r%�bX����D�Kı9��iȖ%�w��?��ӮG��
�����7���';��m9ı,Oa�k"n%�bX���ٴ�K��
���D���ψ��bX�'}���e��MK�Zɚ��r%�bX��=뉸�%�bs;�fӑ,K����T�Kı9���i���{��7���߇~#jˠm��Ս��wcM�	۵vnfw�i�u�Jv\rλ�(�I�W5�u-�d֮&�X�%���}�ND�,K޾�Sq,K��{�M�"X�%��޸��bX�'~�d$�ᩬѕ�LֳiȖ%�b{��*n"���S��n%��s�ӑ,K���~�q7ı,Ng{��r{��7��������umv�����Kı9���iȖ%�b{,��&�X� ș���fӑ,K�����Sq,K��u;�3N]3R�I����r%�g�"~՟�\Mı,K���fӑ,K����*n%�bX�ϻ��r%�bX�ǰ��kZ��K�����q7ı,Ng��m9ı,?���w�T�Kı>���m9ı,OL=뉸�%�bS�z�_d��N֍Z<�.�K���;uө�f�н��{`���fm�Еb����?{���o%��]zT�Kı9�wٴ�Kı=�{���蚉bX��~�ͧ�{����{��??�u����Kc��X�%��w߳iȖ%�b{,��&�X�%����ͧ"X�%��]zT�Kı9���̾�MK�Z�k5�ND�,K�g�q7ı,Ng��m9���1Q�Jx�@(�K�q6�����p�GÊ�"����v��Sq,K��{�ͧ"X�%���r�̓W)�̚aM��B����*!o�vn���K��Ҧ�X�%����ͧ"X�%�釽q7ı,O��d$��u�1�ۚ�ND�,K޺����%�b{;�fӑ,K��{��n%�bX��^��r%�bX�z{7n]hɭN��p�J�T����.��ݷ=Ū�s�ƃu�2~����I�j�,��/��{��X�'���fӑ,K��{��n%�bX��^��3�ı;������B�������TɖN�\/�)ı=0��&�X�%���]�"X�%��]zT�Kı=��iȗ{��7���Ǐɭ6xz�C��{�K�﻿M�"X�%��]zT�K�"{?{�m9ı,O�߮&�X�%�ϻ�-浒�ZMY����K��U��?~��*n%�bX�����ND�,K�z�n%�`x���*'��c4��Q4�"�İT<"� FD�����r{��7������㮸t�[�X�%���}�ND�-�a�]�;�����c�������*
��%�P:b���tm��'Z١��u�n993��0��{=r�M�ǊFI��=�u�M���:��@�X�Ƃ&�6�r-�Jh�����z\Z�٘�z���)1��4�4[���z���V��YM �j`��!Z��� ��u�9ѹ�7�فВQ���Ɓ�e~d��D���q�p�������O� ��u�5ڣ菦|BK��n[�()R�CCd��Li�%l�c��ZΝWf�s���Œ'��[��(�t��p���NΨ�����c�e�۲V����s��D�tqKY�N��J�U�t���6��z����$��ˋ����]2)���ۆW��Xk=�77hS������=<��w!�r�;{0pظ�U�Kj%&�nʂ����w328ͺt���h���[�I�{����ϣ"!E�|O�)j��t�t��,)9h�u:zD��Y�%�㧦�+�u���&�ӕ:�v�AF��D���[)�^�����߿�yS�Z�|��F)#ŏ�p�/[fr�6[��:Y�8�M� }�r��H��I��|���*�ՠs�h�����5����ǊG�@��s�}���i��舝���޹�cAYd��$Z�;V�yڴ�uz\Z�����6��&��9�lv�ݙ�nr�f�nr��ƹ�=<9�c�e�ob���7�I���P�����@7�ܴ��A�52B �����$�����W�F@�_�O�B�K�8|� ��s�=��:"d�C�2~S"j	@n8�*{�@��j�/;V�w�� �n+$�H�<�62\�u�p�������z��8�BS���<#mŠ^v� ﭚ\Z����� �"Ĉ񐤝��A
ɞ��ft�%�2#��ys�D�=�<&ŒC�BN7 ﭚ\Z����ՠ}��c���ǊH7&�W�������>]�����h�YmLO$$Z�;V�z��s��ؙ$C)�t'pbu8��/4KG�'��a7f�;�6�R�@�b�`��uBB�c��A��ω]	��x��=&_	��S������8��]�EF`I@@�CCr�w�J#��>}�hʑ��Y�H&4V'MPC�`c�|h	/9�S��ܛ��a���#�H�C���XZ���y�m:�!Cf�h
|���<r1
I��x�|��}8��U���A<K�X������²���7��B����4*�%Q4�,N��PA� >PNx؇؇ �lP��u��AXB! ��v+�b�� �&!&�Q�w�r��6t}8֤�،NchĚqh{�~^��+|�
�̛P�O��f�77eR��KM�CUwV�N�΍���s�=o�s��]��^yo��OT�f�/G]u�kn��
θ��Ci�x��U�� �F� �i�����D%�+|���b~�'#��D�����ՠ^�s@�wW�Uū}�:�	Odj9&,�Fۋ@�����@��V��}V�}X��X��q�h������u�p9
JQ$B��D�~�(?��&ԊkQ t%
h+ 
$jE�
 �t� ? �s�s�rO}�e3��\����$�@��V��}V�z�h}l�=�{�h���iBG�#��s������{=��wk=n6���ڧ,!rhk#i���H���;�^���[6!DG��7f��� �ڰSMUH�jí�ǅ��C=���7f��U����z�Ɇ7� L&9$4��4
��hW�h����3�s�I#��(����y��Zy�-����h�qY$R(<r6�I8��� ��0N�΍��a"�JH4�B�n�x���V=s�U�sϬ,$��% �ڭ��L���p]p�:��ۉ��[������i���	�\oA�yjIL�)w+���]��듫Z�7(r�Q�I����λZLʷhQZl���r�����%���>���ۮ����<;��N����\�B�gz���۶��e�άk]s�����:��s%�Z"X��-��5��J@��r����?��<���L�MK.��fk ]��]�<�|Qv��*��k!ȃ�;�Gӷ��PI̍I$Ǔ�q������˺��-_������w���1'��!'����@��V���ՠ^����ލc�b�x�H��T�Z�;V�~��˺���]��5���7�-���@�YM��^�WV��v �W��8�0��Z��h.��
���v� ���Ʈ&H����[���6�Dv�;�l�c��h�m�M�ے�[$!�n(�a1�!�|���/<��v��e4��q�b��kX\љ��nI���]�R!Q�"XS����(�s|���I����nI��@.[��"�A㑶�8��v��e4��h�uZ^BR�jI&<�Fۋ@�YM ﭚ�V��W�l��m�53P�-�3������8�k���0�	F�w�߹�<��Ӝ���>��ر�Ǜ�㭱�YƜ�AݹIZ;$��!�x�5w��>�ε� ���n����<�Pi����qhW�h�)���@����H�q#^�'�!]�� ���n�����HI	/�A�v�At�b=�~���rN���@/֦܍�a1�!���@���>���/�S@��q�bi��KEKn��R�M��#��g��~4��h1\
\�#Ȟ'~#�����ʘ�]]�^�`���a룲�r�xf�9mc�@���@�YM ﭚ�V��R䑩$Ǔ�qh�ـ�� {K\�u�pޖ�<����JF���@�������h}cXک�!��$�@�p:�8��05�"�D@H@d$$X�^ �� ������{f�եpy�4�Cl���<�\���|� {�x�-s�rP����޲����)�..6\!	�sr7����a��@;a�؆�X��7W? �� o����s���>� ��&܉��1��h}l�>T�8�k�|�,�I%&��:��FI#�0�@���hs���J������-�c�d�c��1Šyֹ�7����w�zY�p�9��F��L#mŠw��h}l�>^��ܓ�g}w$�O����
E"�����w��?����[w���{|��\0OO�қf��Mn0dk�M��qgB�U���tc����ׂl�Z.u�����N��n�b���Ɨ�� �,k=ض3mu	�3�6�\�:�,�Ն�d;Oc�5����m������Bj5k��i�n0��c���f�1Ju����=��˸G�;-�٬3�mj�
�j�x����cv���hm�O9t>�~�����{��}�������?�E?��^֌�i'�K��;=�μlLvǣ\n۰�2�u,���dn4��L����hW�V��}V��[��}��cj�����nM���u�p�x�|��mL�)2�7�&8������ ﭚ��U�U�+����qh�x�|��t���Z� �74
�61L	$����@��uZ��M��ٖ�℣���3�K%�|�q��i�nѹU��oj�[�{^Ȇ0����ۗ��#�5��H�L�����>���?{2֨��� g�]�b�S��(nd�k2̙��'����<lE�@#�G�UH�A�'k���'{���$��w�@;�ܒ5$�����?��� ﭚˎ�@���@>����ğ��i'$����@�q�hW�h�n���Z��mA�8�rh.:�ε���� 7���"�BP�p��=�ۭ������e��&�p]��wmc6x6NI��ѷ�9���I��f?�o���p��X�n���`u�A36~E���z�� ﭚ�2���Z����f��I&h~���'���� 8��!  �<�(����Ӏk� �N�wvIj������ z�3 �ֹ��� >�f�v[���PX�q9��>��h[ŀkw�=v��~�Q�ssE~�\��ѫG!���{1��{q���W,Sl:q��YV�B�B$�8j�l��N}ذ�n���0mk� ���O�n4��L��o��H�fi�}Ϫ�/[��wu{F�ǎ5��i����fu�X��x��W �i5��CCغ��z�ۛ�Nw�����!�뉅K�R�%K�������$��pL��1WW8�l�����L�=��p�����w���1��n��g��	�ӐX��lwOTV6��yx�n����v��jE���π<�� {Lf�s�>��ץ��Z����1�
m����Ď��h�O�YM�G����' ��#�BW|����?��hΔ��T�I�Ls�q`tD$�{��u�,v���Ss�יXA?Ѹ�D�C@�����~^zn��d����XȄ�IDDH��_�E W�� �P � U�� W�
 ��@
 ���)H� �
�1��@ � �`�"("("(
�1EH"�0E"�1TF
�0@V"�1D�Q ��Q"�0E� �A�� ?�� *��@ U�� W� �T ^* ��� 
�� *��� ��
 ��� 
�� U� U�ي
�2��)A��'��@���9�>���  �    �    �          t7��A(D�P��T���*�U@"�*���@  J���"BD��(
 
� (P	DR� P
()U�    X       � �'e @ $A�  �
gp �%4���n��G=�۟{��Ӿ;�� ���ޕ�ܚ�`A�^�v�W��:�����7�Ω{� �*���_x�۪{;������    �W �ާӗz������x���}�OW� �^�弚��Ӫ����Խ8 =wz��      }��Ws����=R�}�_U�}ޗ��ǽ�N]�ۭ���J���N����U��ͽKx >� (� �@  4=/��NMTŮڹ���[�V�� ���������۽�O�ŕ�p����K���K������,�''^ڸ ���|�{����g�K����6�=���]���o�{��NM��*� �� ��   ��O��:�qgZr˯��Ҙ@Y��w��m>�g�]�s��=Η� )ν7}����g^ ��:q �B� b=so�n,�{� 7SӓR��_/����w��� �   
 �
b ϥY��\[�ӯ6�R� nW�'Je����S��Ħ�� `Q� ��  �� 1= A�PFv tPY�@M  )�4�F@
�����4@4� ������T @����iR�� '�UJ��!���"{J��UC#����)�R�  ���(�C�7������Կ�d|��EqS330��N>v��\| ����
�*�"����
���
��" *�T?�?�����n�g�s�S���9�C�y�8±��E�� F�
��b˞�3���F^���Λ��Ox����bHHFF@����|1 � 1Y���1+�������X��%L ԋ� F4��cp�0�	hEhC�79<�7�2I���װ�N���
c�D�@H�� t���B�I��l*D�i����N��xx�@��m�
�cP�$B��aaB2�$Z�,K߯��*B���`BH¤lxA�
�c�H>Qi)�C�o%*R%C2%�ٔ,��R�ĖE�X�t�&{%d���2@����>.g0����8:Ù�g��$HDx0B�)Ã)��\�cp%З8uy�;,Jhd!��E1��dp `BC;Hz�q���T��)9�;�|�+�W�$��MY���H$)$d ���� x0!��CRPaaC�A��64�R6S"��4c�%�� RO!kB%0�.S�k4mX0�cD�aI!HU�$a@�ɤщ$ֻ,7	�p�����{�r�$%�%��Ct�$�$ ja�HI$
@��n��CaHBi9ɝ�>a������$%Ì��s�y�B�
g	1n�ѶF�>�	���E�F��=��|���9������.:������GTƔ�H�
"B�"��U����,ʹ�]��s��C~ B�����T�BLL���H]��s�y�1naͤ���`D��XłA��@+�=0�X@���22D�uec�A Ye���hK	�a9$�lXA��&����0ZD��c��SRx��0��Ht�S$�댞��!Z9��;)��	@��c�8\���4�$#S\<b����&��9�Ray�tM�@��Ā�F��0�`��{.Isza�BH��#$24��%�P�S��p�-!IL!q�C0�Icᇞ�����!\ �Q���E�B-X,�D`��H4"XHH�W	"�$t��:FK�L&�����Os��|�H�B���XI B��"Jf��!��#B�W=x�)�� ���
�H�������֤n9�*M�$,��%64�F��)�'ghO��S<3}����$,�B䔥��f�;|	sH����o�& ��߮ ��-G���+�O��]�JP�0��䙜����ϼ��>+��a0��$b{>���y�;sy_!<=)L}d�XV]��/�$*B�,��ϻ>��=�p��$�"0X,��B$� 5"Q0cbX���B4	B,���ܑ5�������'=�fL���t�L���	��,�)�
K���|e3���� ��G�4!	w�9�4�>c$j�(īD�jHe�B
d�&�h�?Jf������3�㌎���H�!xG���#��m�V�%B!�(I�)�$��e�<��&�����xC1��+����dL�ġ/�45��A�$�M)0�0�ϺvW<��HN>�5=!�BY!0���aO�����*B��RI�n�w}���F����#z��p��:�|<�iY�0	\ܼ�zĉ�+"{�"H���0��Yg%����E� 0�cB�F�$�J��`�U W�0bЁ�),X2)�$T�	 ����I�%�$�Y�8NM�}ߺ�愜��N$a�1���$�d �1("�\H1Ă�%S!e"�Ӟ�5����jH-z{�	C^!
K�fr���D������r@��x����9sxo&�+��;�g�0�� ���	R���\e#�@�ՖddG5�!D�H�_g�zz���'�����2����Z���B����bJe!����
B F�HQ�X�
H���$H@��3�����XF����!��zx��d�S�0<a@�e�ϼ��!�~=����{�OyO8�{��S��ąq� �b�@�E�E�rT��>����w����/�����g_�|�H"�,I�-���ӗ�x����8p��	!y}!M�4�} ���n	
��X� 1b�h@����<�!�,�X%ɰ��,��@��D��!���S ��xr�!Q2��I0++��C���dj��H��$�d�I!i�>�N�JF��t�x}	
�	
�u���@!���'�.al���cJ�
A�(aC&-��$>�nYx{�}���a\�y�!���r0=H��<摀A�H� ��)�I���,7�K�,�$2L�I�_�#<cR&
Y�,��JSs$2{�w���>����3�bh@hć�ʐH1�$�����%1ՁS7����7�z�	 ������bHG�\\�4eR$03������.L���Icr@�U�b A"P��I�Љd���-�E�H4k�E��E�@���T�����o��ݛ�iL<���NS	�H0#F$4$���-#S$�E"G���$"X�(*��$biH��C7��g��H�DO� �bT�P�����@�������s���@�`10B0��BI"�C��0HԁVU��4!t�wnh@���/6�o�!O�7=��v��66Rg3���;;��g����,0��7�#p���s�0��LM=��ă!!H�l,�è��N��"B$B&l��hf�BT�q1�=�4�H�e1�$�Ba�bZ�"��hj�L5�HVP�X��B#!I�8��l��f��
HK��� R�!p� !*ư!�0#��8�}��g<ra�p�̽p�a��H��V+`�X�4B04����� �(a��ie�g��݁<ä=3@�Ő�(I����3Б>"E��zW�H\�g��a�Wd�S)�y�.�8F-�l�3%aYq�yXp�2e�x@*�D�0$�\"i��sɗ����D��(�)�
f��$a�7�4�5�KO�X���:�HE����sÇ�!C�
XB@�H��^���ԃ�$<>��mx���+
F-������!�]F���!����x)�I��VRP�}v"E�vHl�đ���+\ %LH�xrHA�cNB���I�$*I
@b1 @a$,�bHH��!��B$b�ЃH@���5"X!A�ĉ�|9}�(ҡ�J*�1`���)���.��+�����OOu׃�8�($l(����`jp`�b�0^)�J0����,��,/bH||Z��Č�HRB��#<f�'p8} �H1�y繶�Á��E�%��)��3�ϸR���,y@�R$i	2���e0ԅ��>e�4�\�Y#ZˡK�|�ߛ�>	p�B�T#P�0�	$���z��I�#"A��rHX\=N��o��}�ZB�"\%Lb�+#HX�
R�b�$B��F��E�A�RB0�H$ �H�2F0�B"�0��1B�)"�)� ЉW�D�IA��D��o�,��v����j �e"R%l�U:�,)�J��a+)-$�ZJ�#	YXFRRB���#$��Vx���W.�$`L��<s|ዤ�*����]h^CBO\g
� �J�ؤ�_��QL�C�I�*������    m$     �`��}��     $  �     �h[F�   � �HuPP�X-������⪫���:��g�8�@Z�B۵\��5rI�j�b�"ʵmm lg� �Xvs7Vtf�㋐�p��;(�@J�U]�6:jU
P*�U��@�5*��JKte8�Z�]�,�f�v� p�m	 �a���c:��$��n�;3�넝� hZ�vʂT�`���	6۸i�p�6쒔ֵ� m i1m�\ہm$�J	  ���U�@U+����.�)v�tt��U�RZ�U�R ���;T!��� %�  � t�$ ,1����WT�mJ���Hb��8�v�H�n�(�UU��n&�U��I`m��kX�6�>����0[�ͤ� R�꣨�9�vr��ۺU�!���u˻I�޵�� NV6�ְ �8h ��h�,0�cm�		6���3�W�4�@��/��~�a��T�.����T��
�`m��m�M@AK�WJ�J�J�R."���gF��� �*m�]�f�`S)*]WH
ʥ��uW�
�nU�yݥX[x [@��UL5RU]/�Z����U� �-�jn�NSTM]l�,��'�.��mA֚n������b�+P�k2�UJ�M���Zu�[���,[GdSg�h',qT��J�)��	�Tڷ^��ؽL	b���/TB#��^�ɒ�д�N��l�f��N@��k�`���-� [m�4ȝ�c-6m�   2h�c��b�nZ[A!i�À�U��U$:4UU����` 	 �-
�[[l6���B��N�l��mKW@E!5>f	H��&��J�S��ʵ:L� ˶��k�*t**�JuR�� u��H���m�T�#�+:�U�㨞��Lkr��^� ��ꪪ�R�A��) Y�ͶH8��ƴg����q&�������;��IN݂�Nσ�����F�[j���ڦ��[r� d孩�']Āpp E�K8�e5=�Џ5T�#K��n��˦�� ���G;<�*�5Vy @���`H �N[%h�	 �۶�X���'L����SF�@4P8p p�X� �f� ��E[CZ� m� �b��aD�ku���h,,�$�T�@ ��8A�f�l�m�[�HH-� z� $ �`m�� �m}o�|�[@A$�  $[@ UZ����UmP,�������u��j���[F� H6Ͱ   h� $ [)��b�Iv��mj%���Uy.}J9X4۶l� �a���tإ��ImM����m��� �qm��[@  sm�b-����M���6��x6ٶ��íZn�08�䋵�[xm�m�-�	�6�m�aÆ�n�^�8k����څe�^[�y�T�@��A��]�p Pb��'�j��iY[�m%[v�� C̲^��m�-��ZGj�l[C�9��m��$b�R� n�ư-U+/n�[*�� [����)-U�J�m]����m� �U��-�d���G+�lp��.�R[���T譖�l��4�ʠ�e]R�����.K��N����"Z�e	��)qB��++N�Ƅ�������j�l�FE�&�m�X��]Ӵ��s��[&�P���:-�i��Kd�  ]Ѧ�c�%�IVе͇6�M�A�GKŴ  ඀-�h $N��D�6�$�����S]�-�     m����[s�m�
�*�r�;WT��  �l�8 �6Zl-�K�m�l� �   		 s�ۭ̀I����� m�    86�8d �8m�_V$�v�,K�m�l  �!�j� [E�a ��� ���m�   �t�4���||���� � [FA 6�  �E��x t��(�`   ���"Ai�ƹ+m���`  m$-��nm�-�� |  �m    �\���m�"�  ���6�H2;]1�n�d�[% �m� m�&ϯ�7�D�-U�U*ȭ�(�Ylk���0��R�uF�%ҭv6� ����VA@8Ay�j��Z �u��=kHH$�m��ɺ��[L6�R- BIH��m[[v� e�j-���fٶ����6� ݲʵ@@UU��R�F� ��&tP R�M�m��$���հ	��ěY:٘��.]e��*��cC�u�j�r����/m����5���n�n@n��eNz�:msm&���A�T� ���m���m��HI �umU�˶��߾�����&6��$�)-P�6�UUVl��n1lu�-öYP��-�䑶�H �h��v�(��k��,���-�6��<���-�$Wn��:v荀�ڕ꫃a�-�q�ǣm�YD,�n��k"`kY�  -�"I�km�&�t� ��c��6�m�Q lHrE�A!"���d!�(Uv�hJ)M�Ңi���i�-��+�f[�-�Y1��@�v[�f�M�Vΰ���l�'H N��>�ꥂ�X)�e��&մڠ ��(m��ț��􉜷`W��j��n�����˳+��2�@*��u�ۋjYm*���m�$�6��YM��c��6�lF�8�in*�J��=m�틕n^ee�nfSd
C��
`��u`8q��cIg`�(^�/:�-�^�t����mհ�4c5�� �m��\�]6p ��K(��% l� �d��Q*��`�Z��m4�Hn7Uh��e��!�7mm�^��(�m��� [@  �` @[m�I�-��8 �d� m�m� 'okͳ[v�m _Sb@pWE�WK�U����|���mp��i��퉶�I ��i%��k� -�-�� $8��m�` [@ l�ᶖV�`ݤ�@;m#��iK�#�d��J�8[@�h m�����kXp$m��$am��fC[{l��l a���4���n�h0Srݶ�E� �Cm����llV�9��\��.Y��2]\6��4�䅦��R85�4�T�x͐�]����h��u�6J庺C�:��-WC�]�
�nÅª��uV�IŸK��[/Ꮦ� ix�.���kX �`  m�m݁�5�9�m�۷�mp{m�m���$�� ����z����k0�n� n�jͭ��m���&�M��8[I Z� kA��m����l r�	>���O�n����ut�6ݗ�u�������[9�n���y]�2�ө����g\ԓ����o m[[A�u�Sl����h�[����[����[@ 7�Ͷ�UR�*�<*�5UT��i[�K��a��v�� [R6ہ��h��-�d����m�m�i�@^Ҷ��?}�$�iw��.�˱! �m�  �`ڻ7kl�i� �՚Jm,`��[
�m�n�R�[P;�0�UT�m.ܷR�ʔn�VV��:R�K�h�8H�����^�SU~����Q�˝����;5J�K�����1«�O>���kU�D�n�$���� IۮH[�\m�� �$m[l g\c*�V��v�D�.��p kh�H ڶ�� k7[iib�(0�QEJ���v��(�u��oPk�n׃u�p �kkU`HH��m�e�6�!�*��j��UUWf�:�֊L�A�� R��.��ۛ`p ������M�2Z���  ,]�ʬ�Ͷ ,�^� #�	�. ��o��� 8  -��kY�uI�!%�m�i�հ �[q H�h m���[�n  rY@΃i6-���[E*�+UUR�*��  e�[D�p�-�n�H vSvH�G0&����I'm��遶�m��p�` t�I����� 	gQmm�sA�l� Z-���	6�6��k�Z�lm�JJ��.ʑ=R�UV�[	m���m��J m��H��jZ-��@h�7j�$�;8$������ɫ�hƕ�{S����vl[@�c��� �kh�l�ai�[`� [C!������:-�<,0�v�!'�8�e� uJKUR�+vy:24 PF�Ep���:[@��  ^��v��X�lUtuA0t������ ��lIaҶ�R��v���iT �:�Om 6�m�fe����n�-��[��� ���"��~�@+� ��D�����tOTCE���$bz�c��Dz+�A]$�����1X����CA|GQj��Qq���,:�g�
�u�W�Q�A8����JD^(�$T�E� 58&.��S�r,$Bu�$Ji�PǊ��=$D=��S�`"h�� �OO�C�%O@ �E7��/ԇ§�:�4�qO������0 "�R$A<
�O����@8��CT~:��:*x ���uG����E}t��9ST�SA;�C�@���~ELW����1aĄA�Pu]=A������> |{�`�� ��h�������"���!b}P)�����D:���U�!��Z�8�F �� � �2!/P��(���N�����zzQĀL� `��^U��M����`!"���A�C���z|`"#��&�'�E�	��x���@�h��G��p�W��|X�� 
A=� ��{�8
��$���C��PP��u@SǔU}S�C�����1W����HB�D�@��,hP���"�S 0
C�C�D(�`�p�V&�R5"1��(@s�����&f���`mJ�"�z���赪�,p-n���D\� ���s���x���B&�2S�h����.�I/T����E�ڠ�e�h�x	�@@k�����/\p��AKn�U6���,�II�@ݮWg��5���<Q��Y
�A۳�h�^��Ғ#�Ў�yt9�,<�m;'��mh��!Uuҧv悸8�*��Z� ;(=�z�����n]�a!c���U�M�ѬOH��'�<XC��Ҋ�m)�<v���P����RN�H��K( ��Z����W�[5�Y� �uCav���0��⮖eY	-ʪ�+�b����Ŏ�A59'�ZB�u��s8y�{e���TSŭU��k ����N�P{%q�g����I��ZBR�g��#�Z���e9�Zj��rRtn{:����Ks�6�8�2��ܓ�n60�J���hr�2e�JV��k���lO�SaN䘹�X^���t������\��K�Ąr�*�Av��[�fN��ؑ�3��H�7k+�8��v����Y���g]�u�����F{v��g$Ny՝�1Ξ��#�K&�K��k�wOul�h�vɹ�����h��6f]s�lW��7	�;<1��f�+۶x{AGi�T����ö���nS]s.7+U6�j�	[s����ZA���]�L]���\%.M�_\f��8�gC��R�Hl���F`$�!�Ü�g`���(��Ѻ4�
[��a�b��zaH�]��W.�kp��F��ˇ>M�e���e���]\�'5ύuu8�v8�6^;Z��]85�(�fu���ۭl��Nڄ������[�;&@s2�5�;9�g؞��ZA8�8\��.;r�ٗc���B����b��(��-v��h�	�f9ku�D����d��ۋ.�*��tj�I��Z6��+dML�%�[=�(B,s�I��o{�ܯP�ˊ
�����C�MT_�G�T9�^�{
+�=A>�N�
|��K ��AdC��7l4�a�w30q�w8`nc��m�W�F��=��z���Q�i���<�pj����W����K�:eڥ�gM��MkwkkZ�M/��Knv#�^��r���h&Ʀr�v3ok����̀m���׍wnz�wg�n\I�{Q��Iɜ"�.8����������N�J�󮺪��$�v:�.Lᐓɒ�ksvf)� ��@O3w}���N�p������T1���x���gg��˖��-1�>�sy�r)=�sD�I߽�S�I���h��"X�'w��O"X�%�{ܿ�[��n\7��7v'"X�%�~���'���İ}�{59ı,O��|�yı,O~�p�Ȗ%�b^�}��3.�Y�4�s7x�D�,K߷�S�,K���w�'�,K������bX�%��wx�D�,K�^��t�d��i73vjr%�bX�w����%�bX�����,K��>�s��K��Q����ND�,K������rf晛���%�bX�����,K��>�s��Kİ}�{59ı,O~�|�yı,OȪ�4���&ݞ�Gn��-N�y�	t݊���>9�7CŸݜޓ����,��M��N������X�%��w���yı,~��ND�,K߻�8�D�,K߻�"r%�bX�����͹��Km�ٙ���%�bX>������G���%�OP1;W��'�,K��}�'�,K���s�ND�,K�߻�O"X�<ox��9�Baҕ5�w��oq��%��wx�D�,K߻�"r%��dL�{�����Kİ~�����bX�'�����I�C3����O"X�%����9�+��,K����O"X�%��w���Kı/�����%�bX�}���܅�nt��D�Kı/��w��Kİ}ϻu9ı,K�{��yı,O~�p�Ȗ%�b~  ��|0��0�n��n�
���`-�ɮ����ڛ�ўw���©�M�.�E�D�ci�>�t�#��R+���'"X�%�~�{�O"X�%����9ı,K�{��yı,K��s*6
�ܢ9"��9H�#��R�ݖ�D�,K߻�"r%�bX������%�bX>������\��,N������7!�nk���O"X�%��g��bX�%����<�c�U�%� �Tƀ�0�#�D�?wy59ı,K�{��yı,N�[�s.d����m��'"X�%�~�{�O"X�%���٩Ȗ%�b_���Ȗ%�b{�s�ND�,K�v����5�in��ۛ�O"X�%���٩Ȗ%�b_���Ȗ%�b{�s�ND�,K���x�D��{���{{`�w�[]sr�^q��<�!+آ��Qv�.砳�J�\1N �r��Ls2��͹�59ı,K�{��yı,O~�p�Ȗ%�b_���Ȗ%�`���jr%�bX��O�o�&��.��n�<�bX�'�w8D�?șĽ����<�bX����S�,KĿw��'�,KĽ��m��[��˦ni�,KĿw��'�,K������K�C"dK�߿oȖ%�b}���'"X�%��{�6K�nK6�7337w��Kİ}�{59ı,K�{��yı,O~�p�Ȗ%��~:����M?';��}�'�,Kħ��ن�IvM2�33vjr%�bX������%�bX�����,KĿw��'�,K������Kı>0�YNݱ�$w��m/G]7N^k���7����v�&��T"�t�"���7!�]�.��<�bX�'�w8D�Kı/��w��Kİ}ϻt?șı/~��O"X�%���̹��&��st�Ȗ%�b_���Ȗ%�`��v�r%�bX������%�bX�����ı;�͙ܽ�v-�ܛ��O"X�%���٩Ȗ%�b_���Ȗ?�dL��g��bX�%��߷��Kıo�����*k^ﷸ��{�����߿oȖ%�b}���'"X�%�~�{�O"X�%���٩Ȗ%�bw�}{|�7Hfau�sw��Kı=���'"X�%��9�߿oؖ%�`���59ı,K�{��yı)ʺ��U@��c*�I"��RQǧ��UFt��qC*jU�[ڒv\hv8J��m��2��ئrkj��m��n^Jx����n�*[�<�R���x�Xě���a�(�v*�����2a,=[.c{jx�,��[�.۰�\��x�l6�� �׌�:�h�U,�659-��g��n�[��r�r�Ӹ_�g��o�>�U�8���ql&��ά��u�{���ܺ��P�G�\�rJ݊���F�Ņ��<7j���M{Sdb
2;��s:D�%�bX��߻�O"X�%���٩Ȗ%�b_���Ȗ%�b{�s�ND�,K��nfݗm�7337w��Kİ}�{59?�9"X���~�'�,K�����ND�,K���x�D�,K�}��˒]�L�L�ݚ��bX�%����<�bX�'�w8D�Kı/��w��Kİ}�{59ı,O~��m5��M��˻�O"X�~D����'"X�%�{����yı,~��ND�,K���x�D�,K����˘�snM�7H��bX�%����<�bX��of�"X�%�~�{�O"X�%����9ı,O���ǳ���e�*���ͻV����g�]�H�7����õ�lj&�V�����~�߽�7������S�,KĿw��'�,K������L�bX���~�'�,C{�����Ls8�a�{���{��%����<���q@��dTAP�'W�=�hG�ı3�g��bX�%���x�D�,K߷�S�? eL�b~�N��̓t�fYw7x�D�,K���9ı,K�{��yı,~��ND�,K���x�oq����~��@�p=19����,K?
@ș�߿oȖ%�`���59ı,K�{��yı,O~�p�Ȗ%�b|w��m�۳r��s33wx�D�,K߷�S�,K��G;����{ı,O�����Kı.��!~!I
HRB���5DM�\���U���m<�c�!��8���yw�����м�GQ0P%8��!9Vr��G)����'�,K����؜�bX�%����<�bX��of�"X�%��}�s)��nBm�2��Ȗ%�b{��lNC�r&D�/~��O"X�%��w���Kı/��w��Kı:I�w��a�͹6ۛbr%�bX������%�bX>�����c��$8�J0a$�p�8lO"^w��'�,K����؜�bX�'����ٛwa0�ۛ�ww��Kİ}�{59ı,K�{��yı,O~��Ȗ%�b_���Ȗ%�b�~3�Tdb��7!9Vr��G)���/��Kı=�{�'"X�%�~�{�O"X�%���٩Ȗ%�b}��3'�͹�Phܦۋ�a�{FT���t����}�yO)��׎�Qy��ڻr�^�������%�b}���'"X�%�~�{�O"X�%���٩Ȗ%�b_���Ȗ{��7��??�����`�}��KĿw��'��c�2%��w���Kı/~��O"X�%��}�ʜ�z�Mr��G+p�?�Q���F��_"X�%��w�ND�,K���x�D�,K��w*r%�bX������%�bX�����%�4��33vjr%�bX������%�bX����S�,KĿw��'�,K�r/�j�ߠ�{ɩȖ%�b_��w)��nBm�2��Ȗ%�b{��mND�,K��;����{ı,Oӿ�br%�bX������%�bX�v�Ӎ�����;��܃��/S/��BXڮ�շ���y#'[:��^t���ı,K�{��yı,Nϻ��,KĿw��'�,K��}�ʜ�#��R9]ܷ�)
JI8Ԓ_+����$&k�P�\E��$���~��+ �ݗ�
���JH*q�B:�� m�]k���@k֡�q�U���mҜrX�4���`f��Xn��jR(��Q�Mـۼ��ߗ��׀k�s�	N	��T"t�D@�I��؋2sN�i��$��n�t����k��5�O-�M�8{'={2;�L�1֪ㄷ�f����ج\	X�U�ۇh�vӣu���Y�j�V�qm(2�k�St�lϒ��Uٷ^6u�T2��:}C���l�ͻhT�GNtF�Z�z��f� :Z��[M��N�d�N�ݎ�c;��M�4 ��������c�2m\�]�M�l�����<�e�p�6S�[����msJ'�R����c]�,��a�@�ب&-g��V��������� kn�u�p[w�^�*�l-T�MZ�m���� ����n�365S�:��))�%���U�kn��P�5�hF��]]}M]R���� ����ŀۼ�(T�\����i���(r)$�3u�@۴�l@۴��n��t&�eχ��M���!:���@ݞܩ�ō�8�^N �b�u�ҋ����O�n�nـۿB��9�� �Ng�s$͐���vw��g=@�b��  "�$:˂)� �R�B�E"+}H||}���}�I=������V��E��6�H�I�+ �ݠֹ@kmB��c[W3n(A�um�,ǚ��۫{��`���0�
��I���X �'�� kn���pQ�w��oǍ����e���m8���r�V˻]��=�Ws ݶ�8�5�mPu�zwh�K����t�m��k��� 2�4ێ>N'�dV��,ǚ�m���DOoaӟ�L���T�r�P�q7����ug��]���֞�Ċ���<F�Զ���%������j�
��)'CK����)�<��	�>���F@���������C���>����H���8����\@� ^dBF�b��C��Sc5:&hna�f���V���0�B�A�K�d/��Q�8������M�G����@�����<T}�H��>��*�@A=W
�+���9[ߧa�`�zX܍�J8�Ɣ.���p9%����;zΜ ���z"��gzp��U>���䢩U�����c�DK������5����=��M�����2�n�fK�QǛ�ˣ����%�@.���?���n���&���;���k\�����}A��<�W�~�n(GMTm�$�7j�R��v,����m�rS �k�T�M���EM�� �� �v9â�{�����3��"q'R�D��rU�%
{{� }�x��8�B��	�P�� @��b
�� �*Q�g��ɇ�˫����WWT\��� ��^��IG����w��X��W�Vt��H��T���p�S��g9��w�5{8ݹnw]��u�~{�����u
JqG����3wn���W����@o��`fz5�qS�)wUws�kotD)������׀=����~�7��6�8�Q�n���`|�(������ {Z� 5�x ���Bq�M�NT�+��[�zX׽8��`tOoaӀ>�ɺ���%M��U5wx��8�^��{�/����� �ݖ ms���*GDb��&EF�\� �6y{d�R�Tk/��ָulA���C��`Z&�Vt+�����RmTt��� =��;r����g�����r�
jWj��؁ˑ#]�k6u�������^+���f��hH��ͥ��x��jҝi�&���lii�scF׮�כ��MJ)q���u%���8-e�\�s��$�����'(�67Eۮ�{���{��Y�9�K�x�Z#Tb���7�g�I��|�n���m7��}|�
��I@��߮���U��w_���׾VsbU�$�S(��'%`�i�rQ2t�u`�����:�H��x��'�ԍ:��������8!B�*�{�ŀyח� V�/v3%�76��$�������������� �]8Q
�wu`�/���Ԫ���������o伔/<������`k\�� m*��_E,����Қ�u$��Θr�QZ��G8��\�)�Q'�ޮ\����Ҍct�RW@���~V��`k\���B����b���I3Y�际�6L�o$���s�,F$TD�(������_����8>�X��j�ܮ~�9T��߿Z��)�ƛ����N �x���#�{k�N��Հf<Ф�(��HԊ��^���X���@9m�'5��kD�5Awq3Wp��S�(�@d�t�m��D&�k�.�6��P���ʐ�r�:�=���.8ɳ�.-����<�K�v:��3���F�E�^������`n��X���`z�\�s��W�Ԩ�	S�5%����� 3)Ô��@9��mG)S�)"��!`����{Z�}U�ŀ	$B�A�BLK�^_~>��^����i덥���
9,=Kޞ�+ �{���٥��o���+��!'%F6�9P*�� kn�P��8���Xt֫�*����� ���8�4J\�N��8�Ѯ*����%���x%��\�7����ī�
��ci�:���X��V���z���}�K3��ӌ"�A'' ��,�G�yzp��^ ���r���F��(�3J��������t���J��t�p�u����dq��q��'QXz����ޖ��$�����=P��:�*�pw{�\F�P����� �O�MM؊V�������ֹ�:"%�u���t������s} �Lc�C�B�6�G�9�t�5��3��Ѻ���Q"�V�'!���s�_)9J�iI��] ��ߥ��{Z�7v{��k�+�O[�1Ӝr`�i�z=A�{׀{��8 �w�(�{��n��&�n��(n��{ޘ��8y$�
�����<��Ӏko&�n(*S���$�����{ޖ��j���`w���(�B!�Dq`m��I{�<�? {���k\�H�|����r9�u���.��&�եm�Fy���ں֛��m�n&ѷ �k���M�/F�gS�X&7�9��r�ˡxʩ�(�F�͟;��92k�hv��cgY��]�Ƴ[X�b�J\ٶ�;F���v����5��n���W�{�l���jv��/\�y1FB8�&m�Y�I�4ܦ���[�6HvJ <@øA�;K�]m�ݞ��]ߟ���_�~���m���r5�uz�v-�x�&��n-�۳a˸�#��
�u��2���ڮ8k�0w��� 6��k\����X�j�H���u#�X����6~����=�{ �m�:Jd{O�UMحM��������;k�p�ŇBQ3��# =�zX�P��R�R�a����BJ�������`m�*�W9\^��+q���P���J��`�DBJ{�����8m�X�n�@9FJaT�7�����N,-�<ݤ���M{ ��{��{�r��E��&��R����=�zX׺��ۯr��_ ����b�rD���e6��䓾�{y���	�C1��!��q�!f��_����`m�r��;���J:�(�I�`{��Ձ�z����Q�{׀{��8�m�.I�j�]ڕ5V`r�=�˧ ;�� {Z��\]���X`i�u8�����n�G;}>;�B�8r��ӓ������;i�8��ժ��(�*[�9�(�1��u҅�q��\x~�yJ�qt9��~��(������ŀ?��>��H�����F���Ɣ��7����_�Rv�.� m��k\���S�����
������\�pw]���B@{��dp��D"#�~���<�k��p��ŀ笙��W15M�u��In論�{�`}��V�잯+7}jI#�NF6ܒ�{Z� ��w~_���:pw]�'��������s>N�H��u��|A�k�ɻp86��5C��7��{����h�2,WK&j��wv,�M9��w��9��X͞ED:��D�z��_�D/(J�;�׀{��8��,�
d�ii�u8�c��u�n論��U��*��{�^^��t���V��f����������}� SNp-��>'�>j#��~��g���I=����w*R�RP�Vۛu`{��=������X�5X���m�IJ8�"B��t�]5x�JuiGK9���}�óO�Sv-��7��:)��RW�{���3����y����}u`��������n@*�� nk����ΟJ9��p��T���ZrI"�S���$�=�|��^,:L��.� z����U%�U�%M�ɚ���zV����<��Ӏ����B�DE{��8�_�W%+�-]�n�`�i�脡z!W>����ӄ�w��䓇�;���ϐ_!�4��'���~`����������zM�� ��`�{�����+�@��5L�8%�.3�����=��V��Q1� ��$B�]��*��`�=�"v0`�ް��B19ImW%U�QTP.��"crI IR]U*�uU��6���wD��XB��ݞ�F��<L���9�\;����h>����#��n��7S�*�e���<�h]Q!������dv1�0pEe	8ۨ
��	/,�F�0�se����m�
P)ʅ[\���8���ٻV���"rOx�Og6�;�3�5nm�m��D�9��t���1�m@�.�@����1�ܛ[Uǲ�1�f[��8�uvm'[lY��BH�v��v�Qy2����,�N�aj�U���[:����1��Ѿ>`Z��9jU�V�@u3�Wn���v��#i4#!tlV���jU2+WXp�y�K��FK#�2�MGm�mv�$�9yVn�K�Y��]=�f8-�{+L�F&�J�� ��q v]μ�1ɭ�ʹ2-$!��,kM_&����t��d�� Q�sp�F��{H�@���%��"uY�.p/FIe٩[��"������UT�]F6ʵ�� "L�n��Yf�f�l�P׶D��:2�,�F�>qV\�gkP�N����8琼�D]9��q�'\#HW[�e����/Z
���O^ݴ&GE;u�,�����ac�m��mU��lr���J�]��8S�� L̪*��۵�M�d+ۃ�Aq$h��ڃ���
�ZXG=m7Aft��ĩ�&�2���Ӛ��M̘9V�����������6��N���ㄝ�����#�_}��4s��ݸ�έ��i��E!\�We#;<F�-K����^ .�./3��M�qrø�<Q&�$FG!xL�u��H���:I�V�۝�Q�6s��ۗ�4�si�坵F���t��!^�}^��7�;r��T���;Np�T�9�&`3��B �MmG%�������hVZvرP���)e٨��!q�ؗ��nP9m�� '���j�W7F4��ν���]V�g.��S�k4�.l�:{7j�N.�1C�t�frnl���@ 4OL?Ϡ+N�/�a�"C�������;��8|�!�z#�ȩ���wws߼��g}��D.|�;0>ɤݟn1�2��2Xq��S������'(;��=��Wq��#�����X1xΉ�uNhw��6M��s�,=���[MM��D�Ju��.&����S�5��n�z��{���ۂ�c7��*�NM�an۵[m&��{�0�8�:���g�t�n�� �݀�� �TT��^ݻd�T��&�&��n����˅|@��;����e2��k���nA��.�^3���-�շ���y�o��u�S׆�.nn��w����0�^.�!�O��;��jB�)q��������JO��,��)��]�)�ɽ�7JԧRA9��]Xkͥg�#s},͞,]ƴq�QІ��jJ��η�(��@nm��B ǮfiIR�NA�IJ�չ����ߏ����V��Ұ>��I17Z�4��8�|��Ӷ��"CQ�#Qp!<��m���`��I��m�%��ɥ����Xk֧������޼�z��T�.���E�3g$�w���(v ���Qa
)(����7)� ��x��,�&��"T�HTrJ�;�6��gse��ݺ�>�۫��Vl�:�L�ԕ7jp9)��� {݋ �����B^I����V~~��5!N��pm7%��֡�g>�x�}�75��ֲ��M���퍇F�JS+����dT�Xܳ����G��5��=q̅i�+~�}� {Z�������%���� g�/ÍҎ�6�RU��y������� {����Ş�(QT}�jG)�B��IIJ�=��,��,��u�ҔtG� ���~��'�gR�>�m��&%9��X~���\�9Ȯ~�� �w�`:֧�IB�\����B1J$�M�*$�`grTyQ}������@nkP�̧QL��&ɶ⮞��;�\e6nM��v����l���1[h�%����w����N��V�nn������>�@����GG�}����3[��u8��)"���gse��77�V}���>כJ�IY��ԅJR����@=|��B;��}�����ʺV�]���7h����Q��{�o��� 7�w��D$�"R�*&*$F(��`��`A�`�A �1�`!�E��Q����/��y�NI=�?g���f�(�����X�Z����\������ͺ�5uk+J�'I0�r�D��ky3W:��M�e.k��Ţ6����=p����O�p���mФj�%.�{}�X�۫�ͺ�;�6����dM1)�M�ԑ�څ���d�|�ΟD��v�L��G�lR�*Sr
�%X�����y���F��X�z���wU��)�)���ݬ�v�N =}x��X?s��`wZz)N()J9%J��l�<�{���|��� {�b�1B�ĔL�hʅ,B�S�d�ɳwLsdNz;n�Tj�ъ]����,��Җ������8:5��f�lvc]���q���Ơ-�s��x5�Sh�眽n�ۍ��n���e�RdGg�:�O[�k��ʄMӻh,��P��K�]���öq��u���0=��{�Xq����Z:�V.���%L`)���x5�1��Av��Ru�D�Z�S��{yi��z�ķ-�-E��A�)�M��f�-��2Cn9-�s�#5��H�i���\d7kS�봶��m����V&�)Ґn�m9<~��Vۛu�=ֱJ�K������qwJ�+���.�Lլ�׋?�!L�ϖ, z�X�۫�T�����GCr�RRy�(@��������;�FԎSn�$j��U���Ks},��X�B�������꛺��&n-UMT���;f�QQ�����~�� ����{�PQ �C��ax�%&����6�������kux�p��x�����u�@nAQ>��]X�ڵ����K�޾0�]L����f�3M��9$��t��8������!��#�D~�O�}��I�o�~z�g�B�I(UF����7t�&��.��Z�6{�X��,:!(S?7ذ�������5!N��pi��r�܄�N�~X��,�b�������տ�:��F�����XfmՁ׮ =;����@y�A�UL��G�it��G�n���O��(]�l�u��r�x.n�)#��r9t���dt1�)�%t���t���@n6����!���]�3wnSn�q�D�*��fk�Uq#s޺�;����WW�RF��q8����7wX��X�׋��R�D4�K�(��*����]X��vnM� I�d���B��������w]`rT�=���?6�ȕR1��U���b�:G��W�;z��?n�X�#�K������i��w%�-��Ϊ,VF����=�2v-��v�=�M�����窻sk�K}X��0ۯ�%�C��`w�W�ԅ:�6�ێ������%
d��ŀo>X�Ӻ�<�B^I(�'�t�R��nʻDլ{�� ��X��
g�o� {݋ ��jj�ꪈ�6�6��r��g���X[�vw^,�_)�D|�"(_S���5���9M�I��$�V�3]��ݺ�?n�X�k�	o_qrPI]ط(\z�y"��k���SVLP]m�w���^]֦��ʎ�ܑ8����7#�����׋ {�b�������+�.������>�۫�8��o�������w���$���^���6�IwD��n�`�� �;����G�׀|�b�>]F��R�I$�V�r�u����ր��P�׮ <�e�SvEDq�Q��;�,s��w}�|{}WV�3]��S��%�jDD���
o/�b������ G��{p�0�v����녭��S�8Ǔ�SAd�cF���>]��յ���V]���;ez�����}�4��v�Q�؎ ʚ���0�ÛK�n[��ݞ�-x�M�P�]�kN��ct���.ƄwS[���6\\�l[��X�@\C�b��y�fH.�Q��i��dB�6���ٌ`�z�+�<����߯篭�<s����ڷ�W\��ƻ����uwd�7!���\�c������O\�8���5v��� 1�N뮏�= <������8�m�m�mIVw6�gB�>������I~����|�b�>KwRRI�I�AIR��f�;�L=
&~o�`ϖ,uۻ����f��U]�(R������ֱ`y$�y(U����;�~Wt]�݅U�(���'�}��~S���xpO �`�`�`��w����A�A�A�A�߹�pA�666?�����ga�p{Ok.^��W�KB^�y�V�z6̉�q�����nx}r=��S�.��q*��{�� � � � ������� � � � �������lll{��~�|�������>A���߶���wp���&��pA�666>�{�8 ��=G��E��� ��H�~LG�@FA�V1�@�L�ӄ��
)
@� !##
�+ ��x�(�Sπ�A���}8 ����8 ����Â� ,ll}����˻�6�ffnpA�666?���ӂ�A�A�A�A������ ؃��r9�߿�>A�������8 ���ߌ�����sst�vpA�666>���8 ���s����lll}���pA�66*������� � � � �������e��&fi�wN>A�����8 ��;���� � � � ���~�|�������>A���߿��B��s��;s�y�e����ɬuv�1����A��}�{�����`��!L���� � � � �������lllw�?N>A������� �'�A� � � �~�9�8 �߿��٦���u�&L�����lllw�?N>A������� �`�`�`�����x �s���|���P� �l�����ɹ&�ə�)76pA�666?w��� �`�`�`�����x �x��Q��O�ĨՁ��ބ&����� 0���:O��A/%@}��$�4�ON<G�MU ��*��x�P�O�H`)Q��x�!4Q�"QR��Č,��"<3��dE7�=�O�U�2T�P}=!Uq	��(;�zu%�-q⪖e\*Fh�ӏ�. >�^�ঀx�'D����?����'�!��x�� Qqj.���8+����{������lll}��~�|�����m��źir�3K�wN>A��D,~���ׂ�A�A�A�A�>�����lll{���8 �~��>A���ߦӿ�7p���&��6�A�666>����|���������� � � � ��xpA�6	� �29�o��x ��v�?�9�a�&d�r4ɒr��.M�u^Ktģ�$����qq���}��/��R�f��0�33s��A�A��"��A��������lll~���Â�A�A�A�A���~� ?��>� �`�`��~���|�����?w)�����.����lll}�xpA�666=���ׂ�A�A�A�A�;���� � � � ���~�|�-���{��I�w32nL���e�8 �"E	D��H��t��o�B��U]�_�=��V���NIQ)t���9O��V �����ŀ�G�BJDq�+5��4�F�INJc��ݶ`�������V�w]`Qw��N�ڋCڹ�'&��=2Vn�Am��&��ో���٘��/����e�:[`��B�ƺ@zw]w�;z�@=v��RR�FJ�IV���`|�5�ݚXfm��#�5��q��q�������Հkv�:&~o�`��N��Z6�*A��m�`f����3n�׵���fk��ݦ��J�br��7f�u��<��������V��0���B�JU�|Y3Qwd�kwO\�3�9i�-J�m����Y�f�qˍ�kYwWS�p�W�-�n��ѓr3���M㥞���Vʬ%��'���u�@��r�@F�l��5En]�=�r
�v�V��l��\]�Muy���]�Ѿ�>m�sSӖR�%^�\� ��\�qFKur$��^�N�"s>��q�����4]��N)�F'PO:�S��� �SO�=���nܺ�ͤ۶�ܼv��Ewb�.��N���}:Է��v���[���>�6����jJ����ߝ����`ovi`}��V��֓�TCJGT�� �;��������}� s�]gq#wҟ�M�����7#�=��,�^,?�����<�Հl�z��me|$��!���f�X��]�}�����/g�Ł��y����8����9ծ�Q?7��޾0ۯ�6�ZA!'P���I� �g�+t{-�ݖ4��:�uѕ��\ΐ�d�����&*� {u�� =��w�G�zC���;��jB�d�m�,��.VjE �(I�@�����w��rC��v�n� ��v���*q���+� ��x�:���I%2}�׀v��`b��أm��s�rU�W���Ȯ�]6��^�ZX8�	D���� =���ܒRCI�Q�v�we����f�;��ړ`�MLXI��;#�n!�t́A�n�1Yb^Hخ�m�=�W9T�ĝ�FRS���nO��zx�>�x�:��%�� |�� ��q4�J�d�8X��Ձ�k5�{�,ܚ_�\�RF���JJQ)�8�wv�<�V }�w�$�T(��B���$!b�Xz��?�>��ϋپ��>�։��x�cQ$�� ���m��� �%�C�@g��ᑔ� �JiI,ܚX�f�~_�s��`�7x����I# ��1Yü��/Y��Þ3���ش��Y����خ+`�`�;��ۮ��$��3�����35�@�]�=�����| 5z�^�6�M1�8�%Xmf��Gq�N ���P�Hn�ŀ�z�j��L�&��I`}ך�r��~>?RY��u`��K���țe%9)�NEa�R���� kZ�P��ٷ��nf�`�	R�7R�!`}�۫�K}[��ǾVnM,�J�$I�R�����m�Ԁ�l���[>.�Z[�d}�vȧ]�(�s��+����4H���7վ����^��j{7USU�T�ɕWx啕�$�y(�;�~0�ذZ�y伕Q��⋡]�sT\�]��u��� q���nP���˸m�7%���.�����o�� <�z��Ss���W{�x�9~���(�q5M�8�%Xmf��9\����? ���kŀ	(Z�%R�E4`� ���,ٶf�۶�\��J=��{�E~6�]��m�T�%n�������\���Zpup3����.���7b�UW7j۪x�� �7[<ri�b�e�m�`���Gv{��]��pU�7^n��u8K6�^���ך8��fi�ԕ9��dx����6+���=�N뷬-����٧FXCh�mf�*�6D\��7Rf�T?sv^O<�]���4�.n졕ד5s�8������Z6��9�]5˗P�)!�۔��&���Ł��K�ͺ��͖f�[�INJcp�1�=�����, �.���v��9����	R�7 rf���3k6Xwf����imm%(�r(�"��9L��׀}�ذ�k�DD(�T߿v��(�!�_��`�%NK�ݺ�V�@fkP�F�@laM���\U������C�nku-�NW{x��)wmv��= s�.X�deJ�7"���=��}� ?����I}A��ŀl����u8�㒔�X�m՜�9]�J!%�`6�~�^�0�k����=��2�jq�J�eo��������s�{�X��Հf�o[�JHi:�&i]�����0�}8�7��#���]��9��g�Su\Z���� yZ������x�Z1����{��~=�ۇƳq��L�]�r��(ݺ15�'B�yB7^NΝ�S���x�o�E����h�*���n�(@#]�3P�x�U�޴����N9#t�U�ok6_$�ɻ݋ �Ӏ}�x��"d���J�]V�U��Wx�v,��W� ��P�H���%��X�k��?Ks,��V����fK�X��$�_�x��b����Ч������*��ttM]��7b3Z���v5������K���0�Т��'NB0z��:sż���v��Cպ�,䍛��W�{?[}Xz�Ț������ p���=��@{��ϐfo��|�ߔNRCI�r��$�?|��/B�����b����yEW7}^�G��Jcp�3=<X�^,9z"*��z�~�ڇrU@Ө	���,=UT�7�U�eg�,����b�T"1b�B�郊Lj+H��� Z1F�;��*��ٟ|Xu������rF���� ��v���#����5���3Z��U�h�rP�����*�Uԅ���%���ܝ��ݶ.�a��Uƺ�*���$�����c� 35�菾􁵛�`u{�xdeJ�6�H��٦{�!EP�{ 4�׀~��3��>��?S��`��AHX�� �wva�J��z��7z��6[j�݊iT�QWk�!L����>޾0�v���f����~��SI�qP�G`{P��v�f���t�߾� � "x�H�2Y����8�i�y�x�#�>���@=ce��XS�"�BJ�BH0�Ȥ(�%��`u�V�3�0#(��3�0�XX�(`jƴ}�b�0I!聝qt I�_���N��G���$�@� b�Q�ĉ�^��0�� �+ �HH�0$XĨD������N�?
�'Ą���2$�Ii�		��0"E�Kl��	0!���N!U�- v�oKӧ�q���a{M��m���v�n��n#��l��ý����s���2�F�ëN3s�+�g�l=�=N�5���T�H�=��ŻJ͌P���:˶3��Y��	@��nԏU3Ū�2�1�`�N9Q�0;���L����Z(5I��e��c'm����
�V��z��s�^n�F�9�*���j�؈�jB���$�@{.ӻ#�6m�C��j��$���TD\�$�$<۳�r�y�Ω<B��H@�� ���U��[m��ڶ8X`ڬH�
���� үF=���eC�5 +]\���j(����l�� +5m��@�+��dT-��<��	��RcR�D![r� �=N���k9�lG	��jAvs�]gNI8d\����C��%NI@�G3b�Ot:��f��-��T���Uɬ-���]��^�)�]��H*�(p.;MZD�{Y"W��UR]X�y����8ї���e=amnۊqٳV�F�V3�g��wd�r�[s.ƛ`���T
;L�̕��^S��v��[���e��;r@!;�'��0����%��[�R�VIn�^N6j�&f�׮T$�Y]ř�ܣu��Mv����4���61�.�",�uR�ƻm��vvRdh�l�԰W�q��� L��׬�+�:btB�ldr��+��Ml��n�eP)옢��W	���,ty�k2�A���ۭ���[�ܲ�����Bj��r3���
Իv�	���e۪S��Őܲ:�@,砐�X�Er���#s7���[<��I��$kkq��\�✍���EC�t��5�[R��.wjj�pʩf�2����ZVS�nЎ���4�読�� Jvڥ[��FgMl&���	�����( �Y��ݴ�:n�1ѩ���%�a�#�cf�n�M��ڸ��v[�����W������+@��&�hb5�R�<5Gދ҈t�`��(u?/���b���Q���(l?=�ncQ�m]�����a�'{#�i3�ŕ�W��4��������S]���pa��5f��X�nҗ>��ǫ/v$�s	<�,�lh^[�.�c[�=��;<�[Y5���g����$�H䓥�o4%M�$�;En�a�E����L�u��T����7;�����p��%�s;n�ػ��([�9�v
��I��j���Nv��+�|?���Q��ϔ.=!6F��n�j�����m<� !;���pO��G-�q��9�LbRV���`}��Xέu��_Pk��`�z�����T\�6AWb3Z�Nƺ@{ŀ~�l�DB�QT9ryyLڹU�J�������Hcj�l@fkP���E�j����T��r�s���}| 35�A���� 2{�x�谎4����٥��3}�|-��>��Ձ��U �4�'H$)�RP�/�z"�ڋ=������V�ڥ���?s/H8��)���]XY�����~�W9��s�Ł���r��9�TR���7ka���#�}�k�h�mՁ���Xڱ�QӔ6�ӐN� {�6� 35�@�v��q%���9�LbRU��ݺ�;�۫ ����6M�U8��*bɚ�@fkP�����ܡ���o�����\��&�:��&KTW	�ݛ��8;=�[Â�dh��+̵�4n��� 1������7_(@w����1��NR�"I`}�۫�+�����kv���2�.��&�jK�X��,���HP�D!C_B�fmܰ;��V�nm8�F1I$���@fkP�3[���:'_w���K�*Ӕ
���%XsvXwZ�kj�� 7�TTEM�ͭΝ��m�a%ŝճf�kݦ{Fw�xv�wc��F�qGNPڧNA9$���,��Ձ���~���K7ѯ8�|䪩����ڄf�5�@��~����t�J���CU��3}u`kw�/U���{ذ������q5#Lq�*��RY����,��Հ�*�!�aDd-)�~��K���6���m��t�N9RP���n��؀�֡ n7h7O���ULۓms�<��]��0�g��Q�ݧջs��[�-����>Νm6Bn���@fkP�7���H�Ӎ�`��JI���sn��r���6����Q
g_�� �w��;%�R]ApWU� ���mB��mՀwV�lt��l�nI,=Q9�ބ��� ����R8�9���Nw&��U�r����� {�x ���G�D I$D(�t�	�-�Mwm�5�]��#�M [�h)��2�m�e�l��ֺ��G�r�+I٭�b�M�H�q���S9��(rw'bR�	�nǮ���n�i6����=�P:(��N[��Fuj5Zb榻��b��ix5rj�5��ۛ�n!pܴ�u��<>t<�ʝ�M7!Y��8����uћ�ۘ�[&ڒ�=�����t�7a�n���r��߿=������~��{Ih{W3��=��Wzfa�s���ݸ95�q]��e�՞8�����k�q�@���~��������k�~��N&��rU�gwe�}�ـ|�ـ}��Y伪�~=�!55J�]�5Wh_�րǶ�{�s]ŀn7,�х4S���I��م����XwvX�ݖ��Ө�F1H�j�f�������@c֡�~w�b߆���;d�=�\g=d���<��i�����|/3ܓ��MmR�]x����9����@���m��j5�qӔ6�B��K �����v�U+�dL}VK�b٭B �n���"?�C��O����N6�rX���`w��V�ݖ�����:H|[N��B��D$�w����׀|��=�`�K+i)S���8ܕ`��`~Y����|`|�,�B��*�U�����qs�-��Mq9k��ĭ�ey0�׏S���L[Z��$@�n�� ����zXܶ 3P�7��2YE�VM]UM]���frIDDɻ݋ �^ w���UU_�����N�u)��F�Bp���`�k�3�	B��@D)�0��Т&"67t{�^�u� r����Z	WV�����;�׀�׀}�`z!D��~X���v��UT��"j�� f7h�n���n�(@��`|��4h�i0�1EIT�>�X�c��1�%����YlO�a��n�'��}��������v�cjf�@�����KiԤʃR����r>��ݷh1�@{���l9&����:��`�l��vXwf�����6@�eN9cRK �ww�O=��rI=���I��tH*�j��w���3FFT��MI`{��'w����h1�@z2)��4;�^xN��ˤ5����0�����eы�;��0ݼ;C7=/\�ݥ�m�cv�3��ݠ3� ��S�:%��9,�ݖ����٥�w���\H<�����C���ݠ��@f;b �n�cv�ͭ�RH�9)����,�_� ����}�w��$����"$��w���k¤�=N�&B����vX��������>��0�JT@�"D\.[��������[�޵4q�V��n#nwvx�'E-����l�Q*��X�c[=F�Y��9���nf8�v��kXT����������z�Rۈح3:�ʯBD�nծ"�lI��:{:���5g��^�^�أ�q!dN܆[�M��^FDaZ$��U�^;]�d��cj2g\��v�Y�:0�;�lb㞋��nI�]�Y+�w�N��C��To�����X�c�qO/�gv��`�ckl�]��nsawG�1]�=��H]��M'=U]��v�3�c� ����QmM�8�p��;��~��Fg�� ����w�����4LdeJ�H*���v��ݠ�v�3�˺��F�S(�ȓ��w���;�v�3���^���������*j� fk��ݠ=��@���X)�U^a鄨DP�
�Pr5s$97c�\�刲%圁u�s{=�M�+���f������u�=��@d�t�35���H��s���nK���_+����P�T�| ����'/���}��`��;�։4�m:��Piʰ2q�@�� f7hcj�3��)Q܍S�ܖ��� �we��via��Y���;�(�M!6T��rK �n���3yq���@���������Iv��k>�ƈr%�H��0��N݇=W�r9�"6E��I�����tѧ9�AUwx���@�� �����h���:�ԦQ�'����U)�׀��脢?H}�|`;�L�LtJQ�rX{�,�ݖn�lL!'�J |��P�H�&![�r!�	�
x{1��|b�F/�d������5v-cL����5���`rF�p�(��p�h��5M3�,|�$N�}� '9ѷ�N!Cp�1�{�pL'Dh��(~U/ `G@kC�� ;
pMT$5������#���}�P�}�
�Uh��=�b�"�("��w�����Cnj�]�C������r�������ŀw����^j�;�t�99)���76؀��������Pcv�mۻ;����y��k��x�ڂV��-�n��¾Pѽ���97K����n�`�n�u�Pcw���� 7jeǐ�DTr5N�rXk�V���3&�����*�;�Qz�CmT��۹@�ր��b'��7(c�R����,=Kwoŀf{��w;��>���\ȃ�qq+
>�U� ���y��y}�t�7R�9DnA8X]�v��U�w����ɥ�ܪx6�O��dO�:M�Ssfp�ݳC�-�d��n��9.:c�O�ھ�$⎉@�9CNN������;��`fd��;��`���(m��D�V�ݠ7v؀3��7+�}�L�}�#������rX�<X{�,����V n�_���C_+�%M�J����؃�;�ր�o� f7h:>�q��`f4��IJ���j�F�>Y���n��jcv�q�A����A\)W+l�J���E�P�j�$��ܔ�g��m�l�T�\vSЮ񃁵��ͷ��2FoF�K8y�Hn����rn�������vɝ�{N��ll�jFֶ�����;�T8[F���kG�'NF��ڞ�4;���W�]H��9�4��;"��I����T�]�L��pcJò�8�mv��e�k���k�r�c-��`�̯[NW6�tɶfM3%�{��p��i.�I�Z���v"-��2#2��K���i���j�0d�E�	��>>>�2�^����m�t�P�jcv���@c�UE9RDۑXfmՀw����fk�>����B^I*�e�yR��j��UvM���z�Ӻ�%�̨��o���]X�t20�c��9,=Q脫o����zp�m���u��z�(m��G$vz�U���s����� ���HN��t蚂����;okk��ԍ�N��t�0ay���6y�@B{r���`�8(�q𓒘�n;�ɥ�w�� �:�z"G��|`>WU�J�E���n�I'����hb� ���"D�z+���6���rI�=<X̚X֖h%*"���u�����m������ ����Qm4�ک��'��r�\Y��|`���z)��u`<u*�(W��9��K ���囮�������!G5
S�A!M��r\�]ڤu��0��v��;�z�P�D]bk�V���%(܂p���>Y���M=_ ����=��t�h�c��9,�7H{l@f������=U]Qhn�9#�;=�Ł�ɥ��\�P�
P��E�����M����Q𓒘М,=T�f�X��v-�vw&���oSC��n��+g�� �P�s���0u�p���n_���][�{r�nk�fz��N�7��q����tV���|���4�����y� 1����g����Hm��q8ґ�ܚ_���{�`j�y��5���[eH87��,ך�;�,�%���`g�x�5n��Q��l��r�"���:��s�O{��rO*D��ʱ*�d� ����
9UU_>}U�9_y��X��N0��Jn੫�N�HѼ�]wJ �n���;��W�$T��c!Q�1�(7��ufp�]��뎙�q�'���
d�%	��W4A3W^y��nP�w�>��Hl�y���<��%JcBp�;�uX?7Xӭ���f~��/D+���}U)�&
�l�yo����w������?+:��R�"IdM�`uf�;�4�;�uX{����樽M!��r	��vw&�q�w]�}߻��_��
�{�ozn�6�.l��
�GAlt�͊�%�"��b���v�nǛ��6]��A�v�nՠ�+1�1v�;��P�6S��֬(k7�1cR%�Xt.䀁ٗ*jKkW�ꠠ�f�+<s��u��<���.��v���i��Is����;��9��v�dvgf�;<7�������5Na��8n��#)Cs�+iJ�S�M���[ܶ�{�{��o����krm�q��ۊ��,�ã�9�u��O������n߾w�}�A����@�=�1wu�nl�;�4�>[�iҎ�%(ܡH�]n�^��>{l�5ֹ�D�v�ʕ[Ω�4�v��K��K=T��w}�`�lZ�*���!�0:""=O����]������w�nl�R���8�'5� �7f k�x۶��"���5EʪR5Eޛ��z�M��f�c���Mۃ���5��!I%5Q�ڒ���G_ w}�`����d���y��δ��
T�ffIw7y$�w��8+T�A�!$B�%�aD�uf��0��p�����i�6�N8��X̚X�\��2|�� >�e����,�ƜL�B�Է�|���K �͖O/�f�rI��s�p����f��� ��h^�@f���������ߟݪ9.�'���ۧ9�#Ñ�sR�%_�����o����\�j��J��;LZ�UU������ـk�s���׀�6��CiӜ�I%���K�$w}<X�},��,ݍ=r��RT�PMY�~�l�z�W�/"P�E
�j U���8�_w��=�M,�ڏRNA����X{�"�|��[��5� ��ـ7�-��*qIn�rXs6X�o��|w�ŀf����*ѻq�nJ���N7Tu#��k�<[��vVעW�ۖ[��4���m�S�'��nM,�f���?|���K�O:�I� ��l��p���L��׀�^��u����?S��N6JQ��`����l��Z��vw�ŀ}����8�)�I4��l�1wu�f�,/�R�"���X�� �Ȥ��D>�3�7���I<���{�%&4��D������`}�4��l��l�>A�Z���N*����'R$H���L�Bk7C��j�]���1֥f帥N66�>͚Xw6Xs6{���v���RA���9"�?UUqg>���� ����5�s�Q'7s<���$m���`�zX���׺���,�"�m�����F���{� }]Ӏ=w��I%U��� ������T��m����U�չ� 5�x������	,D$��Jb��/G���H��Ȁ��0�a�	����!䉆�b'O0e[�0�"����`A�ht�a�c
w�����H`���MU�^�"D����>���=`��~Q⇀e_p52 hA�|N�|\��{��ob���\0sgPM^,&�`%,��;��2�HS.���� <��H ��#D_S��̬�b�%P��c_<�CGΏ��(F2ғ�n����͹37]���g���2Hqt��ѹt���;Z��n�J�k��]��TjI��E��Wl�m���a!ĝ�D��4cʪ�u�n�&��Q�c���="r2�e	6�$����԰U�qʰ�΂�8r���	)�G��[B8ѳ��Zt���
� f��ճ��(	ֈ�I
���Hcn��! xA�9:�c��<۰:�
X5��g�f�v؋�=��s�����w<XƜ� �v�7�n���!R����
�T�h��KG*�sA�u�R�ð:L4#�,����T�����Ishꑷ[��Y��Q����ʇE�ų¼Rg�ĒhX6$8����	h!�Xz:� �k���9���	i�Z�\v�m��Be&��bq��q�*R]�%8rԫnͨպ5]*1 �*�I�@4�n�eh�qD��뀝� ���=�P�k-ӮͷZ�-ƚf�rq�1қ;�OE�'���w�ALY��	�D�h�5�)S(\ ��uja��VX�\n(^S��T�qr�;z�'���v՘��Y��F�#h$w7g�h
�xpTձt�2����N�`.�j1������kAn��ӧ[�۵s�h����x�3%ecC�F�yd0]7s�,��qF0��۲�Wm��,gj�h+�� �.p�&(��^U��bd���8��O�yoa�v�����g�9n�k�2i�qZ7aŊ���͝���Xrj�m�kM=N֜�a����<Mnv�,��4��u+�p�J����'XY5�t������s�ۛ��fèl�F�۶r�ז���7��лB<�hC9��,�w:�t$:�k:z	���B���-F�`vj��)N��j�T��V�'m�2���k�v]���<u!n��8��
�6�d+`Z�v[��]Z� f
]ۘ2s����f��R �#�N��l�
�6ل��QU���	��_����N�Ep��X ����ꈡ�Ǣ�}��������o8�/m֓�bh)�'"D��T�U^C0�n����B�,�:�v ��r��7B��L3�	��m��n�{=� ���Bo.�N,m�!.���p�k;;����&n�u�^&��u������۝u�tX�VXv��ڦ��g]̼����)�Kg�2�ɛ$\F2v��닛sgb,n�]̞=n{Ok�u���  �n�߻�z�v�@Ŏ'�	���Ѥ2N������En�
��ܳ��P��$29)�n�%(�9�|���5��6~n���$���W�8��yU�-�NSR���3we��3]���U�owe���w�m/8
�ӧ9�K�wJ]7([v�3[���TS�M�RT�qI��{��3we�w7fD$�E>���'u�3wd�VJ�]���� �_u��wN��s�z��t��$��P�����RI����v�5�R����J�4ܜ@����>�>��ѪIt''@7߿K5���W�������ؽM��u9"N
9,׮VDB�|������m5(u�@����GV�t��T��'
m�`f�yX6� �[ŀk�� 7u�WT�*�St��Xn�1f�5fk���OyXv��N:#����$)%��7]��]M�~z�� �� �[7���웾���kɽl\[�
�m˨�5pݮ�@k��]�5�o�{�q���y��������`�ـۿ��!�݋ ���g���)*q�����K �ݖwv��Ź��${�zxjH!��' �>�6�"��������~؈�s��`n����ȖԤ�N'#m�NK�Ģ�vq�9�Հn�fB^U]������M��u9"N!H�[��ݚXnl�7^�;KscbR���˭N�LㄸcM��8�P������t�{kmMdݏ[�:v�T���4���=�O����g�H9�Հ�R��\U����z�:"&N��X�}X��,��R:Q�NSR���`fn�X-�@cv���@��S.��`�:s��*�Ź������3se�y���? x����}�y��'�����a$�%N66�;�4���`���Ź���쭔0�p�J9Q�8��msUyv�Cur�y�nۨ¾PI���wκ+܍��� �͖��,[����,ǈ�	J��$M�nK �ݼ�L�{���0[w��>��SUM:��N2IV�o���٥��7��`n��V˦:ؓ*A��P���f k�x�x�:%�>� ��UԺ������Xnl�=�n��W�j���ݚX�YG
�~D%F�Nq�c����ue���v�����4S֨C����k��ÃQ�cqW�g :Տ�4�5WUq�>z�͓�b#�1�"Sz$,��� �KZL=�SN�4�4٪��vq̒��
Aee+n�����H��� ]LZ'��h��{Y�&�zu9E�w\��%}��r�����m�b�N$�u�]AZ���{�������=��+	�S:)���t��,��DݳM]H�ңe3H�ue�)�ID��3}����U�f�� ����ܡҍ:s��*�Ź� ��s�����,�Q	L�k���qI)8N66�3��V��,�۫�3f��Cp ���X�v��mBe�:nP9&ÉR�)�i4�37n�[���ݜ ׮������,�4���nH��7*�k-�p�J7#F�7g�$��o3ࡆ&��m��rA8�%|k����{��;��(K��w�� �}Tz�lWeYW3e���O{������ �E-*�e���D=57�$�����y��g �=�`��q�S��r2I�w[�u�0�u�8�wN =�5WtG9MJJ'%���K���U�f�� �����!$�t�N��Htܠz�����pE'i:�ɮ}����Z�-T����뵲gy	��5��̄�7U�^D~�~�)�@��u�/] 7]������8'$V��,�6��Ź��ś����#+i)Q�NK�����߻��<�b�b��"��_�(�=�����g$�����ض�Ӧ�rA8���?-~�;���]�1����a��"�*.l&�:� z��������S����F�8���'��hã�Uf٧�O7sn���,�ˤ���۞�<�wwH^�@7����H/] �R�rQT�5)(���M/+͇������9���v�Z�bI�J�&��`�}X��`�w�6�U��qGOd�*I8�Cq�~���y����y$���I�|IP_DT�޻3f��)�p��q�n;@cmBe�ηH�&�7�'C��iC��O��Xvg�(α��j��prm����&�?�tA����=~����v,e�g[�~�>�w�yQ4�u9 �M�V-�v,�v��,������k�D�R����I���R ��hm�@l�@�⮝N6ND�$�; �se��ݺ�1w5�z�����wh�Q%�NSR���`cmBg5�g[���>����	�����f�f��%�^z�R�5�(��8�Mn�Ǭ`�9��~����vM������S��]爎6�I���%����W;vkc�K�3��jx�"�C�R��Ry1Ɨn��Pt����b�<ۮSuU�ΡNh&B-�����㳊�]CԨl6�v�:��A���OB/u��ml�{n
L�d�h��۵�쵶�plg�����@P�[4����f�̙;y{���Vbwfpn�\r��)�8tpfwǛj)����G������ś��>����UW�3��Ձ��򒤔��n��P:� 6�����+��UI�<1�H����՞�>m�ÔB�ޮ�����7��-*(�)cq��۫��U��7]��7]�޽[I&�u9 �M�Vu�(t���9}Ԁ�ڄ�;��om����8��V�3(��5�J�cH�F�%��۝'*�(�R1��&T��(4�1f� 6u�@cmB7(��U�E�U5ۺn���$�_���,#T�8�G����!6� <�@l�t�d7`}D�G9MJB�;=�]X׺�Y��Y����ŮA�m:s��*��M�g[�ηHm�@y��V�*IJI�ڊE`b��`b��`wwn���Vk6!�R9�#�%����8�m<���׫�Mۃ�XK����CsrV�r�nn;n���u`w^�1f�1uj�n� ��1��m�@c�����g[�e9p�i�S�
Dܕ`w^�1f�T�>�>�� � �0$�!R :$ �E��0�/8�9HX@�RK �*h@`F�l��0��ف�	i��i�k$
��w�}�������e̊��P��$ z�{�ThR�B��Q$w�s�����D׻�R�,il(,"�Y�+
]���BB`
âpO����W��|���A�0 �H��P=P�:5(QSD�}����'�ͺ�s��$ux�^�2�GQA����� f�hm�@f�r�=��]TN6NE%I$��;������XǺ�Y��Uwf�D�SR��GD����p�`yPkT��O����v�����} �:��t� �5)(ܝ~�u`w�1f���|�����ei�(N��q�@f�r��������P�������t����R+ �ݖ�ݖwv���{��\�U$w6x�ʉ�c�"rX}\��URY�zKI%�����I-��,��'�>�����y������:S�%I9%�����_|�[�m�Kn��I$�vKI%��U�kJ���..w�v��l�\f�/��r��g΄��s#�cB\�:�b���~�����|�IfnϾI!n떒K���}�I3S��B�GQR�R��K3v}��\�Sm}�-$�{����$�^�+�Sm%�����Ru9��O�I!o�夒���_|���9�ZI%��O�I!Wk6�t� �5)(�r�Iww~��I,�4V�IfnϾI!f떒It�:���:s��r��$�\�ZI/r��;Ԓ��ZI.��Ǟ[n9�zb�(�b'��ߟ��u^v���cu��9�SF���c�ַ.�l���X��	�X:�NJ3��vsc#�JT��Yy�1��]zmy�<�e��/[�@�S��#��ɧ�g�]�03���q[���a��sOT�Z:u$� ��9��'6�dڎZ�_%��+ӡ`�N��CX���2�R<�R2��f-f��Z�G������t\nC�BcC����C�ߞ�{�}ww�gY9�9�ɽ[�t�6�*���'�	멈�ą�.1:����������c� [����n�i$���W�$�k�+I%���ӕ��	��H[�夒���_|�[�h�$��ݟ|�Y�[�N� ��RN9i$���W�$��+I$�7g�$��u�I$�իi*Hu8�M�_|��ʮW�/´�Kwޟ|�B��-$�ww���:f�w�J�
����Y���H[�夒���_|�[�h� ?]��?{~�^-�<r�!�s�]D�&��\V�vH�nY�e�I�΀k�m�u�I#��H[�夒���_|�[�h��y�m������/{g�w�6f�t�nno-������;��(|'��}�{�ZI%��>�$���ZI%Ӹ�\rP�:s��r��$�^�+I$�7g�$��u�I%�����$���v�$T����NR���M��z}�I��K���}�In��V�K���ӕ�4�#r}�Iw\��]�߫�In͊�I,���Wz�_������.������� �'-=��u������"U.�y��ZW��[CHRN9i$����In�%��Y����$���i$�{�[��N���*�I%�6+�9ʦ�Ksޟ|�G�<KI%�������Ef�2�P�Q�Q(REi$�罾ym�����O��@i @� 7�|�!W﹞s�<�����o-��=Ǩ�T�d�RG$��^k޿�Ig��W�$�ݛ�3����f#jGJ8�ȩ��&�@c֡ kn��v��w���݇���:���T�D8۪nR�-�$ۧH�1��Pu�Yɋ����&�UÒ��늛�����@��[j�n��h1�J�t�RK �͗�L��b�;�b�>t��D���ʚ�s#p�!��u`n��Y�q,����{��`}�5���@$�%MIV��ߖ�]Ӏ�>��YIFV����V�VhĨN�����{M� o]��� 7���.���Wn�Γ�n3�]0M��%ʜp�N���u��P0���^�w]Zۨ�m��h��@�:nPsi�u58�9q�I`fn�X�l�;�uX�l�1fRڒR���Ԥ�r��v��M� o]�7[P��Q4�*Lc�9ܖu� �͖f�,=I{��`n��d�T��(�"����$�g��}� ��s�j���- ?D(A@p�@�`�Ǽm� ���� n��b�xr�"m���̒��x���\�{0mf�m���Gˎ6��p�[R�q�Hu�<ە���IY�qd'�ul�ػky�)ĩ���-WB�;�f�nŌ9B=@k׶dN���ܜ�1v�V�l'.'.�mͷd؀��=���ƚ����3ĂN�	�m��1�Z����$�7ql��].�[ �v3�"^�>�{���e�� 66��t�Ƕ8�S�4b%.���t��Й<��݇���,�\�[l���Zw���]Ͽ/�oWt�K�����n�0P	$�P�,�۫�$>����׀kv�p��OӬ�e	�ゑ9%X�uX�l�3vi`n��X]Ů�$ʕ!(!��7q�[� ֡�����rU��QG$�n�,�۫5� �͖ʰ=�!j�\#r��(�Vn�E+��t�f��͍g�ܷ���&�f�긌��Ԥ�!������{��7se���K Ӹ�=�Rc9�MIVm7+Ѫ���������5�b�jfm4�rRn����7se��M��j�@{u��������˫��7(��@۴�g����|�Z`�E$iSn+w6��>m� 7���npJ��WD�.Β]g��$i�i�#qQ�'Mqv�sŞ_m�z���鐡�Ӄ�:�pR'$��3�����v���H6�,�X�f���.ົ@�Ven�wZ���`j�=A�M���2I,Ǻ����䂂���#����|��|���y$�}��$�^ඤ�� �5)%V�mՀwwf 7��9B��p�_Z���SEW�n� |ۼ�B�����p�n���rDT�$7
ht�s�bݚ���+Z��RV�bq����������j*������ ޻@n�r�oZ���,��mF@n �8B9,Ǻ���@۴ ޻]��2f���M@�D�iSn+��]XwvX�l�3�>ךA*��%'$� �� o]����t�_��)LdDG-�����`mwE�q&T�R�Q�����ܠ֡ cn�������b���Fsp��:0:9�s$/�m�ݓ��4t�tv�C����N6J�H��3�׋ >m�(�� w>�βy]ڛ�SR�Q�`n��_���,��K1� �Y���*Lcs�����ݠ��v��z� 75�B���Q!DԒ�7se��d���ͺ��6Xfij!�I t���>̶`�ŀ�]�z� !)��!AU�C�'�BL
$�I!������ ��3�E�c��/���>4O� �F& i��j>b>� �O��ā�MP�����,�0 S����p��z�i)!FS�~�BO�`�x�=���)��͆�DϏ<Eg�P8�/_'��\����=J?$	�	�@}�y)�O���j�|��F�:D�􃦄#��a� aK1�"N�=�����w���F�p� ��X�/Yћ�X����.yd�b)�=��a�C���A�;��'m<d2J�k��b�@`S!���CXU�%�[`.Pc�xml'�a�����n�E�o:E�-�6u�
�ɑ�!���a�2�P��(���Shݒ	yKl�rضu$�Jr�,Sc��9�^�4�,�${6�����WZ�:�޺�D�Il��[�N;n�J[�H	���02�k���\)�Bm��F��{���������/W['954Q-er��ِ袬�mJ�c,<����U*�2Q]vqt��e����8mc�tTd���d�u4��6��e$u�'�s�u��D��ӭ�L.Dt����^���!����k�֨�Ĝr瓮�d�%t�V	�v3�lC��!��,��ѱ��+Gi瑩x�R-����� B��	�ΑV����P����Q#h���w��Mj�!u��6$�4Q"��lteT-ӧk�d.`�Hsڮc��Ӎ(v͑�r���.�VyV2	g�=Za��cb�E����.cH6�{�F�YuK�sϮ,�(�+ZD� W�n�\b�V]1	�un' t���#���ӹ�xHr��"�҆�;1��iM��y��;<m ]g�G:��z� ��'�7E�:�|�h��K��:��g7���n�9�ɣv�S`*��V�.3�N�����[J�[Y����nC�="��eYβ�#��V�A.6�e��l0��Va�+gi����t�p�K`4��:if$�Kq�:ئ=���J���m�\Ꭴ��e�1	۹�*q[$�Th|�k����XZ;rc��O&�kֶF-�OAT��Pw,Iӣv�v���Zf򚣧���윲�V�ADYG�����:\�ق&U^:@�٭Ha)K4���:�&x��,p쬎���	�U�@�I�,�2�s�&}X؃j���2��WC��8�$��u%������єv��mI��&��J�P>T<<����A����O�>>�E 4/��@P�~:�3d��喹�۲ݮ6�m�����e��i��=2A�R�B�Y�l�Ns�yI��L��z6�b��0 �:��Ȏ�U5��m���۱to[�#Mgul�lձƻ'M�.ɦ�C�\�j�L2-'j�m�B����n4�Hl	��j�@h\���õ��cJÑ�ppv�a�0��We���Y����|齧X���u�n%�� �F����o����G�dg���V&�>;��u;%�+��9���89;t�zD
S8��`�E$iBH`�۫ �3e�}����2i`o^kT�	�を�rU�{u� ���m�ۮ�艑�t󫉰�R�#��;��`}�4��Uĺ�|�����q�8�N6J�89��@{v؀��@�v�=����-�%(�r���r�3]����_�1���m��#��p\U��[r�Ě답7i�葮��qλg��;u�Ϋv̔RJNH�1��A9�}����fk�>̚X,�v{�ԑ�莐�˻��O>���C����?�`R�� �B��3���rI���s��6_��r��3}�B�q�t���1�� n�hۮ�6���mU�B���	!a��8��,���,�v]ݿ秛��N�������h�� =�l@���6�=��n��ήx�s���FYU��2qt��z��=;]�Kv�Fl�H�u֧k���Kn�ݶ 7[Q�DG�o���5��n6J�8H��&��(Jd��ŀ7׀~��Y�29�O*��8���&܅���]Xٛ,�9UU��A��'OS�r������NI՛)9"��79� �3e����`}�4�>�۫��&;�8菉GSwhN��菾���bu��6X���eNG���`�8.
�NB�OT�bZv��g���\�.��ME�ƛdUU�۶��7(ۮ�-�;����J�$iBHX�u_� �論���>̚Xܚ�%Bu8द���>��`un�>̚X�uX��i��P��(�KR��y�7|`�ف��%���J(���^w5X.��q��l�u)���e���mk�Kn��.GU��E�ڍ˸��6�U�S+ĉ�dD��gv;c^7\֜]W�p�o������r������b {:�n�l�nr8�,��W��8��}�`w�<XǺ��5��NJ��ND������b:>�>����>�nm�D8��:p��vw&�sf���U�՛���n���J�$iE�؀�v��k�Kn��l@TK ��;�M�npݚ[p��e�"}��)1:��S�G�S��{ly�e�!��eY�s��	���8�Q�vᩫL������ӷQp��<ܓnXh����tG�ĵ��7fcZ���.a牎x��p����k
�f���W:.՚�l���#mGl�Y�����|�s������	C�ݷd�Vʳ�E:�L0�nfakn��\��Gub�fs�Իkgt^^/m�c=l�����b�8eg�ў��<�u2�v��nZ�4��(�� 76؀�v�f�i��	)�F�:�u��͞,�O��U����5��n�%E%�WwH��@n�bε�%�H]�mI)G�Ԥ���36i`}�\�N�X
D�y�ΟZ��S`�79R��U�՛�������l��Ջ*�1EƩӉ�Q
�@1���.[���ԼmLF�$.���@��tإG�NE`uf�3�4�;�4�>ך���D8����M8��M/�(�1���$S����M�'[�=t��@���*�B��l���^j���K�����������*��"n���k�N�HͶ 3i�@6n�����E�����`gri`w�>ך���k�ܦ�;j��7r�cDOc3:�j�v����z1�dr�r�R��r;;�K��V�ֹ�>�n��P��������\Ԧ�G$��3_�����7]��d���y����1���Xc�W$����'�'���%D	 U�4B�^Q���R1஡��L�����'���rC��cnӃ���'"�>Y���&�s&��.��+w޶)I�G��*j���b7m�mk��[������?���� \���q��V��e����[B���G����湀�u=�k��l��������ӭ�}���Ł����h��"n8Xc�W�rd�}Ԁ��n��,U5Aa	E���f�>̚X̚Xc�V˸���j0Q�nGa�R���kw�������	tA"�#J�$a�	 E�G�)��s����RJQ��5 �rs&�N������9ı,O3��8�D�,K�of�"X�%��^��ٓ���g�w޺�8��������#m0�H�Y團���Íu���r�9�zf������ı?����ND�,K����'�,K���{19ı,O~���O"�oq�߿���響��9i�ﷸ�bX�g��q<�bX�'g�ىȖ%�b{����yı,N��܉ȟ�r��G+w�����#�$�M8��ʱ,K������bX�'�}��'�,K��}�Ȝ�bX�'��{�O"X�%������%�4�������,K������%�bX�ϻ��,K��>�s��K��#2'����Vr��G)�g��t�'S�D�{8�D�,K��w"r%�bX~>�~�'�,K��;��'"X�%���s���Kı*D4���/
�)W�R^���G��*n��0�k��e]e%��ܼ#kWmVM���Ǫ������7#m#���VJb����7l�fϜ�ݝ gm�_��N�s��T�Gbv8�n"[���K��΀�k�Խ�n�����nn^a�vHוyr��QH'&p�b��qnL�:�[98�nn�ٵ��a�(y@��!�D7�bs(6	�)4�"2-�9�y_�U���+��Wnsε;��/d�lM�Ë�rvCn������]�l���ŕ�kkS�e���X�%�����O"X�%���y�Ȗ%�b{����yı,N��܉Ȗ%�by�����5�6�s37s��Kı;>�19ı,O~���O"X�%�����9ı,O3��8�D�,K�Szn�w6�wff�n'"X�%���s���Kı;�wr'"X�%��}��Ȗ%�bv}�brr��G)���u��1��G��ı,N��܉Ȗ%�by�w���%�bX>��jr%�`�"}���q<��r��G+w͍��	*>8��g*�%�by�w���%�bX>��jr%�bX���;8�D�,K����9ı,H������K7rHf�4�f���5.�õ�4��^k7v�L� !sۅ7=uu��k��sfY�����	 ��q6	 �{��8$�H>{���K��>�s��Kı>��Nnrm�����n�"X�%���s���=U�2(Pw� 1�O"X�gnD�Kı>���q<�bX���n�"9S"X����م�\5ݙ�s7vq<�bX�'��ۑ9ı,O3��8�D�,K���S�,K������%�bX=��snd��6�n���ND�,K����'�,K��>���Kı=��vq<�bX�dO���"r%�bX�����6�f�.fə��O"X�%��}۩Ȗ%�a�#�y���{ı,O���"r%�bX����q<�bX�z���_�}�v�����Ғ��:�uOi��z<��p�ӯV%��՗;RlȖ%�b{�y�q<�bX�'��w"r%�bX�g�w8ȩ=��,Kc�)ʳ��R9H�g��Ғ���79&n��yı,Os��D�Kı<�~�q<�bX���n�"X�%��s���Kı>�s%�3�L�q�ə��9ı,O3߻�O"X�%��}۩Ȗ4>�}���"�u"TB�(a�#��HM�� |� ���t]�No�����IP��H!`Ed�I$TO�9��{��D���5�&`��}4�P�Z�D��&����0(uE9j�e)��	׍Q= "BG�!��! ����@t8)�$`I]�	#>b���b�ƌ �}��T4�bH�A0`���2�9�g,~��z�(�a������q��fP���8S�r" }�P��A>S�Ѓ �`EP����"uV(�U��u8x���� xa�o����!ȀtS����H�g��)޸��!�P�蝉����p?�V{"X����u9ı)���y����"p��w���#��U@�?o]ND�,K߻�Ӊ�Kİ}ϻu9İ? �"{�w�q<�bX�~0��nɶni�w7n�"X�%��wÉ�Kİ{��jr%�bX�g�w8�D�,K��n�"X�9H�v�3v��!@�G��Dbq��z��5�Xzk����$ûm���d���nƖ^��[0���Ӊ�Kİ{��jr%�bX�g�w8�D�,K��n��g�2%�b{�xq<�bX����9r�n�i���͚��bX�'����'�,K��}۩Ȗ%�by����yı,�����bX�'��s���rͲZf�ws��Kİ{�v�r%�bX�{�|8�D�,K�of�"X�%��{�s��Kı;���w6��]�sssn�"X�%��wÉ�Kİ{��j~�D�,Os���'�,K��@}"/���`��N�Q������Ȗ%�b{߼�SP�� ���_�r��Es~��ND�,K����Ȗ%�`�>���Kı<�~�q<�bX�'������)�a5y5�d�=vku��=!a�`nkz���H����i�s]��z-��D�,K������Kİ{�v�r%�bX�g�w8�g�2%�b��\���$)!Ii�T�mU�T�ʸe��'�,K��}۩�~U�DȖ'��gȖ%�b~����,Kľ{�w��O�S"X�N�9��3d�74ۻ��S�,K��>���yı,N����,Kľ{�w��Kİ{�v�r%�bX����al�wf�ww8�D�,�������'"X�%�}�����Kİ{�v�r%�bX�g�w8�D�,K�w��I����nm�Ȗ%�b_=����%�bX=ϻu9ı,O3߻�O"X�%�߷�br%�bX'�`�?N_��ֺ]Z�.��-�{t��r��=����#p=��U��j����� ����s��YФJ�rbW�F�����nҏn�,�Z����)�ct:Ep��i�D�h]mi۫�M���?������Σ�����a�l,!#��.�֛��u��GW ɰ&ks��]r�!����6�#����U�+k����]əL�nI�(��!W09�ͽY1����ӧvgq�,�y�[{p�=^��]m��Y�
؆�k�g~�ߛŉbX?��S�,K��߻���%�bX��{��O"dKľ�����{��7��������7%a���Ȗ%�by����yı,N����,Kľ{�w��Kİ{�v�r'�PL��,O�~�L��&L��l.n�Ȗ%�b~����,Kľ{�w��Kİ{�v�r%�bX�߾��<�bX�'ݗ�a��3.���m���,Kľ}��Ȗ%�`�>���Kı/�}��yı,N��ʳ��R9H�c�֊�q҃�n�<�bX�s��ND�,K����'�,K���ݱ9ı,K����<�bX�'��v^d˺��M˔ީ�ݜ�!4�Ð�e#Y�\<����t`�#3��H��A^狀�u��=����wx�D�,K�ov��Kı/�w���%�bX=ϻu9ı,N���R�.���,���yı,N��������Q��'�,K�|�x�D�,K�w���Kı>Ͼ�q<�bX�~�˔�vMɹ�6��Kı/��w��Kİ{�v�r%�bX�g�w8�D�,K�ov��Kı<�{���5�4���.n�Ȗ%�`�>���Kı>Ͼ�q<�bX�'~��Ȗ%�b_;��Ȗ%�b ��Ο�.��4�we��ͺ�D�,K����'�,K��۝�9ı,K�{��yı,�ݺ��bX�'�>����{r�6���ͷ7k�՘��m��ݹ�c;)�8v�ۑ��jNK���y��3��~����{�������Kı/��w��Kİ{�v�r%�bX�g�w8�D�,K���3%��˦㻛w6��Kı/��w��Kİ{�v�r%�bX�g�w8�D�,K�nv��O���)�su��Dh����|��R9J%����S�,K��>����%�Z/��"?�)�࣡�.���'�sdND�,K��߷��Kİwt�Q��DG ��)ʳ��R9H�f}�s��Kı;�y�'"X�%�|�{�O"X�%����S�,K���r�p�v]�L��'�,K����Ȝ�bX��������%�bX?����"X�%��}�s��Kıwm
ʇ
��J�LBCPII,.�Y�!�N`ڮ�շ#m�]�)2�	�V��ә�"r%�bX������%�bX=ϻu9ı,O�ﻜO"X�%�߻͑9ı,K罽��5�iK��\��'�,K��}۩Ȗ%�b}�}��yı,N��l�Ȗ%�b_;�/���G)�r�fV�GILR
G��S�,K��>����%�bX�����,Kľw��'�,K��}۩Ȗ%�bw�S��7Hf\3]����yı,N��l�Ȗ%�b_;��Ȗ%�`�>���K��F'�@�C�7�D��
�t\�O��}�'�,K����	�o77.��˻7vD�Kı/��w��Kİ�V����Kı;����yı,N��l�Ȗ%�bu�{|����g;(ǟ�����]R��T@���5ہ��&&+R��&#1������~����{�=ϻu9ı,O�ﻜO"X�%�߻͐?șı/��~�'�,KG+�/Z�(p"#�R9	ʳ��R8X�g�w8�D�,K�w�"r%�bX������%�bX=�{59� �TȖ'����\5ݛ�Y����%�bX����"r%�bX������%���D�?����"X�%���gȖ%�`��᜹d7a��vffȜ�bY�D�~��O"X�%����jr%�bX�g�w8�D�,K�w�"r%�bX��{{3nk0Җ�ܹ��O"X�%�߷�S�,K��>����%�bX�����,Kľw��'�,K���Rt���i	��AY3�3,۪:�4V{�v";w��!�󂝃�նu��*Z(!_�t�ƕ�%�U8��//]��Ǯ
<�.��nDE^��0�A�c�����p��I){W�����ه��T�P� P�F���Ц�F[$k�W6�bX���G�1i��	n��ۓZ��v��<肄�O��t�nh�LS�E>A�h�p�=����i��5ٍ�nؐ.m-L���"_ǭI�P��gv= �9�U��3q�RSR=ߴ�X�%��������%�bX�����,Kľw��'�,K���٩Ȗ%��ȟ�v���n�̸f������%�bX����"r%�bX������%�bX=�{59ı,O�ﻜO"�oq����?��OEf��}�X�%�|�{�O"X�%�߷�S�,K��>����%�bX������G)�{�ТDj$��W�*ı,�����bX�'����'�,K����Ȝ�bX�%���<�NR9H�nK"9#���9J%�b}�}��yı,N��l�Ȗ%�b_;��Ȗ%�`�����Kı?(�����7i�nK�1�]r؁�������h�͂���Y�tfݴ*Q;Zkpv�k�.l�7s��%�bX����"r%�bX������%�bX=�{4?)<��,K����'�,K����g.Y�m�]���'"X�%�|�{�O!�*{��H���>�+�0E���6%��w���Kı?g~�'�,K����Ȝ�bX�'��s�6�)n�����yı,�����bX�'����'�,K����Ȝ�bX�'���8�D�,C{�3���:c��T0ֽ�oq���b}�}��yı,O~��Ȗ%�by��s��Kİ}�{59ı,O�'�w�7fau����'�,K����ڜ�bX�'���8�D�,K߷�S�,K��>����%�bY�����[��y��=+�V��H�vNoC*\�lY�VD���٥�)�sWF�3mND�,K��{�O"X�%���٩Ȗ%�b}�}��yı,N�z�*�R9H�#��wZC��D�����%�bX>�����bX�'����'�,K����ڜ�bX�%m��_�RB���F�Yvar]Z.�sf�"X�%���{�O"X�%��۝�9����+���`@C��=�y����%�bX>�MND�,K�w��[.��74�7s��Kı/�gv�"X�%�{��x�D�,K߷�S�,K��w��'�,K������݆ۦ���ڜ�bX�%�~��<�bX��of�"X�%�����'�,Kľ��ڜ�bX�'����L.g���1y�6�͒N��ՋS�q��qۖw[��X�Km�ٛsY���w&���Kİ~�����bX�%��wx�D�,K��wjr%�bX�����yı,��5�L�rD�r�g)�r��Y�wx�C���,K�s�S�,KĿw��Ȗ%�`���jr%�bX���^��!���%���'�,Kľ��ڜ�bX�%��wx�D��
�"d�����bX�%��wx�D��oq������1\���9h�}��%��D�����yı,����"X�%�~���'�,K��$0��TB 0�E�!A������Kı;��߲�4ɻ�m͙swx�D�,K߷�S�,K����O"X�%�}���Ȗ%�b_���Ȗ%�b{���4�w3�Єp�fY.�&�Ղݎ������F�X�X.XE��vjm{���x�,O�����%�bX7߻���bX�%����?�{"X����S�,K���߭-��vfn����yı,���NC�r&D�/~��O"X�%��w���Kı>�{�Ȗ%�b{;�^\��۹76��jr%�bX�����yı,~��ND�,K���8�D�,K��sS�,Dr���bǣ����dr_+㔎U�������Kı;����yı,���ND�,K���x�D7���w���q��å*(k^ﷺı,O�����%�bX@?3���A$N���NA$S�s�H$���
����
��@_�@Z" *�� ��" ���@_�DT ?�*"����� �"(��D"� �F"�1Tb(R
�1"�0� �E��D"�1�����B �EEO�@_�D@_� �@Z" *���
��" *�Ј �� ����
��" *�� �� ����
�2��<�`A2�����9�>���     4               (�� 4|= �������APT� *Q�"��(P
 ��AD��H��%E�"A U�    h  @  2�}�w�ݫ�wz��gW��ڞ�y� ��_K��[�o6�Ysjw���w�ޠ�: 1  D�   	�>�  ��`h @ �f�  �   � D �N� X�4   @( � �FE @�4� P��`���	 �E tw2���� ��ԫ�p��yix ��W �  �:@  �{v���r�j�aַ}P ��}�.�j��;�]�u^Z�R� >�  @ A�������޴q�u�'���N�w ����s�����������'����i�,[�>��:� �޷>�[Ň�x�h��V-�U=��M/..��{��>�n����_}���ŗ�v�=S� >�      ��Mr˫nN{z�3���m�o�
H秭�s�|��u��+�n�jz���w����ͥ}��  �x���=�k{�}��|����_O�k��Үp�Eު\�Z_x��w<�^��wJx �      �۠�y��'��/}{����{���6����{Ҝ���v�r��������>�i�ʙ;���j� ��;��o7�S� >�>�NO�<�������rz��� �h�)��X\�����\�zU� 4�Sm%J� h�H��T�@  O��(��F�LD�*�&�*��db41�BT�ԩJ� h ���%)�@G�z	�����a���������O�\��w_*�����@ W@ *p W�� _𪪊� >��=�Q0�����$k��Fa �!��a1�e�F$fg��K���A�$BH�*h!sWZ������A����"R%�4�f��8@��d6�a��^m���Pc�"i�HB�N���X�4�5���f�B�s<��F@ F!�L�$�x�bl:�H�Ȱ��gP3P�8B�YHT��(Q P �#R$a�l�)�Qi�H�)E�kCI�:(�!
��)!	�H��Ba�h�1cII8I$$
ā�ID�Y����I.^\ѸЃX�`A��n2\��Y.��=RG YBR5d$�dedal��z�R�ą�|�rD�)�J�4XBk0e�s4��SE�\0e�L�KtS
FHB�@�XR�)t��V������4��0�bJb¬i9�P�
��
CA+H�ЈE�E`G!!M���\��d��$ a�0)5�$.ow��3�	=���$ja
@����H��5 ����^34h��|<��H@�c�bZd�p&D0H�!B!㭓���&˽]o�<7�!�;&�R!��Ski���9��xI	����0�5Ĭ$����Y�'�.���a��#�u����D#=���0�$���7�5	�m7�l�$$�:���x����
A�aR�4F�nf�����u�����B$B��秩E$�\�0�{��ER!<5��r� ��=5�;10�#C �df����B��[r� �"M4�D��R���z{w���d�Cx�SEcMka.����}0�=׊O-tzH��|1��_�`]Q�>_�.���b�z`ņ�݌���F���f��f��0���$%�$jHB�2@�OH!�,!�Xi�\ ���5�.�Q"R5�d��|=3{�-%,o��`D��B��f�)�<#�@�'<�d.&�y5��hs����7�<��N�	6��Ӊ/7��1cI �5��F8H�}3!��5W�p����G�P���7�9=�I#�	ъE�!Bb�r
�"T#� ��-D� � 0!��1"�=���z��vMS}.J��H��B$G�"E!!�22D��E�6@ȕpcV,p	L4k�2e��� � O�8$�%$���HB,w�9�7sK# �hMl�YL���c	HQ#�Xh�\	r	
b@����wd	R�1cD�
< �B	R52$1�!w�%�f��B�5���Sn3S�d�$���5CRRT�\�7	[
PА,��bF,��=eɫ�D�eξ��#�s'�L��)�r���)�ha�h�(I��I�^�aN�.��f��뚡6�g'/O4�m�k�k=�R4��
a���l�Ha3ۼ�
�4z�!J	�
,�(�)R�)�3l�@5���W�2\�@!�
J&&�����[�k�
��jF�$+
B���<8�afD�/
q��.I���Gz��X�e7�a2���<�<�����0�Ú��#s��&�3zf��A�)���G�7�֒#F$}�YVP�s����k�n�B���@�+	.�S!H`�$��Sc����i�:짔���!A���@�C 6ZR�����u淁���+�Ha�	!��D�"䐄+��v��ᡂ���dB�2A��4kY,��R�p9�h�sr�¹5/��\�7�80)�a!��4B�[7��o���4I@!���lĥ��8�˽��D�$	"Ą��I��w3Щ�DhA`����f���Q�㰖Q��Q���[��x>�oo�).�I�35����M � Ġ¬��VN x�6y$��X$}�I-X�����!��9
f��T��B����0��	cs[=�0�q`F6��H P�S04BD�D,�m�VE��F��J{L%8���&Ķ	�)�E���J���`�w�܉u�߼7d	��g'.�l������5����!X�ccFY!	XX�4&h�Q4��0�HB���S�R��K�r#R4 �W�b�e��k��%� �!J@��.$�<<pq�:W�W� ܔXD�zL<1�%�8B�F��$�)�l�RH-Bvxh�5�������.��<�5�j�X:�0b(��bPLb�X�$��@ "� ��`�JC
�&�p<n8E5\�A�+A�GD��P���<Yw���A��N���#V�$Y1)�Ȥ/��2�5�ײ,���)B�nz�<8Yxq8s��5�zaL	r��(w9Rzf��	L�RB,���h��w32���<�z�VK�r�8f�&0�T���R0��{�3��i�$�)�B�sc3�i��i��B�,�te�5��K/k�[���Ϩ�VJ�ޥ��oRС?V�a��FGRB�B@�0�k� S�>뤥Z18��yJd.1�Y`V-i��#GF�C��7����'�o�]k�l)h�D�Æ˭llM<A������1a��!@�!Tc"���d�"@c���"�@�1H
��A`�jD�A�
H�$�g-$`�$X��{�i��,JH�J�
c��1��#�Q�3�!Lr�eÎ�M�R�#�I��)�MJ*��q��i`�BB�!!,�:Gi�k0�CP�(����\t;"Icrf�ۘ�ӗ7�u�o6j�u2��a(�4���FH�&H�HH��ᤒ\ѳ��HD�I	���Q!n��K0�[`q���j�(1B$K!$k �L��d�q�.���m"PO=��Z�!Q���]�N�������ѾxY����L%�2�_vxn����u�FHS#S�,6<NH=u!A!�cA�,"D��D��P)�jH�Y!Ie��1�#HML�<�@��jŤv
"z��6��0 Y},
�5�cX�a�aHX�4�tB��.�Й�OH2BVXq`@�HQ�H����ޙ�]oV3�q%Yc͑���p&v�s��䏧��d��H���	b��ʹա͞�C�&1����Z5��Ɖ�$�!=�,����=�j0�͞q�x��g5�!��/=4���������g�5�f�)���CE�-aZzā"�,l(@�,a4r\u�+M95�{'����!\��CW0�� H��E�r����׳�c�5���bA�����3�F>�	
Ǉ!�xor^AY�V*�v���^�}B��{���>����H�*�h�ĝ���%��#!\�+][���g�)�sy�!{�:��8эfp�5��M0��,������)��H��BIHH�F��IK!kJB���5��L�e��)X���Iu�$���n����I��]�6ص��7��;��d����������W��=v�E�`�{��ݬ�^��ad�i	I!urI�2�p�H�WC[BP�5C1�u�r��f?F�������?)�G7��I��o���c�1�v����0��H:L�Yᨚu��f��sDt\�]r8�01ӥ�Reg�g�(5R���.��[�bs�c��r�߄�a�ss0s���8���.i.L�����~�{�B�k��±��k���S���@�%b$]�K�|�!N�XG�<�Fp��'c@�G��(B�%7�wА���\��r�h�|aM�w~��o���1�.Jć���0�I0ŅL=	q%�4zk\�'���a��L!�!���4]�L)��Hs��z��e�������6��u{�ם򽙿f�\&��8B5������e0Ӵ!C��)�����ć�%#VI,�� �0H�FX�	�.]i�Fl��0���!P�U��R"�0͓�$�<�U�	HB��A� ȅ�d"P�����@�$d3Z�ZH\`D׆I��gC3{�`,���0�%vI$�Hm�m� m6� �m&��  8  �J�`   �  � *�UumN^[���r�+S$֗��5Ht�&�t�g/Jt����� �ko��t�m�    -�SH�$�`[R6�Z���鶹Rl � �=�2YbZF�  ��ݛk3[V�$8	 �:�m]6f�iv´�֠����mN�6�I�\�8[V��6ۃm& -� Zp��l3�gd�]6��V�w��	���2P+da�l 	  M��-p�����@^�u���L���  � m��\+\��e@��S\�E�ZUV0�UJ�k���	��Z�Ԁ:I6��lm�sK��I	ء�Z�ne-���A�P,�U���V�]�l\�k���]�]��� �i��ꪣ�DF���&����5��-�-LYzl�E��k������j�%�$�� ֳm�lh5�m|�֯f��:I@��y�i6d涠@���p��  _�:������"Ҷ�n����ֲD�]�vm��t�'k]M��̭�<����җ[e�R,�;j�A�� 8@լ�3����e~��]Z�[]�:�j�(U�.��GPN�V�5T�.��e��ۃ���u�+a��8tņY�@�M��T�,�P� Am��R��N��畨��ڪT}�U��i�Wq�g�vjWd�9%k�yj�U]�v�T�	 $[�p7*|�ܭn�P�X6W�����86U�
���4�U�J��U[@���m*�W*ʵԻ�ٺ�X}=���*�#��U�l	 ��H 6�����m�� RYu�m����$ H��%� ��jܲp6�M�e6�dM��6�M�8� ���V�#_k�8����W5���m�mn$���`	y�m��h�!/-E��5���kn�Cd-��֖	V�̳�wgL
�Up \�5*�掳&���5�2tm�qخ�g�( �;a9�YV��[9��4:CIŗe�z��"f������ַ�N ��j�	V 
�*y	�4$gI��m���0  [@-� -��rz[
4��-�z�cgh
��2mU*бvM���[E��YG��n��>�UUPH_G^�ۅ�L�#e�bۭh76� F� 	 	 �I�W\9�������S��Ā�H�mgi-��!  � �  8   � 6� ��i�;ѵ����jL  ��(6�3��%  ml� (l  -�-�m��>p ���@�*���m# m���Z@H�6�[@ h�` 	���i�� U9D&�-W:["�"�< 8�d��)��9�J@�{ 7�\nr �T�Q�wkk�����	L����!���mڏ*ęj�)�kh-7H���_��  ��a$[m��/[vn����+��I�UJK[.�L�v��l��7]fZ�UJ�H*oX���j��u!p ��+�Fv�i�Vi�P��f��`@ڶ�U�Ö� z��Z�R]n���X6�f���1�R�Y(�3��ݘ �n�U�@kX(l�"�V����b�S�q��D�`ݶv��I����K8����;!�br7��S&Q��Bn��U�(
ۦܬ�c�7��.H��p
�t�#�l�T��P
�9�̀]&ɒ]9�Nu���ot��Y�`[VXI�l8	:�\��G&�dՖ�U{n������Ȓ6�a��[� 9,x���I,�����ZRL�6��6st*�UU\�e�v���a�����a��quT�P���?.�ˌ(UUT �km��^���l�H%���^Ҷv�an� � �MbI*���
�uv쫵UB���8m �  uO-�٨nX:��hj�d���#q���ѵ �'�,;HtpA�yJ�����-[:���WvU���[dU�K�\n��P7H�L�7���U:�1�t�җ�Uk)fϲq�(䨜ַ��:��v��$� �'�|�_����
]�檁6+R��Yn5�0m�     q�@ @ � �  �p�l     ���m�  GP�`�[p�Kk�K/���.��N�Wo�]�]!r��T�@��� ��@    �-��h ,0  -2�m�m��Y�k��q�k<T5!5�d-�k�����Ӷ��^r崳�^�m�$ �	�K(:�l4P[@��   j� �`m&��ݶ^�K�m��R��5� 8!�k;P�� A�$ڑ�í����m�u�i����%��@V�����ڪ�U�!m^�m����l(86���H��@�MzZ�m�     -�m*���feـU���M\u#Yr ����! �  m���Il��P��2 ��t����.��ų�)����w�4��V�m[W���8�lV6�Rf"���w9���n�U��7m�6��1��r���!5UTUUU�Wc�]r���\�rF�սi67m� �6�U�j0K!�����6�*ܫ˳q�8Z��[4���d��5����H��rCU�n�K)���J�Z��Ujx&�]۶���U�[s[]oV��ln�^�&Y�t%���'E*�2�c&9�m�Z�HUU])�$�l�Y�WvX�Yy@mc�v�U��[l�P �Ŗh�K���fKh]K]Ė����m��`��L�T��n�(�`���H   ����)�B� �W*�U?ʶ]�,�)mWUUQ���4#_�U�G	]���'  6�ջZ��B�3˰j�jV^M�h��B��*���`1Ʉ�V���V�U�8m���Fq �m�7Z�m�� -X[�m���6cm�@��m��W*ڪ�4�UAā��UBj��T ke�ڥ���� ծ���}3��H��m�V`���q��(��S�e�NL�5J��/,�ô�n:���#ko`-����Z��-�uG=��-�gFn�&�	Zk�z�
�k  u�ʉ����N  �F�P[Rq5�[���p �A�:� f���H*�1��K;�jW�V��S�*�ڒ�J�F�V�Z�i�����h_b�(
�][	��Y[j��<���9���u�f�t�t���t�� �̩wÃ�v�Y�l$���U�X�:��daYUg6�s5�vtdSeeEfBW[�Ͷ�$��Hڵ�F��gC�R�� �@9�մ����5I"�Ϸ��UUUO*���Z�W���m�l  pp$i6�WV �@ m�4�1I[l��8p  H[Cj�� �nEӶUu;Z�����@v��mlm�m��� 8$�$m[{E�d��m[ 6��h  ��mm� nސ�`p�-��e+e��N� H��t ��m���N4� ��W@*�]P���UJ�M������ �6F0i4���M�!�X�5n�[m��V��v�ih�6����֗E��6�K�� 4Ye�6Z��YL���F�蚁c/V�	jع��nSv�`hm�i6l�   ��`6�`p6� Zl�&��ԁ���ZĲ��[UU^˭�u`��8S���j���r�!8��`,���$��'If�ը�kEs�]�윗q���^V�� sJۍ6�=z�@9��l-��`"+N�#]� ��(L����ӥ�0p�nd $m	��L��� 
�ݝewK�$�i��K2��9js<nP.������(���H��V�UUBI$һ-�5:�[E��v�u�������O@
IKm.�f�F_Ļ��l;i�2�8,0v*�)T���|��Uc�F/�(���$Ͷ����$7k5Z,�!m �lHH��m���[v�Cm��6�l  �d��z�m��@�8m"C-���A��t�  W[+��K9��%V��݀�x.��v��7nTUV(�5��PR��l;6�mӶ�`� �H  d�  X`-�m�l��M"-��hղ�h$���>-� mU��Y�f��jѥ����jtN6�,UKŬZk���qu��Vƣ"�R�	�"�J���e%���n�)y3UAD�T�^�P4Q���h��� N��6Ӧ  ���i	vf�>�m,�����m�� Hl  	��M�� �m���a�i���%��m���M�h9\�l[@m��$�  6�m�f��ںE����Lp�V�յR�*���UT�UJ�h��A���w[��Fۄ�h6�Nl-�   H �	��;`��:���mUN��̎�"l� ��f*��h8�U��)	�W2L��UUAS1q?���D��E0���i1�A��b�".�
��D�6)�(�z�X�
DM��P�j�F�¨b@^xL�!�"�At�Ҧ���*qE_q�=UO�*p��)���C�)@`it��_7�"�T�ԧ�A�D4�DO\b�"������1_W�a�z	���UpH�������"(�Y���,V!�G^�Q�ht��B�"�گ�+�PУ�Z!P�S���8+衰@邨�Q�I�ŀ! AC�
W�����V � ��Md�`�8�!���A�D�@t������	㇨C*�bA<M�����.� �t�o�JUЦ�	�E��U�� 04�'Z.؈�
�;L
�t ��_�����J�ȈE��=EO C���AXP� $D�,B3�:z%;�)ā$X�H���:������/|P�q}R�#!1�8h�@@E*(x�u�Z#�(z	�x(�;,����AH ���"0H���ب ��_T�Ar�k@*�$�A����yID���"�"��/
�\Ev����1A�1��A ��:�HAP1E� :�D� �"�b.
 P*��!��SHb��u�@O�  x#��#��A�X�u����Z�(�0&(�C�`P!HZ	E<��2�0��Y�f�jtV��U4s��R���6�u��4�$��-��+��N��D����˒�Md8��H9��R�%�k���N;zU��HE'V��\�<B8�|�E��� Fxˮx��e���tf�N�u��ɨ"7	����e��z7TK��)=��ydwZ�`P����nЗ8:����R`�V�P��ݣ���Z�5��z2I�Ū;<��%�UoA�#Z�{�ɐ�;4]�7*��	[=�)���T7mvNq�q�lUuU ��Yɒ�VЭ�V�[]0(%�jU%l��nCv�(强�1ӆ�sJB]�.u� ЦM�7lh�]��N�,y!�蛌�,��gg����̫�۲�	ֵ��gk��V78*�u@�v賥`xHA�:k:��k��*�pb�M�6��u�Br��K���1��U�A����v���Υ��%k�b���n��I&ٱK@U�����e�P)	�̕mt6hs�6;u¯$Ep�5Q���ۗeY�G(6�� BxC��93p�PR�;WN1�;��ƍ��tx�i���QsY�{�����i�Mr�P��C&]͗�2i�����\"�h����5��H�Vz���P���[;H�Z5����Q�����Q`��v�Q�I�mp��nr��{;��1rs�E�祳�(8�^T��h�ͷ�9u��c���]��&N.�x��WKu��½c���� ]�8��vuP�������v	�\��+Dtlb�޼N�����AU'8�T�-r�+b�-��R�0@W!牸��-��Ÿ��[t����৩ܞ�n$;:�����<YvW�Tm��S�����Z/b	n�n�n�۳<�<���z V��\�ۇ[��D��j�:toI��nY�0�,��>-v��#GkHRxz��r\2!��U`�j�	K���{%hkoe	�,<��T����k5�u�B�$�I\���� ����H+����W\�U�OW�@�"����اAN���US��D4#k ����L܅���3X�j��&p6����Yu�����t�Y.��t�.��{/i���k��'V�ZQ�I�]�^7�GF}�Oi5����5�v"�9�r�4��gv]MF��j�y&�,pm���j9��2]IG4�v�Jтyl�Q${C]�kXݥ��N�Y.1�Kl�

�u�<9�v��=]��U����;Za쾱��sY�L��F[�Y���+E؏sy1�ܲ�K���	K�	������v980`v���7=��,b��1�5�>�W{^���� ��ο�g�g��4b���Ǎ'"X&�x�ގ��� �Ɍod�"`uJ+��dDM6'3@9�f����07nD���t���u�������f,Y��od�"`{z:a�_R]۳@?-�i�O����;V��qڰ�:�>�q��Q�M >�/nTK�C9K��Y�ޔ�QP�fx��#� �i|㲜O(<NV��t��m�?:`E�-��� ���[��LjF���v���w���g|����aM!��%��)�<EP��D)I4�"K��K ������튊�ш������=��`y^ק��o�4
�|�Z\j�F�U�W�x���2wڰ�ڰ>�e4b��Ǎ(��<jE�~�n偓�u`}��,�c�R�	-�͓�8�6]+ӵњ*��l�iR����&9.�[1��\��d��ZӺgti�]?[����LoGLwF�'28�R%�@���h��Z��j���:�P�S!��f���UP[.�7$����rNy�vn(��B	ń$�H@��"D�qՁ�|e�,쫉Q�7X��z�v�h�ՠ~�e4{w4��D�SزH�SK�� ����wGL	[������piexu�^��J��瞓�l�[I9�;p���7F�Gnq��n�+W���2	::`wtt���&�\j�F��G������bE�ۚ�}��~�S@�����q�J8��+��31ڰ�jͅ�{��,�<hAҕ�fLQ��s4�������8���#a8J��S�G�]�qM|C�}���s���534j�5���T��0=&A�7�{w4[��6�c�n5 ��A5�@��-�v%萊���[����xÎ�4�B�%WAt����0;�:`M���W�sޞ4;佉xi�Ɩ6�Ry��7��l��{ ���#w�ģSزH�Nf�{n��[���ϒ�l�w�ۚ�VD-����O��b"^n����,�v��v�iq��pYI��e4}��u���7ڰ3�ڰ*"DT(��A`�T{l������[����w���us�*3����ys[s������r�SĐ�9z.����ʲ���nH��:�׃�(n/XtunM�n���l.y�5�Qѵg[���P�N�'������Z�t�v6˞WܤT����M���r�֧�w]�WV����)��;D'q��vM+\��s7��mʬvhwV�홅�h;Qr=J����8��������n�����R���u�Mq�dN�"2_��|�M�u[�u�.)$4�a����o���oGL�0&�A��:\d����ks4����ϳ/��4v�yn��v� �"�B�f*J�::`M��GL	�-X>�'3U3ʩ����+�
w#�0'~��7��Ύ�lJRP�j�Uv�Y����ގ��X��X�!(�{uU5�̩���8�,�����v�.�t���U��vۦř\�1�m��I��v�s@�{w4��5BK��mXܡi$�rEʊ����s��f�<B�*�₟,4�jU%�ap!��z����ϋ�������3^���AdhxI&h�4�s@������Թu)���2�P���	D�{�7ڰ>x�X��X!åfIɊ6�Nf�y۹�{3���x�3�����M��
�b�V+��M�`���i4�	:1�t*�-]r�a�l�3�s�c�TrDA�E��E�9��۹�^w ����7��S�uD��˵t���+�8�؅2<��`n=�`|��hr�p�46A�m`�4�����-u(�P�O
#"ݻ�V�즁�t�xڃlQ����/;w4N��{ ���;�;�Y]�+�`ztt���m�L	�w4b�b��'2bk$��d���0usö�mԜZl�6x{eu���9綴X�]��������&N��ޛ��]]�cQ�G�$��j�:tt���A�ӣ���#Pq�Vf5�maZ�������;{w4�}�@��u�ndQ�8�X���s���1�`}���TBW0�!E�	JC�Ǟ�[ٹ$�O)Ӷ�[�˄�s����aB��n��={j��g)�~�)�s&D|dN&�>�D�"H�-�3��bZ�j/\zm%m�:�'�ݧ\ ��2�*�Պ���0:tt���A�ӣ��mF��6��Q����;{w7�+1�����Kı;��eMı,K�{�ͧ"X�%�､2Yw&�5�fj戛�bX�'<�}�ND�,K��vbn%�bX����m9ı,N���q,K��{ن���4e�ffjm9ı,N�uى��%�bs�wٴ�Kı;�sdMı,K�{�ͧ"X�%�}���[��k5Ip�f�&�X�%��=�fӑ,K���߳�ND�,K�{��ӑ,K���]���bX�'�b�"E(���!C�t�9����kDֵ��F�t��ţu+D�:�t�Z�Wh�&��`�Y�r�'B%�ו�L���ĸf�!z��I�����xQP���N.��9�Bth�7T�������1�#�Wu�4�;d����aV� T��ZI�j�3��`qo;85�n,���K��I1����M&k����'R;
�K�z�۩��B��:I�2�W1���b.ӚA��[s/.SfMe�D�/�$�F�Nn��m-��V�-�f@��K���V6֦��Ԧ�[L���<�bX�'�fț�bX�'<�}�ND�,K��vbn%�bX����m9ı,Og����"�A�R,I�>�>�}���~�v�ND�,K��vbn%�bX����m9ı,N��D�Kı/g�Ν�Yn�.a&kSiȖ%�bv{��Mı,K�{�ͧ"X�%����ț�bX�'<�}�ND�,K�vޓYr噫�̤����Kı9���r%�bX��{����%�bs�wٴ�K��Ȗ{��Mı,K���sW0�u-ˬ%˭M�"X�%����ț�bX������M��,K��믥Mı,K�k�ݧ"X�{��?��!����f��5��/(�I�u�'�tT��k��ٽ+������`�s35�ț�bX�'<�}�ND�,K��vT�Kı9���|"O"dK��w�dMı,K����CWR�2�3356��bX�'��쩸z���8�W�J8A�*AD�C*�l@�x	Q,O{�}�ND�,K��u�7ı,Ny��6��bX���gun�٬�Թ�5��7ı,Ny�{v��bX�'��u�7ı,Ny��6��bX�'��쩸�%�bs$�vu�k5)�V�5��ND�,K���ț�bX�'<�}�ND�,K��vT�Kı9���r%�bX���ަ�F��Z�j�T�f�&�X�%��=�fӑ,K��]�7ı,O|�}�ND�,K���ț�bX�'�	��yI���ѹ&ʄ�"�V��mlgC�Z ��k�-N���Od���g=���<[��Ȗ%�b{��Ҧ�X�%���iȖ%�b{��Yq,K��}�f��oq����w��~:^D�'(b���bX�'�{�ͧ!�1ș��w�dMı,Kϻ��ӑ,K�I�=���Sq8�eL�by߾����˩n]a.kZ�ND�,K�ߵ�7ı,O<�}�ND��hjb@מ�H;a���B�CP'RT�D�E%%4��H�I�/<�<$�Sd��8�!)U���k$�%�&�d�`)�4 Z��~����C�H�8���Ƥ
w�4{m�&�����N	㉡�R�dD�6�^D�I#�2������)P(�8D�!�oR����[h�U}��HF$��;d���F�Sm
�C�d8����#���YXYr�03!\#X�Y ���4xX�$X�d%%���Z�R�2I�0d����P����Y�&Đ��!7p |���z�z���z��!�E|F ������
H��@� u�U�<� �=� 
UU�&&�}˯�Mı,K���]�"X�%��{L��o5m5�ff�Yq,K>@��=���m9ı,O~��T�Kı9�۴�K��?����������%�bw�߮r��іa�����Kı<��eMı,K������<�bX�'s�k"n%�bX�y��6��bX�'�;�>�sY���$�nh�3W]F��ݞ�۲g]�<�-��ܡ���n��J��؈�j�L�Z�.�f�R��,K������9ı,Os��"n%�bX�y��6���&�X�']~�7ı,OrO����k5)�VY�֮ӑ,K��=�&�X�%���iȖ%�byۮʛ�bX�'<�{v���:��K����}i�&�ڧ����{��7��;߷�m9ı,O;u�Sq,~!�2'��~ͧ"X�%����ț�bX�%=�Ν�Yn�.am�jm9ĳ�  dO~��T�Kı=ϻ�m9ı,Os��"n%�`T<�%V�~",b��Q\�	����m��߻��r%�bX����5�fd���f[.j��X�%��w��ӑ,K¡�C�&?}��$�k�<Z�
B�'\ P���g<9{`zc�i��t\v��ٳ��
"��Q��@�W��_�������B�������,K��w�dMı,K�;�ͧ"X�%��owC�Ișı=ϻ�m9ı,N��2�Y�մ�9���dMı,K�;�ͧ!�G"dK߯۩��%�b{�w��r%�bX���D�O��5���'߿~�a�j�SFY�ff�ӑ,K��w��ʜ�bX�'���fӑ,ș�ߵ�7ı,N���6��bX�%��gun�[�L��Vf�Sq,K>�}�ٴ�Kı;��Yq,K����iȖ%��L����T�Kı<�;>�9�f�4j˚�k6��bX�'��u�7ı,?~+�߼�6�ı,K�����Kı<�����KİOw~h����&V��WgmGn!ه8�$)��)%��>�Z�T�6��85�F�f��G���v^���bC�!����۞��g0+�FR�uz��h�c��'cHT8�G�Ӻ�l�1��4s���V�8:ױˬ�E`�ث\&�{X�m[�{�XH���7&m],$ts��)a�B�N�J�h�[Dr��6���̓J�'A)�K�L̓2k2�\�Bf �7{�Ͼ��1�v��S�U���ظ=ZK��l˹�Vc�ٴv�������g+Z���D�Kı?{��M�"X�%��n�*n%�bX�g{��|�șı;��Yq,Kħg���u��2�&�֦ӑ,K��]�7��DȖ'���fӑ,K��w�dMı,K�{�ͧ"|�TȖ%=���/+�S�1X�}����ow����6��bX�'��u�7���)����߷�m9ı,N���*n%�bX���������n]a3Y�ͧ"X�| �2'uߵ�7ı,N���6��bX�'��쩸�%��"{���6��bX�'~��I,�Դ�9���dMı,K�{�ͧ"X�%���^���*yı,N��߳iȖ%�b{��Yq,K���G�	*�s�� ��؍*��=�<m��Z�]Od�(��-�	ۣ7�w��~~{��c�L򭸞D�,K߮��7ı,O3��m9ı,Os�� ~�"_"j%�b}����ND�,K�~�����u��]j��J��bX�'���6��x�����J��P�DȖ'sk"n%�bX����m9ı,O;u�Sq?"�SX��b{��~��]Jh՗5��m9ı,O���ț�bX�'��}�ND��	�MD�~��I��%�by�}�m9ı,N��Zn�����g{���{����{q�;߹��r%�bX>����q,K��;��ӑ,K����ț�bX�%;�>>�Yn�.am�jm9ı,;��&�X�%��w�ͧ"X�%��{�dMı,K�{�ͧ"X�%��;~���jf�˗D�j�r�a�o\@uK#�E)��[� ����v�Qt�fK�̦e�Y���Kı=Ͼ�6��bX�'s��"n%�bX����l?	<��,K���I��%�b~G߿~��\��շ.����gȖ%�b}��Yp��G"dK��M�"X�%��w��Kı<�����O�L��,O���Ymޥ�����k"n%�bX����m9ı,罺Mı���
1#@"�@�"1� � �H>����<2&D���۴�Kı>Ͼ�D�Kı<���a�j�SFY�ff�ӑ,K>T��~�~�Mı,K�u��iȖ%�bw=�&�X��"{�������b>�}���A% �H˚�Mı,K���ͧ"X�%���o��ȞD�,K߾���Kİ{���7ı,O�?t������5VD�35O\&ٻi3A���1�t��[ιuJq�0_٘-Y�ߣ��&4 r�:%�bX����ț�bX�'=�}�ND�,K��n��Ișı<�w������{��7��~��Zn�g�O����bX�'=�}�NC��+���`�Ͽ]&�X�%���o��r%�bX��{����"�eL�bS������u��,�5���Kİ~��t��bX�'=�}�ND��T"}��Yq,K����iȖ%�bS����ɗ�e�e�Y���KϕD���iȖ%�b}��Yq,K���iȖ%���W֐R�b��WH�4��|���]&�X�%��{����,�[r�	fkSiȖ%�bw=�&�X�%������M��,K��;��n%�bX����m9ı,O�/Ś�,�E��E9�ɞ�Wmy5ô#]pݪ�52��v�gsC��\��ܛ��}`������d�,O~��ӑ,K��{ۤ�Kı9���|$�&D�,O��k"n%�bX�{��95.�2�2�jm9ı,�{t����uQ,O{��M�"X�%��?~�D�Kı;���H���K�����n��]k%֮�q,K������Kı;��&�X�E�%5Q?w��6��bX�'響\Mı,K��vtɬ�d���ɚ��r%�bX���Yq,K����ӑ,K�����n%�`~?%�O����iȖ%�bv~�sy�ra$F�>�>�}���^v��ND�,K��+�o���Kı?w���ND�,K���"n%�bX�*!�"���,ɚ�33�ˆ](�F��TU�祍¸���-v�&��m`�A���\���"er��v�zs]�nwA�k<ray��J��ek����
,�8��n���FF�w;uUֳ�C\çzÝ�����̕�vn�W����tr�4[ǜ,ֹ��7>�������c)�tu�M��ﾎ��غE��<���v��a�Wt8W`��qVl�@F������ߝ������Br�Yz�������M*]v��B*�.B�n4ֈ|/=vi�{�5��Bs&Y.f�Ȗ%�b}3��q,K���iȖ%�bw;�d�'"dK�����iȖ%�bS߯�5rfd���fRkZ���bX�'|�}�NC�X�L�b}�}����%�b}�~��Kı;3�����eL�b}��Y�\��շ.��f�6��bX�'���ț�bX�'|��6��c��C"dO�w뉸�%�b}�w��r%�bX�����w�V�33Y����%����D�߿zm9ı,N���*n%�bX����m9İ>P����ț�bX�'������-�kY�ND�,K��vT�Kİ�X�����%�bX�������%�bw���ӑ,K���d:';�s�	T�]ٻVW������=Oa+�6|ձ퐞?}��{������`�ԩȖ%�b}����Kı=�{����%�bw����� �DȖ%���_J��bX�%��}>sY�d����u���Kı=�{���x��c�����hM!����J�4���h� � NQH�>����'9��6��bX�'�;���Kı;���r'����;�ow�~��Z�J�j�K;��Kı>��p�r%�bX����Mı�~�������M�"X�%��?~�D�Kı+�/��f[��0�S34m9ĳ� dO����n%�bX�{���ND�,K���"n%�`|�L��{��ӑ,Kħ�[�̸fk-�2�Z���Kı;�wٴ�Kİ������ȞD�,K��~��Kı;3����bX�'=��G��-؝̀���cVf�������mӠ�#����_��/�I�f��<�bX��I�_�k"r%�bX��߸m9ı,N��n�g"dK��߷��r%�bX�v}2���Ն����k"n%�bX�y�xm9��+���b~�����Kı=����ND�,K���"n'�TȖ'��}pÓR�a��	��ND�,K���n%�bX����r%���@P��� �EXȔA&Ǜ?����O���ț�bX�'��}�iȖ!���\x���Rb�}�oq���BD�߹��r%�bX�g~�D�Kı<����r%�`|!2'�]��n%�bX��i��Y��Mm&kSiȖ%�bw=�&�X�%�ʱ�����%�bX�L��q,K���fӑ,KĽ��u���d��)��08ی�;�m>u�mҩ8�k��.{gi���`3�~�ww��}~�Clt͚{��g�ı=��p�r%�bX���n&�X�%��;�͇¨�"dK��;��&�X�%�_���Y�n�0�e��4m9ı,N���p���P�&�X����M�"X�%��>�����%�by���O�Pʙħ�[�̸fk-�2�Y����%�by���m9ı,N��D�K�'���j'{��ND�,K�Ͽ\Mı,K�'�����˫ng�z2�z�O"X�~RD���k"n%�bX��߸m9ı,N���q,K���� b��@�t��lWI �.ݝ���9�s��r%�bX��O�+-�MXk��f�&�X�%����ӑ,K��~
������%�bX����M�"X�%����ț�bX�{�����?���E�[R�\�.��m�vꄤK8שrX�ݱ��+���~�{���<��Űіa35���Kı>�߮&�X�%��;�ͧ"X�%����� ��2%�b{�~��Kı;���k.�[�e�Z2�&�X�%��;�ͧ!�(G"dK���ț�bX�'���ND�,K�=���O�C*dK��;>2k5�)�-��jm9ı,O��k"n%�bX�y�xm9��U�DȟL�뉸�%�by���m97���{�7����h�{T�Y�﷋���AZ�����iȖ%�b~�����Kı9�wٴ�K������'�������%�bW�o��s-�fL�2捧"X�%�ٝ���Kİ��
���~�ObX�%��?~�D�Kı<����r%�bX��S��"v�f��nĤi2jK����A�	��
q<�J�)�z��8�@<	P�:&�ұ�n�m�G�x>	�����Ry�.�Y�tN	�����0ָ!�l�C�b���/��D�@6)�����M���s� F��;͡���ٷ�@����������p�E]Tmm\�{mbȹ�W��T�N����,���&���KYkn�\�P�R�t��e�tJqF\�@[t�0s�<��.�l��:sN��Y��<�X1kA��iZ��KPzyv�X�� �s�yI;Yu��j/���ں;=Am��,��ugc��Z��k�փ��g/b��&��uefx��d�0��wW*��jz���u'1F��mNx^�'{�۰������⃎&����9�E8*�#Ɉ��t��/�|o���s7g��j���L�3�6�J�ґ#l���(R�*�<M9ū�z�w1�>b��X���ñk� �F���c<��a�0�s�����b;\�\��2�lht�x�k�7���p���-�kshw�mժ��Q���d,�77/=�� ��]��� �u.��K�v�C�/5��3�5��ܵtv����`%�������J����V�b��c�-9a(ڕT
%*55�;m��Ep3������?}WKQ;rE�)�AW�-m�Ņr<��Ŭ[7e�h�]u+�9�u<c�-r�`:�%n�%��%K��TM�-&�I��\Wa�l`��
z����ΧR�^	��N�6m�H��e���lig:i�M��2�6�[��{]�\��)#�u?KC�d�s5�[�0s��򝤴vW�7�X{!K�:.h2t�
ics���N&�bDM!�\�Nu�-D��Z����W�K�`X�c=q�Vr�9�#�NӒۋmU�.^#���Э��1��9��'&�0�*�Ar��.��V���/TY��C����yZ��FY�ݛ�����n^�*j���جm1tf6�-���L�!��қ�͛t��ޏZ�8���,D�/vt��I(�3�]a5؝7.AȹU�Hs��{J��1b#D��	�������ۍY�1� ���ӍpC����;T�[erMq�]��'&&;m��U��"�^p�7�܁�����#����`���`*��S��C��C��*s��}� =TA�补LU\�5!u;��Zզ��I�Wlg�(ĥ<���n��T�O���Iv�N�&�y��*�f�Z�{3�wk�v1v�׎�R�j�և�����%��6
 -烂�a��j[���[:+���l;r;˹�W"vd�^ׇt�$��:��0G���3�5���N獞9�p��<��nt�t�.��gP�<P���v�JF"=.�]HX�:��cVy������)�~P���p3&��I��Mf��X����j����5�h3]��u����xM�w��{�`��n�n��MkW�,K�����6��bX�'s��D�Kı<����|�<��,K�}q7ı,O}���j��S.][���r%�bX=���7���Z�&�X��߸m9ı,O�?~���bX�'<��6���S"X�v}2���Ն�̙���n%�bX��߸m9ı,N��n&�X���MD����m9ı,����n%�bX��aɩu0іa35�iȖ%�!"}5��q,K��߷��r%�bX=���7İ>&G;ݾ[�~>�}���VV/F�H�F'�.�q7ı,Ny��m9ı,�{t��bX�'�k�ݧ"X�%�ٞ��n%�bX��Yۙ��L$����n�Cd��[n���vױ���Ŏ���i.K�s�_�kt͹�kY.���5���%�bX?g~�Mı,K�5�nӑ,K���{p?+9"X�'����ӑ,Kǿw����z(�T^ﷸ��{��y�{v���qT4 DiP��Hb��\@��x&�B <dK����q7ı,O|��6��bX�s��&�X�%�^�};s2]e3�fk5v��bX�'f{ۉ��%�bs��iȖ%�`�=��n%�bX�y�{v��bX�%<�5s-�5mԙI����K��"y���m9ı,��]&�X�%����iȖ%��W�u��߮&�X�%���~�9��2�L�E%�֦ӑ,K��{ۤ�Kİ�#���i�Kı>�߮&�X�%��;�ͧ"X�%�n���~~=a�sF+��]=�#r��a�uP�j��Ճ+��y�1��;���:7O�&f�t��bX�'��]�"X�%�ٝ���Kı9�wٰ���/�5İg��I��%�b{�߮r�%�	�5v��bX�'fw�p�c�2%��o��Kİ~Ͼ�Mı,K�5�nӑ>Eʙ��N侍F��NcR'�i�#�G؏������Kİ{���n%�C�OӦ.�~U��ȝ޹��r%�bX�L�뉸�%�bs�Y�Κֵ�K��e���r%�g��������7ı,N�_~�ND�,K�;ۉ��%��Q�O=��&�)���'M�,�QΨ�ݷ{��?����n	"�E=���O�X�%��}ͧ"X�%���n�q,K���R���~tnc�&��k,ݎ:� r��u�K �s�U"��h��d{����]�$��&f�W��Kı>���q,K���6��bX�s���	șı=�]��9ı,J{����ᚶ�L��j�n%�bX���Ӑ�B9"X?g~�Mı,K�u߮ӑ,K���{q7�r�D�=��쳚�ɗR٢��5��Kİ~��t��bX�'�k�ݧ"X�$2&D�g~���bX�'���6��bX�'{;2���Ն�̙���n%�g��%D�y���Kı?L����Kı9�{ͧ"X���E��Ap Q"aF�@�Aj�ЊPp+Wi�HLP?X?��]&�X�%��ﾸa�L�4L���fӑ,K���{q7ı,?/���~�ObX�%��>�t��bX�'3��6��bX�'���%���3.7k�^�j�8+����cK���%�0vR���i������Hi�����oq��K��]�"X�%����ț�bX�'3��6��bX�'fw�q,K�󺳳:f���f��f����Kı;��&����MD�=Ͽ~ͧ"X�%��g��q,K���{۴�O�=�����~�WL��G����x�,K���fӑ,K�����n%�bX�{��6��bX�'s��D�Kı+�/�e�ˬ�ar˫�ͧ"X�|2'�_}q7ı,O{��6��bX�'s��D�K��&D�]���r%�bX���~5s-�5mԙI�j�n%�bX�{��6��bX������D�Kı<���m9ı,N��n&�X�%�bE)A���%H <��̗2�d��n:ӛg\�;=ph{V�f�qs@q�0�8Dy]sA�f�����m�X5xnLk��C��#"V�ʫ�����م�m��V�Ɯ#t����h��jU�*tvwhL[8톶���0���$h�Mŷ5�Y�닮mY�̇�q�S�ˮr�7F����d��=Y�6��������~۝,�L@t[f�ՓS�.��n�K�p��eԙ3W��P��o,9.��乕��$�^I�s�7vL�Z���S<��*�öw5�u�|��^�`�o����{��'���Yq,K��{��ӑ,K�����1_�yq,K�}��iȖ%�b~��ee��[Mc����D�Kı9�����?�"dK�}q7ı,O{��6��bX�'s��D�O��2%��{�\0�&Mh�&3Zͧ"X�%��Ͼ���bX�'���ͧ"X�0ș���dMı,K���~��؏�b>γ�V5Dr18e֮&�X�|�2'��>�ND�,K����Mı,K��{�ND�,�dO����n%�bX�gg�>ɭ]e�Fe��jm9ı,K��Z���%�a�E�_w��ٴ�%�bX��~�q7ı,O=�}�ND�,K���s�s����۳8LK/i+�
�'�3���׫2UǕ�OIgc����_}�q]2�E�5�9ı,O3�}�ND�,K�;ۉ��%�by���|�3șı>Ͼ�D�Kı/a�~ɩr�զar�fk6��bX�'��쩸hq�R݈(���Ȗ'y��6��bX�%��kQ7ı,Ng��m9�/�P�&�X��߻�
.`-�����7���x��o��r%�bX���D�K�R"y����r%�bX������Kı=��ܳ���Lնh��֦ӑ,K>���ț�bX�'�߾ͧ"X�%�ܽ�bn%�`|�̉�{Ϧӑ,K���S+-�Դ�9���dMı,K��{�ND�,K�{���Kı<���m9ı,N�{����%�bq�]�K.gr0��Y�lL�����A��ݫX˙������K��%��foyp�p�5�d�f]j�<�bX�'�~�17ı,O=�}�ND�,K��� |�NDȖ%��u��i���������@i��K��x�,K�u�nӐ��U+���b~�ߵ�7ı,O~���iȖ%�bw�gmM����,O���d֮�٣2�kZ�ND�,K���ț�bX�'=�{v��c�#�B�P�KE0���"#�X���>�7ı,N���v��bX�'}���F�Y��WZ��5�7ĳ�H���ӑ,K���ϭMı,K�u�nӑ,K�n�~�ߵ�7ı,x�ߛ��MbRN^&>�7���{���Y�Sq,K��>�}��<�bX�'�ߵ�7ı,N{���9Ǎ�7���w{���7��m=��]��w-�Sh���K�r4	W<�k�n3�67=<�t)�5�mԙK�թȖ%�b{�w��Kı;��Yq,K���n���"dK���_J��bX�'}����]��K�
�����7���{�{���|�"dK���ӑ,K���_J��bX�'���ݧ"~Q���K�����nl��9���dMı,Kߵ���r%�bX��벦�X�C"dO{��v��bX�'�ߵ�7ı,O|��pÐ�5�d�d�k6��bY����n��7ı,O{��v��bX�'s��"n%�`UC�	�T�. GH��j'w�����}���#쬬^QD��RK��Sq,K���{۴�Kı;��Yq,K��{��ӑ,K��]�7ı,Oʇޛ��2�k��l�mv`��:I��Ŵ��	���X��#'Y����u;���Hk�;T����,K�}�Yq,K��{��ӑ,K��]�>Vr&D�,O{��v���7���{����z(���ۉbX�'3��6���$r&D�>��Ҧ�X�%��u߮ӑ,K��{�dM��(��Mbj%�~���Y�u�u��.[��fӑ,K�����Sq,K���{۴�K�XdL��w�dMı,K���fӑ,Kħ�ze��kSZ��L��ԩ��%�
�!c��p�!I
H���VӍՀ�8���lM�8�jcĤ�@���b"!v��|��,�c��D.Wz�~m�y)z�'t��F�W[m��3����8�V�mb�÷n8�X�aŗ�OV��i1�mn�E�ӱ�U�-�A�Ol��ZJL��}��3��g�n͡��˩mm/Gv�NUz�۳4Ϲ�ҫdlr�N�bQ�^w\R�$nѵ�kX��qk�VK�)q�]=������:o�:�,/GE�6M���֘v�� �`�\��ɚ���V��^>��Nn,��m-���˳l��sͻ7E=���#V;p�������+�t�e�6Zk˚�k�O��ߦ�y�e�ܬs�	B�@�����M'�`�0`�G�^�S}������∄������{�{ �'g�ə8�b�'$4�|��٧���|�����g����#���o����;���;/v���Xz$��=�����Ƣ9��G�H�ɠ~]����ޟ��̀���Т3Vœ��Jp��]MG8�;3����v��B*�pv�i�}���1;	mbRN^2C?ͷ���r�̀���DG���V �+kÒD�5�Hh��[~���3a#0��HI��$<S¸�@#>2Ghn`:`1�!�iRY
*`FF0���SDA��8'�%���7$����^�S}��m^Kbl1Đ�<jNM������q��З��U��x���0$�Q|$��X_֯`���-�;8� �c冨P�soK�ښT�E�()Q\�X3��5(��oy���4˶��ÿ,K�<����%Cr�b��]���ݷN������S<e����{��r}���#��H�������ye4���P�]���<X����s�Dԍ�#�ɠ^YM�����h��3?���;����E�"�|�����z���YJ�q(�R��)FP���UaHQ �b�1X� e%Y|�V%6/&�'����i����4�%����kG����6
mO8QCM��D��R@�0@�@��!���T����y�D_ ��iEzJ��.�z��9�^����Q�"(`�*,5H�� H� �B����Ň8xD�x{6���g��B$L"��x3A�������#&D�Xz!��C����<؏Qq���hH�M��|U�����$�pp҇��D���|W�( �p*	������*P�b!)�����K �ctpM���D���gً�� ���^YM�k��w�[��b\�`��T(����6wv��Jg]�4ږF�~i,Ln`)���9��N�Y9��O^Gi�Mŵ��:2;u�;��w�}�q$'2c��留�k�/{)��������^�L�Z��O8)�MC@�����h����o�/��R�b(�AJ��*��$P�kw��<��������A��0P� �w��M�<���������A�lllo}�~�]e�Y�d�Z���؃� � �7���؃� � � � �����A�A�A�A��}�؃� � �(PB�"�"$Ta��`�A�A�����A�A�A�A�;��}�k2\�3Zֲ�ֶ �666=���lA�lllQO>��]�<�����wM�<����{߸lA�lll�t��.����K�h�OWWY�i�n�]�n�Y��.Ջ��;If��l�;��_||�%-x+}�������7xk���A�A�A�A�����A�A�A�A�{�� �`�`�`��{���A�����~uu��̦e�f�Wb �`�`�`�����b �`�`�`����y���6 �666>}���y[{'I���f�YrL,�Z�y��p؃� � � � �����A�P,l|�_}v �666>}��6 �666=�o��,�[e�&�4lA�ll_��� �߹�lA�lll}��߮�A���ϻ���A������6 �666=�i�%��%�]j5sSb �`�`�`������A�A�A�C�0@����6 �����<����}���y���.�^߼��	)R�T��� ��@���f�˚��ln����lo��,��M�GO;V��^2tUQ���o,W	p[L���X�^ެ�����V�Sh��!���f�4�Нm<g=
0�����EK�,��+��!����U5��s�TV^N��I�;u�ӵ:&zl�\���&��e�t�&�H��%��]��As�K�;s�ն߽��ww���vUM󅮦<�\���3WSZ̙��5�1���1%ֱ�KcX��]�un1�-��2<��ɭ$�2�Wb �`�`�`�����lA�lll{���b �`�`�`��{���A���ϵ��b �`�`�`��'�/�˩&��3Z��M�<����{߸lA�Dlll{�w�؃� � � � �����A�lll|���lA�Tlllo��C�˩r噭k5ff��<����}���y>��]�<��?�Tb!�A� �����y����<��������L֦��Z�5u�[�M�<�����k��A���ϻ���A������6 �66
�=���lA�lll~��ߝ]k5s.��f��j�A�lll|���lA�lllN��p؃� � � � �����A�A�A�A��}�����=|f����|�E�9��'kW�ɫH8z��f��������v��(LIAJBy��m�;�e���a(��9�<h��[�q$'2a��w��t�|���D�4��>�� ����Xo�X��X�(Nf���R�N��נ~���ٟg٘�-��{g���<y��2W*�尒�J�ޜ��;�\
�b����\^�@$�qD�^�遻2	�"`ñ��g��v��lZ�r�5�.���ܽ�c&���ȐC��\���ݛ�3�_�����۾R�&jc/�����}����_�!%􆷶���ndQ�<X���x�Z9e4�������31#�=W��G�rQ�<�M�����y�՜P�A���D
���e1��G�c�E>U.}�5ɹ'���w$��q�ڮ(��R�n��YK��ua�
'3oK����ͩ+�2'2a��s�S@���q�����Ɓ�c�`Z�Q�(B����JͲ�l�-%�#r1i�=�U�M�F��+�����y;t1[�6��۫�|e��c���y.�7�x���Ǐ4��O$z9e7�$r�nh紐����8���*÷�P"�dR$�Z���h�����@��T�ڂi��Cs4=��o�r�f����>B��!".7Z�>�j�'28�y���/�@���Oy~��s@�l��s�,_u	�$�%:�,���.^�!idQ�zY��s�@o�}��ߵH�N,'�8��?yh1ڰ3䒏�;-�X���U[U\�*h*d�96َ��$�F������Xt�ߗ��7w�53jjxL�\\B�W���x�>��V]76َ��=��)-ަ�j�P������*~T����~�zl��B^�[��ŀ�����2d�2H�Wj�?�Ͼ��{����XNc�8�/�B�BxH�E$C`P(���c�Ϳ���mM�]h���@bˡe����i͖f�����uۅ�v�ѧ�ĉ?}>�>�4�bʛ�"/l����ݝ��W/&e0/N����������#C�Í�2.nն�^;vx�8-v�d�U/>
�m7j�`cq6����c���Ft.�v����i3M��,�Վ�6�tD6�u3�g�s": `,�ê�u�����{������n�.�ű�5��u�D�F�E�6�K�tF��1qImt=c�m�����L�`ywK`l� �P�,�[i9#�nf���M��1#��=�~��?w�sϒ=��Ndq��I%!�j���6\������2�W}�4�"�b�G����=�r�nha�#Тg7}VJf�UW����V�fb`{�:`N��t��j�ּFU�j0mH��"dwV�>n
�M�k4��:��d��3��{��~��C�MAbNc73���4˽�@�vϢ�B]���Z�<��U(�������M�9}�������	�q,�c��;��X���J"d��*V"�.M*9�U��[�`}��Y�%2��M��=��QH�q�l�N-숉�{��i`}9��=������<���_̂m�䌍��;�)�fGi���ٰͭ>�v�DD(x��ep��B�ihn��b�e�n8�JڽY��i���8�wz����e⧂��R~�ˑ0=�0;�A�Wj晴Ɯ$XLQ��Wj�g�|��}��[��@�����g�YҠm�7#i�L��&��{j��|e����""b P���vVM߾�nI�s�Z{ړKD��9���}����BU��X;�����O[ߕ��v���D���p�?.���>�識�����d�\��
�J������:To\�z�B����34���nD��v���3$�Zx�L2x%"�|��~廚{e?� ��@-�z%��aTrI�M��>2�B^J*��zՀ�wՠr�V�}�$Tue��I���������K�!U?W�6o�����Oq9�G��X������]�zI����rN{�vnH8�6��XT �VU����L��� �fs3����M �W~�Gp�a1�9V]76�DyDFo���7}�g2���f�ppk��8܃x��4�d�۫����h"�eq�n�4C�y�ɑbi�aib̶�d� ���/�}��A��y���4�I�X����C@�_z�(�2[ڰ2wv����B�/}�`��'�'���o���k�=	B���i`7�����u4�X�8����*��B���ڰ:��X�������]v���/D��L"I���L��d���5I-��-$�4�^�&�� ,X� F""�&�Z�\GL�8@�=*ȏ���CH�~t#	��JH���FE�!�v�bsŉ�s��@�0��jd"#��&_4�kDT�1#4>���"J��N����↗ł�Y`Ec�ȸ������j�I$�Z
�(X�Â&�mڣW���iHZ@�B�[-�Y#HD�8��!�r�����Z֮��ejU����R[�5pf������7�6�qܫ�v{+�4[v"�-�k$�i �a��/F��U1n���b3��P,��9�9v�%�ڮK��M�q1�
�CL[atka���Rk�.%�=��j�R�d�,*7e�E��ݢ�sך ๮U�
M����*y\�i�C\m9t��r�ѕqq��Y3ŀ{t�����x���[j�d:��*�Ύ6y�i�8Na�;7�j�&YӚ��T ƚ�a09��7-�0 F�LfZ�[Cm���]V�ᝤ�W�
%�ȦUY�Mlj�����M�Y�g�{�]6��j�lK��*���$�D�W9䝙Y��]�u���*˲-r�՝�����*�ΠX+vrg�t��iS>t�$<�-ո�]U�I�Yc�h��:�{u��U�TV���`9x�na"y7[x4v��]�<�u�Y��bb�s������)`�eh��:n͵�DQԫ*�l�m�a��F1�g���VѪ�j���������ڍ�5��#&���ӕ�FK��t�I��6���˭��Wm.v���k!�k����Z�pA�x"�j���kv享\�q]�T�7=�.6ж���X��d����k��te�%vĽT���]�X�R�I\��8���X�Ͷ�o<���mK���u�Ћ�q)­�F��D���"g3q�.�.�a�&]�h�u89K]��"��m�2=qשZ�V�;��; k��\GW-6UH�K �tu���+�	�v�]ofSr��审&�5��r�����%iแ3�9��۫{�&7P��x�dU��.�� ���v�vm��I]�oF�6��2gk��`��S�a9B��a7JN��w6M�kT��o9eYiD��[W���)�uv�ݧA��lUP[Y�"�(e���I�u�*]m����a��*����KT5����I&���Q
�%���S�u�Z�OD�D���OP<@:�H
*q���އ�"�Eا��������!
5�V�����lť�qb��;u�՛�����n�m�{Ocb����K�\��z�@�;]@�6+�8��{0�R�WN�t��͊�g3�R���*�82�\�fv,q�Qu�=�㎷k���]:1��T.���n��9���H�n������/M�J@�����<M�\[.���k���P*hx� 3�;Ad3SV�e�&����螈���P;ￜ�	ٳ�i�\�/F�٬D&�7`�@%s;�1�X�\V1˦ro7~�����>wB�W9�9\�������VO[�DDz33�;���h����'28�qȒ�-������u`}���:�ߡ(��%��z�}��q�	r=��=�L�e�L]�����We��v�4���{3/�Ɓ�;�qw��{�W�y���4�I�X����C@�s`{)���s��`}���3���[/��5�jx3�;<�K�m�h�t�\UX�{r����\���~y8��V��O�d��`d���>��z���ͧ�`w�ɼy�4&�I���^���
�W8����Y��_M�>�>�h]�zmQB$�6D��@�`u�9�R�3��Հ�7j��;9Ҷ�&�NH��4Wڴ.�����}�����=��d�m9�$��@��k�=��_}��_O+�[��?��~w|0���U��ynNB�+���L�U����q��i�<��8G�L���*�s�`d���>��Xu�}	yD.0���z�?�6/�i�Ģ��c�/ДDL���l����c����M-dHI�xG!�r�x�8�����i ���0r������{)�r��IlqHb�p��}�)���-ڰ>t��z"���z�7�4Ƃd��	#�9�ܫ@������/�����@�L��P����n��0%g��v.,b�[���=/���ɧg�4��!��S�B%$�6H�ȿ�yh�e4�j�������:�,��YmfZW���`t�z�	���[�f}�E����72(ۘ�I�h��Vr��f�*���M����`���<�8H��8���ϗl��|��s�]���*1�'�����Z���Џ���'����߽��C��'sA6�x����Z;e4�j�9�ܫ@?^�dm,X��	�Xl�@y����hy��)�e�]\t�,��s��w}1���c�s$�_����v�V�ξ�Zk�h�����qHb�W77���EP��zl�P���W���9}<h�����L�7�$zOSu`}-���"g5�K�{V �ⱨD��Ȓ���.?{�@��`d�:��Q.��V�%3j�rj�Ms�H���7�XQ
2�v��3krO<���I�(��H�H"A}}�댰�:t�S��mF��H���]�Sxq���,;"����r�X�^�d��^�U���Or7�tF��Yvخ�E��ήh!��p\�^�^Wb��m�m�fՔ����k���X�9z���P���ىb�&Hٺ�1n�Gk��cP.ŵ&m]��F�Uٳ��:4\)�!�<���{)e��6�Mϙ8W&��q	 f~ϖf}�O��ƋÇ���N�8�������ٴ��C�z���d�'�)nu�镔��m�~~�X=�Ձ��s䗡v�=�x�����I#N,#�G�us�=�v���g���y(���=TL��T�<J'�-��@岚w3��P��[��0)X��|���/H���߿[K�&��Lo($��2C����נ{��|/�s��Z�S@��>x�h�I�1�� ��ڱ�t�CZƤ5-��on84���m)�[�k�� �r�u����s`c|g��/��@?����5��`�n@��j�E<X Ɓ�Cn�w]�f�_}�@�}�������l�<���k"i��P�@����4.v���*�9�j�9�׬�'28ۍ�܆��f}��.������+�`n܉��2�WT�cNǂq����*�9�j�?[)�qrנ{�����3�f����4�uvv`4'e��v��X�ΎՍj��;\���q���qc�������YM�����k�-�Zb�C���Url�񗰒�Jd��ڰ2qnՁ޻V��H��bI�4�!��@���f�_�7߆��@I�@.�6<s;��˹'<�]��y�Sx�Lh&L��=��k�9�j�9�)��>]}���v�/D�AI&W�j�-��r&��05l��յ+�σ��&�b��Ss�nbG}�l������sk=Z60m-ٹ�9Ս��)ЊNH�����x�8�k�8����v���z̃s"���i�h\�쪪H�Ւ��"`ñ ����7q��n=��k�9�j�9�)�qrנ���������z{Ḿ޾2�������BI �  SK|��nI��w.K����H��@�,����_}�����qڴ#8���2i85'5�B��<\�>a	�G�j���������G���sd�ư�-z2נs�ՠs�S@�7�4Ƃd���5mIlۑ07fA��} �bY ���6�G�~�ՠs�S@�_j�8������V�O�<*�6�����=����XjJ"���Z���Gq�Ӑ�;�ڬ�Su`|鹰;��X��$�P��F* X �D;�9d���c= l��7aaUM�U�y�R��_'H'��s���ru�6�9WV�Qi^�۫\��}0���j��ۗ`Z���%98[��W�N��)��f�h�x���n�8��tD���`�6�d��*/�LZ�ϭ��\ݵ�^91��s[��<���A�'Z4��2�s��nv��N�t;�.�P��M�F��OQ��UD�ޭ+�<&�����̉V;��ۖQKeVL��g��\��69����ƛ�5�'$ZW-z�Ș� �ղ[ ��"+�J�4��qc�@��}�f$w��4���@��Z�nV�����xŠñV�l[R[v�L]�"q�Ik�qrנqs-z8�Z9e4[Sx�Lk	��"`jڒ��"`ñ��&}�{c��+���v��͞�mg%u=�ls�'�*6�/e�[lenn��[Ț��]�e:���r&��0;��`jڒ��YJڂm��S��9�)���Y�db�u���j����7��.�:���@�]�@�-z��s#���i�������Ș� �+�z�i��YrE�qs-z��Z9e4�����*#m��i����X:nl�K3oO�n�́��Z�}�.��yB<�ژ��8&�M#�Brn�9�v���`n�'!x*��u����}���������;�ڴ.e������~��:�<D�L���@̬s~Jd�ŻVv�g�#���|��<�5�ɂm)��̵�����] �	E����*3�c"FD�1�25�Q6�0�:`5p�D�� XL��g�N*	��\�8�'+jB��\ �H:k�ؚi ����-�o�ڑ	������Di����X,M>0<xI"����=��!$�T �<}��m
j)�7�f��M�'� �NJH��2q��V�t�r'=�2�BKI�8�Ͱ�"�K*D�h�F @cm�������T!�h �@�h1��4b_@^	�!���==8*� }P�� )Q`��Jh��h-E�d��L8ܮr�=���ٰ5�i`fV9��7ZŅU��܍�qh���<�C|{?��v��76͜��<�:m�E����v��Zv"Y�kj�E�+���7�孹�t��[�����Su`|�Ԣ>�����tnM�ƛ�5�'$Z\�^���V�{�M�}�}�ؑWJy��r6�i�W������`N���&[R[�ܭ1h!�
E'��>��wƁ��~��v�w��8E")��}�� @�L@		���u�P���Z�zP�'d�Ơ�4���-�-��r&��09u�/.�qƗK�ҭ9��n���u��J{-4�a��nD������w��g��'k�ͷ�����=.D���u�LH��d��L8�����V��H��Ɓk�Z\�^�f}��w�/6���8)"�=l�w��i����s�z<��w9ۨ�)28ۍ�܆�޾ՠ9�X:nl<��^����n��28�q&�$�@���@�]�@��vnI��n�M /���?����Ol�Y]�U��ә��7���ļ��%�lu��sl���F��{J-����V1`���$�2��kg��'ڸ�z�Ilg�u+UA]�p,���{Ec(����Z��9r�t���' �:�]���Jk��7[�9���(���%�v�')�h����m�j�U�V����VL��Z�" ԙ����֤ˣ0_SkG7��5rԇ'-̴��u�\v띹�9��Z�%���]�pڳ�y�����}��Ti^�ç��ٰ�2�̬s�%��i�`[s�1�dhPd�@���{X��s�:�>t�ިIzUF���DN4�!�A8h����*�+�����fb#������,�:��R�yD�yɰԼ�%^���3��M��q�z�V�[QbY ���6��������D%�o�:�o��s�:�>m_�nl�ZZX�z�b���MM��cq���1аɎ]3�==�v�K����M��q�ec��X�����ݝ���F1I�ĜM�h��[�ϲD ��Q9��&T�  ���P��%

>�����{6y�h~�Yc#�7k"NH�
�J��76jP�gu�K�{6 ��:��r6�hq�=�Ͼ\�����Y�@̬sa�I)��6��ښ$���� �Z���?�2�|���z��Z-āM�%��LH69�=7i4u�\Y��y�.7�.ܩq�v�GY8�4��5�w��hr����f}��g���g�Lk�LƔ�@s�:�>t���`fV9���CwR�k$�`�Lp�@矼�{)�P$D!$D@��ec��`��:g*��&ؚ���C�fb����-w�@���@�]�@�s�Q��dQ'�rz�V������矼�{)�s�ܹ��M5��s�&H��9�f�=9�YŪ�v'�l�ѧ�����˨�L0��5�'$_���=�v���h��Z����6�r4�����Λ��&��t�l=c�3�if��Ab� �Z���;�ڴ�%��z<��;҃#RD��PU��̬s`9�X:nl>��I(�~C�Z��S!L����m҇7����w�O��)n���uɰ���.�7g�7_4�3+�����߻�����Cr��"�Y]�v4��&s�n������$&x���!ӱ���8j���+�g�ޛ��,��?�Hl�V�;���lMH�Š[�M�}�`9�X:no��˜�rH*�И	��?-��z�ՠw�Қ��ܱ�Ɯ�k"NH�
�J��ڴ{)��l�Z���<�brEe��ٖ���N�0;��`E���������}���Mf�V��Ax+)�2a9Ҙ��]�]��r�j�@歖�Gql���=M��^aɺ��a�E�9�fչ�z�̶L8��ʽu��/��.�ۚ�!�T� �K�u�l���
}���;5��<�K��]�8��5��l����t�Z��N0�I,\v��h�s'�'WE�y�R]�9�vv���oWOI{6�w^�� k�����w�M��Y�ݸ[��Ybf̆]�r���	�e�����,��Y?~�o �BD������@�_j�*�+�?Wj���F�5$L�5�fV9�����76y�_��C�L���5�O�
cJE�+�=�v�����}�@�{��yM�0r&9XzDB�g�ޛ=�Z�3+�-�z�9UoD��G&Š~��h��l��VΛ��"!f�ZW^uٞ��I����^2�ӛtf�Pti#��^���9���}���t��8[��"�����!-��d��{�e��4�I�#�G�uZW����o��a*DV�S��O=Ͼ��}����qs��^"�M�N8�48���i��:۵g�Jg'Հ�tڰ�i���d(H��Zً���f�Տj��lua�"S�㹰d�+�F�i��h\�z��}������]{�`u�j��c\�"��ʒjy1Ċ�ړ:U��l����U��5d)l��'ո�1�Y>�X��`����x��?qڴ[w4.v���+�dq7$�Ș����տ�${�x�:�|�
�J��ֱAH�!�0n-��h^{�ܢ�U�D��C?5��4Au���C �U#�"��_��~z|���/s�p���N&��BQ9X����j������j�3�Wr��"JLfE#��v���K����=�zՁ��:�3�*��\m�6����r�{j���ו�`{Xk�9���.5�:Μ��F��f�2��m���6mڰ;=�Z�}!��ڰ7^���jKK$HN-�w7���H����<��=��|�S����9�q��+'Հ���(��V������*�:-RY�P�32�t%�=����=�ٹ6 gtbAb[ � �"0]C�'s�s7!��^֠�nI��i�=��@��t�ս-��a-�N�:^]%v�:�5vk�O���<�wn�)C�9-����1�+vnϖe���b���cN!��}}��qs��\�����������s"�>5U\V�%X���i�`}�nl�w7��9U��"JLfE#��=6��M͞J!L�ݵ`d�ڰ���+x��&6G�~�h��h\�z�}����=����,q%ąx�H遫z[.����[�h����*W�6�]�	x�$i�-�����F��$4�b��0��� �xW�:5�a���`$`_S��Ri�}Kd�|4��}(C�
�'`��!��|c��������=����P|3�1	A�Bl�X��O4]�b������@�iCh��
���<"B%x�{��� �y����P�k��C��6�#�yxav���F�����&�Z	]!��0X�`�<'v��������+�u]S(�R�\�ء5^q�5���N�`'6�2֭Ӷ���P�U�u�H[v�:[#s�����c�iM8�Z���ӷH��7h���5`vtO%��[�����R�G����ˠ9��ȏ]���Z.��*�O�4��5�j�2�yul%�f�F5L�ɐ3#�%vl�4,����=���^�DRv��M�'���C�(�	^u;�@��v����n�b�.y��Ʋ�)5��,bь�E�;�y�R�K�����gr��r��U@+hV�h�HBQ�p��*�j�꼤�	ʢ�M���Et�r��f��q��@촷,��ڳ�.���0��R��!\�.;i,�Ż�2���.S���ܜn�ͷ%2�L�-�vR�h9�C���l
�D�tz�"㲄9�Q�881���ʞع��m1�	+�۳��O/6v�Ctܰcc�.�v�
uԋ��6��UU&Ā �2��Rg7:�]2��S˳˰U���7-���G��U�΀�b����T��ٶ�ZX����l鸹�Mtd�:�Z�y��儻)�ek�٣c�
�Ҹp.��б�U+��v����8�2��H��c�tv��Չ�v�b��p�oifEi��>L$㥘ڬulĴ&�q��fDa�f��c�v6Ր���=��n7!�y`^�Ŋ7.B�����]�HP�
ŭȑu�t�Ў�R�3�h��U���,N.�vM��*۠:����B�\c������C*f���Ơ��Q�Z��g+fќ��mL4v��� e(mJ�V�e�"�3b�lI�+�fw��瓳�D���ɌSeic�꫏cb5;�6��܎��B�;�;��<[=��鴼��Y��y��rl=/N��a���m˹�kT��k9��Q�	�\!�l!�[�]\�[�q]�5b���4���`1�vI�-<�GEm�;r�;r9�q2���^4+@Q&v�mlg[v��{����N*`#�x^/}��A�q �Q*$PB�SOP��Aqሏ^��_���v]�9R�XM���<�nmu^	̛v	k��h�\u����Wi�m��]�n��zS�������n�;Zt�4qYmx'ҝ`�w��9w@9���SO�$�g�%��&���]]�e���ECv�kH�-A��c��k���t-a�Ճ&�;ؗd9���f�x�ǋ^��L�g>aefӺ<�ڑ��I<�j�qۛ]����{��o���gk-����o��\Ƶk\�ձqlE�s��KBA#��G�s4�����Ձ�i��Q�]����V�L�+��ϲ��������N��\�{�H���jPq�$�ț���s���������l	���t�����8���@�s@��k�;iw4���Ͼ|��z3�|$��H�PkW���u`z"P�M�|g^Ձ��4gٞ�����'̄��6�p�.��<\v9u�-,�-�g���=$�;��w��>�!"JL�a$��ۚ�{^����B��{V �$�3���W&���%qXK�W�Q)J�-�O;^��K��[��1h�8��q��ɐ`rޖ����:[ �Z dr5�N)���@���<�K`l�tJ�0-RY�P�39V6;V�B��k����Oqց����*�b&��0$d��B<�@��DJ���Ѷ2�7Bm���MA0�]���I��{^��e4�v�}�ߐ_x��S�y�D�d���z�[���-���t��-����	+��-Z��+����:B:g�U�R����!� �`����7$�������9	RH�$�h{�����M�X��V[�,6!N>=� �ؗ�����h�mz-��7��`t�t�դ�T��_Ⱥ�
V)Xn�n�X �FGY�uSO��{p��3�֕m4�$�Ĕ#����9l��ξՠv��h�mz�� dr5�O��r���#�6Ձ�{�`u�1���LT�}�,���#��Il� �޾���ȃX�]�̡ee�����-��d��0���Z��D��7�rI�󷹖j�kX�^^�-��d��0:B:`yvנ~���24�O�<����v�� ���kIqAqmD���hv73�qV�aj��[%�:B:`j�-���h~��(�$II"�H��;s���S&N����O[�؉��R^cNF�45���:�|���i������/��s@�֚Y���J��q����:�k�;s�sC�.�_= ��x@��jƜRW-zmtt��:[�d�U}��S0�f��*m))mbͤ �5���hJ��m;�����pV�l��v6����}�w�i�����;'��s�����8�krz�1����������ڠ��w�on01�p��!�����$�מ�7NY�; ������vPA�n2ÝɫŅg"���DlI��=lKvD�rp�{*���̗���[���md�v	���w{����q�U��,���d�[�sG)�B�$j�-4�sh{r%�	�[(�]n���8����8�k�;{)�urנ~�R)�(��L#�&hW��y�X=n�k��IL�:n����Ǌ8��<h\���۹�q^נw;��w�5�9��l���T�l��`�\�9	RH��8�����8�k�1�`d���5(�OuIei�T�U9�ݞ�ʋ���d�$�-T��ϭ�4C�y��LJ6���������uz�����:�k�}��Y�@���Y���KSY�ˬ�nI�}�f����	�Q��*P��8�L�����;)�q^נmKW#��N)����;w4�ؗW���}g���\�"�(0P#�@����T�l��`r�-���h�,X��fP�*��`j�-�Ӳ[%�:Wn��\�DcĈ࣊9�ɉ���	ٸ���Z�a5��ХXr�L���{�Sl�b_Z�e�:vA���&J���{^���b1	�R4���4��l�����l��`i�B�	RH��H�����:�k���Ͻ��<��R�P�
�� �����4.��@)��*�N6�*�)��t�N�09N���]0/mi���N4�r5zoe4���+��)��jR�`��!Rs]�����ι���\V�Z��n%[m�u�d|z��8��G����4�������t�N�0;�R�X�K>�`,�`t����#�� ���埱#��Z,J8��LK$��u_y�; ��:[�tt���]�.��J+��q�K�V5�Ճ�!��1^��srOO}ԅ��4����^`��}�tt��:[���{�˙���XǎbY$�f��;$����+:z�V��t��ϑ�Tr�TX���Ta���Һ:`r�-�Ӳ�ڴ���$�i���73@�-��2S��6WGL	�Z��Q�Ɣ#����;�)�u^נr�n��{^�e�,k+��pmI�J]kڰ3U=�%�:ݫ2�~�/�>��4��@��ڴ����v�����(���@�!BI7s9�ZyY��na�k�9����<%e��Y�K�@����K��ݑ"�7�m6Ը�"-��7&��>	;k*c�Q{c��x��[��]����	P"s�{mq�8�p��u�ں�=���;M�\I:2�u��f�h�7Zvi}t�C��}�̴ZĐ�..ɘV���n�I0��K��*��@=C͛&z��Ձ���fI�m.���04��8QO{���p�#���-��+0�cKЈ2��̺������t �5�랑MA2�H�L��'�6}��:ݫ%��
>���-ʞ=@6�>j
8���VK�V]���x��$���Pe�E�D�6�hz����z{>ϒ���@���8��YI"�%$�řlu�[��l�09N��)���'O�!#�:�k�=����]g��:��V�,���݀��:�u�G=f�<�yhXklF��n/F7h�<;"2
4�Ȅ8��q�zyn��t��:[��l��U���t�5���Y�rOo}�o=�>��@ "���D>�d���'o�|����������<��0��R=�Y?[��l�09N��=��1(�n90Q$H�=�}���_=����:�k�9Y��ה��X6�>j/-��#�)��,�lS��=�_x3��Ɠx��0$JL����6��wJl�9%s��[���Մ۬�D��7�ng�*���9Y���������8wRE"JI)���נr�-�ӣ�)��4%�J��i�8s�`d�u`c�j�D,_B�Q�`Ec88���	�L�3Đu�:�ڜ)����M�=C�:hB�А�4��`ob�s�2�9�T�H1#}8�Ѣ(vh�p$0�S �Ā�ǡ��<���N��7meee%��HR�҃��MBBt ��%�m�6�2)H�a #F�����T!
RZI[cm�a#HR���B�[F���m����#�HF2YHH0Ȗh�����"@Ѡ6G	�F��B�d�P�IHT���@�$H/�F��"��D:&�=@�T�QT�W�/�������m:%E"
���Q �ER ����99���1��P�M{�4�U�N8���&��/��4����v���� �{[!�8��q��U�V:1Ձ��Ձ��a$�rwys��å��-J����Ӎ��أR=k����7�\N�q������t�O�a�j��x��ǎ��K�:�����J8��Lđ#�:�k�f$__nhz����z��To����e�:tt��:[��-��t��V��rC�3�WY���cs4nN"WZ���=�%�BJ5>��\P�s>��3�߽=��yx�z)�%$�	9V:1Ձ�!:׵�^ڰ2^:�9Ι1�ن8��>�E�I��l�����΁v�m�N��Ƶg���k��ip2�k��3-��t�N���K`t���9mI�Y��q5	MǠv��o�Q�G:����K%�Ԕ%2v���Ӊ8Ӊ��*���;s��{����/��4S;�
bS�#If[�vA��t�N���K`{��u(�n)0S��u^נv��X/X�q�����$uR\ �@���A���,ɫ��32��˴��m؝oƺ��NzӳtWX���94��r�!sG)Rs�;m;�C�3�՜k�������le*���j�:���dn3Co�>���c��Em�[W,��]�ƻ��T���glJA="̱RG`yG��n��x�؃�^��3ʹ\F��GE�gMԴ�#��Zl�a��Yܮ��c���eyL�m�Ƚ;��w��콷}�`�:������>Ϸ&�p�ݦS���nZ/i�cr�f��e���W��V�Yy~~��09N���]�`r���p�r`��ɹ�U�zevA��t�N���\1^U�Z̻Tf,�`t��09N�������z���*�N6�c���ϳ3~�z����{^�۝��9mI�f��A�H�n=��s@꽯@���hW�������0��Acr�<qmd�Ǟ+�q��i�ub�݀ȹnS��m�K���q���u^נv�e4���J#��mX�q��L�9 �S3�U��gt��"�)2^:�1��:�k�?w�R��nI���G%�;Vl%2�^Հ�M�`<�krLX6�1�(���.����^�zm.��{^���v�qɂ�+��)��$t��:[������x��k�QZ�m6:��\\`ɮ0�ՙs��-�����t�����^�O9V6�X/X۵��u�X{��%��q��x19�U�{��!)���ν�v�bd�ݙ�%[m���&��/������7��ϻ�8��
��G�6��b����yv����@�6�IƜNf����U����ۚU�z����$�B����b
�If^4�]:z�䒗}.�I.�=^�I
t�i$�W��������g���љ3�Ɋ����ɪ24(/fv��$6�p���酫�tnL�K��7�$������I
���$�v����IykrLX6�1�(�z�K�����y����5$�/��7�IV�[�g��K�3¾���73����Ԓ^�=^��UWw��~�i$�Oޯy$���!��R5#k"�)�/f|�/����$���ٛ�����9m�� ;ljb�V��X�b���n�m;�-�bW�j�����J]��i$��z��%�X�I{��{�%�Y�f
�el�l�a����i�KΓ��M<��ۀA��d���A1g/X-@,� ��������K豤��I���J]��i$�wK�8�q'q9��$�_j��K�m���$���v�Iot�{�%Щ�!g؂��Y��$��OW��R��K��w�~�{�$/_9�$�w���,�&�I��3�䒗}.�I-y$�:^4��뽟�m{�IW��{&,i���DӍ�I.w��~���\��f�m����r�{��s7m�����+Xâ �LH�0G-�p��/H֬	�p8�"��ԋӹ굞L��؇r[<gk$�0P�^[���ã][md����.�k��v�t�m����GKع�6��t\��]lgO���*�;e#r�O\�q)���ƃ��Ѭ�Q]XnHsz��L�u�F�W�$����m뙞zSǇ����w��ۣ��s� �e�.FyU��P�m��f�[X�g����[���%��2�MP�>��ٳ[��͵�"vM0�p��&]s���YqAqmF�%:�g�8�mb�f�,>￥�_�~�n�o�|��xy���߳>E�e����~��^y|�!��R5#k$�9�$��z��뾗m$��OW��B�/U|�Ie�.%[I�����s?~I.���I%����$��KƒK�'��I#�(��m�$�"I�ޤ��{g��$.Z��I���K��]�$��]���J��e��y^�I%�f4�^�=^�Ir���I.w��~��]�#��JLib�F�o:�M&fzzuû\��]u]��cJ���y�7Gg�� �>�1���jI/ݷ�~��]O�[I%����$�[&cI%��T�U���5�kF��S���n{ۛ��LB�ē�=^�I%:f4�[#������_���x�G"i��$������$��4�S����\����Kn���j�`��Z��y$���m$����&�D���f/_{�h�_-�cs���QI&���u�l�ڰ���؄��c�~�C���MٽMš+;V85�B*w#�u�39���h���=��[��v�̀�V �>5�:g fq%F�7P�F�4w� 9����h�ՠ~�U4�$�R4�&i$�}�$��f�Ea�Q"�X
EV*�$`(4"�
�1˚�z:`l+� 1>���g,����s`<nՆ�3���)|jDq7$�L����h�3�}���޾���/[��Babnym�l��vn$�k-���Mh�t(�g1[:$d�O��M���w4�٠^�M�ڴ,�܎9�9�ol��f�k�Z��#���n"F�m���@=}�`I}t��RK`9IK��m<nM�}�@��s@���C狗j������}��'�[�off�İ�I]�`wH��$��L`w_j�?.g_ɤ�T,Lra�ę�_'ogM9d��H�M��v�nݸ�#��0+� �e�e0<���6I���UU}��ۚ|e��i�O��8ӏ@9m�u�L�0<��������3(̬�����:`yI-�l�h�VW��i�����۹�yI-�l���05PBL3.�����0<�K`$���L�6nIé�]o�F¡��#'t@(PJ�_`�c��cGkS>�_�`��Ob��}4���a'<����b�Q4����=�L6d `A6�`i�P��������O���G1�b��}`���S��`&�:`�+�� {֝�M��Lv���Ѩ����M��R �Pо��Ni`��<5\8ĐEښ~B��<E������,c	�Dͪ� 4����0������c���	Y(I��"V�XHDI��@�C	�EB!�TС�jbl��I�i�ѵ\�k�bH��̺�-�		8��ŷj���a;6f�-&���I�z��7��Ե�5���89�B�-�uT���*�h����`�7B�HΑuÐ+(N�پ���R�3�pX�6�%m��Xy]l�4���0ObX�+h��U�q]�k��pg`�r�gi4�b�oj�;�8��d�h�lIYp�B��N���W� ��9u�3�tpl -Oon\mKq���F��j�+�/͔�Ʈv�V��+a�,��œm�%�R�R�Ɲ2�u����@j����t���AX�8gnj��T�mX�Q�e�� =�m�$�i3������v�m5P��j����0.iR�v�3=r�mu�mkr.���3�}��9v��k��v��Ŝvۧ�V���9Yl]�*$�(;N��P5�+����7"�5��<q��i����	����/a��6+X]C��i�N��F^z���3�{,�O�ґ�X		���v~����[! [u]V֫��L��4�һ=M�s�l�5P�>6�!Jv@�GYͣ�]�K[��UE���d4-mP��:z�v9̹N����u�4r��i��n�cD�5��Ÿ�ܫ�ێ����*=:�^�팛��(p\�`��J̆��
ְ]��a@K����Jy��/2=]X��$9Rwb��R�1��h�;]�m�q��l�'+4d����2s)�k�I�5�l����):�(-�F�^y�9��&�����r�jRy,��JQ�mH�m�I��b�bz��L`���@��O(�Y�d�x^N�kXHa�n�݀�G��2��Wm���6�sR�0Rڕ[z���3}��f���LGb��̘�V2R�e�=��z��q�VN�m��S�2]S�<+9p�u�6��s$Ӣ�X��$��U��r[��I�M�MZ��m�LAYi���p�k5�vżt�l��)$5�;[#���أ�AjS�j��ej�n�#fA�c�hV�uc@��]R�j6��A)� �G��61_
 ��Oʂ��A	��D��x�Q1��@v$I�<���bQx�$8�ܹ�@��D�Ly!�������8)���������W��]�F��Dm0iz��-܇Y�Kd�ƶ��8��cL����nƤ�s`.we t����nkW2���0�c%�2/G�xԎ��ų�=k�N�m\ 	���*9�MN.֤���쁺݉5�qR����Aw�WcC�Tp,z,�rH5P��g��ڲ Pj�8����[a��u�kZ�z8�����8�"s�n�j�зe�$�	<�O�꺸hEݱ��n|�z�y���+*��l{������:`yl��6*]B�$�i���94q�������^�v����>�Խ�g�X�iBD�W&�z�������aD%2={�2���{[4Q�$�R4�&h�-z�L`n�D���a]A�e����= �h�����ۚ\��m�x�翻�a�d�L�/C�+��2N�әt[����7l���[����aj�'�I?�g���s@��� �h�Օ�hx�F�mŠw��k��>�zDF+�P�E��HE�T�'�)���M�Հwsy`w��os�ϳ:�</{$�A������`$���L�0:��T)^D�M�F���}�%�{�@�]��;�w4˖� �X��V4�i��Dqh��0;�t���-���LwB�yn��i�g�\ƨ�����(��J����-����<<`�<U����f7j��z�Xt��Q	}!�Of��l�G���M)3@��k�f}��ݛ2�́�ݫ�2f��б�r����r��ݛ��sf
�I!�J�j;� '5Ͼٹ'o��n�ˢ�8��a&D�Z8�V�����[�2	�ʥ����+.�]�&�GL�����ll�09�ڴC:֓$����r	An��M�<�X�rj���Kd�������XN��t�Eb��3@��k�9]�@�j�;�w4�:�S�$mA�(�z+�oR�2fSٰݵ`}=n��'�e�̵t]���ݾ���#����Wj��R����Ici(��Ԣ[��X�ݫ������
 xU'�`�E�*� =�v���i�I�ȓ��~\���D����GL�*�\�)^Z��J�%k�5ф1���J6����k�k��ټ`Ǩ0�5��qǠq[^���S@��ˤ���Te���3+	�*��gz�D)���Ve�Ձ�m����hl��n{n���uf�
&rwv�o�X���+���v����`yt���܉���9۹�s9�2���j�F��?q�6s8���j��q��>��+D(���ϣ�~��`��j{s���O9�c�R��ѫ��8#=b��X��<ݬ�桔űv����W�=��bgi��0ݹ��5�'O�\ٲ���W��7C�Xp;��U�Y��#����z�֡��ƺXkN�[\Bh0��'�WB�:ƎItҲ�6�M��̕�s��֔�26
u�Y�����m�LY@��e�<��\���UG�����{��wo{���6vs��؛Bb�M�F1�Wgn`�#:�u�6�.g����x.A4���]]��~�������ˤ���Z��W+x���KHR9۹��L���Vr�f��gz�IL���F��pr$�&hW�z�;V���S@�;w4�3�SW�5��qǠ~�76s8���j�TD(J{Ov��� �&�&(�Z;�M����?.���v����1�m0Ŏe������7d��>ݭ[�bx"�^�s�q�ݛ�n�̼�r49ȜI8���nh�mz�;V���נ~X:�E�lK����uyQ�(���M���u`s���3�S)�̑���n=�۫����(�2�� {�� O'[m�#O��Ǡu[^��۹������;R�ĚjciD�Vcv������ݫ%�V�~o��fݰ=���6���h{�f�Pֺ��ua����W)�ۙ�WZA�@�V��X��X-��3�z�!f$_~�Z������NM����:����� �&0=�Ti^+/2���<�X-��3��Y�Q	H�PBB�(T60�&��M��}�U|æL`j�-��R�ZW��D�IǠw�S@;m���{�ϕ~���k��D�)�5�Hhm���$�)%�;�A�+d�J��v��4���Ŋ1�x��Ԗ�a3i����.�8�ǉ�	����H�PmAI4[uX-��3��G���X͗F��NF�'3@궽�}�E��4�ޚ-����v��Cd�Ҋ��� �:I��:`r�[�ճH�M'"LN�>ϳ������j��mՇ%'��!��`�>���!w���;�(�3u�rb�jk��>x�X-��3��X6�`lv3n���8�=qq�!�v:������4dhP^��-�Hv�3�L9�WS]���߭���� �&0=�:`��.F�9ȜI8�s�s@;m��[��u[^�1#��xO�"oƚ�ܦ?~��l������tt���nC����6����v�hVנ}�v�6�J&^���d�UUS\�M"�$���۫b;�~_ =�����f�"���Jx��>�<�<d�.�^)*�u!`�t��`�ι\\�n&{v���-<ܾ[�r�Nm��c��6�l�d�kX������s��n� ��g�Y�j�v���ʹ��z�d��]�Bٖ� w:�3���3�1[S� RNWL3�TVI�i��0�7k���ST+�5c��vl��M��&d�ν��\U	�����z=U�e�%��-�����<�}^ks�<��!�."�ܥ&��K�.(�W8�EU<r�n��<;���&<M��J'�{빠���;w?� ����9o�4���pr%���L`{�:`r�[����]A�3�_]�W���tt��$����hm�@���Պ<Q�L�ILRK`{z:`$�����U��� �'N=�;w4˶��;w4u��e�J�x��@��d[]�&l7"8.a�cuu�K<�C�f2��4��v��!R&�Li�ә�����w4u�o�ws@�-[���8�!Ś��9�ٺ$+��� B��V���qڰ>�n�T)�Y��mU6��<$����-�;w4˶��;w49ԮTǉ�ciD��=�0<�K`{z:a��u���'�H�CND����@������U�z�v�h�브JLib�F�j��'b��&�v��ݮ���E1Ss���tvq|Z0�>���^^[���Wt���s��ٟ�q_y��^ǫx�y&E�����-������[��� �Ϊ�x��"q$��?s�s@��k����o� h��x���78"l��c	�P������hvT|<(��{��G5X�#�za�,�
oӄ#��<��M�H�M��� #!	�B}���Gf�]���WL��q�P�	"�1!"q��c��@�#Ly�;����ʓ�b�8j�JJQ����B,mqC�|dkC i�}6���!��p��=�	LF� @�o�&�=�0K����D4�
x�@�M��^�z�z�U`+�� lDB �UJ"x�b�N��0(��pت�@<#��H�$L�%U����M�ݻ����.�=֒�d��&D�����=��Vq�����aB��o�f��|�!��$q�m(�z�v�05wK`{z:`yt�����3-.�[�]Z�� qhCB�K`L���a���CD<a�p��F��{; ����?��ʰ>�;VӍ֨QHwڰ�gsɏd"�҉Ǡ~�n��vנ~�n���נ~�kf�8�ND���IloGL]��ގ�9Q��ϲ�����`{z:`j����ٹ>|��\@��⦨XJ�Q������?s7$��꿱��(���4.���;v�]%�=�05l�����
����d��D��I��k���$ZldUԆ�:���2$�(�x��"q$��?s�s@���Xw�D(��2[ڰ��Zm�*Q�ɩ���>�n�T(ID��{j��w�@������o�ndQ�A��q�z:`j�����ˤ�[�"��NF�nf��31u��{�ی.��z:`�����]^+Uv�+�`M����[oGL]��U��w�w2�p��.��uf.����go���6����-͵��է�;=��: �C�q=B�RX9��HZ�廵z�����ܵn6�ڷg�5��Z�Nj�&5��x���J9e�/4����L�����=�;X���m�*��5m\���;�;������t�<h�ht��F���sY�ر���c��D1�2R1���nX��Μۇs�Ͻ����N����v���?�c�_��-�OB�8l`���ݺ�6�b���OE�4���V,���̊���Q��s(_�瞁y۹�qw���~A��nh�a��Z��z�n�����}�j��q��IBJd��u=X����rf��o��y۹�~]�������U��� �'N=oGL.��z:`j��ݴ�t��5�4�s4˶��s@��k�/;w4�̹�8�k��K$��:.N��N@���y%gOU�݇=������ZX�d�rm(�z�vS@��k�?s�s@��k��
��M8�x0IHl�����OP��R���F� �WH'G� y���7$���ٹ'9�M ��+�1�7X�Q8����`yN��=�1��z[����� ��e�2�S��oL`rޖ����XQ	�F����**�S\��;�y`d�Xw��x���	%حF����j,��#�C�j�pt��s���̆������1���+�l��.c�3ĺ��?)��loGL)����05�e�a���W�+�`{z:`yN��������׷�ϒ-i,�d������qXK�V��2ɇ�%BJ�BMBO��#�%�����ܓ�~��rN��7�9��A������M���@��t��-�x�Y.�Z��WE�S�OqՁ�Qǿ/���ڰ>�q�;�)���1�`�i�d&9�)���ג��]��W����'�ݧ\ ��Y
�K�=�0<�K`{{ ��/@�����)jF���@���`rޖ���t��ʏ������-^[��-�loGL)���\z��l�"�W;^������9{�sri�aaʠB5$�����B�����nI坝�k-�r%�8�q��۹�g�fq�����Ɓ��נ~�u%��F�Т#Y�c����������z,�l�i.K�w)�b �FIȈ�M9��{^�����:�����s�ۚ�� �"�B��Xw8�'������XK�W�bGt�<�M8�x0IHhv��ގ�S��=��`ڔ�wWv]�L���Mr�6"!B��ߕ��[�`}��4.Z���m��!F�j��7nD���A��d���� ����!�Z�N�@����n�\4+3��j�N�\�n]ur���v�qʹ.;Nؠ�bTd�9��{=kWS�t�hS6[r,f�2�ժ{i�,��[�<�R1��L��pdB�{c%>$%L�:3�`�͆ͅ�����:�0���(���\nyǭ��i�Vܘ좧N�	y�������}�<.뺝U��p�Iusd3�z�Y�f �ڔ����*|�tj���|��s�=a�Vx�R洛�7d���<P&KL�mp�vo�����5�k>M,6�����=�c���v�&�[D��$ȣ��~�@�����}�@���h�ƱD�K"p�@��t�ݾ���� �Ɍ�IT#$�dQ&�Nf��>ՠ~�e4�-��v�hy�L�s"�B��@���X�o���j��k��
����g8�]�6G��i����8��gZR9�6I�j��t��]*#*���<���0=�07o��^A�3��3�J��Ƙ�icjɠ~�n���f��٢)M	��L@� 	�RcUM�@������@/�����zx�ܶh���Z
F�-fZ�/)��}���ގ�r��a����e�&���&0=�07o�`N�U�Q���+X�^�&0=�07o�`{{!�w=t~q���,rC?��k�@����g��bx"��Cr���7RJ�휔�CB�X,��:~�:`n�D���A�{d�z�YJ��2"&�Nf��>ՠ{{ �=�c��� ��eaw��/0�U5\�&����X�o�(DBP"<P ��A�X�f�ϼٰ-}������NF�0IHh�L`{z:`n�D���A�V�]IB՗yiU���1���遻}����@�3��|���P���D�Y��{�㵞�dz��Z����G�����S��#:RpJ%1��s?޻�~�e4-��ގ�r���tb0��w�������W%�=�07o�`N�U�x��U�^-��ގ�UW���Lod��Z����]2�~��oOަu�Ɂ��R��1���B"B('�Th�R����ܓ��,�_�f���2ڼ���L��[%�=�0?��������ػ]�)�U���Vݓ��=sc6e�׮�X��6�sV�f�r\�beb������[%�=�~����Zç��i�O	)��}�}T��?:`w\����0
�K�(Z��-*�U�yloGL����0?.Z���I�"A)�H�#��ﾪ��ݓ�`oL�0<�K`{z:`I��Z����lJG�~�e4����'��F���y�nI�UUE�  *��UUE�  *� W�  
��UU��  ���QO�"�`� � �"�0@��V�F"�1
�1 � �"�0"� �"�1"(�(��  �� T@?�  U����+�UUQ_� Z  *�UUEª�+��UQ_𪪊��UTW�*����  ��  ����e5���0=.� �s2}p��{ �@  �   @         � �@PP(� @(��EUQT�( �(	�PT�A(H ����( �� X   0`  ( 
 ���ʧ��y^s�{��n�N[��� ܯm����c�o��ҬwJ���{��o7|�Kż� ���vn`���wT,�k�s�iӈ�� 3�r�MO6�7��ހn��x<    U  &��)�}rˬr�tܞ��P�}樂�o{x�j�Xu}��>�t*X�
���@ U��R����M�R�0 4    � P  @@ �   :��hR�� gT�bj�LZP�v�Ur�*�8 (AA@ �`	t*�ZP�3J�\�
�t�� ���ҩVZ��n�J��R����3ϥ��n����}n[�nW���|�����������x�W�����z�==]���9ׯO&{z���U_ (  � ( c` 8���n1����k�|������7�ח�]��������7�O���f���y� �����qg5�� \=�sr���n,��&�m�� �<�޷���W֮��UV-U^ <  P P�c`
+�%gn��^/����]��0��x y^ۓ]��^����w��־��{�B��,��nm> ^�����{���m��秧{w���g�{�y�W�y�����/����9��s��Z���^��ܪ� 4�2T�IJR �O�L�IR� �D��P�T D�*�"T � S�BS=J��  !HCRRD@G�|	��������3��������u/g;�e��g��q��aPAW���/�A]�����⠂���A_�UeQ9�?��Q�Ѧ޷ksA�BH�:s����.9��M��7�\沠��0�Ibq!1d�Xe�RjJ�YV�:<�w1���c>8��R��4H3�� ��a�{�ҏ��j�bHPi`���chgc�0�ӡ�EPU����˯8�1��"��|ûE�oF��|��7�oϬ�5Ü�L3|�E��,�p�)3*d�Y�0'�0#�ĕ�jq�p�0c��ć�0���#�Fi�l�Ze֜�X�:��3V캢�����5��FZm��lDL�N��	l�0$��pB@��
�0�B��Lf��U�f�I�t��w��_LHDE%!+-2ؓ��o;�E�4q����.(hiY�����lѾ��v
`ܓ!! L$9����[<<'4l80T�2�A3���]:�7B˺�P�^�{J�y�6����W5���k�s�~㇆>�,0�ٟa���1��l>KԘc ���DX�D�����==�a�n Ø끽��"*b	]R�J���V/��Ov�{7sL��p�H�;�4X���"�0���Ӫ�m%�I��9����� �$�%"D���}p0���O���bz{�X�O$4bh�Ģ)���e��M,��决`Y�6���u�Lta0	0;	0`�r�ő���z#����2��ؐąp�5;c ��5Nkm�����< ��	%�:c9�z���'͚�vJL�>[���h���KS�� �HI��6j�،�2��QX�d�$������ݭx��Ɉ�A���"�&L!\]$b6;h"̵���ܘI��u�<Ҥ\��2gC����gvs����p�f�S�ec#0���5�3�1�;����[�k|y�l�7�,̦Ň����}�}1�m6�WD���`�K FF������I �T�.B8)L�02BN�6{�Ǧ���Q��b�,b�#	���  d!§��Fr�\��5��oe����턆T�ѧhh5��> t���2!�w�¼~z���P�h�R+�:ͥ��j���y���D��va��Y�u��P޸�����Hbj �A`F6�f���Z���i  I��H���HC �JIQ����	(I�$�`��CJ���$�)$�$"P�dg �e(2��LuT���a��6i'�� �L�c���g��P�8�lpޘ���' ��vh�D�l����<,Z/0b=%�i�Ƴd���jj~���s~yk�xk||�TE������3;�=�;�	�3Ph彻���Ň|;��	Ǩh���B"�ͺ���;ĆG��� LY �"�)��� $�A���鉁���%.�n���8h�FKQ5��8��ϴZ],�Xh�O�>��8��Af���K|`�l�[>��٨�D��
s#1�B�_]�MJbC�1�#����>*60�8�غ��>a&4fx�}cx�p�Xj�Mk��2��n��!1���u��0N�,$�� ��C�&��$!J$qJ)����B&�Y��t�931!��1���,1�`K8�驣-��V��*�of�D�3�a���Af�&j}�,3�.k
ʳ�2$�a���
b-G�mȍD�,�HXj�	Z��hV�!ZLj���_�\�VeV:�sSSf���1,�ݜ��c)��U�s��9p��
d'C��I�%:њ2Z�4Z�gv�� �K�X3�`�D�:���>7��*c�5����Zѯ�n��3���ׇ�(>��{�0�� �Z"H&F��XBVRY#�h��N�a����B�	R`��D� z$,x��A8O<��<Xi�+LѠ�ӦLөp�a���}s>�,ղ�F�:d��'ƈp* �����m#��ޝ��tI	Lc�dh��)()"#ȒL&I��	�d�pᰌ�L�'I�$;P��\�<���}��}��������y�{l>�~c�q�a��	fc4��h8�kv��߇3 �,�Vh�I&Sm%�+-}�o�"�Ah5���#
2�9�aI�ЌH�&��.A�Hb&��J1#������66fY�`K$��HHD,�d��,�E,0Á8KPĲKR�K	D	&F4FI�8�U��,�̆b`�����b��)��,2�I��6�E�Vi3DF��N�hmK0����U�N�0���5��5���*��I�>N:rOC�ŀ�l4e0Υ2L rW1e�$JIHX��� H"BqHR	�O�81�����ji5�|��Ȋ(��}@�$�H�ŗ
fA�q�F�p�l-pt�*�0����dDZj!��H�!a�ֱ��z���^��´��9	),�,��XG��y��k�;1xld���qCA��+��.Rh6q����8s�W�%��P����l�?sy�՚KX�1a��fV	�Qi�'ɝf��}湣W���F�b��H�KA�&���D8��h�
(4�8C�-�I��N$K2T��bk���'�g���ﷇ���H��i#	�6MH��5nb%� �ў�ϹE����~_Y�d$D�%a�}���q϶y��g���f��Aa`n0�B1	��&C��Z��&��-���XU��a�#L��a8Md��l��݆��:���#,|��a�ǀ�%&kw3��>��sE���%����p	g8'ϡ�+l�4�}kE����h������o�6Z8d� H��$�����LT(eX����8h%�,�d"�T�.��]��e�$�LH�4�E2m�i��vm8�8bI(h���8��!&,��!+1�Y�SLfIq�1!$�pq$Y�*CL���d�9)�:�%$�62L8Z	�͘��M[������1��c8:4f��g7�>���v6h]�A,b�ĝ�,�������[���l�2Ιd�8��o�H����~z`�q	�da�~���<�5�5��J�
L�ADA�a���h�BH��!0e�a;�w����{�� �$           m�                    � -� ��   ��                         6�p                       ��                            m        -�m~���b�݅J�-Dd(n�n��h    <^���[l�Lp �������ݬ� m� f��)Vk�m��8!�h��^��mT��	gk��� �   ��m[��:��ۤ;Z�:r@5�XI��(�jՌc 6��YL�r�b8�leYjt@W.m��6�m�:tK:�$�aaߩϾ�ܾ�Zm��F@t�    m�N j�lv�l^�f�8 ����%��]�np�L���$pM'#k�l 4]� u[R1lJ��iej�W-�� hh� �6� ��Ŵ [Am������I�햗L�	�Ŵ �kh�+j  �(�j۶�]�j�/I�6�*ic4�[@��M�4I{j����\ �ղtI���&�8  ��6i6��`-��m	D��e�� �e�L�CZͳUU�Q����eU�ںI kY�l� ��&ăZ���$ �YA!��6��-�[Hu�e[�ZWq�S5K��oam$ p��UR�!P�A�\qp�;#-���=��Wi .�&��Q�հH :�g'L�gkz�$ m6�m��n�[B@�[�Ć�@�P	��� ]�Z�ۭ` �����m�m���a#��K��[��m��mӀ-�@[B۵l6ؒ۲���^[��l���u����v��2�9{E�$�9MJ��i:��JےA�m��GZݐ���L �@�m	 �� $X���k���YW+���@I�\�$���[� �C&��[x�� �l�Y,�F4Q&��5�j��&�4�ͳr�T� �e��n�[@�  y��m[m���MA!m8��SrA ��lH*����LU��Uj�շ ���۶ֳm�9�'Y�Η�,Z��-�5� ^�X&��0&F��^ZU�*��VU�٦��-�4��n�@n�-ѭ�}�t�-�i [W��m�n�Lm��m�-5�݂Am ���&����j�a�*��bU�mm۫`e�$5�!#8j�
#s*�P��s�m�o68 Xc��
I@��h  m$ڶ�m�l	:�lm6[�����a����-�10=z��sZ�0 J�P�Ӭ�$��K۰�e�ے[B�Y��M�m��`hm�kX   �cm�$�Pʀ����Uu�,�&����5Rխe�Z�%YUr�ʹ�V�F�-�l ;m�ml�x������@�`�[\m�lp$GP:�o��ﾕ8n|�V�@E��J�� �m��6�?�o�|��m&'D�h��m,���iI����X`���y�m��ӡjN;��t�+��^Pv�*�tTjKZ�]����b@  -�kRd����Kl�5�����m�k���7#Um� q� ��`  8=m'mu�T,]�"G)��m�%t�j��&���m�5� �v�H���h  �` �ۂYC�%�f�ܔ�vU��J�2��UU��k���[rΖ��ɀm m��� �  H��#m�Km���Ŵ   �    [[l l�F� ղ@�A��a��vH*M�֦��D�IS[�� h6� l � ��  �J �m� UUմ6��^P5
u+�-�      ��d� 8 � ��Ā$� ��@   ���I�m�k�l8 d �`���s^m��϶�}��yYu�Æ�K`�W�V�`���| 4����1�������lqͻ`�[p-�� m� �Y@  �   -� �Ā ����I6-�  �f��;,�� ��UK�˲UT�T�)j��Ka����@���z�^�m� �J$�r��՛� �� �����鴐ڶ5� �m,�@si���k H�[�  H��K�����V8�7/-m[r� ٖ�� �������:-e[��mX$6�nj������m�p[r��u���P-Znk`�r�]|��I]�L
�f��:*��5��dg�Em��!v��q$�	 m��ͮ���6�[y� Ӥ���2 �`p� $ p [@��ے-�@-��,J�s��9��[�
h����6[�M�KP�e���PP*�/ʵ
�@U*ԫUR���4�(d����5��L[% ���7L6؝���M��n@��l�cY-�/`H k[$�V��6m�$ �a�i�6��aס�m T�U[�`��������� ��M�J�@����תLk�-6	 ��-�mm];i 8[B��h -�l�3�TAt�P �m0����f��@z�m��t�6�UT����uU�6[�6�%���[R[v[��H m�cf�H���� m6[����[A � @   n�#� �v�U�Z��)V^[�P6�m���cm��������O���l� ��im 8  H � � At���[PJ�TK@T�*��PU*�P> 0 -�h��mm$ [@  ���մ$ �� 6�m�@  H ����[���m�� h mж��e��` [d�  ��� "F˭��i�  "J佋[mm�m �b䭶 6�H�of�6�$��L�   �Y%���L���` �� m�[m�j�t   �^3mQal�j�m��e�0Ts�d Z٥��	U{HV�
x,1-nZ)��A���P:w;�f�mU ����]UVݐ�'YUk������>প�p ���E�B�Žz����Ym��Z0�::t�]� �sm�  m� ��@��m8m�� m�E�����H9ml[@m�H �eknUfUU�lp lZ`[����2���m��\඀�@	�-��I5�� -UR��UJ��/6�*��ޓm���! ��n�����I	$�`����6�ko[C�h;vZ� 9��v[hm�m���>8
S%�U�B�* �Y� F�6ذ���o���0�6�$6��.�P P�T�UP�H�m( �1m$m�j@m���	e �`�l��5�  �	�ܛ�j�(UVҵ�r@��5�
�Q���َٻ`�a�ŵ�������Zl$ Mlmխ�H    ��q��r�]���H mי�I�Af��+`6���$���&9J  � AR�v�ݖ�ښ��դ(,0�E�l�`�f�X��6�[��։  	 6� � � �� 8��%�7m�P6���@���� p[Am  �f�$  @ pR�m#m�K���͘:U����H5J��tqz�p l�l 	   	��8 m��m�i��rD�6�j�����I��ӂ��8)Cm�U�[@��$-�6���~��-� �	 m��Am-�ڶ��"M�8BIe�b�n���[Vl� m� 8�a#����l�H�`:�h8��R[Ӡ
�A6� [A�� ��m������z�o�zt8�c[�� Vݚ�Bj��UUU�z
�i2�:�����,�V�Πm����u��Փ*�$j���ٶ-��m�  �5R��iA�� ��ۭ�f�6���p � �Zm��.�U@T �;` �� m��v�i��m!#v� �|Hl�zF��W�  .�$ 8��v!��V�*հ@C[�1��SS�m���d� I'\	��X�L ׫���ٶH}o�|   � �ۂݔ-�� t�Z��6���@�mt�WP�ob���� %�k�F�  ��S��}�e_ ��f���Wf��������TJ���P���$@�(��?��!p&�d��x'����M8�;T��P�DÏ��0�ꪏ��~_}@8��=8��M�����"� o�*x"�<C� Kx��P> ��> z�Q�v:�(��udS�~ ��5���C�| 0 !�v�*� _Q��A}O��A�(�T���TN(�����$�}���N�@6���E=8*'�x�:���/S�S��j���M����� � ��:M���=Pd�(�+��=E� � ���|(�@t?"|'z����S�Cb�2� ��p@z( ���}���Ὀx��<N���(�.�}:��8`
�/�
َ*z�8����B�(0x|�P4 `��C�hE` �� р���;U )����A^(����%`$>���.�8�,�ዀ����!���Ot�~��- �   	6ۍ�I�l    �    �     h �ҝ�M�Խ皕i��9��<��Z�.�r��ڲ��..�[M��ڠ�\BOl��zG	��*eML�C��sHI�0�蛫4�����9U�j#.��kfy�r�m�YSs�����/d�y���;4�#���i�ڮ������2��{c�L�Ȯ�:�1�gn��WP�B읃q7�d!p{�v�ە�6�0i���"᳹�;vuܓ��и{c�n��w*]L%�(�98/�ι'bwy]��F.5p+����1��U�tnb �eM��HmR��]mm]�5%�9�Z1oh���gm�ۙ-m3�d���:	s��\¶�l=�_mW$�j��:v��gk�"Sn��yZPr����,�"$��� ��F���H[�[R��6�t! �bMId��u�vJ��j4�e�\�&kx6!�P��U�V23j���b�ʥ�Cs�i@d%�ë��#n\c�vїH�em�P��r�  �[nv2�6ܤY�TJəҝC�n;u&J�VWA��m�]� �ud�˸�їi�*\(gc��Ɲ�Y����.�l��'I�`Z�%��K+��u�YiaZ�4<� �Ժ)V|�S�����:8��*�Wu��Z		�h�[v�2��)�[&����G�Tŵ�ls�%�r�Pb�F�X#)[�Lצ��:#�m��rnqhVwc.;ۚ.�D{!*m�nRWgv`�Ypf��D�N)xn
�R����$!:Nf�eG �;\�-�5ִ�J��)���x�(�Z[H�ѓg��bA�e���q�6@@���W�$l:�9y�H낪2;\��i�Za��Ip7`@
���n�wj�i5=�U�gMҙ6��r�+ ,J������v�l�_.ܖ�:6 kiM:�]��[U�v�+�-�۝E��~G�T��
iT�����x�z �Pv)����vxQ�v� �v��ֵ��ְpl���+��Y�^dU&�]�����06��ǰ�d��S��5��+��y�j�u�$\m��b�����%�y�ꢋ�(��g�q��㇝i�@S]i�ն�<�n^}dN�r��ZP ���lRV��M�������t1������R��ب1���y�SI�oZ)��8�6ۜ�6�u�{�����t����V�̲՚4Yf���۱��{)�]�v���!��k@�HM,o���B,�of0w^ۼ遻qK`!R����E�̡f,�`�1�}U_$I�u�W��� �-1Г�6�K$y�	�0;���6L`�1����ƛ���0Ć�π����� ��'�����D��J��Z/2���1�zt���^�
�J��|�ݻ��n��8,�t���[4�27g���bح'<�V�q���Y2<����q��=}4��������٠}R���ǌ�H�rh�w�4'�L	T�x�qլ���r����h׶h�v�ǢcD9�-��&ɌӦ0'tt��	,i����hq��y�3ʒJ�9���=��X��_uy����y�"��fP�f0N�������K`�ـz��K����ZhNƢ��,�7D���v�1��Rs{V�)1ķ��@�qlp$�<M�����}��us�^�^[4��4���cM�i�bCO+�Eҿ[ �&0N���������#֑����<o"hrdz���@<���/O�IکJ�� ��{���Z���]�je���/1�zt���[ �l�>������?�)�M��s@�R��1�zt�]�UYt^�Һ������b��k�V�T<������b�"lpLa)�$s4�w+�	�c ��	�0<�D]Z��M5 o7fyU�s��{wذ�w+���ʜ�"�"�h�n�{�Ň����W� {����V���6�i"H������+�����U%B��9�K7$�����6�F�9�$Мπ���= ��4�Z���s@-*�)�MX�M�7Vͫ7a5rU��x�ɴ�	�:�,\�G;���X񼉡ɑ��{�@��@�{���_�;~��y{T�M1�5����`r�-����T��&Ɍ��?`}��+z6!��H'#�/-��9{կR�����L �� �v�w�la)��4�w+��٠^٠^[��|��<j���<y�N�Ӧ0&���}Q0�}�3��mh ����ް;m�9M�Hkl�c�rE�cF��ѺN\O@:ӭ�����̛8ͩ���[���`z�b��-@�B�>��|����=b݇�MrTS�Tݬv��t=��g��D���=b�<����ݻtۥr�:��-��U�r�nH�������>8b�n�/`l��0���'l�ny���9�YV{8���}���9�\ٻQ�g�蝮�˞��M�9h�[��!�"H�(ddnI�qI��I:�o��6GL�ꉀN��*3t+���2�dtϾ[�-�N���4׮���ǎ`��9�Wm~�;�0N���#���Z��lRݎEԪ�+�n�`=��廚W;���wl�#ƛ���=:cl����[ ����{����@�;WIue�Nݣ����6��2s�]
��U[r��l�kv����C�Q%�����b�;|�׀���$�������m�I�!QRf����u�P�@�4��u��^ov`��,�vr�ޱ�~���q4<��`�~���z:`rީl.p���1)0RG&��3�\���?t���z��	�1�z�*�f`��w�����ގ���[ ��׶h�%SŊ��4��70����m��%�ۅЫ$=]2�gX���.֮7����l�`��Ng�U۞zy�4��4����;j$����ɑ��� 篦��}��us�^�}N㭦�Q�v�r`���{�ńUJ���"�� �_6��k<��yl�>����K���&�y۴��R�ޘ�=:c����ҳ11E��`rީloL`�1�y۹�}��V�1A�ɘ�$q��e�9���qQM��Evv+1N���h�@sغs��&��1�����h׶h���W;��\�YT�c$R`��M ��ٞ�Uv{��X�uy��0��BL��ۃY$�@����:�ܯ@/;f�}{f�s��4�ǎcX�[��}������ݘ%U��w�����3@��jI���&�q�x����J������ŀv�կ �~�/�:y�ۙ�8"�t�� ��m��ݞH���f�D�z� ���t��[Q����fc ��	�09oT�7�0>����1?�'�M�s@��r[ ���L`v�Wv���� �e�)��z��	�1�zt�ގ�*Px�[�<ǃ�#��٠�1�7��-��*V�Ȳ�*�jLJI$��l�=��}�Wny�}���J|����T��m߆W.o���� ��;Vۗx�vzn�MlIDK������ns�y��
�)�ݗ�nf���&�y��zڵHB�^Q�cnA�jpc�k����6"�u�h�[qr���)����QQĭ��t;	ܹ2�+.�k�\��]q�����բ�v�y�6�U-
�W=5ڴ�tY�\������ܖ���aɨ� ������w�u�.��܅�6͵f�]��慷v廤u���Mk�'m.h�=�ɒ7m�k��?O����K`zc ��ߺ��E�'�cX�'3�*��= �����n�z�jI���&$䬶7�0N�������K`�q��#i�$��l�/;w4�:��m*J���0�kMmcbn�⼼�ގ���[ ���Y�vڵ�y?A�ӑ'X�X��-u\0�sv���⡬�Ƶ�D��qե	^�h�-fS��K`zc ���y��ŀr�x;��F���ƣ��{�w� � � @a��8�+���&� = 0U�9�w�9�w4�w+��²���F�Ħff0N�������K`zc �.QА#�ۃY$�@����:�ܯ@/;f�}{f�}�ח�,�<s�t+��t����S�c ��	�}��~~_�{�^��=[z�=�\��&��u���0�7m�v�\=���B@�+���`zc �Ɍ	�05oUz�^��D<F�jI�r٠o;��_:��|�U߻�����/W�[/��Kr��0w}� ��^�*�/�`4�N�QX���k�x�j�I���L���f2"L^Z�`�2.���y�'5j��S*+��1k�O%َӯ��O% ��H�Q���b$��Ï��^xb��先�
�l�����d�ы��iB-mC��90@���%9�L�>�꧃�:"�EA�S >$B~ 6��>�:*/�(%T�PG���o���W���xyݶ��l$��q�X��W��^x�� ~�����_*O���Xo������.&�� 7�ـ{��~_��wذ�:����v�ְ�K��j�tm���u�l���ۆ�����rP�{77�91����O�篷4��,�έ~_�w}0����H�ۃRI3@����bE]�����>����H9���� ��,���π�_< �7fU+�{}� �ذ�c�&�LȘ��#��ff%{�M����^����a��6(�b*�JB�T��RUI~��qq�=�G	,hj�&�I�~��,�����R��~��W������7�ukk�L�Ĕ�ttEb�6ʶ��7
K2�fNϖFIb׿;���MJ��;c�.G-����� ��^ ~���T�Xs��X�}m���Ie��9!�v�կ=Uv�0{}� �;4ϩ}M����:w��F���ƣ�8�T���}?�o�a��}�ŀm�W� gs�YTr~�H%$�h{1s��f��_nh\�W��@>˔t$���I"�9��X�T���/� =�}4�n�g�{[nI1�nI$dRI*������+ή�ą��8�n�/Li�hd %:���ݞ�y.����zY�Թ���\�tu�tS�F)mnr*�Źm�D)�c"�v��H��U�KKuƭ�s��ƵFl��$��j���[�C6�ͦ�gfo��ڲ�N�iU��<r�,�9��P����]8x�#��4YY���ʹjϻ��w�����������!�\<�F�[��.���F��vf��p��i��Q������~��8A�!i�m����� ;�ـ}{w?� ﯷ4V��MD��yr(��ݙ�9��,��b�;|�מU�/��9����ԓ@篷4ow�*_$�S~�������mi���lu%�帰=J������0�����ݘ��UW�o�,{�[�ym��)��έx��������9����즁����`�H�&�B5�p�;VS:���4��=vj[�o=�g���Ux��Ӽ���q48��9�z`��� �;���%��o���qt�z�2;p��I0��Ŝ�U
ꤒ⤨IW�W��^����� ~��ϕ$��ë���	4��,�H���� ��<"���l�}�o��X���~Ni�Zwn?��J��� 9�z`��懳_o���c��Q,x�D�N8< ��ـ{��~_���|��;��?�{��~?���v��κi�a��b��V��m�;T[5��(y��t]�ww�럦�gKv��' ߽�,����;|�ԕ%���}�|��R߫����v�N#���o��*UJ����x��� ��qg�$�������[vIe��[��}��\����|��p�e	!���W�����߾�ʾ���~���N��#E�����T���z`����u�z�R�����s:VyI&2D���I�r��h�������v�z�-�Ƚ�b������v���kS��I����gV荒�Kzx���D�{���}�����tj��[o����;|� ?svz��/��� w_���9N�����I/�$�w~�`��ŀr��y�R�v{]�C�Ǎ�M$��wޚ/n���UU�o��m�|< �5=�K���n�w$��$�����v��xo���x(����NBo�?�w��}�Q�׃���Ӆ�帰_;� �%���� �}�s{���R����+Q>��sI	�N�c�%�с��k�F�]�����<�]�ws��
�cl�{o�|��7f����~���|�_���.��Ƌ��� ~��ϗ�ٿ{�X���v���%J�Ô�ͷ$L���$�@����8������]���s���e�:x�dD�L�8����7^ ~����U|��}ŀ�����A�qZwn?�m��x�U���}8��4.v��߿ffu�u��%$�d� K�;J�v^$��m�.el���~���A�̠]Gl;�MÓ�Z�r��0$	�J�V�b��oS`�K:%�۩�f�.�ঢҫ��9x���N�A���5Z��a.Y5ڝ$��殞�%U����I����8�rM��j�5W�lڔ�tA�.��/7c�.�k�͌[m!r�NP����w�tq/RX��e�w���t|�[���/_�.H��v�ɛ�%����:t��6���'����g�ǉ�M$䎀z���@����8����
��= �{��#i1I4owz����|���� ?svg�I]��x<�m����dq`������ԒUvs���;��,�]�mٖݴK*܏W�%I=��� w}�s{��<��J���|�_���.��Ƌ��� ~���<�%I.�}�~����:�k�-}*Y1㉤�?s��,���+H杴��v�Н�Y-�^L�u�%��ww���q��$�H�s�|}}��qs���n�RUU_�wޘ����$ӻf����������Ao�E��4�C��S`��S��g�=�*��o�s{��ԩ+��w��p����8�����< ��هԪ��b�;}�<{���DX�<�����{����w�ۚ��u�y+��y�zo�m�;j[M�&��۹�{�o��U�y����jK1a&L#�4���68�]f�4s�]
�j���oh2T�kv���}���|ؤ����*U]{��6��< ����W���s@��M�jm<"1�H��n��+��}�w��X/�מ���_���.��&��0�������������H�B��+���~��(���s��rD�-���LUR��}�`���l�ʕ�;�L ��x~	<i2"I&h\�z�e}���߿cgGL����R��+I/�]�6�mNK]P��oWHv]Z�h����;rb�*��~�/�7�q������r٠r��g�� ����=Z�I4E�[R�v� ?svg��%Tٿ{�X���v����IR���v߉,i�n�$�;��,�����_*UI�^�����L��5�ݺp�$-Ł�J����x�}���0%W�).�$�J��V�+Ԓ_��U���V���۳-�a q1܏ ��u�U$���w� ߽�,����~��z��q8�Q�
�&ʉ���IkI��X��ج�&E�DXמ����̘�kDx9�$ ^��@����9_j�~�]���\�g�rc#N���`��,�IU��=��}�� w��<��]�W����M�%�I�=���n�=J�]��z`�� w�,�8�v�n?���%�UT����x���r���>K�Of��}�~��ݒ�VԶ]����ݘ�K�U��|��}��;|�xMb]E$$%U�*F��GM�`x��� \H��b?`&��P4����},	�}HX�m�Ӳ�R9�fh�`ٳe�В@fN�@@͚��c�9���ξ����t������h �   [x�@    ��         � �v�Uin�B`(yx�b�c�Bj5��2ù�ģe��.��m�2�qđAD��;g��ۍ�a<�5UU��9Ο��>6.�����2�aȻ(��:0bY(q�z͜���cm�A��X���c�,�6�Μ�
�78�s�W�N�[E/2�rJ�<�I9Yu��S�i(�76�F�(�S<j�;c"GX9X��g����o���ۍw2��ux ��i̲����J����3��-�ǖ�6#Y��������r	u���v�H�,G t��P�7XB5�LhxL&NՋ��3���F��i�E�8ӭl�p5[g��Zp
�Q������7@�hU��%6����R�5KRU[9R�U����U��Pq�ԯ4���Ф����L`�;I�lmJ�ԪO�Re�Z�S��K{�b�[�ғ�gQ�v0j-Q�m���̨�!����@CQ�\��1����$M;�"�iմ*��m�[=��j݊ոիm�D9H$J��a�-�@��k���3�cv@u=q˸�ѳ�ez�n��_rf�S�T�$�=���Q�0M	9+Q%/]��I$]6k��ۚ�R��յ-[R4�I(Y�ڪ���Э�Y�:@@��v��sn�W`�.�B��w7M3Ŷ�je�)���BvSﺾ��`�]�l��a;kd�ݸ�r;։����NMG�r��)]�R-�+ZM�D��q��j�`ںۻuJ���K$P�@Pu�oUn�K���V��o���r��[T��8:�#
��PP�ca�	��Y^���9�^�Ƹx�J��C`�H�m���r��4�5.��_}�'����*;A�g�Pې{�M�:����g�e`b�r�UR���m�W8�r�_/5&�%�	B%�dK�[M��^�������w���wGȾ��}Nh~E���*�ǿ��=�N��C�z �����w��ۻ���w�ᗋ�� ls��T���:hY6�Q�S� ����+�NF����\�h�7����m�5�ڑq���v/OZ�v�<F;k���>6�*մ����Hpq�:`��7�.�q%��)v���r�96�<{vqz���J�Mh���5{k����h�G4�k�U᭗Қ���䌹ش �
���8��`���&�{���������k�l�Nv��\Xh�m�W=��-u���8j�z8s���X����Fy�A�g�5~��l[���K`�1���k�c�t�rI-ǀv��y����l��� ;�����^z��w�۳-�a sԏ@�����l��yz��v��*e`�[�<ǉ9��3篦�����w^���龼 ������ncrM���g�ٙ_o��{��h׶h������a���Clݫ�l��WE�s�[��ӓ���㖺�v��Iec���ӻr��$�������x�{������|���},�pc�e����y�:�R��R*]�LB��(>y]���^����U�{�y�T��k�=`Դյ-���x�o���ׇ����������^ qwS���ƚ����T�_��� �����n�U$�����;����tऒ'���נ{?fW�y��_M����խ�$����1�&�K%�뜦�0�sv�.�&��5��Y�+r�����~F���ƤW}�^٠qou�UUW�Wz��<��`˿���q49#��ݙ�I]��o�����:�k�ffbAΕ�RI��8$�I�}���\�����LM� ��o�����_�И�<i8%���$�UT�����z�� ~����򤪒o�� ?���|���Yn[r~o�p%J�W��������ݘ??>�x�"��!S�m��{=�����']���b.�8��V�y*��y�X7���� r�M��� ���ٟ�>AW}���dM�<���@⽯}� 徚]���}�٠r�+kV7��jI"q���W-z�{f��{^��t��jm0�9��I������x��L��ׁ�Ij����P	"Ȱ��`����҅.�J�_���Lo��c/͢4\MH��{� �T����9��urנsjK��Ʊ��Lq�1M�����z�砮�7UB�ӵ� ��ː�tG&24�'0RM��� ���@��@>�l�e�:&G�'�z��[%�wL`j�-�������	�ܟW}�w�hW�����P9Ls"Cc�= �t�����L`r�-�z�J�8BcǑ4�rhW��˗ޟs�ߵʯ~���Y�e	0 3&�
{�ww{��ϭ���n� � W:�ܽ�ȳ�d��u�Ur�ͣi�^�s2Q��lԹD�l\l]��U�%�!c$Tu˻��;tNe�]��;6��m��Ru�U�M�J�0q��.�l�Ӹ�n1)v������I]����담�O'H��$ͤ��$�r�a1��7D�F5��ϯ�K�,ˑ�X�ӻl��mӲ��8��粖m�����4�ﻻ����������O�y�#J7'$Q�&(�E.��S�˴ĝ�vet�^M�D�^uhnIn< ��f����w�
UK35�z9ڛh��a s�@�[ ��S��t���-U�#�Lx9#�w�hW��ݶh\��s�eRI��8	�I�S��t���[��]'�`^^�(�N���ǀ��0�K��|���� ��u�gzm�bl������ۡd��7jT��܃z.��n��j4P'�f}������	8���/��@9�٠q^���>@r��@���HqB'�q�;ݙ��U*��%IJ�%�K0������0�7^�U�J�l;�|��%�i�n�qɀm�� ~����$����������6��M�V�ێ<����}��L׿|����$���o��ﭼ����jQyWb��-���L`j�-�{��ξ��"I�cB90�ӒF���sd�4Z���Gntѹn5�j��X��w{��g�����SH� ��z�m�T��a��y��O3�$��\���`����UT�w�}0^���w�3Ԓ��xO�Q�v�w��o�9W��{�[N(�<A@�D���;w�@������pc�$�O��I+���< �������U%w��M���!�	�dX���;�4%J��o��o�0��^�UK_u�T�<��z5ع�"��B�0�&�u=��J��.�g���9*�Z�z�r~o����0��_ʩ/�w}0x����iա�� ?wvg��ٷ�����`���R�����w�[yݻ�&�r`����w�0�Uz��/�4�(�X�o�1�܏�%w��Lo����0-*�J�g�ag���gzy�RI��I�pRM��l�&09N��7�c���l���������%۪1�뵅G��F��s	Ր��c�%�<R�]K������]t����������9�ݿ/�}�� {_��8��]�rI���L�*����׀z��xo��?�}T��;������D�v��#� ߟ��o�ׇ��IU�y��}4�v�QȲcǑ5�G/�$�ϻ�AKN��VH*����R���>�%)N�{wZ�Y����f��)JR}{��y)@~P'>���┥'߳��y)J}�������[�������o��l� U-qVb�
9[��ep���&�
v�2l��c��h4�7iU�l�긝��'���{��3�jpq�(��������8wi��eL�.�> P�n�=,4qͮ���u�w���#�{�R,�Y@n'�T�<N�2k�@f��rZ�~�����[�$J+ei�t�2ƒ���$���lVn}z{ hM�n�r4/\�������w=�>��l`�jNݞ,��\��k��j]�����y�]�{��}�H;]�����?JR��o�R���>�%)O��w\�˒���w�%)Os���m��ˉ�nI�H*�R���j��$2S�������%)?~���<��.����JR�ϯ�w7��ս��fh��x<��>�{�qJR�����C�H�K����)JR{�?~��U#�tOB(�N�˻���R
�$#$�s��y)J_~���JR����C�R�T���߾yT����y��pc��n[�W�R;��ʤH)~>�t<��>�{�qJR��ﻡ�{��������0?��^���'��2F�*�[fΝ!1GM���㣳,Z�٬3Z���~�JR}~����R��=�u�)JOo����~���)Ew�����4Էjӹ�*�U.�7^���BEJ�s��M �	 $bI�	L�F��2���� I#�L���$��R���y��)~����JR����C�JS���o���Cm܏*�U �ý֫
�
^���S�@d����C�JS�����R
����#��v��q1��*�R��w|R�������R��=�u�(O͒}w��<��=��me�y�֌ެ٣Y��|R�������R��,�_~��)JR}w��<��/{�w�-�v�����߁�<��O��%kXe-���g��3ӹ�m�]�V��`�^�uf����ۛN����\��$j�H*��}�H*�'��wC�JR��w|���ԤR��j��AT�/��"�4�ܻ�=�\R������y)J^���R��_w�JR�g����JP���Ͽ�pM�;n[�W�R=���ʥJRy}��y �|!��µ�\\L!6p���"�Y� �i ��Fd��z�'��0V�p�N2�.�a�=�)�H�@А�.�S �I�����H����"f �v�H 6�v�$����PN�|lШ� akr�0&�v��G�$ �T�������P\^�R}P���қO��u x���01 ��r����qJR��w�ǒ���k��fk7of�kֳ3{���A�{w��%)N�߿k�R����v<��/{�w�)JU��N��Kj[�N�j��AT�|�|R���ﻱ�){߻�)_�J���o��aT����wuh�"�d���!h�pʽ�NY�՗�R�q^4-N��n��v;�M��*�UyP�������)����┥'����^J��v��<�AT���}m���ݦ�Z����R��>�u�)JO/��%)Os�)I��wc�JS�����[���\N���R
_��XU S��{�)O�$�����)���R_�u�rH�%Ȯ�	#U������\R���߻��)�}��P��F�'5'���
�H���=��;�.�G�H*�'�w�JR�g�)I��{��)�w���)?�k3?Y�F~�fNӮ�����T��n�t�H�b̙�tI^�����W.\c��n'v�n*�U �[{�k�R���w�JR��{�qJR����XU �_���ݎ\���[m�)JR{}��y)J{��u�)JO{�aT��v���}wT�V��;oėhѼ�a���<��>���)JR{�{��)�}��R���w�JR��]5�v;lM�v�ʤH)s��y)J}�w�┥'�������*�U ��wm�v�dWn(F�y)J}�w�┥�뿿h|��>���)JR{����R��6C�_������m� 6֖q�M`�N�ض��2��4�L�+����l��B�:Ĝ���v�Pn�D$�l'I÷!�f���4K\c�]��B{U��6e�ݢ� JZ"�����;��nx��[vQ.�C�8z�gE\���t�P��50��h�	r��nv.�sm���k�()Cr���ٌ�ɶ�n7z���9�l��NX��~{������?R���*l������TM��ӔW�q�b^�իil��5t��e��*��\��y)JN��hy)J{����)=���y)J}�w�┥��ڻ���j��{37�{އ�����xqJR�߾�ǒ����{�)JRy}��y'�UH�գ�Eiݹwq�U �AK���JR�g�?���>�|�aT��m���*�U U�_oX�6�٬�e���R��>�u�)JN���%)Os�	��O���%)Ou����.D�v��ۏ*�U ����O%(�?k���┥'���ǒ����{�'�J��(L���(J!(J��30JT�RH.��]ڒ)d�)�5��v6���ce�]o]!9�4ގ�v�����v����fn޷��(J��0J��(H��(J���(J��"��(J�~��^x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~�p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bw]��^x%	BR�	�%	BP��%	BP�$BP�%	Bf`�%	BP�����pJ��(O3�(J��J��(L���(J!(J��;���Z��vؚ�7�ʐ*@��
��(J��30J��(H��(J���(J��?w��pJ��(O3�US��>:PM�&BP�%	BP�%	��(J��(J��(N뿽מ	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	����8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	��߼<�J��(J��(J3�(J��(J��30JT�RH.����F]�n+�!-�IBP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bw]��^x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'���pJ��(O3�(J��(J@B��30J��(J��(J�߿xy��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP������%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BQH.?;=-��q:v���RH�(J��(J3�(J���B!�߿lA�4?~�������v �D�%	BP�%	�w��y��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP��n�����j��{37���8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	��߼<�J��(J��(J3�(J��(J��30J��(O���pJ��(O3�(J��(J��30J��(J��(J������(J��(J��(L���(J��(J���(J��?}�߳�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP���fg���i��]F�q;]\��XM�.��\��3uu�/Ԫ��0O(�N�˻�H��RH��(J��(J3�(J��(J��30J��(O�߿��(J��<���(J��(J���(J��(J��(N뿿k��(J��(J��30J��(J��(J3�(J����~�	BP�-	�`�%	BP�%	BP�&f	BP�%	BP�%	B}���<��(J��(J���(J��(J��(L���(J��v����N��nb�
�*@����J��(J��(J3�(J��(J��;����<��(J��(J���(J��(J��(L���(J����8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	��߼<�J��(J��(J3�(J��(J��30J��(O���pJ��(O3�(J�(J��(L���(J��(J�����ٙky��٬3Z�k[ߞ	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	��~����(J��(J��(J��(L���(J��(J��_�~מ	BP�%	BP�%	Bf`�%'"rE�>"��(H��(J��`�%	BP����8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP��߿o��(J��J��(L���(J!(J��30J��H#V�;oĖ4Էw�T�R!(J��(J��"��(J3�(J��J��(O����y��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	���ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	�w�����%	BP�	BP�%	��P�%	BD%	BR�&f	BP�%	��~���(J��0J��(H��(J���(J��"��(�
��Zy��v��47$n?ߕ T�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&}�߷�P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'�����(J��(J��"��(J3�(J��J��(O��ߵ�P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�& ��
P	@�{��~O��\pMطm�@T�Zι��5���A�P���"��u��VŠc7)��5��lݼ���(J��0J��(H��(J���(J��"��(J;�߷�P�%	BD%	BP��f)BP�%	�%	BP��%	BP�'�����(J��(J��"��(J3�(J��J��(O�~���P�%)BD%	BP�&f	BP�%	�%	BP��%	BP�'���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'��v�_��ִ[՛4j�o~x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~���G�(J��0J��(H��(J���(J��"��(J�߿xy��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	���ÂP�%Ȩ�d'��P�%	BD%	BP�&f	BP�%	�%	BP�������J��(H��(J���(J��"��(J3�(J��?_���v�:�2w��w�N�I�<���(J!(J��30J��(H��(J�����x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B~�p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	A�����JR��ߵ�*�U#��ЊA��˻�H��QI߾�ǒ�������)I�{���J�@�_��xqJR��gٝ5�֍kz��e���R������);�u�y)J{����);����R��~�??>�x�XԊ�V��6x�]7���i��2uF�wbf-\܆kY�k{┥'}�%)Os�)I߾���o%)K���|R��վN���j[���*©R������Lu)I����ǒ��������)I�{���?��0u)��~��sy�֬�Y���l┥'����JR��w�┥'}�%)O{��┤R�;��Gwn�"�qB[���A�eU��M�����)JRw�_��R����)B/�������%)O�����[m�2�i��ʤH)o5�%(�R~�����)?w��<��/��w�)JN��0��6��t�u��ŷ|er�$  W�[��n��{r�<�-@�ʫ�u+
k��ֵ���m�p�-�w�X�hܖ�gmt���#z��F��V��b1p#��jQ���m����(�����pW=����K�7�˨�����_[��jk8g��a���ڒ݇�u�4��s�*�R�@��[�=-��x.����g���� v5�]Z{{��%ŗ���5��h�q���{������k����] 6瞠��y��.�D��q�l�����tt�fo7�n�)N������)I߾�ǒ�������)I�{���JR����"�4�ܻ��*�U ����X/Ȳ)w��o�R�������R�swqeR�%J��v����m7]��[JR�{����)I�{���JS���8�)I߾�ǒ������f�ˁqKVݶ�ʤ^UUBVR�|�*�)��߸qJR��}ݏ%(?��T����}2�R^^�;o�4Էy�7�y)J{����);����R������);�u�y)Jw������Q���4�.9�����i��Oj�YGE2�1'g�0�ڷW�����q��3o�)JO���%)K���JR���]���3�JR������)I����r;�wmEvℷaT����ėPB\�����a�){��|R�-�v*©R�zt�m��ˉ�f��)JRw���R���{�)O�@d����JR�{����)C���6�2;�]ˑ�VH<*W�{�*�)I�����)}�{�)B~K$��?
��AT���?QF�ۅڗ$�)JN��v<��/��w�)JN��vJR���w�)JOE�/��;+�v��H���u����H�⁺f�+v��RM�l�����m��l	�璔������)I�{���JR�wfU �AK{݊��AT��^�wp��ټ�Y���R��w��<��/{��R��}�v<��/��w�)J+�����"i�n�K�U�R
�s{��)>���y!�	�<M���߷�)JO�}���R���۶k��fk,�Yf���J_�d��ly)J^����JR���]������w|R*�R�7m܎���Q]��-�XU �/>�w�)JO;�vJR��}��J�AK���XU �Z���"��D��N�c<l���i�i-ut��N�,a�%"nƤ��De�ӻreR
��n�������w|R���ﻴ�y)J�o�2�R\Zk=rH�%Ȯ�q�y)J{�}�qJR���ǒ�������)I�{���?9)|~蟂(�N�˻�q�R
��w�V�������?���ߵ�JR�f�U �@��z��"c�n�qV
R����┥'}�%)Os�w\R�����!"���!��@mI�}ݏ%)K���vG`ӊZ�]�2�R
[�z*��������)JO���%"���ʤH)i����[b����7E:q1l!Whl��5 $��Ká��3����p������\��*�U.^�^)JRwﻱ�)}�{�)JRw�z*©R�E���6[�Ƌ�n<�)JN��v<��/��w�)JN��vJR��~�C1JO��~ַ�ff�Z�fkf��<��.�����)I�{���JS�����);����P*�/N�qB�h���e�2�R
]���<��=���qJR��}ݏ%"���ʤH~Go��rEd�"���y)J{���┥'~��JR����┥'}�%)HX�B	=�8ʦ��@�G�S@QJK S	��N�)�e��bY�֓I�Fp�@`� �#�Ha2�L�
������F掰�0	1⯧�0@'E�&�9�3FF��݃� 1��&�����o{��{�� �   ����     	i�         h
��N��r�����+��!�m���B9�j�����㣵��j;]����b�u�gӮk[6�NEE��%�v�uu����M���W;Gi&�t�AR�<�-n�6�^�. :�m��=[��[$Rg�x�#A��;iW&�y^�2��[[�T� ,�q	-��a���D��EE�2�j�X�m��s�wF�P�	͞;l!�#�Z�[�*%�ՒAz��i��E�LR��!�/��V$���b�e�V܁�i<Y6�'�n{>kT�X�$=�u�լ�Iq��L��2L8�Ѷa��{���G��ю�*�tU���� S�бAɴp�T:X���s]<ٽ�$���8
ڔ�HtΨ�M��1�ޓ�� -6��L�,H6�� ��]R�m!�:�jF"A�+9��P5mJˤ�<�uӫ<<���V����]�*Rݲ��2�`��Ƥ
wk(�qr���u���'e��PA���v�����7ct쑘��GkBnjJ-ci띜�t�� �l�[XS����u�m⣲�>��n.{nW�6�z�z]��涐��݉c�a�5�`@�릂ېBV�t����lM[PmJ�&�*���z�R��T[eK�� CQ�<���R��Sʝ��k�.�dM���.c<�=i�u�t�'<�E��m�;Y'���n
&�[\ncgET�*�$����y�@��6��`�6�up���x.�A���7X)(f������H`-v�ʽ"&��.�EJ�j�\ml2T��5[K������F͹I����x��j�^�v���9�ٚ(��.����'Q��঑�<p�k��B�m-ѕWZ�P�S�+�9�J��HAdu[5<�,׍K�	��%�)']*��]'5U@Fv�'�����غ���=��Ƞ@����==���T�������w��?V���ݶ  *��	���o@��۲q2��:!'��#���Qң����u�$4]��C�AU�=K�Fbt@f�$�)<�*�Z���&ݝ�L��Ud�n�M�U�n+.�Ep=u]�9���q�u�t&
w��O�Ms&�[��%ITx�qJ����,W[�����nma"NS1�Ƒ.�j�A퉖r���Yţ�����wn�wz��~��qˎ�]�\�GE���i��ete�7	uٺZM��W�qK6�uN�7�Y��Y�ַ��)=���y)J_{��R����쟒�R��?w���U U��Y"c�o�ۙU��AT������)I�{���JS�����);����O�R�����̵��ټ3Vf��)JR~���C�JS�����);����R������)>;���XD�R��.AVH*�/{�*�)I߾�ג�������)I�{����AT��i����챢�ۏ*�)I߾�ג�������)I�{���JS�����){����+{٘k{��U�pZ��0X-�f����ˮ��ۊ��Թ�]���]p7Z��{ݷ��������)I�{���JS�����"�U�H){wҫ
�K���ⅶ��5�5��JR���]���(�SHi
SY߻�)JRw߻��(w��*�U U���nI$��܀�R��;�u�)JN��v���/��w�)JN��vJR���F�[6oF�5���5�qJR��}ݯ%)K�{��JR���]�����߻�)JB��]�r����̪�U �F����);�u�y)J{���┥+{ݕXU �G4�궭�eݗ%��b���ݓ���j�l��HLQ�+���x�̵֩h�kf��Y����)I�{���JS�����);����(%�)o}�H*�R��;�oŨ�j[���'����߻��VrR��{�k�JR�߿o�R�����<��>�;��dl�e��<�AT����*��AI}�{�)Nȁ�	�;���yU �\�AT��8�]����dWof�涼��/��w�)JN��vJR��~	�E,��{�k�JU��(]��2�i�I�H*�R�k�<��>���┥'~��^JR�wveR
����n��2�tXԷ\D�kɯNn�$ֺ;bS��N��,�ʯ#��	���ղ\�&Ir+��XU �]��yT�JN��v���/���R�����VH*��Ή�"�D��E�n<�AII߾�ב�C%.���|R�����~�������\R���k;��Z�kyY���k|_%)K��~��);�u�y!�)������)I�����(n��qKV�rL�AU�IP��~���C�JS����qJR��}ݯ%(8�� �τ3�|FT�s}�┥'��j�f���fn��JR�g{�qJR��}ݯ%)K���┥'}�%)K�~�f8[�����Bzp�z��a�DN�,�H���t����H���:%�n`iA��bZ������ߟ��伔�/���R�����<��>��yT��.qn���۶�E��-�y)J_w�� ����'�k�<��@�N��ߵ�)JO���%"�r��.�Wq4�$ʤH)o��a�)�w���);����R���ݙT�������rH�%Ȯ���y)J}��u�)JN��v���>���┥'}�%)K�ߣ]��7�Y��f��޸�)I߾�ג��T�~��)JR~���C�JS��{�)JRB� ?{w�ֵ��{���c� 6��L�.v;f�mu�/3S��n5�Ӌh	�Y:v�s����#��&$��۪�u7#xK���S����i3�j�i����h�y3�bWd�ʲӍ��gqG�I�
<ݲ�Z�9��B����	̚l��Z�y�s�U���N�W�*�N���k�ZN�]������+;�&C��Xg��������J��H)�������Ӗ%��:m]v�ƌ�̨�j��4vj�=MV 7c�o�neW�R�{ٕH*�Q�{���JS��{����)I������AT�{�yhi�-[�ʤH���]�������\R����wk�JS���⟑�R��j�f�ٺ�F�Y��{����s���┥'~��^HB����b=����c�5�2,-f���~X?I�����)�߿s�R�����<��>���┥'���z�fk4ke�ٻy��%)O���R�~���~��JS����qJR��}ݮH*�8�^��6���9ι�\[��Kv���D��u�0�4�VT�X�Vlӛ���)I�{���JS��{�)JRwﻱ��JR����8�)C��\�&Ir+�aT��m�u�"�ꁚ\q�JN���y)J]����);�u�y'��K�	�Ewn"�U �AK�{�O%)K�w�┥'}�%)N�w^U �@����T�m�X]��neW�J�L�����)JR~���C�JS��{�)JRwﻵ�)w���44▭�I2�R
[�z*©�ϻ�qJR��}ݯ%)K�w��T�������=wi���q�m�El�l:C�ac�[<vX���X�͇i��9H�ma÷Q4Էw�U��AT�{�<�ATRwﻵ�)w��|R����a�T��ov�䱦�E��*�U"N��v��� Hd����o�R�����VH*��w^U/R��AK�^���k5�ff�n�kk�JR��߷�)JN��vHz"�T$N�7)��{�)JRw߻��)�v������\M7�T��-�aT�N��)I߾�ג��߻��PU U��Y�$��\��FGXU S��{�)JRwﻵ�)w��|R����a�)�zo35��.�Z�YX��m��V[�����j6��^v%J�M��TQA��(ӻq��R
[��k�JR�����)I�{���JU��וH*�*���z�Clr�����_%)K�~� E�);�u�y)Jw>�u�)JN��v���.��t�h�ټ3V���R�����<��;�w�┥'~��^JR�~�w�)PR��n]�i�n�XU �[w�┥'~��^JR�~�w�(N(�"���Rw���R��v�X��!��*�U ���ʮJP�N~���┥'�k�<�����וH*�R�wn7v]�"m�J�-e�WG[5�ݨg�I��Kqz�v��QjW:H�w��m8�qB[�XU �F�ve%)I�{���JS��{�)JRw��©R���c!vڸˉ��*�R���]����s��\R����wk�JR�����)C��ڻ���j����FGXU �[}�yT��-�v/%)K�w�┥'}�%)KW4OB(�N��\v�ʤH)o{��JR�~�w�)JN��vJP~EI^{�<�AT�W=z��D6�,.���[��)J_�����)I�{���JS��{�)JRwﻵ�)�>�y�zw�{ӽ��t��[Fv�� 6�ݧ8�}*K=$����Z�p.���zVyG�@��RG6�61u;��ȓ�� ���v�=nd�x���&��z���D�eB��9�Y�㑛4g$u�k`��c$�;.Y�����9�v�I�v^�)Q����঺�:�u�����B�Ͳ*ګ6ӝ�؎Ī��mg`�Ժ<�d7���y`"#0?�{���v�{�诰9�l۲�����@x�nkrl���sx+��v��u&�wlѮ�A�f��Z���T�);���<��;�w�┥'~��^JR�~�w�(K�o�km�0x�&�R]�����{l�>�S@��Ԟ�<a�6�yl�1��2�K`n�V��&<s�B'3@/m���hvנw���8��u($�(�1�yy�	� ������0	�c���~����S<��� �y�Du��Zgr筊I�\���3�(ˢk�#bk30`E�[wd�1�6d�h��R4������8��)Kir�U+ sL{٦��׀T��G�lqO�=��_zh�Q�Ilِ`t�(�Aun�TYy��ِ`E�[vd�1�8n�m�[���;��6������}�> �����YMݵkh�$�B�9��6��U�m�^����˓IHצ��N�'�1D��x�50m�����ƀ^�4r�{�W�z{��Z�I��`��R{l�9�)�U�_�?~ϐw��4�_��m��<n94{���]ϻ�r�q��|�0�+"Q9$�G_tx��b$�i}5�/������6AB�6b��o�'�Ԛ=5��R@�{��!ѱ>�GX�D&�\҄���A#,U`8&3k��C�
6&��<7��	%�#���	�&�`��<VbC���v�����UH��YDC�l_U4�@��s���W�}������6�L��\��T��}�w��0�٠s�S@.s(�L��I�i�`ñ �&07fA�IlF��v�ۆ�m-k��ۡL$i*���,'BI���M�!�<۵�+�}��yg`ܭ�@?�cvd�D�ݙWQpQ!���h����߿f$z�yh留 ��h�\�ۉD<yQ��ڴr�h�@�,��y��=���j`ۑŠs�SB��{�U��nWD�Ή������4���Эk&<s䂐�	�cvd�D�ݙ�r]���z�<��ɚb�=�,��+�`�WFֺ�N���Ug��):��NӋ���m�2	�"`ñ �&0BY)G&27�j8h�ՠs�S@/m�9e7�� �C��L��I�1A��߳��'I�ِ`E�_＀�ճ�&�q�'�)�|�����@�����RW��<`~�y�4��e�f0�1�:GLِ`��W�m��uC�Ю�fw{ޕˀH  Z��m��E�u�uRp]U�l��Ҋ�k9�6���f�	����-΍F�)��[5#��u��pm�;r�Z3�M���:Ϧ�a�gk���۵�m��i��'�K�Zܯ^Cp��W���V�:�-�5�h�ٞ�d���wiܴ�5<����̹X����Zh��TJCr�ݠe�Vq��L�5����������W�ҳ�n�z6Ui�dl��Ԁ�Bvg�A�L�>�F�FۉD<yNG'@���h���g�f|��}�{��=���5��+�`ñ �&0�1�:GZ9B���Ŏ`��R{l�sva�]�*����ߗ�;�O/�kdJ$��1Lm�&�s��������{l���.(��F�IȤ��07fA�N�����������7Wnf��	�^s[7	[f��#�aK6�ș#�����+)��2t��7d���W�~��:`��'��av�-��=���H@)��(9 ��l@�T�����s����遻2R��C�29$�r٠^۹�s�S@/m��n����M9�߿~�^��٠w��4�٠�@��I�m,x��I������{l�r٠^۹�yڒ���n~jnv7�\t=��Z�3C�Z���N���F��Nt$kI��9 �4�٠�@��s@�,���ڲȔI��b�ێM ݓ�t�ݙ:L`���LdnD�"�h��h��p���I���0��� ��B)�����s�S@/m��[4�w4�u+�x�`���> ��� ���z~��b�9͚`4���Xs�����:���k���ʆ�7AqDìR�Z�e�ŵ��g��vsU��w~��	�:`ñ �&0%I��b"<���rh��h���f�s���'���BF�n'3@ݙ:L`�ct���%�m&,s䂐��f�s�����+���Pȃ0dL�]�@��Hs���r������(�k�1���[4�w4r�h�@�_J�Ll�I�0jF�pܝg���FB�-dn"�v�5\��\��q�pe�M1��!�@��s@�,��^�4��h�Q�ɒS&()3@�̃ �&0�1�:GO�}���~��+`�n�!�{� s�p�ŀ}�e4�B���29$�l���#���0	�cT�+S��@�rh��h���f�s�� �WUT�b�UI��m��&�E b�����r0��\bWg�Ruo8�2����/IkJ'N��3��������v+��N)v٩�PxC�˻vl���e�(��ݍ�bL�4kiv���i�``3f�ڵ�G]�ug�l8���cN��VVnx�vn�ۊ�a�J����9�Լ���5(��@�A5ب]"��r�a�g'd$� z�Ӂ�^G�w{�0:���e�PJ2�Ƿf��l#�Z�qv*�zn���sv��:\��������^�h�@9�f�{n��P�kbic�'$��^����#���05tU3�&�FF6�@9�f�y۹�s�S@/{f�}Jˊ91��s"�hUU%~��� �}<`��0�ݘ�:��ɒS&)#�@�,��^�� �7f�{��yUR��Sͷm]�48�n.��Cq�+��Ւ�΋�,�&]W��Ñ��M�8���v�.f ���`�K`M�vd��a�]k{��k[��W��{�GIB	 DdRA!N�:��w�ʾ�e4��h��1@x�&��Ǡ^;V��YM?�f$z�M����/3��lM����8�r�h�l�5l�þ����N̉��Zwb���y�,��N�[%�&܉��3LԒU�ܿ6����@�!q�ꧬ��C;q1d���i�y�b\�N\�I$�(�Ǎ�'�uw�z�h��|�����g�G&27�iH�	�"`ñ ���K`NT�������Šs�S@/{f���_?؍�T7	H'�]�:���>��h/X\s��O�S0�$�+�������ݼ�٦����iBcC�X1�&���^��w��>�����@��,Lx�Q��]Rr�F�X1\A�Ů�]�b��j��Kv;F$�1�&,���M)�@��s@�,��^������;^��47$��l�=T���۾�o���7���ԕR�;���e���-���"����5l���#���0<�Eq�$�)�1`ۏ@��@�s@�;�ܫ�@N � M=@�К��?~� ;���(��F��)��n�͙)%�5l���wbJբ]
����J��6��0�[�%��xQ�m:�*^�$b$Ǔ&H<mL��Nf��YM��� ��u��%��}�b��Xy8���v�����?��^}��o���;m��9�)����#�uy4�1��,� ���xww*IU�{�� ����KӢǏDґ8��w4sw��ׁ�+�����[��� �Cm�3@�-��:��@��@���U������$�u-���ȚM���X�:O�x������-A� 3H�G@�!����I���#$3&Ll��Z<��C(N� b���!���H�֊��B��83߁�5���ۢ�㠆x�(���I��<8"C�_}@�����#�5��E���-h
7 <��Ou�����{�����������$  �   ��E�     �           rJ�[!R��J���Gf� �*�(\acn�Y���T���v����,j��kvͤb*�!5@WTQ Q��gkfmـ��R��î�5=&�t�1
�v$ ȧ0khݢ.mu�Gm�;n8\��JŎƦ��.(ې�h#3GIk6�g���� PA7V�+S�Mo-'�l��rK�[�Rf��k)�4q��+f��7�ϥAՄ\��������pYEv`���e
�;R]���luc��|�]���2s��j�� �&[��ڍ�B�Z�n:�QÍ�[v�l��s��:hC\��iv��P ڨ���*���.҂�D�]U���n-�g:�j�	ydvn�(�Z�#i��4��5H4êl�^�8[�!Jqm:��f|�%ڑ͠��=W�L����]�Ur�f�I��c=�S]����_5�ݛL��ƆYx"�`�U�ڡ�ts��j��Bc٣/�֪rfN	YU���.����WF�5=U���X��..v����+tk<lfw����X(���@l��7�+������yF6n���˭���SX�!�YU9���j�'$l�A���P@n�+;,���P6���k�m�KԱ�����̢�O-sHR�ݸ:�!y��}�b�O��N��NSe��)X��j�|�u��70���+��jΐ��&��5\���h6M�v�PB��O�۶זF��k"�u
IG͢�C�b�]@ ۣ`�d�B��:�x4�)�� ��U)@�K٭+�d25�� �:�`�j\�,�`2u�[K��S0&V��uP&�Xwi%�u�&ո������i����p밹�7-V1�IJ��@@r��#�%��e �g�B��Y����e��i�N�;[֭Ff�k[ټ���P]!�'��Eڞ�`|���)�� �~AN+�.(���Ϫ �'�]��mh ���Ky!��m���p�)An���^�v9�q�����VRNv�k����S�����;c�v�%�q�AV�g���/8�mYF�+cM���n���ř�ɵ�]ZɘN'�*έ�.ځaq���Aew]h�I�i�X���F)K�N�F؆�u˔^lLd\WVaes�fv֎�=�`(�Y,c�[f���{�_|JlEv;��9�k
�1�Mfy�P�N�M98�s��$���줠㛰Ն�ͷ�rנ�@�v�g�;�{s@��y5���1�,q�9l�;]�@�,����[�߱ ���{rc#p�Ƥ���׀s��������޼ �}��V<�2A�jd�$qh��;^��9�0%UU/���=����yH��.��3�m��x�J���z~|���9͚`T������ӐD��6�Օ:#u�O<�]k��ܧ7�r5�z� �wo���֭M(Lhr�q����v�V��l��U��o���=�зoŰi�n��r`׻yڪK�I% ���m�u�9l�;mI�`�#Cm��͙)%��1���L�ӻI��rAHhVנ�@�v�����-MU��1�,q�9�0RJ��޿�w��0��W��]bGS�����NH�l7=j#�űI;I����k�l����k�-��RM�ڴr����������_{&H�ڙ1H����s@궽 �-�m����$��O���~o���ovaĥ%T*E+�U�]������X����7��m��&��Z�;r�>J�+��}0��� �7qh�ՠZX&�I�Ǒ4�NM�GL�09I-�nɌز������"f�v
��U#�/F�s!̓�i3�4;,�z*�i:�9�۶;�'��#���lvL`{�A��Zwj�l���q`��^z�%v�0_O9n�VR��4�)�1`ۖ�7d��d�:`j��=ˊI1�88�jI�}�)�s��h^��w\�^��H�&��9��·G�&H�ڙ19�9n���נ:c�#��z%@���2��R5�ܗ^�95��Miƭڶ�I�It�[�6���	�`�BI��&� ���z�ٌt���:`vܸ�,2���
�����ݙ�Wg7�ŀo}�X/�מ������v������ ��ذ�05wK`:c��[�
U�V;MȰ�w��u�7�0=IR\���x�f��"NH'3@��e��1��l����R����ˀ�  u�^Me�t��N�P�A�m��䛳r)�[�ej]U�a�lg�5J�^�K�A�v��᱂4�;�mi�a��\��X�Ztv�@An]�ã�9���=@�.u��ij���w���Xv�:�y�hNg[]Wga\�ni�Ӹ��FhS@9�n�E0�r�K���Vn��ڒ0�s�\Gc�[����C�h`�k����=_|t�ӗl�<jㆺ�����
�z㊯1t�ݪ�ۊ�
���)�l$M7�c�X6�����>��;�w4.�� ����c$y,���`{�t���Wt���?��UU�o��הR;���G���L]��Θ��H�t�	Y�$��	�
Mπ��@9{f��n��[��^���R!��,h�@9�ـwwq`��,��� ��W|z�/��˜�<�<��pd�:y몱r.�Ԁ�iݩ�n��3�Fƞ���Z~}�b�;��Xow_�~�;���7�����Z�Q��qŀw���R�\E	䑂`E
�B���:��٠v۹�w��S5�4�q�q`��x���<��w��ŀo}���)וF�x�#����h�0;dt��[ �%���2�̻3Y�������#�����٠quUR��3#y rH��0��	E�0�=�kf�+vn�I�IzH�����Rk����Y�����IlgL`wv�hoX\y!"$HO�Rn|���7d�wGL�0$�2��b.��Z�ǀ���;��,-ZIҪ��|�/�H
8�o>���(����-k�Nb`�D�q94���vGL)%��1��Ev�,��6�Rf��[��|��@9�f����h^v��,$�JC���\X{v&lsG>���mK��㊺]��z��*,į/�0<���7d�wGL廚S�*�&�FF<q�/n9IL��GL��?}�$��R�&2F��rh�nh廚�����hs�\�#Cjd�&h��,����ov`wREURI$�g�����[�f�}��q��2D���#������6t�wGL�0���8�������.&�q<��tdfU^��Af8��UvNe��(��ɲ����L����;��_U%_�9~����G�q9��yN)&����h厘RK`:c����
U�VZ.�e0;dt��[ ���0;̦T�lM&D�q9��������?c���l���pX%j�Y�]w��6t�l�0;dt��;^�UJ�UU*�6��Im�$�$� �h��1m�䖲��4�,KhZ�F��t`í��z�o)���	*u�����xm"Fm;�oH���(Z53��J^��R���t��#їI�ۯL���g�Ӣƣ�KK�諡�O*��*t����K��.q���T�ZC�{$��÷]R.�ك��m��"��n��2[��5�k�ãTv�G7����NoY���5�Vx��3ώ��T��S��Ѱb/Z囶.Q�L����"y1����x�;�q`�K���o� j���(�v;YX�K2��:`yI-�l���Y�J��o�����2K���ɋ�����7�0����wذｋ ���P���4Ǡ��@�{w4����mz�>㸤�����������#����Θ�=$Ә¥��q���۵�[�{���.��T��wi9�յ��F�u��+�`���IlgL`wtt���ce��K�n8�׻���J�T����Ēt��ـ~�w�n��*�:��~kdmn= ﯦ����h廚���>�e��	ɎH���g�m�٠^�ۚ�����hr�Ǘ&H�ڙ�4�������ov`�w�[�y��N�����pݢn��q�����\�9�w�9]tt�F�3I=�H�ж]��}߹'������1�����GL	�&fZ�(���U���`:c���l��+k�/0q�N	��qI4���*����,~<Ay{�4��v+(�m��.> V&���8�)�H�L�b`,)s5�Vq0<�a�3!R����"L���Ä�J��p=֏(""	!u��H�B!Z� �X!�"� ��)�BVX&Y �`�K#����U�)-���d�!4���
Y���Adj�B�� ؀z�&�<=8��\��@M�C��
b|x��
?=LD} p �
x�����/ ;��ϩU]��z�Ȯ�B(�m˒��~t��� ���0;~�L���dI���}]�@9{f�����#��b�t*Aw�°��([n�z�;T����E�#�8)C<k^c4̪7�spPI�Q��	����h�n��[��}]�@3�V\�I���㗘��l��/�`:c �1�ɒ46�DE���s@�v� ��f����R��]��Y�$D�9��.L_���I_�}��}��7�� ����T�����sf��p���E���6t�Ύ��:`v܋����~Û�����g/\y�aУF�u��Ɇz��� ��v�v���a��-^,�`l���#�mȘΘ���ݼ�ըE��r,��Ş��J�޿z���L��ŞUJ���x��[I�'Nf�z��r�S@���yn�՝+ʠ�X�#h��; ��#�l�����+ЖL�I�����4��h廚\�x9�Lu��*�Q
����Ͷ�8 kw]v-v�8���q��Y]�1狰ܨd���1v�"���=v�g���"듳u�ٸ%FƓ86�-�v��*�r�ـY!�����ͥ�N7g�]����+,/)Y�*�^h5R��S�6d������&��m�(֮΋��ٳ��I�ۢ�\�
�5ԩ5bc!S�9-� ��y{d8�z��tsvjw]��w��L��ێ�p�	$�.��a�8#7-ۖ��ۜ��髫�]�!"G��d�S"$:���4
�k�9�)�^�S@9zʉ0�c���%&��yw�z�[4�w4r���Ydn8� ��R= �-�I07dt��$���J�V�v�r`|�%W���,���`��x�[4��=��,����jL�9�09I-�nɌ�:`oH��A�{������k� Mf[�	ɵ�D���l�WW7Z���$t�w�o���� 9�ـo{4�UJ�Xw��,mx����j27`�G���ͪ��J�^���9��0"�-�i��ee�2<���M���yn��ؗ|w��@.^����S"$4�06_D�6t�l�0�j"@�d��������- ��Y�w�S@�-������,�1��LcF����ҏ&/]v�\����;M�h�2r�#m��ƚN- �zh��;�w4Wڴ��wȘ<��#3� ���e�Lv����Xg�h�E��0'_D�8|��}�˾n�|��}�ܫ�^�1kI�ȓ�'3@�}�@9�Y�^YM��s@��.���ő��o ݄�l�0;dt��}V���-�����j��sWC�NK���s֣Xl�.�b�-�g��!mZu�WZ��qa���l��l��7a1�}��<�2F��ȆI��s@��� �)f��n�w���I�F�����6��< �4ه�Uw���`�{s@�9c��<r#�r�$t���}UU^��$��=��wȘ<��#$�;m��;�w4�k�r�h�k��A5���
,�8mG`mS���!��f�ur7;���u�k�{=RF��hn5&h廚U��9K4�w4��
�֓K�7)��Ilv� ����Atu$�,��x5#�r�h����W{�{����4�E�BF�+ņcwd�:`E�[ ݄� ��X�̑���"$4����y���;����L�]RUH������=�����Ow�������8 mm��lK�ON�'Y�-��+@���nh��l1R!�[o��%zl����� ����H5U�Г�]�󹽵�r�@ύr�.�e��Z�Q;t6��QY�:�����on���'���y5�O/=v1�t�R�uS�ϳv�jkZw\�۴��T�Mc����fۙ�c�2��Я@e[��C{L$��2�ܝ�{������8�Ā^];\ۭy�Ji)duQ	fzd���$,6����|f�H����˹1h���� �*��_{���ݞ=UI~���ذ����A�!i�\� 9�6g�UU���� ��ذ�n��J��S��U�-�R;r2L{��0"�-�n�cq*<��Xg�h�E��0"�-�n�M��M��B���ю
G��uoK`������GL�}U�ټ�f�5p�����C���L�4m�t��OX����ы�bx�Ӟ�O�m��L`v���#�����	fU�"d�En\$�9��,�>!.�~I%��`j�-�n�c �9U��̴]���A�����ˤ��	�w�s@;��C�QG��Rn|���s��~I.u�ũ/�����ϾI#=��� ��,h�ԒK���|�\뮓I%�'��I-��ƒK�W������ue�.�6�p#tS���l�u���{4dI!�8w�tN�}�&�g�u~�bK��t�I.�=^�Im�v{�]���m���rllC�L��bԒ\�w7RK׼�i$��&{�%�q�i$�k%o�'3�K��Y�$�9K>�>SH���B��x����]ũ$��g�$�t�شI�YƳ,i$��&{�%�q�i$�d�{�%����$�R�b�Ld�&'$��޸�4�_����~����]?6$�݇��� �?ÝӖ��K[k�������Tu��:�N��,lK֮�q\�[���ͪ��A���I.�=^�IoF���[���K�wqjI%�V��D�c��%��u$�~lI%�	��Io\t�I.�g�$���#jx�4(�jI%�	��Io\t�I.�=^�IoF�����B��&$i��>�$��w�����$��F��Ͼ�꪿����SO��}�I[rklC�L����$�yo��$�L�$�݄�y$�H��I%S? �;WI[Bm�{ .#]���0�s'>��a��J��z8�j:��5��y��w��]#`�I-�L��K�����諾v����ϾI.����&�FF0���[���$�)[I%�'��I.��i$�R�d��$Ln(I��%�n�i$�d�{�%�6$�݄�y$���<�$hmdȂG1�I.�߳�J�J�I$�a3�I(�:��Iv�D��K1�$'�)79Ē���jI%�RϾI*��s33>������Ξ��X�?	�~'&,̠��f���T����s1��&�>����ﯸ����C^h�A���af�F	�gn��߾��O]H�=}XR����xc��:M��ӨdqD1_���4��������Q|�b�_�*�����&6��.R!�   ���"��x�A�x�{�w��?>�     [\mZL     X`         @ ��ͮ�l�b�%t��y�Zn���0F�j�dݜmv�=eݗ��c��,��T];g!g�I꺷�L�����8D�i��Y2k�^�=�ut��n�T�\�����M�4�Y1.JmU�S��3���{Ll��T&�u�C�kcEU��X�L�$�'�M���qڗ-�mā�*ڴ�v���-�P�v�)��i�x�M�1�ӑl튰�x3�q���7Z���2�l�±�x�!��9�NQ��]ͻuP���m������>�5�g0x㚰`�񸝳�X;Y�F�6X*�2��[rZ;m�Ѡ��dqq��U+���n��[C$"�s���q��IJݳ�4��k����l�T���0@E�U��ZPb��.VP90\��U*�W[l�9�p��H4S�i!�4�G����`�u5غGhU�i
vZ��ܻ�ZwXu����+��W�6�]X-��nv�;
�*0�����E���Etq��j�j�j#����PU�S��+-�X�9s� f#m��1Vٰ�д��m+[m��܁��� :
C��b��Wa7���[�U�<�;%�6x��/V����+J1R�+�	�UD�(d
��)vC4�f�`$�U�|$��z���U��e0�z�V2l���Ok�C�zV�\e��A�S�#s_Gn2�L��IFEkuDt4�mq�t(ngM��:�u,���Ɂ�n��5%*,*Vɰ�v`-+��7F��q Fc%�늩nVz�d�s�m�pWP 6��nf�H(�<�Kr�ϔ�W`X�N�	&N����g9�ra���-������(�ՙ��ű3�ڛH���6i�f�T%�!n��H
���t�*�ZR�!´�ʖ.�ݱ�H���@#�
A�i'-Y1��v<��Æ�Q�̎ÖV���V�,��(
�f�ݫ5n� ����E=�
�� "�CI���~N�!�H~ >�S�\���+� �� i���ȝYG�y��F����*K��Kx�� ļ2QX�\�/�دM�q�u	ιֶ͌���wj�L3����Κ��A=p�θ�lJ���C��Jv�+s����Jg7�n�p�W!��x��!d� �IE9�4{�բ�wil����b�[�c%H-<tv�Ql�6t��IA����L9���!Y�b���������.]������K��\�Ԗ{]T�m���*��DF��A�+��5JZ�5��4� ���o�{�%GV�Iv����JvdI����.�q�&$i��>�$���z�K����䒽���$�9K>��3?cmv�&��<���ڑ9�RI^��g�$��-I$�a3�I(�:��K����YuxR��W��$��ȓI$�a3�I(�:��K������V�ԓH##H�5$�݄�y$��4�]�z��������_�~/mČk��Z��̽�uF�!nV���Wd&�%���훞�ؑ�Gv��ʻņg��F�CI.�=^�IodhԒK���|�Ig:c�2F��L&H����������:�ߑ~U<�4�	� �:�����g���2�ffg��]�|�G;)7��3����I^���!�q!_�n�����$�݄�y$��jI.�߳�K���n�F� ��0I�䗮���=�:g�I.�=^�Iod�jI+��w
ƈ��F����H�d1����� ���n�c{�$��θd��i���[�vح�nu�d����T�M�G��kqts+�ֺL�5�۶GLwd�&~����d��	ɞ=i�ӂ�����g�ý����@�-��f~H����ԓH##rC ;����ه��J�$�ｹ�s�x���o <��P��=�1��#���v�z&�)�ڈ�K�`��, UJ�����n�c ���u\����T��95�����..��z���j�G]��E����d�$��	�	�π�l��L`ޘ����}����2�����+���L`v�t��v�h���V$F��4�d��-�ގ��0l&0=���,�5��nL�U�wߖ��`�i��g���� �s����*��]UB61�$�s4s�s@>�,�l�����Ӣwt*AuyXV��ܴ��qk�y�E�vd�
F��טj����Q$�,��l�f�}�Y�s�h�n��;)���o&&7$���7ؑ{}��s�x��K4
����#�6�$NM����=��`�L`ޘ�;e�V`ff���x韆������4�;�Ƥ�<sK���K4�;� ;���?s�L�IUB_;�����m�( �q�Ft7/<1�\�T����5��4'ey5� �o�j�].56gA�H����[ڝ�m�>lJz��s���9�*�ƥ3�ʠ�OX{L�h���n���9ͳ���f�Her���׋N�5nxXz�����Jptݮ�m�y���7�P��Z��o���r�aN2\F��d�r��ϻ�7��q�ѵz0�[������Q�c��q[a�b��j����Wk��7����L�#N����?c ��	�0l&0$:S˰c����jI��l�>�e4�R� �����bE�?/((�"NG��ޙ�`�L`ޘ�;zc�����&�FF6I ���@>�l���0=J��W��x��2'L�E�U�,3��0����t�>�,�9��$6�Ƣ72LQ̗Fݰ�l�ЗC�X��c���O8��$�Uː޺�=]G�mL&H������v�hݥ��;f�w���I	?�Ԧπޟ�:*�}��{	���oL`���I�x���@>�,���0��ٽ�L �w� �Ӿ���[�j�,�`ޘ�;zc �������͍�F��RM �;f��ԩ+�w��;�� ?s�0�v�W$�=�Z�i�Z���ӝ1�f�Y(��]zn�%���",YG�0��m�ޘ�=���=�1������W�W���m-I� �m5� �|zh��ގ�ގ�ZH��Yuf]YV��L �����0%��!*I!!x��0�M��#h`�Q���ŀޛ0��ѭ�F�n�2��0ޘ���t�=����}�[���kȐ$��#�MJl�v�q�{a1�{zc ���A%�fRr��6�ēT�Β3	7<���7 �b�#8�oXqi� c�&4��a�bnf�}�Y��ݘ�wgԪ�Xs��X���~M0y#RFG�s�o���s�ۚ˔�@�9ܕ�mymI4��0=�0<����0;j�	qۻi��[�Ԫ�����r����W����P�!
©*EUZ�[T�/���=��=�>w�laYv�e�0<����0ޘ���q`*�-�뻃Q@��BH�+c�.��l��]6t���,�6j�y���S��5f5�2<Lr(G�;}4������>\�zY���̑�S"$NM ��oGL�	���mKE�I	?�M�>����S�h��yl��{cp��0ı7)�l:c ���6La�_U}�R[���=%�h���mM ���@�J�����w}0�wf����YT��o~Y��~m�[@� ��뮊������i9֜Z�D�
�U�ɝ�e���Gmp��e�{/\p�6*�h,���ZŻC���*(A��<a�ݛ3�rV�d�g�m��m\��V�7��Ag�j�)�g]Wd�yv���e�u�6,�k��מ�,,s��N�˻�k�n.E6*uE��jG6�m�Hqt�s��l�;��*�F�3ب;���{��_~�҉+��kZ-�X��l�;[wG]�שc*JF�ZJ�n3��̻)���T�P{��h���v���v�h�2������INM ���@9N�`ޘ�&Ɍ�!wi�H0ŗi]�c ڝ1�{zc ���0>\)rcQ�#����rM ���@;�c ����:c*�*�ef]"�ee,˼��&0oL`S�0oY�<��bǃ����bn����*�wnpڬ����Rc�oO6�����k�j�"G�M6l���gy٠s� s��hs���ӄ9�PrM �^ټ�����RRs}0�}��ݙ�%vz�,K�<�<���I4����[4�v� �^٠}��J�F�wk3l��=�1�mN����}Io_M�)��<b�������4U�{}? s������wn睌�Duۅ��v5���Sy��V�T.�W��ԯ;'�B�c5MG3@9��h�n� �7g�UU~�;���9}<yD�<dx<�َI�s�hyl�>�n�s/l�*�tǖd�ڙ1Hܚ����W�����A;��Bi� [h}�a�����V��5��8h8�I8�Y����[�,HI �C �H���If$f$G0���	��0eV ���Nsg0�R�0�n'�(��y��}ޫ�@#*��ڎ���l2,0ʁ$#� y���&*�˚���h%N� =H�("u@��s���S�Q<�=AW��{�wi��>	��ߎ~��f~��{�h�1�$"�$��6|�}� 8��0��f�T�]�}��3�p��0Ę�� �^٠^��;d�oGLЊ]Zʻ���-s�Гo[B�
��W��i�K4p�(��6ȱ�

by<O"i�RM ��� �7f�wqz�$��`u{}0/j�i��F��RM �-�y۹���4��4�:�x��8'#�ɠv�t�6�L`�1�vɌ�!v֤�j6�nf�s/l��l�|��߿o���4!�&sBi]�����$]�y��*�~��&6c�h׶hyl�;��� �^٠s�uT�7��6I�rG@n[3Δ��#�=u�Km	Вl��Ư!�uܲ���L��R��4��h�n�s/l���ϐ����3Ȑ�L�4L2d��}�>UT��ë����`yl��tec��0Ę�� �N��=:c ��0%u��������i�0<�]����z`�n�s/l�>�ܕ�c<�����L`v�t�6�L`�1��������w����V������  ���KK-�mŝE������uJ���#Iux��aEsnM4�@�V�'�ODW[f�ӷ.�;ve�I��2��1UU�� +��-<�r�t�e��s�� �H-+Pc�F�z��Su��4�$p�]�Nn�c���q�������nu�tl:�\��sQ�	����1��j8����ӄ�\M�����{ۻ����ww��~���v���ʛ�vLF�c�.	��>d�ֺ�ge���oG-E�v�Zy�
H�r|���ۚ̽�@>��@;�f��t�mjLa�jF�h2�� ��ـ���;��,����������1����cf9&�s��@;�f��v�h2�� ϩ�,���F�"���&07z:`S�0l��;���I����͟��nh2�� ��� �-�+IT�b���5�\�hrth8盖�����V�*%��:����ǒ'�a�1�� w=}4�I��L`n�t���v
+��J��f������{���P����"+��'ޚ���s/l�>�ܕ�c<����[4s�s@9��hܶh�t��x��8'#�ɠ�l�-�� ��ـ���?�T�]��c5R73�篦�}�f�w�� �;��R�\٥��
�,��%a{a���u`�jn.b+�S��Z3�&l�,�1����cf9'��4��h�n�s/l���r̎Ldje1fc ��0���I�f~��_Lt$�I�F���fπ�o������-'����*.���;���o�0s�l�5%��ݗyLjt��l�����s��p���<o"mc�hܶh�ĕ�}���}� 8��0�f�ڍ;�\󂇃��[�6�:�j�����P;7-2�WtyH�A9����#Cm�&�w���GLjt����V�ե^3/�07z:`S�0l��;�f��t�c�1��������L`�cw����R��c�G�ɍ���-��[4�휠�4���b�"��
8������� �S=��$���)�@9���>W���u{� ?sv`Iw���UT���w!A�랬��/Y��z��՚�L��W�M��g�;$9N�G��<y�~���1�{d���hs�ycK$O��I4�e�@?sv`9ݘ�wf}J�U��އ����&��&�s���s�i���h;���/3�,��yn94=T�*��w� ;����[� ?sv`�R���I�pRG�@9�٠s-���L`O���U�ʞI[�˭�	  �.I��m"����sI�HLq����J�/���vmO��:Ws�-�f�@�k�̗=J�:�O5��������µ��mA/I�Un�uR���=m�t��g��t=Z��x�#^��\��e��V�K$Wn����ݎ��n]R�E;tu�e�Fw�}�&�D'K{$�[���WP��ˤ��Ϋ[ukZް�?���O|�f��1�պֳJ��i�N���t�U��\2]�⡤3Ƶ��͒��1fÝ��SP��O�`�1�n����[\��x��y1��I�r٠�l�s�h��f�g�˖2I�qI���1�n��������9Lt$	&I?��6|��M ��&0l��7zc ��,�����b���1�{d����L`*�U��z��i���DW�n�u�{:�����=C�ݷG긻;p;Y���M91��;�M �;f�^�� ��l�;s�,��yn94����A� �:�14����
p�`TOk����ʯ��� /-�9�����8)#�ɠ^��`ړ�1�n����-�� 8��������٠^٠^��h,�o&&<y�M��L`N���z��:��K��~;Bs��f��F������z�ۆ���[]�fM��8���u�N��0N�������K`d���B@�d�����g�z�nh\�W��� ��� �w�����0ć��ʾ�~;�Uw��|��Q�!%��=o�4�k�F�x񼉡̬�6L`�1�;��-�����M0����qɠ^٠^��`�uk����?�Is�������]�vX�i�J8c�Ei��ڦ�),˰�ϖFeb��4���8)#����ۚV�K`d����b��Yv�2���[گ���tx�=:c��s@�e�x�OLǃ�#�	�c ��گ�J_GL[�-�T�\�d��"�h׶h������u�ރ%�#�S@,*'�ޚ��1�$�I�F���͟�}� ��^ o7f ~���?�U/?_�!֮ܖ�IDλi��4��7hvF���7�vZGi��8�tmg���y�pdn�t���&ɌӦ0'tt��V�	1<o"hrdzyl�~ă���������znw#��#Cn���L`N���}Q0	�c딭�m?�
H�rh{�g��}�h�W��&ɌӦ07j
�e��h$s4��*�"��|�\���9W�������b����"� ���� ������*�
��*��**�� ��*+"H� �� ʀB��� ȩ��B�� �H�� ��*������A_ʠ�����
��A\|A_�U�TU��PAW�UA_�U�TU�TU���d�Md�| �[f�A@��̟\���   � P �        �   �  � �E   �! *�"�R��ET�

 J��B  �P� P����R��   � @�@P� �4�����^^�w�:��=�����l��{�����n|Z]9qW}� ���������x K�ݗ��ʧ�PO>����U�]����W�y��� =/(�ھW��/N�o�x��JP�
@ 1�Gz�N���}_�L��M�/M� 4���<��5{��=���Uu��/� :�d��R彷��Ž7���z�� ��\[�g[ŝ�O7K�   }X  	�{���y�l��MJ���@*�( � �4���Sw�����v�.u6��*���7zS�u��wU�G��}�S�� ;�Ҕ���z.3�@ �"�E/������ r�i�ER���ӳ  ���  ��� t� :1(  � (

(P�R���zi�,�@=�(l��N�s=4�N�(�3�� ng���P;�N�0 �iJ�����e� ��K����Z}��T=_m�=�Irk�W}ܫ��U� ޞ�}n���������qeO��� �
 H 6 �If��t�a��r-֖����V-U.���j�i������z�='�Y�]/=��� 	���������}���_isoY\Z�7W���t� Gs����ڗ���|���n��ʞ =AL���h��!?�S�J�H��<z�TOTj� фOb�Rl��  �%6JR�  "Be%(P�2hx�R�������\E?�_�r7N�Qt���$�Q�7���
��DT�`W�`W��X�"��� D�ԈX�`�a�F��	 �܅?_��3dth���R6HG����2�������K-��>���� �������s���F�
���n�ٽ�� ���@�>���oE`W�z�k!!�,\	q.��|RЗ������BcDHD�Ft�a��8Ĩ�	� ��$H�:��Ł�@���Nsi��y�L�rk�RvX�0���5�R@x�,FH#��
��JƁ��qSB����H�`�!#!H�B�"� K
��HD�p��HaR� ���@� h�%i�1�#B)�#R%�X@�"2BE"��D#�0*ƬkrRp�Ȗ%���O,(Z�B�8A���3!�[�q�rb\�Fa%%�H�a�Fb�S[#�vH$"?!
a�B��K�d䄺���Kؖ$�H�b�"Vb	cI�^�с$6QM0���J�F$H��@H)���>�V��
 �@Hu�I�)P����p(��R�\)ডr2���3V��I3	JIBB��$a�@��jB�7Y��%6`NO�'L%��4\4VP�'�R}�T3`��J(m`WZ7�d$a����h��k�����v �Xt@�:�#ą&1�I���@(h�J��4I(|}�J���B"���
|Ƅ�
8C�IeōXĈ%	!�[�ѭ�d���&@����ZĲ�<`˕�0��=��H$�2���\���vu��󗓁]�Z�ۢ�,����ؖ��H��%aR�I�!�i�֌��d��8ɘ����PR%J�DS=���ۭkXHh��&��4Sd	���w���� B�@��, %�#R��V0"H��"�`3A��1'
22	
$��X�FB�e�YRS�1"�D#0R4��`I �@� H(@4l�U�Fh~p�`i3G�+
Hpeb0H�>��\7��{<@b��!@�Cd�$�*��@F�*BHI ���܄l$�u�a����� XVP!6B�D'�$
a��<����'���E�X��D�2,l�a�B\�D��
�	�D�$+8�N|��T�Y����m��5uV|=n1��CA�0��+E��,,��]�}��{��!�$`%�$�X�`V@����r��M��`�(ƃ#d�ы����&f���8HB!R1�`�����D������I9��M)�`B����*H"�Y ��)y��k�99 ip �4tHE�����RdI}���!A�.�����cRc,+��p��m�ec��s	B��WC�J@�B�р�ABFFA�H�
�B�h�"�`Pb���5�I�Q�B��
�D�����)��T! � h�́6d!��D62�HU�V\ ���X!�J'T�0 D�hY1��`�#�
�kW����� B0F�ͻ
���$�RE��ɦ$�IH�������ᭁ��4��JD٘�l����iԍP�# 2V�$n]o����HI$(�dB`q���$�$B2z�BH�D$B$�i��Ʉ+�Q�D��RH6$"@g��H,�C�>��p]m(�q��'	��!L!�4ˬ��D0�&z8B��	a5�++aA!�P�mvFF��<v��x@�I	�,�d#
���K�%i�F#�f�
bԺ	��x�KJ�
��	l�t���*Ƥ�n��Sa�HGCb@�JB˛��R0#��5�Ml�!��	a"L�,9y�|P�͛7�ܑ�d�mԡ'Ƃ7Z+tBP�FX��%HP�m�d��k� I	I��a"ȑ(�BB���sI�n6藦e��`D�e�p4I
��@,�$H�I�5x���G�!���9���׺�ΝB��$�	�H1A�B(V"�!B!	!�f�zӘ�I�.����042wA�1!ƌ@�ҁ# ���`�!B	 �IH\!�|�4m!VHЍ^H����zk���]sL�־c����I�s�!�b�	B4�	 B��rp!IP�HX����n����3�v�WS��)�a
�#ą�X����������47߭%��5?
D�x��X]Y08(C�.�2�LcVi�Q����y,
�xH,J�������
��+��6L8�\%١�XWи�
jB!	$�$GS�!VHQvmB�#a #����:C����W�wJXXx��k�ጻ�
��F�+D)�A�H�F�(B�!�H�cJ�.0�W����	/�}N8���S��tp���Hh �4�!F0b��ϴ����n�f�\%�LX�p�CaHaC"����%3@��!L$u�E9�����Yop���H�/M�e����i���,n1,s��'��II��Rm�a� �B��D���)�	61�c���Y!#���$�I��J4!B��#��2Xc�I,��@�)ah�)��l��7�dHD��$��B�U}�XL3�.1�
A��1*�b�"���š�$qXH1�]6N!���ب�f_|y������Á�q*�$!��P��'D]Sd��FF$|��RM��f��fSi���d������0���Z�K������2nr�A���^}����to飄�G��$�H0�¦:6H�r1�$��O��!����w-�wt��G�f�u��:3z6��j P��-�p�5�"��L	m̧9p�%�c!�I��G��!RP�7�%�o8k4�|���t��� ]�Ӛ7N���[#��bG4ҵ�a�\p� HF\0>$%04SZ��N�� ϩ/,j�dLk���$$�G$6G	p�[HgӖ���v&�d�E\��M"@���cK ��S���f���F���B�J`|B�I��c~3P�̡[f����Ɵ�������T��ļ�����l���1�B�n6IM�27S����aH}	IH�R�JD�V#YH��KJD���V��R5aX����SC��B��Lx�B���Xv�g+.� �"U�0�1�c�"P��
���1�B��e5a�\b�"�"�$!�݇�z#)���G����]B1$�D���ٲ P�P��B�6�\4B��H\ U��ۭ�$h�L��\H��
D�:$cXS�)6wZ{�5~$����.da-r�@��%Ʊ�08�pҰ(F����P�]� I�XĚe!�H����k�,�����~�݆9�}�/MK���Jc�+�h��F��B��\2��CaG��# �-n�T��u�J�;�x   �    [A��А ��                                                          ��  6�             �   �  ��*�y.�e%iU�PWT��+&\�e�`((����v�R�p�fG ���#m�E[��mm�-��n6�	 U��3�F��4v燚�W:j��$��b�k�m  -�  m�  
P��C��l>���֐2*���A!"�m�۷7M!- ��`�6�6  �č�L��$�X��  �s�8 it��`H[@���:e� �<m�դ��pz��vۨl[@q��m�m�`�Q� $ �� �����M5Qzt��t   >�� pH��I��p 6�kX$.�m� $p�m�m� �;l���- �I� �u�M������͉�[��$��o���6��m�t���&�bL��`  �lk�g@ m���M�ٶ��m�m� l  �m�-� ��Y`�gIEb��f�
ѳm��P jv�kN�iШ3I����� �m�����{[�6ۀJ�S�l��6�%�L�%��־�!���e���\[G��a���l� -�m�ͳ[v��:@[\�i+۳m��8��4=�kh��U�Y�3u<��\PR�J�6[��Ay%ꀎ��t�Քj�M�[T�HJ�e;gm�ඌ�[��-� m� K�͗[��Pp���9�\ޠڔ�S+����2�����`�����@J�H:
ꪺ���Y�	PVV�����(_Z8݋v�g3�/���r����~����=��ӋM4�66� �`�dN�Y\aU�ppY3 ����u� >7�&���vTUwFժz�������$n��[AmH��� $ �� ���ζ��A֭�����g��$Y&�km�]&��M��    Jp�[�8��  �K9�6 ��W$�:��`n��
ۗ�v�t��.ݪ�U ����V1�m-�p�z�6���ZM���z� ��  �lk�m�f�%v�#n�� 	  ��5�j�;m�^�[@	e���̯�h)iYZ�Z�% �.��I[a�  �n�,�;tJvH�`K��T�T���R�5V�����U���^��UUݪ�����2��c�ֽt� ���S�B�j��Ml� �J��UUP&��Ғ�&@L�J�U+j��ʵU9#mf` �tӦ7mnl�J[v�	EI$�8�v�l�n�	��l��mmm�)A�� /*�=���h�i�2*ˀ-��a�k�m� kv� 6�m��6�L�2��np*pF���o�2�YZ�m� h-[P>UK��e:��@ �u�ˍ�` *�U��'f���$�Bۀf��H�dt��W,ҰA��$m �4��@ �X���ͱ�j�bڥ� N1�
Z��VV�A���hH��zt��� ��f� m�� m�$,0m�  El  %�m��Mְh�hm��BO�}���E� ڪ�eZ�s�&̵�8Sm�L�U��e��` ���6��a��Ӏ$ m�H6��������uc#,��ݕy��e-�K�� @v�ӲC���ګ���U�����  �6m�� *ڪ��@VI��U���z�v� *�-ֶ�I�KL�m���Wmz�� h 	9m�[M���長���b�\�\�#u��:Bi3)�Ӎ�@�I%�y��z^.��� ۶��N�c���H�b��{M�(- $�m���k������콡�ڒ�H[��I�{�� ��Ö�H��v^��}��� �m�       �J6�ͮ�֓E` t�����]Q�Bѭ�ʫI9�cG.�Pk۴����p��s�� v�v�ڐq���Ͷ 2I�Ͷ��Ț� ��  m� �fM�H�   ��Iv[&� m    	 8��a -�V0 Hmp����{I��q ����m�gm��֝%l[@	����A�� $kX6�f��@��n���(��P�*�UR��Ҭ�*R��*Ωj��'��Z� 8m�kn�l��8�,�am 6Ͷ�UUHV�J�����F�[ .�]m��y���m 9��i���ͱ�tM��E���&l.��z�m ���"GL��P)��p���R�h	U
Tv�vizɲ�m��p$-�m�`�6��l�-�6�08sE<9�̋RF��o�|	'�����ݳne6  ��.�m�A�n��Y�m �Q i��j�������U@��	Z�g( +[]mn�����m l���ڬb�vy�eY�K� Zkn-+i �%�I�h  m�ԭ�@���  d%�l$���$�V�m2$mpj�M�Jm������96�[ 	  $   �qsÖ^Z�x܍Ul(]e���Gi��$�f˫k�WR˸�vr�@-��n��f��0��s����s�e%��^$ݘMIUQc@���*x�'7UN��jW%�;u�mNl�5�b� �mmCZ�I&s�K��Et�R���=t�&ڶ���^Zu���'�P)� l����[�!��p+P\�m�)���	r��\�oR��2�X�Y�  p[@���   �a���:�˒�  Im$�  -� [@ ZlI��  [A����$����Ůl8�l-�J I'$ m�� 	6� ��� �e��)�n��  p -�Z�$ �Mm�h ���D�@ 8kkm��6ͳm�5�lHB��%���vۀ   m����nI�h�am� �bݗm�p ��� 6��ko`��y�Vܴ   >�}��ඤ8�ޅ�F�m���$��� 6�ש� p �e��h��`�j� 	l[@�66�P[Jܨ�h
l��F��M��&��Ͷ �� 	n�s [Z�o�'�ڦ�m��� @�X���uT�!5J��5\�RC�F�6�IN�!!"YF�6��Z�-�,2� �	 ��U��%*�( ۶���$�    [Z��H,�kav �4^2[N 6��.�|>��3gZBٺ�[��s�M��bpmt؀ 		�28&�i�/�O�vp}JU��!�<�T�ۀ-�57E�@j���  h v� �`` -�l�UUʠ@�6���8j�Ef��V��  ᐐp�%�  F� m� v�$�[7fۀ;e6  ��bKn�Ė㬗Edݶ m�k��Аz�h� 6�M���m��� ����� i6H蚎��E �/Z�9 n��T����8 F�ۀ�O$�6�T������ڵ�UYI��j��YZ�U��{���FݎH2Hm&�L���["� V��G`�[@m�m	  �@����ҭm��2�ti�m���E�[v�9��
�5U@C�����g�W�['^pɭ\6r�YT6RwKv�uB퀨�0�T��3i���i��ꪷ�)���Okm���s��A*�U]P 6�tA�H��mm��KoM��m��@[G6�.�t.�@�m��tl[@8H��ݲ@m�m��]0��m� 7m��Ŵm���  h6�l�m����p�l���ְ�D�:8,흦dv�l� �a!! �
�[gK�j��H[���p[BF�d8�n��+mS4�mٵ�H(x��jVyyV�e1�W6ܐ�m[p �����  �������
ڪ�zp�Ҭڶt���}���p8�^۳-kj  ]6 ����t�V���IU]\l��h6�ˀl�R�T�0v�6��*0�Ͷ=$�P l�&�Xۮ����&�0�v� m��$ԃm�P$�v 86�\�<�ԦPx�:V��$��� l� $֚�U��J͠��&%]�C5Ӂ�!m ݷ6�X`m[  ۶[EWEYD��MR�����\ [Z^vi4U���Xר ��d�֭��f���@����uȵ�P�û-,�,u�m� �m�kũ�vm[ S�)VIV��h� ��lD '���Ab�J�8�A�E'�|&DQ�:�F�@��H	�t�� �\I�&& �"�(�C�:���G�Pz��@�<R�� ��qM!���'��x�b�u���x"���u�(uء�X�<��gH*���ث}� ��U� $!��V|���<p�m0j�� ���*Ux����ς �`�Bh G���
	�^���<�!���:�4bmZ0��	��6�â��õDt�iS�*�# bE�E/U�?|����So�� �Z p����GB��z��"����@v�@D���Q��Q:"�` I�W���@�A�'��>C�4�U� ���q��a�C����Z*��P"H"�D­�t�������.)�"�"�Ci�=`=t_�	��"`�� s�E�Ax kh�P�M�*qx*�#�`	 ��HH�C�M"�H�Ҩb+�"QOiA��'¸?P�u��>���
��?�����$Ũĩ�8�Ei�\ �����"CE� R.4@Ϯ��֮L�H�           l�  [F�$�;mo�n"�V+��J�J��I�eP*�'!Q��#�c5lі���u��x��86r�pj��)����k��Erm��m���ld����[Gdyym��V�c��FP�P2��[uƹ ]gp�];i�*6E[`tP猱F�Y�,���`��&�$�������t�F�I9,�1�\��.T���l��ң7f�`h;$���u�Sn7JN�6�j��#���P��םƴ�#P�ۭ��sbûu��d6��$9ˌp,,��&��[:7*cmm�Ę�1�s�n�Vl��Z2�&j�U<\�� EN@�ۜhr����3 @�A�ƛ��A�L5�OR�N��n;C����5�j�������V�s�#Ty�Vs���gLK-�l6mc"�-lnQ�mNg��t��J�:�]�ιp����᝟F)�l�3\$5U*� �Eʑ>�!�\�j�:9��T�K�$$Z�h\�i��	��T坳���� ԮqV[�JZ������Ά�8�OOX\�8��U���sO*��!��@V�+j�t�*��Q�F�v����}QimXճ��C�M����I�F����'R��F��YٵHB
���L[3�< 2��J�$M�eUX6m6Y�R�6cHܣ�U��*B	�8�1�c�Y,�.W9��]�����:�r��ziѪ1�`��GZ�#�ha��ʽT�6�tF��]�#ur�-N�1��:�7s�A�dTU]�H��dv�d���j�5�-��@���Cͨ8Tx�m��8��ksH�x��m��������$=m��:��6'ףx�%7�)�4��i�k�u�V�(�T��ŕMLWRD�Qk��m�Z�u.B�Eq�p:�fuD�&5�,b�����u��WZԅ�4���v��#�ҼQ���>@� �~Vi
x��x��Mu����{ޞ��zw�wt�ww�O� I�p�W�J�ۨk�G8 D^�I@����(���q�k����tl�-��t��u��)W�+r�==�e��n���7 ��j^��N�n��י�<����͖W"R��QuKzNn2nx�ƞ�c Y����i��c*�c�q��.*���C؆�B=��s��=]��α�^qx	�]f�j[�M[j�Q���v#��n7�/+�����q�g���*�s�9ݹ8=�&ܞ&*C��$�7
�n�Հ}�pǘ���ϐw�X�'���(�
�)�+ >�]�I$�!(��v�g �i��H遳�J�J�KVa�fcK�0>��H�}�1�ˎ�RX�0�������0>��H�}�1�r���=�`uw9��%D��B6�Vm����xt��r��T(J������\��s�]� ��c��:�m]��ez�8{.�g��Rݧ�^�0�j� ���"`}�"`I#��m�r��r�I�`n��~�9^��E(Ձ� �p�ӱ
�̭s�=�ŀs���̼*H��q�8Xu�36��$w7���<X��"Jp|ljE`fu��J(�u��ݽ05%<���s��8(ܡӅ8�X�͖۳K���`ff�X�9U�c���$JS�㛰�ڱ�y��]`WCv'n.�$�y���u2�{M�m(�Ҩ�e4����;�O�z[������.�)R�W�VR���Yx�-�l	$t�>ޘ����9\Hś�:|�r�P�r;���ܒs��[�>  '�Z �HP	A1)D	R��O' ���9(ݧI�y�G*�>�l�7^�>]�v��Ձ�nۧ)�m��)��cK�0>[��H�}�1������R��n֗��5m�I�K�Bl�4P���V.@N�s��t�mdћ"���-�l	$t�>ޘ���L	��HD��$��9���u~�����}����w5��&�ӂQ�8*���s����a���'���6���v��ZI�Ҍd"RK�٥������;��f�򸦅M�{C�Yʪ�v��,Ũi�T�*I�>[%�$�� ��	.D��)޴vv��D�:�V�:�H�m�pբ�����:��A�.ٹ�Y�3�ٽ<����埀��ŀ�]��s������ ,�y�|�#@Ԕ�%X{�,׺���� �x��BJ&Fμ�V����jJr7���U�����r��{��Ձ��`oMKlh�pi�����/_{�����L���$���v��f��*���ŀn�{_�[�����`R�^ޜܒI$�IQ�q�3Hh�4]�qg'9�$8�5ڷG;�	ݴkb�1�loj�<�QT���U{$�>y�b��EƱS���X�\��hq����]ò�L�ƚ=N�'kh깻������+�՜F��M�D�:6��ښ�Nm�h�-��0]��837m��U�sGV��7*��n�9���v�ha�wj۫�r]�/`�ՠ����^�wow��}��<;�5a5�t^ܘ���E"�2󆽂��A�u�Od��GV8(ܦ�
q��^��u�Wd��:`}��*i+�BYH�]�[�nr��
����`��X�u��1m*Q�R��$#���wu��0ޘ���L[ߥ�VV%yY���-�$���L`Ir&�d�]��	�y$�V��������u�w�x�I(����mYjU��8�Q���6�Rnƣ�j����0<�/<�����y��WI\���m�~�<0>[%�;�:�W���`OB�2٫3S.fk&�jnI�����+U�$��"2Kw�,��]`7l͈�$n��HD��$��7�����5wK`}&A��l�d���^REX����N�{X7oL����t��eJT�Wj��������dl�����W�yI�`wL��Wa������{r\�z��0a�4��'0l��Du�����[��W^�sNup�O������lwK`}&A���]�fr�"�n;36���W<�|�y������`��`�7��nDJ�6����=�����Y	��T(S3�\U
e�պ�o ��n��A�F��qX�uX���	$t��}�F%�+�����y�����:`M���%Ș��"n\�bQm��t���]�^��٥�Y����n��]�Y���9�Ʈm��쵰$��m�L	.D��}oB�l�(�
�)�*��y��ʪH���0'�y0$�����#�ޯR���@��bWx���&K�tt��}���)F�eJR��G���U��x����Z�B��X��N��y��H!�d�8�V��Ձ��o��|���`f��`j��䈩*E��':tp�	��|��릺�X���cqӱ�]����9�I'%|���S��L	$t��$wfU�eٖ�eb�����L��0$����L	�R�KW��������L	$u`f��`n��`w�*D��$��K10$����L	.D��}fj�"J9B�
qʰ3^j�?s��^���{8m��>I%(Q	+��;ߝ�r�� jӮv�m���"�8ó��8i�S�]��,�j��.ڲ:'��cQvܴ�D�v��1����eh�9h	X<�X��mГt�M���) Nn�I3�[Ĺf���xz�6�O`Ŝ[��g�ߪ_�:qz�l��A��N��lmzu��nZ%�q��.�.չ�6�@[����n�[7afƈ�ݖU�Y�6H�
M��J
��#K+�EW6s�w�����7]���ۙ��G�];7U����cg�"�ڶ�b��u�;�� �Ƹؕ�(��L��0$����LY�iR�8ʕ�H�ך�܎�_D���&�O��+0E�Y���f&�0:_D��r&��0�k���r$���ך�׮p�pJ"�o �7���Sdq�Q7��l���y���f�X�5X#15�(�T5*F:gk�%��d������A�s�vn��<'�pi�Gu���u`n������w�Ł����"Jp|l�Ea�����}�0 <D�A`$r �1(F ���� 8'���.�w���7^j�;��t:pQ�C�
qʰ6_D��}K�::`uJ�)�+��bWx�/�`I}�GV��V,Ŵ�F�eJ��H��p����`�\�u�8����7�����룉�[��[��OC1����M�P��V�DD'=%�v��nu,���Θ_D��}K�՚�>o#BNB!�V��W�H�l�n���؅��{�ϡDB�5��J�2�8�"n+}�Ł��U�����d����D�iE4�DSjي�"�H�4/D4�|�;XNo�M�K2� ��B�l"B3O�3���2��n��3���I�}^ :^��zQ�K�C��	��`��HH�!��	p<)�=|��?8�J9 T�!�F�|<��(Q�bp�,�Ęx��k���֊�M���H0B$HBv*��j;!�O�������|�:"�t���)�
f�����S�<��E�*�jbQ�$�Z���ݭ���xJ�'�q�N��7���o����Dy%[��� ��>�R]�����.n� ��ŀj����z�L��Vw5	;�N�#��%>�na.y��`����{u�k��;!X��쿽���}���`��2*q��y��Ku�� ��t������J�2��]�`t� �u��׋ n��5/*�gv|�Li�T���������`f��Y�����X�,���[	9L�I����J%�ߖ�Og ���bA�@"�d@����~�(�%
Ds��}8 ׶�5�����䫵�7]s�|�(Q��i���pw����YP��T��%2>$�n2?���n�=��%Լ�a��ָ�n)��������G��Jd#dq������`n��`f�ũBK��{8�eN�.�������Y�7]s�����,v���;e�9_�پ��S���5���UUC������p�D��ޘ�=���2�NR�ȩ�*������X��,�p5D�^���n�ɚ�A%�.f�� �� ��B��}<�}� n���O߽���^����'��� �+���M��ϱм�SmOIg�n��Cm�;�4u�q$�e-�lD��xF�<��A%���ib�M���@�v�8�k}v]��ت�+���������Vs���`�[�$4N�ܜ̞2F���-`��-R���j4s"��r5��814�/X
;<M�dζ9ާ�kv�#��A��]ME8Lru���y�r���H���	�3�%/4̅�jj悂-�YH�J�U��&Ln�ujh��3v���d�`(ӌ�Q��I���Vw6���y���秋 ��	9L�fb�L�?W�H��y0'{<0$��~�9Ik<�O��hI�D�`{�}8�v�?B����ޭ���`��ۧ)�m������W9\]�_�=
gޭ����X�
"����5�K�I�6�8X�5X����UI�� ��}8�v��pnB�����W\b::=�m�)���{Y��OX{GMtk��T^{*��ܮs�w"��S���dR/��{� n�� ���脼�!r�ޭ��w�!J����J������Ƣ!,A��$�!$��Q���/� ����9μY�
<�BUF�{��f���ԖIUs�u��`�\�)B�	DUw�q`��+�h
4�*TdpRB��ʥ
wm����Xu�8�IO;�� {sт�d��I���sn�r����v��:�p(�דR�u]�$ke�7n���5�4��&��_T�CX{.�K�D�9�\���t'��hI�D��?O�Հ}�l���ߤ;׸�$�^�/��NS �#�8ۏ�;��/�RG���y�-�ߪ�=/:H�/���E՘�{89׋�䈈DB���H�C(B�>�W�竕U7���`fl�`f=Z�(�NN�"�Xz��3}�XY�;����ܮr��o�������P�¢��<n���w4�t�ps�������\��f�ml��<^�W�+`Mq����v=���eA4݇�y����Y]�_�o{<0'_D�����l�b�
4�*TdpRB��y���s]0"�-��2iߦX,���ņf,��ݑ�-��� ��} �����4$�"qʰ5wu���0��I7
b���Wj������71k�NS �#�8ێ���4�k�ps� ���(P���S�����:Xb���I���m*I�vi.q��l�v[���9a8�9�+=��ͷ쫞Lގ�l���fA��d���ʼ��̥���0"�-������ښ^UUW1��N	G(U'"̦)%�>ِg���*��y�6�B�&���&�v�٥����ps��W��Հvwg�u5t+WEՓwf ���p(�{�.�~�d��{^��tE� 9W�,33�ֵ�;}��N��5�	��Z��^^x3; �E`��퍦�C�&�k���s�w<%�	K]�`Ҝ۩�x(2�ۖ�Q�îе+x8uA�n6\���`��7	�]�b}���R��!k'Xӻl�%]���t����Ѵ�u(�[��awl64���=p�u����@��;��v�@�ƂP�<�P���bS�Gsk(�];��J�)HJmέ�S�V�%Z��\5�j���؎g>�3�?�%�ԡH2I#��Z�]X�����	}!�S���sH����&j�&�� ��~^�G_���U���ͺ�W*�#��4�Ӝq6��)����>��Xl(��{׸���� �t����*誫�]Y��P��D$n�����`��`l$�S��i�7G�*Q��7R;�ͺ�=U�r�������`wZ�vWR��4�gc�	�/1��z����u�(����#�\�Qs�n���w���>~����7�Ew�cg���|�l�8�z�T$���q`}G�i6�D�A6�>ܚ_yL�U �����H��
9񽣻X��,�7]��[��i�T���NB���}l	�3�yw�lt�iߢ�affb�/�l	�0"�-�'GL�f� �h��x�rrU��d��0'Y��tt��|�e���cN���=&}mQ�v���j��%��I^c���^zvMۋn٧��+�neg�!(�{��t=���X�7X�ۡc�m�"r��f��~�l���,�����Ś�L���̩�-U��*�们u�,��<�%iB��	���mz?�}����Ձ������Rl�(�
�*)*�b"v��X��X�u��w^���3U@IjK&�����`�Z����������`}�6"�dCq���{ti�z��f�(��� ɬ3f����g6׸��t�F�eJ��D�>�O|�	�0"�/� �L��=��唳$�G#�7��W�������=�<X��v��:��$������7�^�7Հy�`�v�8�Q�䃍��=Kٷ����|�I�훟������
�ҩ�qӮs��������~��U�q�8X�u�����qpK�� |� ���r~s���h���g�N����mSh�,\�X6���zJ�+�F����6���Fe��y�-���!�zY=l{k֛m7)!¢��]�w�H��L]k |oj�����ɚ��I�������fk�ܪ����Ձ��>Xf�J4�*Tdr7!a�$�W��`~�,��/(J+ۿ~,����)HBI#q�;{�u`y$�%������ݿ�u�QW�h�l�%���ҋ�DjI�H RCm�� <�V ��
�E}
�� `�|�0Gb!��t�0���~���m^�7ۡ�����pP���>0�v8@�!����n!���2$I�>|{>��b���?�u��l��`           @  ��$Ӕ�F�X��D�H���ь��ٰa��Vv�E�`V4:f6^x�l㓠S^knkV.6��UM/+�KP
=����gA�ϴcYz8;U��`�M\�Ҁ�6Ί�*����n�-�U��gHe*�:�tt ��/�uQ�k�[��*��e
��B.�X
{l�B�)d�r�AuM����&�)��j����0i^��8L�)�(��N�oIr:3&�Vr�� U��t�����n۵���e@V�+��f�Bt�^�E�t�خ�6A+Ud�#�Ň�$�h~�}��뤵���)�E�)�2�n����n�ȅE�\ٲ5v�KKd�*��'�}*�,���gZC���m!F� 9���p�ꍶ؂m<p&���*�	�P��n�Τ�.�Q�O$��kv��Z6c�r-ӱ��p���+����yn}r6ȩF4����An��zTr�p�ZRPɼp��U�R��j���&��0ŷU6t�N����s�B�3��m�r�M1*'<g����QՃYCSEr�fU��``)�;	����D��iq  *��ݞ��
�P
I�\m���Kk���m̜v�'p-�����+n��un�<���\]b��Xsj���j8�0p���vUٙMպj�AL�Ń��3�P�llBH�v����X�ev�iu��2ڨim�s�L|�}�Z�]mS`���%�v�j��V�vC=�ԛ�sﾷ�B���gn�e����Q�<�9e����ܥ���36-�^^��`�ieg�{�m��b��ٞ�9[�xp�jAG��]O@����؍Yq�w(d�7�nsٶR��r�	�N�+������4�!����T�N�F/2�d���I"@�#&�$��V5�j�,D��d 2AD�:%f�YM���ͨ�X�:����iՄ�F�[�#�h�f�Ҡ��u����(x67z���h�*��@~;����L�x q�/��@< �����߯ݻ| ڷi�[sp;��;��ܔ�nnc�Gc��M��uzi�g8�f0�Y��۵�$.�0��Z�X#m�w�����׷cq�N���ᷳc%�mN��%�u3�P�"�����gY���p�P5��ݿc����\�]\5���ڍ�Xr��X�^���e���^5e�&x�d�nh{O7m�竅�G��3���-5h&��ݭ~�������������ς�����[�×��?]-�0�^�1��rk��XM��z�e��SF*�06}�V ��f �G]j��7���{���N8�drB%#�72i���t{h�V��b��͙573��*�q���N���`own�����}������3��h�)��"$v�GL���'vA��{����<2�q�ܤ�
�J�5w5��nߏ��3|���Ձ��9Cp�)���q#����n�H�A���rZ�i����u���/%X����M��۳Ł�fk���K˔������
f��j�ֳ5��'���f�"v6>b��&�~W
"7�o�ŀv[��{l��9�R���"F�$v�v�����g�/n����`|�F��b�S-�l	ݐ`M���������j����Zd�6G$"N;s&����O_�{��L�����bW*)	�`�s��ڶ��pn�-[�U۔�H6�:������:��v�3���7�=��X ��~����ݿ����d��:N�$v�v���$׷�kw� �G]g�z*�{|aTU�MU���W7k <�׀>�هJ*#�L��(I-�	W�:3k ���ֆ���*f���U��y%�Q^����F����`qjP�UZ��K�L��)�q9#��3�� ڮUow~��7=�`nd��ŘkCq��ے'BX��v����3�cT�C�=&kdx*���xV_,R��$`�q�?��{�V�͖�M=ϐ{�v���O��hJI75uk :�6"&Mn��7�=������I���L�r$G$���g���b&w���z���v^!J�*誫���0<�=���`~�,�O}�kr�D��D"����ED�A�HI8Z��.%	yw/φ���&�TIJ��.� |o�%^{������7��vfj;�!���>am앷���fI�Nz���	��n94�l[<��9Wi7Mʉ�eE%|��Ks���Ծ�����z�XISV)�������{l�G���}X��� 7����a�E$G!N���������&��H�Oc�g�8��.ӌ��n2G`own�{�,̚Xy{!�v���{��'!�U�>u��Kۿx�to� |o �X!	��(!����~  ��i[�M�r�l��iN��on�mӶRS)�;l��r����$��-���Yy���DOW�ݡT�9�A�N˲��U�ʎ�ٞ;t�*���}��}��٧]ђl{�!���w`����+�ܬ�ͮy������5�/B@#Ns@��g��g��5�[�-�5�:��ݶ��9�6Rۺ�x֚��iO\�f��5��L��kW�j>M��,���K�%�Y�ؠfT���}�hl�)��������bYE�s����}tx�s���$�w���(��IB[�{x�d�R��ێ$�`oY���Uq#��]X�},̚X�V�IFJ�C��Fe�&��M��K�g����`n�m��m7*'Q��a佛�`y�� |���5DN�w�4�l�HUX���檪� }� �$����ᾮ��b��� ���e��)MIj��qP��6���Y��)���QE�X\�Ň��\�n褢r*8��H|���`>7� :�b(�C[�0X�n�j20m����ݺ���8Q�G9T
���Ђ=b ���$߿}��o]�>��Y�IyD(J�;�h*��u$�]�5uk <���{l�a%�uѾv�޺�7tSS'$N9%9,9T(��i�����>7�ވ��o����?s�'�M�1�I��޳��&��M�	ݐ`}��bu�#��󞍲u����6r(W�nN��7:�4����{�}n��	�N3ˣS������λ�{l�
>������z"�ꦪ��+�\ݬ |���B�=�~0:7Հ>7�5(Jdkt�*M£MDےXݞ,�3]���+A�c�s��D�X�'�C������7w���a�E%��Q�$�B�a(�;����ŀ�w��$�u���i��m8�H���$v�v� ���V���n��(��w'g�j�Ie�F� pZP��+s0=���)��˝s�`1s[�m;/�I��݀�w�>�ـ>Q�Z�!B_HowqX��9 �q��I`nd��UIBS&����owq`�]�%
=	Dq��=�~
T��qĜ,��~v�Xl%&�����w�&9&��M�;Uq{=��=���72i� �|�@�����&�f�׾(n6���U�`��`nd� }�����`J!���4�}�Mvi{�/WWZt��:v.�$�S��^�� �e��UJ�wE���Q��m�:�z~,�:� |o�_H׷�rY�
n��T��E!`oY��ܤ�g�u`Ƿ�>�ٞP�z*��lzꦮ�.�*�����<��X ��xl%3�ޘ���`V����	9�r�=\�K��c�g��:[l��z[ĭg�7���v�M,s�����޺�5wu���Q�w�ճM�I$�I*�eqJb��t��t!�n��Ō[�U��<A�˃��n�G0��lc���i�h%�G�#u�qB�rL��u�[���*&��q�c�}W�k��l���ۂ.ͽW;3���Euf���C���F�Ԟ9.;q�����\Ԥ�Y�(\�	�L�Z�7l�Bv����d"ywx�캍��mí��&xl��L�vܷX{B�^�{��?=ﯾ2��ݬ�y�Sm���Rj�m:o'EX�<d�=�������_mJ�cn9I8x������Ձ�����|�۳Ł����(�Q�t��.p��f6z��D%H{v�`݇����J���F�j���]�x�m�yB�޻6p��,�6J�F���n;s�^ݿ�a�`oŁ��"�o}XgM��M]
�թ$R�!���+��}_��`nd�����R�{�r���r�jP����չ%��=Y�v�9P@��v�����F�̄�m�E��z�����`nd��9_ �l<���`�=�Г���*�=~�| ��H"ԁ#,�@�1��$"@H�!�T�&HD`AH1�E�"A�B0"@ �t�(	T(�����D/G>=����zp�������g��$��6������>v�8z<�EW��� ���`3�)Sc�m�p�>܆�{�u`vy�X��y� �M�n�V�f�UM�s�>7� ��k�5�� ��5X���D����JShpn�9�T�7#�݃]J�\1ql����s[k��?��y����q�ܥmTRW�j��72i`}�>Q	y$�(<��X�������J���� ��v0&���z;�U�~�r��1x��)F�eJ�Hڐ�;�Ӏ>7�B���p�B�N"P�J�@�2���C�1�R�	4�C�U�	o��7����4�`0sB$.�  (��X��R��P��$$O���>R$	��lU�!��
� |�# �%�A�a�4�T����w�u6�P�S�o�`>\Q��G���A�+��N�����C�� ��u��Uو� u�Y�v秋 ޙ�JS��6��r8�{�����`��`>���;���O��Гr��s]�ꈅ���vl��P�����,���7��V���u7It���o��<֮.�k�J�/����ݍ��{�|	y�N����p9
�w<`�f� ��-��DGyo�;��/�B�ێRN��D��#�-�l	ݐ~���$��y
2T���ڌ���{�V.�?s�����OŁ�����y���d�ڑsv�5B�]{X�z`>�����(� ���{��=�[w,��ԙr�+��`N���}���y���v��r�r�ί���I �n&��;/V��1V�<=��A�Xf���RY#.�{��k�)(��	�ԇ@����`own�]�~�W�=�<X��y)N2H�m��dt��z[wd{����t'�q4�nP��`yf���4�ԗ�a�`{w�V58⍪���7u��W���y힜�� ��`oM[t lq���$�`or�/{w�\��Հ>;fq(Q�����{�_���@ ��\�\i�e��p�ȡ)���U��J��Ҷ���ujݶ�Kt*�$��]��.�qّ۷qu��9gC�y�^H�͊����U��M��K�
����6�*�\��S���3f��Q]�kL˥n����A��F���a�p�V7l�qge�Q��'iۦ�v8��(�a����4�7nm�Z�>:������_绽�Ӿs��e�Tp���n==`��xW�+,=I\<�K6���zg6W��v��vU�uv^Y��H���ِ`or�܆�q�ܩMS�U����?%2ov��9�͜��jS'V�R�Cp��Q&�v��Ł��j�ܤ��� �o���h�(��$nSWf ����x�<���S����=���Jq�FГn2+s6��Ԣ!mu�|�oL���[rwz��:v����>�����S��j��8d�]ζ;.M��6�c//#�� -�k��o�����>;f��|���oq`vu�l�q(�GN)��٥�UUUYʨ :��� �>ª�響a���09l����(�U�^YwqĜ,�CU���ufs��*����y����:�nҎ�R�N�j2+��$�)��X{�X���B�<w�Ձ���C��ܨ��� �����L�w������v�]�̬�0�W6a��#�]�Уփu�X&�'p�+O������q�p}���D�*�m���y07{�wG^���}�c��z�H��(��X�Vٛu`n�>ǚ��ă4�y)N2H�m�\�oq`�n�Jȵ*R�J ����4_�D��׳���x��2��>=�I&ܢI*�>��`}�5XǕ������}V��߄����A9,��ٳk��;��s���$��$A"�@"��\�޹.�WWZ����%��G��ѫ3�r-&�م�*ܧA�]!�m-;,�Ғ��1�'�g^V��ǋ >m��r��[��=.7�U�-Z
�j����f�Xٻ,����s� �{^V|�����8ې�� �5��v�~<�eC����	G�E	D���{��<����O{�i�s55&\��u�kb �`�b�`�����b �`�`�`��k���A�A�A�A����b �`�`��)�P!�@M!t��u�ߵ��A�A�A�A��ݙ���fk$ֳ5�Y���A�A�A�A���؃� � � ؠ����b �`�`�`�~��kb �`�`�`�����b �`�`�`��?~�O٤�{BJ;�ۧF�F��z��VqIq�=sgf�(���G��8��R�@�>y���6 �6667�{�� �666?�����}���k��v �6667�?�%�?�����5�h؃� � � � ߽��؃ȏ�
�C ��A�A������A��������y���yO�!�A� � �]�K�Nj�d5�4K�kb �`�`�`�����M�<�����׏�b �`�`�`�����b �`�`�`�~��kb �`�`�`����p�Md�d��f��M�<���� �ʢj=����؃� � � � �w���<���������<���������A�A�A�A��y����h�&a��F��A��������A����*��kb�A�A�A�A������A����׏�b �`�`�`������F
�{��kZֵ�kZ�n�,�
л��-�Vö��=8�����n��xwk��p��tn�b70s���c7�[)y��LdȻ�����^�1��c����䨷��D���r�;-7��Y�n^��ؚs�8��ag��I�g���9b�2\��1�2�ג�u���Y������d�7�RH"�m�T�$��%<���m���w~��{��w�������F6������'�8u�U�źN@����!��펞O��?}�B�4f�3Z���6 �A����w��� �666?����A����׏�b �`�`�`�����b �`�`�`�����&]M&]\��kb �`�`�`�����lA�Pw^?]�<�����{��<�������kb"`�`�`��h��[�ֳ֤5ff�6 �666>�~�y���y��~��A����o�؃� � � � ߿~���FkSZ�as�5v �66�?���6 �6667�����<���������A�A�P���{���A�A�A�A�?��q��-�34j�kF�A�����ߵ��A�A�A�A�����yw^?]�<�������6 �6667��Y/��kY���t���e�� ��7�ĪW0=+���� ���\��kN7:Q��w{�;�޳������6 �66}�kg m�/���5����;���1�I��μ�V��9�;\��v]� �I�	� ���R�2�������s�>����]ᰔ%3��� }{^V�ݡ��q��H�#�a��M����~�y]Np=Q��q`��R�������K{�K�����oq`Ϯ��Q	.�fY54�-
n�h�,K���J��b��=3Ľ�V��.śR�����u�`E�ұ���m��ey0'tt�>�1�6d�)�Ŕ�$��n���۫�W�},g��a���v����?r$�n4I s^� ��z-
�D
x�LY�-�����n��[t��8�eH�
K��	/W���l�� |�� ��[b�m��$�`b�5�����5���ـw�r�eʪ�3���V�n]n�1�n�TQ����f����ڵ�lu�r�:%:�B;s6��>}w�>;g��[6�[[������Wu2]ݬ ���o��?_�gt�`��W���I��e555��oL�ގ��L��ŀ׷�}�]�i��#n!�qk�<��}urI�w�ܕQ_�"+ �������	�h`msj���gŀw1o�9	#t��B� ����<��w�����`��u`�P��Q���s���t� ���h���R��=l�[j�Si��7�5$rU�}�������Řk�9U��޺�7�^�T�I�����ɦy/(�Tl���`Ϯ�ЦN��+L#�A�������t�>�۫<��2s^� ۽0�v)�.�j�U*���>m���]��m�
��y����cQ���C�`nm��m�g�`6�`��.�H��oɥ�`-8��������*w5}0$� ��0�C�fou���0$�$�FZB�T�+``'>�
�?`�� 0R1�	��$0	 4�P�6� I4��EBH�6
8����$��d� ���� B0��	�8/��>����F1���I�@Ӹ Fn6&:��Ou�}�;��>[v���]��            @  ��f۴�tɯ5��9�n(�wO�y��+J�J[)�:,��q]h�8�'u\�������2�lY�� ��U��ev�gIۇ,IzJ��=u�i��l늕j�Mٌ��hj3��}�J��l:�ήX�e��nd�NLVʦf�Pk�ړ
�T��<�y�e��jz,��M����C���kN7&Ǧ�D��mȜq#�t[Y*�횲n�3@&w$�U���]j�	zU��g�<��u���m,t��*;h�zA5ge�7I�uC��nV�:�[#�t��������8(N��3��C=�Ɋ���ZA ��R�:����D�*r��^xK*+v˛&5�'S�! Q���.\v��	��qpn�@�Ӟc��=�)�Z��*���h�N�i�h�-pn�1mf�gE�vFn��i��K4p/T8�둶�-΅褠���[r<\a���U%���d�mRd�S[B�j�6z6�f�����b��.mgg�v�e�;L#��V������T��Rt5���e�"ؘ�NJ6Ѫ�S�"6�T�M�\��J���FJ�,`��n�rP6����U:qvˎ+�K��RTk��S7V;M�E��s �[b��.Jt �H���f�/H�]�����VҔ��pp�@]������9IyQR�N,�>je�Ȁ���՞[Y����'N�W]*����k��۵t���e��aVt�R+n3���vۦʰ�坣�
m*�;�K��9���2�֊�^eg/T�m�B���'/ uT�8��G(q�nu[(�ey@�7����\�\��y;��y{Sq��kW`�`� �:��Rb I�KH$�bBz���T)[��L�	u�Z�e�s� �x6g�:6�gk�Y�q@�' ��U��m��X�I�f�V��GL�RT#"D�.sr�e̹322f�t���: ; M=|B�w�]�(E����v)�`�~D8�����<���kZֵ�kZֵJ��R.Qև
f���ɞN���\�,)�΃�P����;\�b�{H"���k�䭝dz��Ԁ��ʁ�S�,t�hz�j�O*m��u�6��GP�5vi��*�bn�5�c-;���E=��	73uN�
@��F��r��0��0JUjq+�=��%��1�8՘��p����d��yR4��Xn�u�;)��y�[y2��F�5�E��kD<]j�J��Yu.�%I�x�y.m[S�\�_�����e555�秋a������<�@w���<�o�5SSsr]U�.�.�[�#�����_�s�����ߗ�5�$��n������}:c��]Ķ�:��ylm���=Ļ���7vx�1f�<��{�7�^�T�I�����{l�=�6��w |�� n����Z�۫l-nT�cG�'CY�n:&�j��^a%Hvw-m����}�}��=�*U�5g�9l��>�x���~��(�C�����TGD�CN�ddvٻum$���Ģ��>��׀>�� �V�u���Ƣ��irU�}�1���y-�+Ɂ���07d�L���������ɥ��<�Vۻuaꤻ��`{o�M�����Sr���`}$t�>���� ��p�d�����^�[�\��� ڮ9PB���Z��jɬ�s��5Je1v&�GL����0>�ꉀ}[��C�D�jG$� �3e���RF���<&�GL	9GJ��x�Y�p�32i`}�4V:�.QʩU�!(�(W������x87�E�)�.�faI^?��O	����0ޘ��D��L��*�E�-R*iUTݓ�}$t�7zc����	��&���S�͗��Du8���@�p�Ų��;I��k�kl�UrrKԂ5�w�07� ��o���A��t�������䦚 ҒX̚_�U$w�Vw޺��6_��H�:�P�MEQtUـs�����꡽������>镢��D���i9`}���s������$%*<��A%ԎD}��N |�iMIN.f����̼���ݐ`}��L���Ǩ5FQ8� c�M�#u'�D�ӷI��1mp�}:W�axs����ܹ�q|d��;���π�g��}��H���ݓ���=�T��H6ӄp�>���!G�Q�{ذ�BID�u���z`�Y��ȇBN�������X�4��Y�<XǾ���v�5�*��SWk���[�0��'�x�~���+)�Ph�I���d����[�zO�q���{l�2!�����w��׽��i4�� m�s��������[v��;k�+�T�q� V;q��wT%m���e+���tI���E�R;�ֺ|L;�H�v��ݚC������a�%;۵g;7`�rV��az2i�oI�N�,v�V�\r�P�-Y�mJ��a�K3؇5S�a������6;Sny�8���-�jma��-��՗�]8������}��`ը��$�/V�DV�"#�2A��CiyL�qṻ
$F��E]�����u�X9]s�.P=��`���D��6�r
��7n�	ݐ`ovA�6�	�U$R]+E��$�7�ʰ1f��̚Y�8�Vh�f�Ձ��I�4�)�Pڀ}��,	��L�GL[����U�t�ڒN�y��?s��}_�7���d���Xf�*Co����#r����������
q��iKg�ql ;��:3�WWw��0>�05oK`ovC��͞J�����cQ���M9*���mc���w��v���[ŞIDG�����J�q�� 5#�7ޟ���Ԭ�GL[��n�v�bŊ�e]�J"^U׿zg ��ذO:� �ɥ�}�+E)8�`�jH����t�ս-�����`U~����~�U��S7A5�.���/������UWa�80u�kb<���tl�f���M�����m��m��K�=�X��ֆ�J2�
E`w2i��Us�&����{����؈�U��M�)�r$'��~J��7n�����%�Ԥ�j#3v�' ���w����ȇBN�q+Ի���`{vx�;�4��\�/fߒ�6�����nF�H�NJ�;�4�?Us7o��nl�Vٻu`}׍	���Sl�5"�Z��']�ag�Ӕ�A��	��F�V�/oOe�Ź��,�`%x07� ���0>�{��3�<X�[�i����,�ȓ��~��!t��; �����H7璔�$Q�m�"Vw޺�;�4�;�4�3�5+ ��&���6�$r�=�Y�n�w&�a9�P@�`��_w��ܓ���o&]9�u�Eݫ�� �{l�<�>�ٟ���ŀsri`�k�#�6M�D����gk���&`Nhu��c�f9����t�2n�Ww�����0>�06vA��ɥ������t$�1��>͎�; �����$�I���hj7U#I�%X�,�&�w&�`}��V��YN:�1��$�a���L����w��%
�]������P�MDH7J1HXܚ� ԣ����;���>�m� �B�	~���������5UUT
�3,�2r�q��:7u����פ�z3;�,h'�,�Z �aԝ��Unv�a��:�Ѷ�`������c;۝�ۮ��@f���Y1��F�5�Zvvݺ̘���n݅�M��S�q����N�H�U!Uq�	 �ꃰ��b��Um�a�U�^D��'F�n�.�K��v�����2���A��e�z���7��{�w{��|��6:�v�!6�ѷNnLI,�f�!A�޹�<���nW�נ�5��*�%�};Θ; ��� ���0����g�[�&f��u�I��%�b}���i�~9"X���z�7ı,Ow��nӑ,K��}�I��%��r�5k���q&�I*G�|r��BX�{�ԉ��%�bw����9ı,��4��bX�'���6��bY�G+0�e8�JA$ڔ'�g)�%�߻���Kİ{�l�n%�bX��w��Kı;�oR&�X�r��܅n����$�1�E|��R9J%��{f�q,K�绿M�"X�%��{z�7ı,N���]�"X��#������!����"nݓ�{=KE����z�������Nx�sf��,j��\�Z4��bX�'=��m9ı,O{�ԉ��%�bw��z�9ı,{�4��bX�'�w�/!�a�Y1�njm9ı,O{�ԉ�E�����>Q�<�bX��nr�9ı,{�4��bX�'=��m9�k��R+��}Bm5 �)MH�8X�%���s��r%�bX>��i7ı,N{���r%�bX����q�r��G)gL�Jrpl���_	bX���Mı,K���6��������XB��j^Jl��x]�"X�%�a�K�g�5r�3W5�Ѥ�Kı9���iȖ%�a�G���ԉȖ%�b{���v��bX�(m�XB�������Nŗ%��O+��e��� ��|�}�\�z��Xd{/k��nzf^��wg���%�	֫��������X�'���ԉ��%�bw��z�9ı,{�4�NDȖ%���o��r"9H�#��/Zb�R�I6�'�g*ı,N���]�!��ș�����&�X�%���o��"�>��,Kwr���$)!wnV�t\���SS5�WiȖ%�`��٤�Kı9���iȖ4^"z�Ge"�bD���2[D��u���s��>~a#T1I=ݰO�!]&� F(����<�4*��0 1����4Gb&��3�5�����G9�8D���0�!�sDӦ���vj��0���0�wSH4T�kT��uՌ�8J @����)u�+>�Qx��v ��B(m_�C��8�8�W�b �t�k@�SQ>���z�7ı,O}��]�"X�%��;=rd�#�W^ﷸ��~����㺉���M�"X�%�����H��bX�'~��ӑ,K����I��%�b}����3Xh�&:-�M�"X�%��{z�7ı,?wܟ���%�`���f�q,K�绿M�"X�{���7C�r�|���ꔨ���C%ي�v.�ŵ�)����7�ج�7aD��L��˭H��bX�'~��nӑ,K����I��%�b}���a�I�L�bX��~ޤMı,K�����4f�2f�̳Y�v��bX���M�Ȋ!Q
H]ךd/�RB���w,!n%�bX�����ND�\��,K�i���a$Q�	ʳ��R9H�g��m9ı,O���D�Kı;�w�v��bX�{�M&�X�%����>cS�%"��p�W�)�z�U3����H��bX�'����iȖ%�`����n%�`x��
�T 	 ��D�Т�5�}ɴ�K��r�E��N4�m&�	��Y�G)D�;�w�v��bX��צ�q,K���ߦӑ,K��}�H��bS��W�Ws|���HT���RP�Dܚ{h���v'1����YxVٍ�;i�]��������.�R�ՙsY�~Nı,K����Mı,K�w~�ND�,K���"n%�bX�����ND�,K���f]fj��Y�5���n%�bX�{���r%�bX�﷩q,K���߭�r%�bX?{^�M��Aʙ����B�t��&j̅�
HRB�{��Kı;�w�v��bX��צ�q,K���ߦ��G�İg��M��$��Q�@�Y�G)�r�6��ӑ,K�����n%�bX�{���r%�bX�﷩q,KĽ���J!�1�mį���G)�W;�H��bX�'���6��bX�'���"n%�bX�����ND�,K�� h"�H����	��ֵ�k@j�gm�����D�ZWIm��]�5�49��Ѵ\(\�
i�u!�A�㶠��H��z��Ғn�hܫ�E���eq��ЮgR�v{3��H��z��8.�$��qճdN�lej7��ݗ=M�����5�/a��;�VF9�i�q��4a�k\h0��&���[@%�æ���uvu���򝂷�������'n��j��;�n�Ddض+i�+e�d�,�C@��9-�Rn)z&�9��Fۄ�|r��G)�ݽ�ND�,K��z�7ı,N���݇�}"X�}��I��%�b~����58�Q�)*7�|r��G)�緩q,K���߭�r%�bX?w^�Mı,K�w~�ND�,K��������a��}����ow�����9ı,��M&�X�P&
��?M��,K��oR%��r��G+��nҌ��MD4�_D�,�@�=��M&�X�%������Kı>﷩q,K���ߩ�������ow�=���2KJ驤�Kı>�w��Kİ�1�sR'"X�%�����r%�bX?w^�Mı,K�����-4e��4F�����z����M�`oNh���d�=��.��rk
]C5���a�-�M�"X�%��}�H��bX�'~��nӑ,K�����~ g"dK���o��r%�w�������ȑ���%m��{��2X�����rE$C ��_hϓDB��Ȗ}��&�X�%���~�ND�,K��z�7ı)�Y�[ĔC�c��#��9H�#����zi7ı,N{���r%�bX�w�ԉ��%�bw���iȖ%�g)�ӧ����A�NU��r��P�2'߽��iȖ%�bw߷�q,K���ߦӑ,K��u��KG)��1����IQ�_+㔎%����H��bX�������%�bX>��M&�X�%��w~�ND��oq����d�:��nn�.�W�m���	���i�;�CyLtա�3�knN�.3A�uf��m�R\ԉ��%�bw���iȖ%�`����n%�bX�����r%�bX�{�ԉ��%�b|wW�.�j�j\��nkZ�ND�,K�צ�q,K���ߦӑ,K����Z��bX�'���6��bX�'|k�4L�t��Hؤ��Y�G)�r��z_+㔄�,O������ r"�UdL��w~�ND�,K���I��%�b}����3Xh�2�Knjm9ı,O������%�b{���iȖ%�`����n%�`~I�?w��6��bY�7{�?���5vR�0{���{�����ߦӑ,K��=���ND�,K�}��iȖ%�b}�g�Mĳ�g��u�w���d�L�9�׺9��[�Lb�$U�x�dG6�r��(���#6�Lԙ�k56��bX�{�M&�X�%�﻿M�"X�%�����7ı,O}��m9ı,K{%��eֲMkWS3SI��%�b{���iȖ%�b}�g�Mı,K�w~�ND�,K�צ�q?S"X����g,˧5n�kWZչ��r%�bX����jn%�bX�����r%�bX=�4��bX�'���6��bX�'OK��0ɫ5��n�5"n%�bX�����r%�bX?{^�Mı,K��}�ND�,/��P��H�F��U�Q᠑.�}�q,K���_ߋ���Z�,ї5��ND�,K�����bX�'���6��bX�'���D�Kı9����Kı?)�e��I]k�6�Lѓ�ӵ1ɑ�Ζ�4��]Rm�2Y���ȷ]���WJ!��׻���K��;�ٴ�Kı=�oR&�X�%�ϵ�]�NDȖ%���zMı,K�����ְ�,�5.fk6��bX�'���D�Kı9����Kİ}�oI��%�bs>�iȐ[D�{=�e�,��̷PI���]� �~�&��'�s>�iȖ%�b}�g�Mı,K��_6�5����0�֮ӑ,K���ޓq,K��}�fӑ,K����Z��bX�'>�}v��bX�%�����2�FkWY�]kI��%�bs>�iȖ%�b}�g�Mı,K�k��ND�,K��zMı,K��cNAI����=׺ww��{�߿ɧ� U�_j�1-�[�<xƳaٖ��\ԣ�P��M��۲**u�+����.��:�A-��&܌�u�A$;e��������`�u!v:�+YNpnշA�W�u�/`�l5it�J�l98�ۦ�p�:�X��m�Mˈ�����;f���+S�m���� ��E��Ѱq�^�y�\:��� �c����!uW�(4r�c �w��mNv�����z�����ct����ŵÊ��$�:���5�s&@z���,��ֵnk:��bX�'������%�bs�w�iȖ%�`����n%�bX�ϻ��r%�bX����.5fk2ۆ��j��Kı9����Kİ~���7ı,Ng��m9ı,O������%�b{�73�њ�Z�.������Kİ~���7ı,Ng��m9��0ș��~�7ı,O��~�ND�,K�5��,˫��ֵ��.�t��bY�U��>�}�6��bX�'}��jn%�bX�g��m9ı,���Mı,K�����ְ�,�5.fk6��bX�'��z��Kı>ϻ��r%�bX?g}t��bX�'3�{6��bX�'�Q=;���
cU����F,�G��h�f#.c��@fJ��&'U����"F��:k5jr%�bX����m9ı,���Mı,K����ND�,K��=jn%�bX��z��蹭ML4fj�k6��bX���]&�`�F"b#0U��`�
0XC�?wq,L�����Kı=�oR&�X�%��}�fӑ,KĿS�%��e֌֮��Z�Mı,K����ND�,K���"n%�bX�g��m9ı,g}t�9H�#��W��o�58�Q�)"N;�}ĳ�"~��jD�Kı;����r%�bX>���7İ<�ȟk��m9ı,Oz_n�f]Y�̶椗5"n%�bX�g��m9ı,g}t��bX�'3�{6��bX�)��,!I
HRB�Q	=1��L�Wrnh�k�nn�Ka��e�.:�\)ƖJg��L��Ns�ٰ�6Y�{���7�����t��bX�'3�{6��bX�'���@�NDȖ%���fӑ.��ow����d�������,K����ND�,K��=jn%�bX�g��m9ı,�}�Mı,K��='!��Dɖj\��m9ı,O������%�b}�wٴ�K��q�*X1(Ud�1%0E��p<h��ؙ��f�q,K��{��iȖ%�`�/�L�\��Z&e�5��7ĳ�2'u�~ͧ"X�%�����Kı9�{ٴ�Kı>�֦�X��#�����)I�A�c�H���G*İ~���7ı,?��߳i�Kı;�g�Sq,K��>�iȆ��ow������y�S�Mn����
� ���8�������n�1�C���ז�F���e֮�q,K��}�fӑ,K����Z��bX�'��}�ND�,K�ﮓq,K��}}�2��[���֍[�ͧ"X�%��u��7�r&D�;����r%�bX=�~�Mı,K����ND��2%�����L3Z�sY��h��Mı,K��~ͧ"X�%��ﮓq,�dL��w���r%�bX���z�7ı,Og�a��FjL5s4e�k[ND�,K��]&�X�%����ͧ"X�%��u��7İ<�1vc>5��\!q�{y����$'�r�T��\��3.]j�7ı,Ng��m9ı,O������%�b_�ﵴ�Kİ~���7ı,Ow^�.f_L��2�-rme듭�z��᜴�ۨ6z�5���!������ɭ���&�����oq���X�wY�Sq,KĿ}�kiȖ%�`����~'"dK��;��m9�q���~g~��dH��gi����,K�Q	�wߵ��%�bX=�~�Mı,K��}�ND�,K��=jn'� eL�b_��6�5�����5�kiȖ%�`�=��7ı,Ng��m9��!�2'}��jn%�bX�������bX�%�'��<�]h�j�Yu���K��"}���m9ı,N�Y���Kı/>ﵴ�K��U�;�٤�Kı>����4�̚�֍[�ͧ"X�%��u��7ı,Kϻ�m9ı,�}�Mı,K��}�ND�,K� �7����� ��!I�bKG%��C��S�Z ��
A<�P�#���ޕHQ`a<h�Ձ0��$_!�
v$J��n�]B;ZP�0�
:��z�(��M��հ"@EB3| ta ��Ő0�Q�;�1���F� v4�H�h@��ؑ]�M��ee��G�N�. �C��8tC�
 j����! �0:�@=����??vݶ��Z巀           @  ������f�JƎ�v�"Ssfq��4�Ueeh�X�-��Tvz��"r��m:+���s�͓q��$芧e��E��5ʸ���ؤ�k�*�/Ul��+*��s��x6���j��yAW��vP#����1V�D��=���;��uF�m!��Ʒ�YvV���cĖGuc��u� ����;	�Ĕ�M�R���swV�yvڎ<���D������6rI���%j3֎^�Qv�;��[tF�b��b�� �3�Q�ln��iu��h�&��	L��M���J^����7e�k�9��{nR���6^�[��n��DId&I7��l;)p����!8�k,�jAv� �]��&��H����v����kS�6* hu��@ܲ�]nk�i6�]gU�l���"z�*,I63u,�x�!+m��3��U�J���i�<�ivv�'2��>�]�2Ӎd{���5�rV2S�n�.�R��v���ζ�4(!b��3����T-�e�
Y�	��Rj�ukd[���U!�s����[�l�2Oe�����͝6�v�pt`�sU�N�qMIm���ʑ�ݻT�Լ�N�3�#����9��́�9,P���+��)�5��^��+���\�Uc]��	�N�Se�L]�wc��(T6+�U�L���[�UA4X0V�<�QOV��@�m���S\�#�M�����8��@Իl��:B�@H+Q�^I؅�.�UDh�<<��z(�h��M�*d��ڒ�A��L�t�.ݣ�vV��K`^N�)��Wk�W�=�����!`�=n�&�Y� {!�YCHp��Ap�T� �g�ɴS��92�RA��Y�j�H�͛]"�dnyy�(\��,jU�1�t��"���:n�xΰ�#f�-[n�Pء�m:Ԃ�љ�`Q�ڠ� C\�C� Q4{^�8@4E�
@8�����o���ִ ��T�ݚձ�VA83i쬧dh����M���9+���W�뭍���\�p�KC��MR�8�֮������^nе&�β�� v5��L�g�����ӻu��rDL�YrkU��:��y�K.�Ӳ�����9!w��8���TH�R�й0m�w`�+��Y �w5x��<k[��m݊6�`����2;�5��R�$<nVt��Ȭ�ͱK[t��^u�� 0�h�f��N@�����{��7������bX����&�X�%����͇��L�bX�������%�#���"��)�ur��K�|r��G��f�q,K��>�iȖ%�b}�g�Mı,K��{[ND�+��{���������ʪ%���7���w߳iȖ%�b}�g�Mı�!�2%���kiȖ%�`�=��7��r������@l �q�+㔢X�'��z��Kı/>����Kİ~���7İ4��"Q;��;�|r��G)��P�ME��a�թ��%�b^}�kiȖ%�`����n%�bX�g��m9ı,O���r��#��R9_�fh�zt��H۶�Q��V�ř�{iJ$9C�<i����G�W*����%��6��V�r������n%�bX�g��m9ı,O�����9"X�%���kiȖ%��{��;�E߾���������D�>ϻ��r h���6�'"X��Y�Sq,Kļ�}��"X�%��w�I����L�bw���p��R�.�u�V�iȖ%�bw��֦�X�%�y����"X�%��w�I��%�b}�wٴ�Kı<z�tљur�-�5�թ��%�b^}�kiȖ%�`����n%�bX�g��m9ĢZ��^V������$-��V�j�f�d�0�ֵ��Kİ~���7ı,1����ͧ�,K����Z��bX�%������bX�'��3��2�b��ӌ�=�m�^-��$�ᩓ�8{k�j��\�nCO;���}�̑�^D���,K��{��m9ı,O������%�b^}�ka�O�dK��{��Vr��G)����¢��|9ı,O������%�b^}�kiȖ%�`����n%�bX�g��m>9H�#��VݡƓq�q�q.V�X�%�y����"X�%��w�I��=��Ɛ*> }��w���Kı=�g�Mı,K��{%�٣5��4fI�ֶ��bY� H����Kı;����r%�bX�wY�Sq,K��]D�}����"X�{��?x��D�﨧SIE��{��2X�g��m9ı,O������%�b^}�kiȖ%�`����n%�cH�-�@���"��5)*��]p�Nn5և�ez�#�v�[�v��_��������u�����'�,K�ﵟ�Mı,K�����bX���]�NDȖ%����fӑ,K��~��lӭ��m�B�jn%�bX������? �r&D�{��t��bX�'s���ND�,K��=jn'�eL�bwڇ��N�b��I%�9H�#���=��n%�bX�w]��r%�bX�wY�Sq,Kļｭ�"X�%��Mz��U�J/w��oq�������m9ı,O������%�b^w��ӑ,K��:/��h&�T-J�(�sf�a
HRB�����]�3$5nf�ӑ,K����Z��bX�%�}�m9ı,���Mı,K�뾻ND�,K�}���(��\�gRU͹�hI3eu�,=s�$;cզn�G��`��4��e��w��o%�y�{[ND�,K��f�q,K��}�M�"X�%��u��7�G)����	D99M�r_+㔎%�~�I�r&D�?{��M�"X�%��k?Z��bX�%�}�m9����[�oq���]��QN��M��%�bX�����iȖ%�b}�g�Mı,K�����bX����&�)�r����#d�J������ı,O������%�b^w��ӑ,K��w٤�K��Y�;����7���{����������<n�bX�%�}�m9ı,?3���ND�,K�׿]�"X�%��u�����Y��g�w{���7� ��]�{bn81����r���ʥ�ۉ�e�&۝p�w]ѺpB��cHl@��4v��E�u1��L=��y��`��J&����9���\�v�K�b���5�Cq�@������"�8C�!�{]�cit�*�f쫏�|_�n���f�!�F�YI����l�)�N�5Z ����)�SuSvTL�cv��0��֍�^��������o���u�2�h�{#���p�Z[�<Pu׌tVـ��Ӯ{v:E��5Ͷ̙���Z�S�,K��{�i7ı,O����9ı,O������%�b^w��ӑ,K�尿tZkFjK��˗Z�Mı,K�뾻ND�,K��=jn%�bX������Kİ~���7�2�D�=��O�d&j虒�3WiȖ%�bw��֦�X�%�y�{[ND�,K�ﮓq,K����ӑ,K����,��H�ĹVr��G)��n��|%�bX?g}t��bX�'��}v��bX�'��z��Kı/��Y-�r�l#��_�r��Eqw5�U�,K����ӑ,K����Z��bX�%�}�m9ı,O�9���nz�IY�u��Ar4i�`��­Z+�q��x���D���8�s��H�L����bX�'}�~�ND�,K��=jn%�bX������!��5İ�{�XB�����{��*�ɺ���W���ND�,K��=jn���+d�T

�h
"���'"X�|ߵ��Kİo��i7ı,O����9ı,O>�ݺ,֍j�m�\թ��%�b^w��ӑ,K��w٤�K�Oঢj'�k���r%�bX�����7ı,O���Y�5&jf[�3Zֶ��bX����&�X�%��u�]�"X�%��u��7ı,K����r%�bX��׮�Mh�I���Y��i7ı,O����9ı,?﷟�ND�,K��ߵ��Kİ~���7ı,N���g2Ƒ�G2]�uyy�h��M�8��5��<�ɖ{WJgN�'6vb�v�&>�r%�bX�wY�Sq,Kļｭ�"X�%��w�I��%�b}�w�iÔ�R9H�a[�Z#n1A�G�\Kı/;�ki�~�DȖs߮�q,K����iȖ%�b{�ޤK9H�#��R��QA��r_D�,K��]&�X�%��u�]�"X�'M�E��A� B*
sG�,L���D�Kı/����|r��G)��U�l7�)$�=k4��bY�@ȟw�ﶜ�bX�'}��jn%�bX���m9ı,�j��9H�#��W�f���B6H��ֵ��Kı>�֦�X�%�~���ӑ,K��w٤�Kı9����|r��G)νA��n@
r�J�v9���Wc��v)���y�W�c���c�r1�㬏�=U�R$N�Rq9�|r��G)�y�ͧ"X�%�~�I��%�bs�{�ND�,K��=jn%�bX�d��!Ӏ��Q���+㔎R9H�.��� ��I�����A;��֡"�'9�t���+�S"X��5?h�֌ԙ�re˭]&�X�%��~�ӑ,K����Z��bX�'��}�ND�,K�ﮓq,K��;��W3WRfI�e�m9ĳ�5߹�֦�X�%������r%�bX?g}t��bX d H	<P���D���ӑ,K��;�Z#n1A�G�Y�G)�r����9ı,���Mı,K�����"X�%��u��7ı,K�{ڰ6�Ol��;��X�:Dt�\p�M��`Ȏu�\lS�i��?��8�.֬�S��%�bX=�~�Mı,KｿM�"X�%��u��?�"dK��w���w�{��7�����2���)�R��n%�bX�}�p�r%�bX�wY�Sq,K��>��iȖ%�`߻윫9_��S9H�wM����B6H���ӑ,K�ﵟ�Mı,K���ͧ"X�%�~�I��%�b}���iȖ%�bx����r��Wn��֭Mı,�A���ٴ�Kİo}�4��bX�%������bX�ȝ������%�bt�?�Y�5&jf[��5��r%�bX7��4��bX�%������bX�'��z��Kı>ϻ��r%�bX�TO������kZ��$�J�<��SC3��ܣ���o4�F�y��2�onW��y
����]��zp���њe����v�k(=�fܨG�̇wi��5�O+<Cs���'9�.����B�+A�`��&�鶔�X{
��=�W �e�)N2��2۝�Ӕ�-��v�n�l�n]�m�O(�*U���;j�*S�<�-�;]H\�UT �T�n�ܚ�MV�Z;�Nw;�ڼ��+���Zx�X�]Dv����*�v�R6m��&i�����ou�{���ӑ,K����Z��bX�'��}���L�bX7���Mı�G+�^�2��Ȫ4�W�)�����Z��bX�'��}�ND�,K��f�q,K�����"X��#��n�h�8��AK�g)���>�iȖ%�`����n%��򚉨�����"X�%�����Sq�r��G)osX�)I�BA����_	bX���]&�X��{f�w;�]�v�Z�l7�)#����v:`}�"`jޖ�ݾ�����e�U�s�=�cZ8}l6�ۧ��FVϧ��"9�9��Y�����syĔWI]����?��V����L�GL������f[��3Z��}~�
Ў���\P�_%]u�η� ����d�[�y�Ҍ���{�`}�۫<�q���ś�`f�V�� N���e0�-�{�`o_�����7z:`w^���C�P�!IV�{����K`n�t��dt��WzS�"�Z�yY4��tb��wLk���Z��=�=H��u\ؓm�tDF�b�N �/�ś�`n�t��dt��nD�&��HYi^afawif[w���#��r&������F4ےU��wn�Iϳ޻�5�B� l ���(���R���RZKb \��=�����R(�b�bH0	���O/�(�]�@(� A#�,H<!$H��XJ Kg>B��!�B"}g��g�@�@	�Ӏ�9
�f	�c♇�D;���8��m�447�I� �Gh��|K�bFl6�Y��0�`��`�AZp��T����1x���z, '�";��;�ܓ�w�7�����NrD�R'ԕ`w������GL�GL�����v�^~/105oK`n�t��dt��nDͿ���_�:C��n-����Ԙ�ZC$f懫5i`Ӝ�;\˞�''��6͔2��-�������V��h�V�� N�8�Xwv����D�ս-����e��E��.�,�`}�"`jޖ�仧�07��O�Us�����R�F�b�N �+���B��^�޽ŀ}��`R���|뾵`�^�
4��$iH��6����}_�~�`jޖ��dE�ˬ��fա�qn�ǜ�����n�j"��8��`��l���Y�P�8�	N7��I+�;����V���GL�.��W�����j˩�Xܦ�?BJ!~�T9{���b�>�x��&F�ܙ�(�.�n��L]=lގ��&0>ۑ06�su�Ҍ���*�f��罌��L[����H�/ WV���>�1������]=lގ����X! :�Z������ �ʹ�IQwvĲȕ»�.�1�F�X�r�0c�������WE�6��M���G!�]��!�xm���&;l-�t�ܰ�
č��1�
�tgN��ܚ&o��>�[�2�k�h�Cn���r�b��a��Ȳ\�c�ذ�����U��y�R��9���ε����ӗ�v�M��B���2�s����I��m�{��bM�?e���u����Ym��랩��"�A��	z�^���7k�9E6P�:p�ӓ �?j�:����6��U���K=�ԭ���2��L[���0>�0>ۑ0���(�r�m�#�;�۫����܉��z[�:+��̻̻Wu7v�?D(IO;���9�ݜ�κ�;�۫.��Ӝ��H��5%X���V���GL�GL�+.a����.�ͺ��#���nͱj�sj%�Yl���n+A���D΍J{4}��'�u�s�x���-�I(��9�ݜ�o=�Jp`�v{�uwK�9T��7���޾���z[�tH$^�'Lr������g�ıf������B�(qJ:���˹=������7z:`�cd%&����aj̣/V�lގ�����uz�A�<!?(��H�P�a=1Ыtb�Ὂ�T18�=�u%�ں��sBR����m)�����;�۫��`uwu�#r��0�#r9MI%X�:~�������{�������#a�ç9��r�ԕ`w����!ب�(ł(P��LZ'ɕ�K[~��7}�Vf���#iG?��z�.�����<遻#��r&io7Q)�plQ����mՁ��t��nD�ղ[�U8�Ag�+e>z�9,ϴ��\��6)9�d�w���q�����N��t�I �0q���z���nD�ղ[w����v��WXRY���nD���9w�l��L�۫�8����V�یPi���1g�lގ��K��t�޿y0"��ڥ�NB��v�������z������W�C!D+X�+ 䏩���˼�ʵ��L�0>ۑ05l�����Xf [
� �%9R��T8�����}���R��}D:�#�t�w=3��g��+W��]�|��Ɂ�d��GL��Ձ��m�I�T���Ȭǚ��0>�:`}�"`m.��,�x]�/�Lގ�I3��-���u�0�:`�`l���nD���U.�敏�\�U�r�#m�`}׺�UV��/������'=�krN {���� A �`�PG�$�����kZֵ��ݹ˧��m�1nܹ3���769�h��v`��;Ua���ծr =zQ꽁��\3؝�sl��..%۶�)��+���{��Q	��G��+��ѓ���W�Qn#��Gk�q�WF�V���HE]��P��c �v�n�g�2*N�6�SíصV���1N����%k���tP�tf3*�t�7{���s?'�=��Z��i�nc���Hn����0R��v�닧i�N\��DF�b�L�G�ߦ��s��f�����ԒQ�;[��9�s�)�SWd$�HX�m�����,������K���W7+x�	R7#�ӒU�t�uȘ&A������t��i��SnK�{���٥��ͺ���`w5m���T���Ĝ���2I1��\���H���V��Ɖ��=nL��FȩԭgK�H�����;n��v��ͳe	���ott�:I���L� ��XM:a#�`|�u�U�|��W�ʡ�D��2�$z_�v�SMM8�������K��u`r�[�"$�Ņ�2��L��s�x��n�6"'��g s��hJ19'!`w3n�7vXc�Vn�,qn��a������%×E���El)6��F�<a���ZGk��v�y)EJ�9"���� �{����3vi��͕ ��t�S�b�INnF˹`ݜ06tt�:I��F�C	#i:�5#�3vi`w3n���Eb*@@dA�U"g���M����䝾��p;K9��dC�iF��X�۫ ��x���TDO5��S�RU�`'LJI*����`{�]{�?��x�;��V٩h�ND�T�D��R��ѣe��X^hY̎gg�M�)���t���y��(l �q�,�vۓK��u`b�k�3t�XF�b�L����rA�������ˤ��ԑ�^��br$	����]X����n��ɥ��77�J*TI�A�$��κ�>��X϶�
P�$�J%$�9_W+�1�Ձ�����rJ��n;��[wd�0"�-�6���Lq����6[x)��#��L��W8��V��2#G"9�c[T��Kwd�0"�/�_ �=�`uFV�Q��M���f�X����n�s&�iY6�>4I2�l���t������0>��@����DN;�����ɥ��2�K`}!�.�,XZ�+�'vA��2�K`j�-���:$p|PK�S�� 6���B0�aH@a��6)я�,'@�
v�@3J�����ba���$ ��T�lT~3�F)6�T�A$7�=޸�>���!zU��'��v�?W�!�Db��2Dc�Y"�!�*�l��hE��l���H�r��HI��3f�J��z8l��}�x};�nfgu���� �>             H I�ԑ���RF�5Z�ɄK�s���Rrv�ÑW5lі�b8��v]a�ص�.7Dַ �R�P�Y�,��Ĩ�dm���-si{DN���d�J�%��6��>a�}�����m�cb��m�@��J�dv�����-%���䃛�%��lE��[���4��VZ�nL��QmD�v�F'o"�%�ʐH	��nV�d��@82�J��rs�*�;#����۳���ڛ�����m��N�:���ﯤĺ��1��hI7k;ka�P�\����v�ڗꪡ[�m�v�]�n����M�-��d7L�8�60�\�H$�Mf݌��ʩ
&:9v��KՂYIKi�Y2\��Ȼ�F���UvrԦrYժ�r��;\7=��9nCL����]Ӗ�n���	��CT���i���ö�D.}uGn�-q���Y"�UPt�G�v�cm�v=A�g����1��Yn��;4����"���2Bv-�m*M���`�b,�a��Ћ���t�.U�ԯl��zD圵��UREh��*��'P
@&U�jU�1�z�v��:�ذ=�+s�ɴt%�.[ڞU�^.�)eӷ�8�v�ԁv��۔�s���l���݅z\��!!�u,�gi�yWjwLvJ�F�ꐷKb�eH�� �i�R�&�N�i���ifs�خۖ��8[��7۪��WM�g���vx�ջv}���LR7	��Z�Ga.���qW]���U{&2�]"f��b�����c/�[�=�ٜ�컟�\q�o��+On\��d�R����$.�;X��yMۉ -�;���D�c�L���Ih6$桴�-ΐq��F��8�P3�:@�pM�˧aı�[['Q��ɩ�l���W^`���c�*V%bA��Z��*�[2����L�������HuU��m{��Ͽ;��_�*��|	�EBb||�U����F��4ؼO{ݻ�߿~��������  [V��:v���C�ó�6���8-L���$Q�8k��A�ĜE�3�@u2��m֍�&:[V̀a�+ԙ
��X��6��c�N�8�Ƹ��uayX֣��Z��eXNێleZ�Ӷ�zh�RI,K U6�/E&sNs@����2Sd�m�e$Ƹ��n��ٹ�lZu<놙-O1n;K������r�~�o�wu�x���]v+�l��h�p���j6T�x.1�&�Ȏcb�9��:w�a��X���v���&Ɍ[%�&d����ĥ*$䊚���7����d���07fA�u��^~�G$�������72ig�K3�Ł��3����!����v�d� ��d����]etK,�^ie�w�{��[%�>]%�72i`jĳB7���������t��t�:k��*�d�/j#���v�����j��e^ ��K32�l���t����s6���2jN��� �q�.�ٿ��D0\B0��6�QB"d%=�R�����q�q`�w���9�RF�Ǒaq�2TN;۳�{��6L`|�K`{��(�e%�H1'��Wg�ŀ{=�`uwu�y{v�XF{���D�����M��KaݐƒKv8}�Io����V��h��V����C9v���r�ч���S�7\9#7Ol	�X5oRn���$��Y�5}�I�Ii$�ݽ=��z�Ig�%���=����A)�$��4��q��g���$�Y�9i$���������^笈�pi�Mȭ$�{߸s��/��kv�:�� D�ON?�f�}�I/z<I-�R�2�+��J��Kwd��]��_|��^���K��}_|�[�-`8�4�ԒZV߾�}y�mꂹ�f�7m��{�9�m�sd��Y�W����F�JS�N���w`��u�J@�6z&G%�lj��d���[J�ddq}�I-͸ZI/���}�I%��ZI.�f��I-OM�%)9
B�I%�w~���q����KI%׾���[�p��_3sx�
�ri�+�I)�1����K��S����ݎ|�K����9#EI%�Ii$�����$���-$�����O�N�����}����K���HJd�D�r����Inm��I}�>��I!N��$���/�Kl����C\[���H+f�b�t�r�I����̹���ꀌ��j�	%�t���$�:^4�__t��I%:<I,�K�L���1�$��I!nk��P.e�g��9�m����7m���s���m�N��� ڒKI%�����%�1���~�Ww�{�����ƒK�">یPi�����If�-$�����HY�夒��k��KФ�'!fWw�4�_lp��Ix�Im�K��mｭ�v�|!D�����y�Zրm�m�\xٖs��I8GY�p���n��0�ew!��Om��ķ$�}�u�	��Y4��!)q��n�����Τݭ;��__B[V�U�k*��Vܳ`�]�n��Z��"Rlv�%VcN�c��p�v��2��j��9���h��5�U�cT»��(uӨ㶽�\��ն3l���,���ɳ��4ZIIH5�_�����.��֛��T��v�r4N�Z���}���Ի���[w[=��k��` o�]se����c����o�%��/�JH�4�_lp��:,�Uk�Q�E%r9i!u�5��In�-$�����I-ݒ��)��痾p����%A��$���tZI/����$�[�%����k���-��ID84ێF�$��>�$�$�i$�����K߿~��{���K|x�Rd��$�6���$)%�I%��/�K��CI%���I.����'��y�l�v}e���z�����]�Cg��v�!M�� ��{3r&���ƒKoz_�$��$��>�$���ZI/�u%�F�b�L���Kr6���W�W߿~廩k����$)=x�Iu�5��I�))I�@R�i8�K�|�B�/_�����z��$�<�4�]y��6*$�8���}�B[��[����`}� �4�Wuk���Y��
�-��z[ӣ�����,;�7�F'$pm(�"�h�b���TӲ��؏!7ca�9f↨cs�%ie��W�������[���U�s���^���pi�RB���x`N��ս-���B)Y%8	:cM�Xۛ,��*�9\;��B `��"� s*$1P"A1#a�=0 �dcGZ��XfM,ݚ�����DR;V��odl�0�����7��J�6�d��vw&��٥��-��z[��E�<��H��*BN:a�֎Z͋3�튺a�����{6�M�u����r�J�i����4�>Y����Ur�A��Ł�}�I��Q')ř���t���l��0>ِ`f�7�J&�9��vWs]���K�����n�3sm��d�D�wb����J[y����6��_�,H��#�h�'�|���}��nI�߸�i%��n9���vi`n�9<���ـzI6=��雋�R��y�i[p<��	�e,77&�-���I,���u��1ĥ&INN�$��[�v��l���GL�4WE��f*�Y��ս-��vA�����}����{�+یPi�������#�m�L[����E%��®�Vaj�`}�0;o�`|�Ka��\���m��:�����D���I*���ꪪ��z��3�w�����@�!�Jk��3��� �m�*�Z�;8ڇ89�ӈ!26�鋮#ړc�kV���q:Y�ťn�Ӂ6���Ee��[�krf��7��o?-N2^8���'�hT�_b7�6\n�\Xɯ5�_��8\l�vs������N'ed��ڑ��� j��pU�a{-l.�d�aۃ��8�1�'%\���c-ShN�`"�H�A?sտ�W{ޢ�d%(85R�EOZ�fVc���}|p}�������a�\3��M̱�M�R�2H1Ȱ/���������sn���U|������{�ܦTmJMG!I^[oGL���ގ�-�l�im��C�M��U��sn��m��-�7��B�R���x	_륗��ߪ��{�`j��`M�釖��������t�q�S�U���k�7::`}�0&���nKP�3.��.�lV4�7�*�����X�<���n]=���Щ@����%E#�͕ ���Vْ���;�%)9
��K�n��󮳑	v!|�Gc��w �{�`w��V�7U$�Q')�$��ݑ��[vGL[���7�J&�9L�U����;�۫�����wn��vӔʑ����%#�7dt���]}=��:`|�K`l�R~q��Ӊ�$�XI�����݂6���Y��	]�_����N��#6EgSSV��oGL��~��_����L�z�INO�����۫I.�l�GL[��RGt��ux,��.�ʺ��rz�`>�X;��b��]���I�:� �R
Ȳ �>@O
�D]��Ӱ؁�B���d�H�>5�1�%	�@��]�R�@��*P��&m��abB�J"��X`�
p#WA�@y ��'�Q&� hLҥGL4 q~HA�m"ҤcK�a�֜!�a ��%�h���`���� @�B@�� �"�C[SeAk��Q(0J*�)z��G�F�H���� `�� "��}8i' ǅ�B,��x�T�P���d�5!��C��ҧȽ�"|��|�!W�#�3�"y:�'C��>@�=�)�tl��x?���Z�>����DD$����ذ�z�.�U�VT�j殰6"y�~Xg�k �:�`j���]y�;V��)(�!N����V��oGL��l�GL�Z7��έպN���-��բ����\�weA�.ݯMizZ�М��9n{(��Hw�x������ű	B�C�׵�7ǩ�|��rS���X.����05oK`n�t����ʲ�-b���RY��ݑ�V��쎘-��f�m��C�M�ڎU����`w��~D���߳rpR��4�"�؅P��O���=��Iv��f��/2��:`|�K`l�遫z[6�{�����=]��I"k����b��D�LűN⋤���y -�M)�g�Ȫ.U]Z�Owk ��ŀry�[��7=�=^�Y���%D�:��f���׵�>���>�7Y�#�o����:R�b��Y�v�v���wu���V�0�N��r�"���`M���[wGL[��f�7ͥ9)�Dr��w]���u`ry�X�x�
_-�����|��n���ջ�n�T����o	�nކ[74�
�t�f��K���l�� D!�
j� l�L<��Ԧ�<��y�i����il�H���us^ή��;�f����d펰�ⶫ��o����9ó���3��� ����t[���%ŕh��i��͎�eE�[-�\�E�]�`t-�Ƚq������a5��Y��0���浔�P�EW�X����f����Q�q�u�f�
v�s��5WV���n@:Z༂����'q��Ԑ�[����~ŀry�X�x�G�������$�m�#r���{�u�}<n�μY�B�2nѺJ��U�W��/2���L��l	�05nk�7t�'N
7(l��r��w]�;����l	�:`l��wW�^���yl	�05oK`M��廮��ٱ�:��8�U)��)<�e�-��-ud��&��mқ�D�7L�um���],Ff,����'tt��l����u`|�
��Q'*E�#�7��o�W�ء�*���^s��'�{_��uw5����Ӥ��QSpr�����z�fA��z[wGL		ٕefZe��e�'tt�ս-�6GV˻���9U�︽���n9���z�dt��l������UU����Ѕ!願��G��.x�8t6��U�+I�i#���v��������˯3+�=���d��0&�4N�nP�8�X.�z�SV��U~�Tʐ�w��¦�W5u�|��9μXbR�����BP�,Q
�TBQ_n�ذ�n���ݢ�#��J"H���sn��۫���`j��`|�
��Q'*EǙl	::`|�K`E$���l���ږ��WtxX�#�֔�v4k�n��ϊ���8P.n�����]'%��9L��l�K`jޖ�����m�r�Q�)�%#�5nk�:����۫���`gw�ؑ��n8��`jޖ�����d�S��$�tT�)�I�r;w6���wu���r|S@@x��U?
��1�I%��ok m��iU�uV���Uլ��u�yB��og�;={X}y�m����`ߗLu<Rs��\H��5l�2S���l�L�ՓU7�\�ܻZV����yl	.D�ս-�$���]�;V��)"9
t�$�8�����`O��nsaDL���٤+V��"�c����u`|����r����XY�v�մR|ڍSPr��D$�"y]{X�n����ŀ=ն��db�HSN;u����`n��X.���]��U�4��$��� ��3�:e��XF#���A���P6������V#���s{v�7^2[<se��Fڠ���'h�C �Ѩ;Gl�ev-iv�:[�Q�ۦ�b���g��u�v[Yg��E�+ �c��cxʗl�r��Xaͣ��7�))�T:�,�N��yf�t�]T��b�m�n���'E+n0n^�Z����ßS�O&��6k�T��@��qG�>���K�����n�<�MMUd��!�dgQժ��	4S�vn�]p({VȬ٣�m�?���o������c�T�S���c�U��{�V˹���{�����V�*h�8%�0��U��ޖ���L����:`l��SIYiaj�Y����L����:`|���Xf�ID�*R���8�����:`|���$�.���}�k5&�r4ND����>�晱K��z��ϡ:�=1qvHoO>��--]��~��Θ-�l	.D��z:`j"�R��5�L�f�5�7$�����tP����x�G@$QQ����g��������ͺ�7um�r����j��_D��z:`I���-�����!���pn+���X��L����"`IgAR3*���e�e0$���-�%ȘoGL�UW��h�t�� ���T�G;p,�q J��l����uײ%clr��͇�ݕ����WO[K�0>ގ�H遲�P�+-,-Y��2�\����t��GL���.:QIb�²�����\�s� �x���Ӆ
�%�
�V "ql���f����]�>�µ��Q'*E�p�7wn��s]���U��ri`u�*O����r�/)��ޖ���L��	$t��������߽kFa�5��\q�#RNɂ/i�Z�6�s�[/Y�pݻJY:9�y�t�e%y�_��odH��ޖ���6ƈ��q�Ȭ��K�s���$���-�%ȘY�T�ʼ	������o���!D%2�;V�ɥ��ʚ'N	G(T�9V�κ��� ���`M�B��!$BQ�oBDGP���
�
9\�r����V�ǩU��҃L�JL`Ir&���:`oL`T���;?�s��G�x��6״�͖҃v�]	0����\�WM���bd����W1[�o\�`I#����|�޿y09M+Ο%D��B6�V��Հ}��`n��`}ך��7i�|�F����0��0$���$��E-2q�#�1	�a��OyX��+I0ޘ��D�-������y���܉�~��� ���;��0?¨_��_� 
���Z �*����� 
��@_�QE?�TA$@@��E c�P DP,Q@D � �*�� �*�����@U��*�
� 
���(
�� �*����� 
���(
�� �*� �*��b��L���{�� � �����!����B| @��ƃ
 @P� :T+E( ��Z�o��   9A(((P�%U�J�((HB�ڈ��Ռְ�l�T�����P>| � 
=��FAB��J�y���}kۀ�����4$���mo�݁������bY{�=^����0��=����4� ��v:���/7�P�ѐ��N�h
 )�B�����5`6��A���ßx����tr{����m�nǯ�H��A���կm�;��n�m`���/�QE��B��C����/�4Р>=�i��\`v����>��^�-�G@�op<�	!��ެ;��}�:�$��6�����7`4>�`���_<
�������>�`hz���s�/���h
����=WwS�[����|#_}�@�wt
}�<w�
ť�U����n���=5��R�ž�9tY��[���Tx> ��(�>���&�Z��� 3j݁l�*��	*�n��`��p6�Ka�}Q��`����n�	>�=�F�:�`���m���;��݆����RB�  R  0�JR�S�h044ɠ1���R��Ҟ�h�    تT�iOT�4      ���@���M 1#&�2@ ��H��Bbi6����h�S�!��)T�0 � �����|L|��}9�s���������P�6��F}�T)�H�}T)��BP�����[_�de���T�1�9[~�-�P�Y+�s�b�
e����X��-|_/�}}[������������������������wwww�����������������o��{������������������{����{wwwwwws3333wwwwwwwwwwwwwwww3��fe�f���������������ټ����������������������������������������������������������������������������s���������������������������������ffffn�����{�������������������������������������������������������������������������������������������<��<��<��=�YTOY��+�Q^�����S�����d#���z�^���z��X�	� �`^��	OY%�	�^���)^�����YIz���}�Њ}(�@���*��ң��� /�}*?D���z�OYT�Y�*K�Q=`=b/XG��z�*����J�X���=eQ�z��Y%z�C�A� ����W��E�=�n���fM����D������y��z6f!�+��:�,�֏;����N���:�ug%�']gQ��������};���a�-�O�&v��x�a��K����Hh�:+�q�/��Oz���A�q�z`��F�w�GD0�a���u��Rw��!	�K���:�(� �
�z�.A`՚
��X�K3�']��r�R*r�t:���	�T> �.��v���[��bށШ]��d
TX48��������ѥA�j�$�޵�/"޷a��1�#<.ι�O.��ލ���P���@H���A�C+�'(����� ���� ��E�SZ��W<�'=������ֈ8&h�#;#�'��������۽w��8g��$�$�aPN$8��bF�Q�Z�3�	����0��E1@HB��\8Y��N@x�lYLa��h�:$�N�5����|���d�i�s����];����5Le�ބxaw�Q�t`�֢l4d�4w=�t��IŌJ)�(J�;<lߝ{���4��/Bkt=�X��I������3C�p��o��l�f��	�g8fNz��I8YZ�2 ��m:�0�)�aM:�s�q��u$�Nh�p�tлn9a�g�Ƃ�R���ZBI���!"B!�
�5XVdy�לń�l�$8$&,��&��Nc�s�,�j�L"t�vsFaI��H�F�(��c4��l��:$����7I34�3AK#	3�v�l�u|�'��ׄ4+��y��eͮ��c�Ņ��q�,&,d����{;[����;8���YM�������޺�p���u8K`3\ B�a��,2�д�z��	`��AI�
��0�09I�a�d�}x`��q�Q�����OK��`�E�8f�ݫ3��dA��h�ވ�0;[ǚc0+F:�l���CLc&1���FfLR�aui�0�&	R�6���L	6I�D4�$KF,�΂
2�X��Ĝ,v��RA���cK����,8h��9OgD�DE@F��7����S;xy�K�Z�#X�y�ai�`t�@@�˅�����6���]�l��9�#ck��y�dӤ��Ĳ�NI�c	���C�F͜5��I\�Q��j�h78��8\��N��0� ��h�AkV��!������&���d�x��=	���#;�c��3EXe�VL����� 2I0���$4I���2J��3��r��a�Z�5�G��l�oηI�4�	�(����&�x,�G\�!$6�a�z���ltA�$h*n!+)ZsA�k�0Ұ�F��1��6����tn<����4����a��1F��#��XSjѬ�:�7�.��Ef�I���� � ��c]9�����sٶ�{�d
���G<�f��ò7�o�k�±�j����]�³3ABaL��Ƶ��:칪M�c	�t�ދ4��M(v�3��hq6TXh�p�������E�W�����A�E$����5&�Û{<��h�Sp������N[���z�;C���.���z�5�%o���A�9�1��0�o��&��ܖ�j�8@�ҠiX쳆���]����zFD������;�Zי��᳢d��	�a���|�9�a���m��	 �㢸(V^t`�2���M��R��̄�2u�\�l�D+�c &#5hԘRJ��3F ��	p���_��`�`�X$ȩ��#l�4l�a,�΂�#[����H�#,�h�,���.yΘ�")�M8ʓ�!�N$Ac�$�F�ǝmގ�w���.���	ł	q#'#0)�	b0�
1l$��2(��	� 0#4�������1�F�7ˎ�	��<u�Nt��iq�'D* ����Kut�o)�;��A�T0^ز89����*��|��;��� �i��w�w��o4�Ͷ	 3GRh*\*�qwL�K�T�BG	��Y��cF���+G�s)<=NH�L���M��ĪtE�Ԥ&�B�}�E:����ã��:D���q��1&p$ �x�+�d�	pcL L�0�b�a�S����S{��';�4��!��U����xK�r��b^bK	A���}�Kz�RnG��^s�[p���r�'L5T&D�yVh�&E�F1�a�5�s5kF����ͅ���q��1��0��H��#%�:cã��9��F"���}�TZ7Vk��dJ�n�p�K�YxJ�2E"a��G���f>�f0z����n2�p��%BV[�� �p�	a�.wa��fp��|v@Ǧv0D��d������ ���$(FX`��&@��0���p���P��C#1#�U��V֍..�6%�Y1aF���25dDV8f�G5�LN[�:ٌ��Z0'1�,����f�t8M�d�0���Y�Kt`�a��f��	2�P=굧������5���mHZ�&�U8xR<I��q8�b@�t>��ϋ�.u�B��p��d�� �z��h	z������ѵm7O}8
.�X�z�0��]-"�5��|�(�u4軮��k6%�wua��
<es�����n���g1&�m��K����9��}�Iq��.�nuuɋ:�����&��!�ڲŔ�2�)�]|�E4SMl���ޅ�ajZ�%~v��Ծ����wv�����4�'o���u	�I	�����1sQ�:�p���|�@��iȰ�������g�����������~�����I�����ÿ�;����        @-�  �  m-� ����  ~�z                                                                             =@                                                x���۶��j����Ug:F�@-�nB��U����]b"J�F����"���wHH年�n� 4V��%��	�[g��]�m�b�k�v*�8���Z;0�i�P���U��J�J��!I���]m��[pI���*�U��Z���3��n��-���[[I���tͶ6݁Ŧ�m *�TUPs�����5�� -�h[@6� J�  �pm�ݻ`�iת1V5��	����XתN   h�k[��EЛcm�� �W܀�WU�W�  ��V�lH
P$-�6�m�l  �N�!���LH  [vZ G-���5�wN�-��	6��i^ٕ� ��WH� '@8	��q��!�$ 	 ��   �b�Ӷԭ���� h��kt��	Ij�� *�
��=  [$�66�@�m��I)Sn�	 -�ݻ%K�̵��I�;gH�`֊�)�,�UJJ�P[U�-��*�=���S��I��4�G[m6 �6��v�ko\�-����H�T�3�V���a���b�< �g��D��k�vk�i8��M���-s�m���Mv�76��uV�ڶ I[ ʹ�,��r�4��l5U*�E�c�	����L5*��+���YnZְl���B���JK*�MYF��j ���7l;7Pq�;$��X�.��$�w�_|v��WIq�e`ٽ[m� �-l���k` ��8��[8��țŹh)l�%�%�v��;v���F,[[�h���������m]T�'/Z6���f��Kn���[ +UJ���Jiy&-��qm-���m��I��i� m� �{��6�\�[pr�u-[J�\�A�@ ��j�h�om�+m�m�$m�9bl��-�9�� $  v���  m  �UU@�;UuJB�<l�   �`�a H�͔�]k�-���N�zY����  �`5����-�����U`%�����T���1�A�,G*���l]4�g   :@R��I��n�m�� �kv���)V���� �mm�*ڐ�mUb�r�.�
|sU8�h��$��N:��;��2Xr�m�*���c�UҒ�����]�m����������	,���;`�I|�$� m��h ����@r�͗Yy��l�[RR��)Ai��"BNm�-��t����m0[B�L!Pbݷvjݜ�Z�9�  �sI��7k���ڮ���B���mMiB����][p5Uŗf5pqn�	�^;:0�Iqׯ[N�U�9G���m������h-����:�i�hѷl�p	$IoP�$o]&�֎� V��p��ɥ�rlohl.MӦv��Uj����@ o:t������n��	�j۝l����v���	�6���$gjm��h/pR�D�g0&�u�4�^:�:�'�}<���&�H�q�-���k����C5V�!^�j��ᗲ�h��W$ۮY��z�(�I@8��ZKkm��+N��� rҕ�Uh� 8  �۬��[��ج$It���"���q�+VNj��秠�y�7��b٭�EuýC0��$�j�hO
�v�5U��Vݶ�T���ζ��-�9�� ��I*z]�j����I��K��L5��l F�f[1V�7�:xtX���R�"D�&]*�?��u%[��$p�k�5�Ŗk,�h�-�w��y�����:�������@"����0��$תN$��8�wCj���+X˓gh	84u#�×M7W��h��f�-JX:p��m�m��R�^�ɲBKַY]@jNpm�kn5�5Ӣ�/Z�j� -�k�� 5�E�v�탸[*�ۊ�0F���b� Y�타m[淴K|6���z��ԖM;` n����+�z�һ2,�M��mGI@���-�ʭ���L`.�o�Bg��`zbu�U[r�Z�	]��Nf�V5>�m�@j�6n���t��9q����v�;�U� ��s+*�uR��U�T��lI!#��0[d��$���M�r�ZrE)G��ۥ�!U�p*��?`�t�z�@^([@H$lUJ��U�R�e�Z�U�	�j����v��̖P [@ ��� � l$�V� -��:l��^ɚ\��  m���   p�6�ak�k)	.�[@@�6�EX��]���Tӭ�B0a�V�*D�UV�$��ڙ�Z��h6A�C�T��o� ~Bb&e{eѰ�����������Z��ݝ�
��ԏ��N�/9;,䶷mj�N ��m�٭��ڀ$6�  � ���e���,�u�m�p m�  
T�6Z�$��ɬ��:���6Z6.PةvPB�T�uU��Z�#i���[�kX B���   Vڀ� (8����P�@3��]z�6���mJ�Qu6�cj�ͩcQ%���ϻf� q��[�N��Lv�ma����	ޫ0(��	$�J�ѮF��6�&[A��z��[[m����[p�)N��[P@\V��=T�2��[UX�S)iu�[m&�` ��  ��"�qpBm1EP<�C�y첤kV� N �kv���e���[Y%@a��@B\K��� *�`9�@]�5PSͶ�  �m�[x۶�\�8m�d ��J�6�-���$Hp  mpm&�mږ��Ҙ�5SUJ�T��KW[G|:�ZԒ-�Hz��-�,���lf�jN��[BEO4����&�/]��]�n�Kר  ,0F밐$ #m�kF��K{[�����5�eT��ӏ7*���y�|o��)�a���͜q=�2����၄,D�D$�g��jk"���
�2j%(ʖ0�(*X�̈�h2�,
�� 2������T` !�U�Z0��"(���(��(�R"(�R"(�R"(�R"(�"(�""�(���"*�"�(���"(���(�"�(���"(���(�"�(���"�((���(�"�(���"(���(�"�(���"(������(�"�(�(���(��(�"�(��(��(���(��
(h��(���"(�R"(�R"(�R"(�'̎9�G�G�T���*8����F�ړwF��XZ�:\�Dp-c�DC�e��#��tr�U\����j\�'%�R�R�s:�]Ӷ�����9�m�<�i�4I�.R��Ҷ��ݹer��깮�|ԝ�S��kzet�jo�%p[V��.�aN.	r��:�7�y[*'u��fh��In��K��T��\I[��e�\wM�S(���͡m���6^&�f쩔w6�(�u)ۺqԗ0�Z��N2u+�4p��K�5M��4�X�g�sN2������i�UV]�Ա<��q�ә&T̕ٻ�-�ڷ)��h�Ժ^T��V�LҺԋJe<ʮ�^W��GO+r��U�����[��<�Kr��#7q��`���	Ў�-�ʃt7���bX���Ÿ�jO6���q�+�R�G�Rh-ռ%�B��<wrG:H����l�jm�m��ܾ�//����r���yyyW�yN�^U�^U�^U�^U�8PU�^U�^U�^U�^U�^U�^UU�UU^UT�v�  &�nrm6�&�nrm6ڞ��)����#�Mu�[m�����n�  ����o����9�rI'�4(�2��P�H�ih[Jٱ��d�ص5-V�VCcB�CMSFB�Ze����<���
�C�cʙ�h����g���`#];'8��$!�zIK-��I�#Y��d��� �t�f�              m�        ��iuw=�1d^ݬl�q�JM��๧�<��m��*����i���(T���B�Պ�\*l!8�;bȭ6ڙb�]~?/n��eX+s����ճ\B��*d���q��`r\�Z��MpV�n���68�k����¸: Z�=p�(5P9��GfZ�6ffV�P�	y�
J�V��c��R�۱�h��4	��Ycj`� ��UR����9ɭƝp�#q��]nlm��n{0��K��2�!����z��}�Αi^jUT�;��r��:�-�h7gD��t��ÇڃR1���5sP�.�`�ߟ����nhͥ�1��q;�'T�s����;�?�l���#�{0�P�i����:���~���z��`���� �2�72�<��jq�[�N�t����u���t=�D�ǸR������P�tP�4ڣ3m��]��r=>�y���YS����o\I[�]X��$���%�g:�lG
��oD+��i���[��2��0�r�VYp�d$$u��ַdB;6�
݊�ms����0�{:g��!�ѳRT��+4����)m�9�6�L\�beqۭ��kg)X�l�Q �i���iBx%T��κ���7ecHUT�I;�K/��96l���8�$ɒ@7F^�'�.iIyƎ�سԗ7-�ܐE�%���UpW���-��&ÍD��qoJ�e;�ץ��c��/ (lR!bE,/�=�Z�p���}6  � �-c
qbe��V�1mA���������:��Ѫ.]�ΘA��ntKqu��i 4�a���Δfd����@�r\�9�Ě�	k2p@�������o���q3��r�{뾺��5r��n�Г���ծ7Q�G]��֛Rʐ�9v���99<Qt8�lRGwֵ�A�挣B�;�M��.��n7b6U�6l���w�'V52A<��H?�?f�I�a���Z��8I���j�b�6RY�Hh��$$߬�� �i��c����!'��8Ow9	7�$���.@���6�W&�d$�2M5��I���,FX��{�BOo ���{��H�섟UP�礉=v��"6zõ�xy�-�f�١��S3���s}�G��BM��x���!&�0o`'you���Uמ����~P��O��8F핾�f�Z&����W� ;�wd$�o9�M��	+�1Q�
&7$�l�9�!�l�M�A	���!!D9��< 7���A	ʠ�=�I�����im&�&+�pBL��o�9�h�!'� ����]�����є�mm����G��x{6��Ԙ0�I��Ǝ�����%�!$^l��lǈ��6�F�L����	9y�$�.I�;oQ�ď��ݐ���&����TEt*�s9�$�ې�vkc�BM��|$�l������	;��p����a0������b~z�w��~|����<w��G�������O㏾�c�'9�p�g��w���z&��t�&���No�$�d����I��!$�P��A
\� ��Uu�y�O.���m=��@�ߑ�Y�Mj����$��>+�HOW�o!'=�E�n$��<W{�	7�!'pd��(h���@t�ʠE���K�iOQF
��xI��	9�3��͂n�	���$��ڳM�i�@��Y6����4�n�Cb�	jʣh7Q��o���/s��y�z8I���W7�!'0ף�bfF��p�y�!'��!)���w.g
#���"d&'	��pBOo$$�d����!'���F�M��	7�%�{�9�M�ʄ'}�Ķ�wg�ORR)L��|���y�I;��D���	6x^YA�腀}��  J�\	nH��i�s��[OM�v���jˋ�bq]�:�]L�M,#��H��-5\]j�È�<�qY���<���Ӌ�ѵ�SpU�=t�Ц��=n
�'��Ge�m,&nۗ�^���lO �/n���=�ޮf�a.�cf@�n���s�a�.��ϣ�1�:v��JPy��'=pBM��RW�6�d���"cEcq&�	J�i�`6o6BO�d$��w�8��XS�(�L)A�I��	9�!'��BOz�NǘD�oQ���
^��{�$���DO}�o��<`��.7�Os`��� 1��}��C��I<�97��USZkT��ím���ڱ&y�oam.#y�GCh�ﺞ ���A<��p���¸����uo�F�O[��������b#�_;��pN�k	�ڄ�ߠ��� �B�D���6
���O��	=�o������:��b
��(���R��'���!'��	��I��#��QF�M��^qI��	+s9�D�6I���I[.�!b�
�K*r��Ѵ�dNd�y����b����!'3$$��J]���Naz����&�d�>��	9��o�!6�b���p7�Os`����ڡd@+���3��ucW�#Hްu�1!188mu��o�!'p\�"{�$��b@�I�f1�M��I��@�Ϙ���{�t{>�XƩ�B�^.,]mŐ�@�k2�bݑ5I��=6�u����/3���܂o�D�l��Mb"'	�`��)#crI�l��w�sd;�<�(n$��'��!'��x��39	7�����l'����\$���9xd$�6	��U�EN����x�BO2�-�J2��R*�BO/ �;���C��^����Uf\�ƄZ�&��+��%�-an�ws]A�lgn����S�:�� w>�{���W�Ka�ᠠ�΀���F�L����!'��!'��ŎF�Q�F�d$�d���i�|D���t���3�Q�ݐ�y�BO{�@��T�<f�u�Qe����1�3s���~�p�c�'���@eQ�Cj��/9l�!$�s�<<�7��Ҫ��  ����6�-��e#�����Z2�����b#��-Mq�� !(��n3�]�LuR���,�[��y�flhf�:J�5Ԉ��X���ɍ��v���%�q@R��HM��Jݫ�LU#h�d��ThVU|�ܒB�(Kv^.9��f�>W���}���[i,����:��:�g�X�J�ꐓ���D�6I��1`P�	j�xgZ7�BL��	<��	<�:x[�(�>^���A��r��@�_iҫ�7t~������P�rw�凞O���s�opA	/�1p�{��/`�����%��gGFx��������m�:Ș{�i:&�bI��M��	��������U>�w�$�G��׹�f��U��o{�]
H�ʦ�(kCLi��F��XF&X"�q�]I�YIۮ�n�b&��8��䄝́��d�"NbF��	7�=������HI���h�TL�	9�$��HI���>b���J2�Yѭ�������y�I�npp��0���¯ݪii6�ֲ�S*�Zi�$��ݽ�]=�ј�$$��x섞^A	7�_w9�M٭X�䑳#|$�6I��!'���g���(RGu��<biFLN�}{I�O�O�Ͽ�|��  �}�s��I$����n���rI'����*�%f dRf�@�}�#�4(bh��J?����?�����!��!�Ǡ詴&Xa��d.(i|;�l�ι"q�e&*���Co�D�s��]��v.ð&fJ��Jsa��a���k���;�y��˭~�}�!�R�^�����J|(�)���:TM��1t�µ.!��n�������C��y�z��M�7�{{�qn���*�{m�����$���Z��"�#D�ۋ��3��	;�ͳ��O���>��BI�G�a��(DN�B���'HAk��W���~X�7	=�'x����ǭ�B%�nN<�Z���n9s�q��fٌ��F���v��wΜl��}����N,�5#���?~�U�p{�'�����1q2T$�_��2��x{�8���D�����ȼ���I#�x�߾����b��G�}H����E_ц�(�qΓ� ��.������7[=�n%?��s[��2�Q=�u�G|׶��}��V�}���"z�b8�I��2�~� �ذ����[d�r��҃d�ɞ���w���!�m �ڵ�^m��I����I	�>��{�BR��BM��g�����'!�C��TjA���Ͼ�>��BC�􄟾a�{�|�����G��~�		J�I����3�gц~}�y�	=�a�'��)���G�}��'o �����p�v������9�?7�9�GS�	?~��3�]�#�ސ��Xv�?�rzO?�}՝�m�z+�UUUT  "�Hצ]�ؗ��kqق�I΀�[�>��؄��ݣ����^���vQ��#��� mR�v�NK�D�Wl��N���+�@0bgj�f�کK+����pX�WF���B�vZ��s��qhge��F�:��)��Ħ�$��yq�]*���kc����[�9@>�Q� =�z�'8�#vP8�\������xm,�&�~�>�q����%�O�k�%���&���>���%�s�o��P�� ��yϻM��G��+�7	q���2Ox�ÿ�P 	3��	>��@���
FBRc���T ~������W��s�D���K�UUP�_p2J��b�b1��r.�E��p�/�S({��?�a�J��O����<{rI��d�B=3���2J������$���Ӥ�P�g� ����}����@~�UW�&����I��02Sdn7��U��)�Ї�B/��H NǦo�$�~�߇�T*B�w�?����C���ИI���P�ƨ}@�{HI��~��'���@`<Ծ`
��/zw���HI�d��UO'ڡ'�0ׂJ	�����$��=��}D��\$��'�߅V��H�0�M��!�d���6۲��[)J���9Θ4g[l������������?u��	�~��U���$����>E~�l��{�ā;��޶~���6v���*F�m�����'�����NG���K���`=d�N��;a�z�ꄓ��0�)9�w�	������I��P���	?f��l?�%N~�=^�C�o}�d�P��߇8O�s�'W�
j�����H�(�B&��k�u�4(�bWFjY�Q��ĩ1z�ɋ=�*/$$�˟���L��B~F��B�BS\$�����]���HI��a�G������T���k���΄�:I����|D�Xg��UUrb�$�}�8I��X̑�����U}B�~���8���?~����D��3`�7]�bp���{��p���$���pt���Bu,_mo�ݴu}���I��{�m�$���0��A=�K�o���4���A�>!�B��������BNe��'��>��W�y"Qy�ks�'�~�{� �r|�)-/,�K��'�� ��6Jmq�As��y�I��Ϩ~�~�$�G_︸���!��F�e�k��$���}��Gsd'��s�d���Hk Ȋk�����H�>��ޒ~��I���u)��P�� ��̰3O����{�   ]du�+-��ӂݎ��öۂ�V5v��vO9�V^5a.7:��Yv��u;�ظ���gd��kD�)t&�zu�T3�gg�Ђ�Ū�����Q�rm�N��a\Y#sY���nR+Z�n�]���W������Om�z��չ��e�L��V�;�yߢ_d�+인��^[����:I��ﺺ�K�d�..���O}�	7`�3����G�O=�O�W�8�ᄛ��1#���v�G4}	DT��Ou�x*����-tU ׆�H�=$ط�j��bJ&�<-r�� Ug޸x���z��a� B���\�	'�w^��A��t�/{y	<
�BO|��M���ެH������U$14u��d����䱸A�z9��� ����(q��.t�牆O����zz�U"{�!'�Z��Z$.@�$ߞ����\�W�*PA�  ��v�k�B�O��:��=!'���8�!� ��dp�~�ː�$���$�ϦZG���zPH|'�P�}�a'�a�g��')w�-#�5���mX����0��o�@N�~P?{����z���;:k�.�a$�.�p�&?A\G��(��6�I?U
ߧ�=�g~�nG�T8�[�0�9����m�xI����k��u���$���($O�n�&6�$�	>^�	'1Uq�J����eQߣ����}�2�??�޷��J�f$��'h >�$�<0��zB{�@?n�}�y��rH��G��4�ʡW��ubOvBO��yמt��:���U�˒b�qRKW6�CcC�k�N
�P�O��)���j�_��un�K^�4  �;0��/F�IA&���$W�O�@ >�a�o纸I���s�UI�&-fBڑ��I��d�[��*�W���$���'�D�J2�%�U��0ovBO��'���R��< ����BO|�����..{���H����{��K���bބ�s�s���w���b�x�MCA����܎7��d��˰ŷ�&苺1��?{�P=�LW�^D��/}�Q��1.s�#�a�U6q{T%���}�&Ф����RI$iq{�|$����.� �n�z���$���A� ƒap�
�7���q{��;�Ι?
��  o�a'��0߂Q����}�!'«�BOz��A><�z�b_����$�I$�I#m�$�I>�9�I$�IϽ�߷ww��9$��B���� ����]�qU��(s4��22�������-kn�X��ː�׃�u�ӣӜY8���+S�\�e��5h�XS��t�U�ړ�wl^����|�:�/v}o�;��u�v��M��,5�M�                         	9Q�3v�+]6�]�OU,�X�`�;A�]1�F9��(Lƅ+�I���ݝ�ɑ�^�J4����A�'�m��N����;K��]Wg�\ �3lJ[�� ܋l�:7Ms5�̶�}1�c�s��;gG�\�-�K���q�,#Im�K�kH�&K�)aM.[��q<�^.΍�!t�[l'g������Vóg�+*�X'���6p�.2�c<�申m�R8�sgg��5mGc��f��Z�t��A��VP	e�UcYvp�v��Wq5M�n͖��nQ�9ڮ(%�ѶBۚ�0�'��/��.5��'���1�sW=�n1����:���	mA�F�-1��#�Dք�*9�rO&�$n��W�UK�m�[n�v啹�[(x���WC'S�ҳs"��6t�l,�x@.�.b�Gm:����(��YӮ�{K(�Jpt�-�St� Y#�$��;m:e��6���. cQ\���s�fͧ��i���Wظ�v��*�� ��q�*�81�la��X�$�lN7mf]qRj1��CК�[@�F�kY:�"�'K;�M
ҭ���e�(�an��v���gSl�]%�M�Ku����-v=g&��J��gB^�&��k�\�ɿoQw���a�S�J����<O4�s\�o�*B��TO�)�❚��^a��ZsZ�{    sy�mX��@d,3��s�x�/1�����G���ʅ�,�"]�z�ح#�V:u���V.�ϒ���iAE��U�{㱄�yȔ\��95dX�1��-l��e8�7]y��w0[y��v�4u�R�%fa3b�kB����ܕa;��T0�S���'~u�盥T�0�����"u�,9)ߤG���cv�؊�K\g��G�5	�@�=�鄜���UO�L��y1蒉FZc�D�8g�H�vBO�l�����FżCf8�m�	7�HI���l�v�a'�T�zbDA*�79�x���BN�<ѻp�O;�s��"Aŀ�d��S��k�S�-p�w����I��ȪR)��ٳ8ƌ)5L�Ё��=��=�<qQeufHa'��w2g��%}���'�|�dL���O�C�V��t 5�(Pٓ�}�2}ԏO�^�y��J8�p{�Ѭ�buW7�������Ԏ��d��Ug}�����h��;��ID�->k�T�B�x=�s�m���'���ն�p�Z �Ź������e�fxr����'HR��^�y�+��}C��ث������ I�o�� ��b�-Q�6�� ��X
P��1�k�{�P��
�{�;@
�HP�|�����cDrHY\��_P��x�c�߆d� �����sR�%
I�}��ڪ U�j���;��]�k�$,$i�P �H�ٺ�C�����N.�۶�w���
޾q��Cq��D����ޱ�+2�U�C��;����JIH��?UU�^�&/��(Q��z$�F$�,�PG��hz��o��\V���Q5j����1������T8C�(���^Մ��`4�JĊʤ���? ���?&k0���� �O��k��P����,>#�τ�M�$�\>��̢���*-�8qe"�f!�Zޡ\Z��ߴ|�vS����O^r�>�1�$is�Ӡ���=�xG��@o�p�I����'m���{�Yo�a���̐��z=��_��p����<�{dϙ������&/���7�����{��w�)���4�qP�I	��C�t�>�D�7f�    �k��[�d·�
�U'�R>�v*�p�쉚;��$-�©�PlnS��j�qV���9_n�>
[�\3N:���,�y"�dK�_M��.Ûe��<t�soW�؝�	�NM��ָd�Q4o���ӮNNnNs�Rs��j팭�խ����\�f��~�]�ip��iċ$���.�����@
�[��0�Z����r2k3���y �y��u�!߈��ȘB�A�o�	�^�y��y��I��9ıƖNO�������N�������[�B�}��jbO�U���F}������.ڒI��l����kpKI@��-�D�<n507ރ����i�}��̂;��!&��ٳ�u$+�>�9��2 ���K�aR:@5^��kw?g��Ǒ}���+��
F�H"��'�G���c�	���|'װC�T;��� `�>�(_O��g�5�}��`7�P��&�m8��>���¡$���~����7ʮې.��H��Pu��D=r�˗Ɲ��� ����zO���D��HOz�Dz� �$�K	F��,����o�W� �~���\��}�A���'�/�cw����)�u�����TOUd!�#����܄���y����'��	���y��Y��d�Q&�7�>�>}����vFuq#�����|������h<u�#u!.���A�����[ܒIxI0�yE'8��~f#޻0�ןw��fM��//!A}�'1�˄� �r��>����C��c����jM����	�%���n�,���y�"B-����&Q��	<^�_��F�>��П#s��s{�2����h���8w~b�;3_���qÅ~�U����ݡU�蝺::��u��y�T�<`8n�w>���I*�	վP�{���d{=!$x,�C����%߽�N^Hq#�������r��b3�TIIMs��y8A��Q���=����Cފ�$��d(ےt�����Y��w�~�j����p����"3n��XޑQUf�{-�$}�1�P�-w�f�5U:	�:\�I    �I���N�9W��bM�ۊyݧ�o,��5=���v+��^�����%]j�m�$Wr�q�i�x��˹�H��S�5m=��Xm���jv�������^����H@6ݥ�XJ�ͮ�CKl9�$�I�kҪ��sg��l�9nv~]�����s��ۯ׽��|wŒ�Kj���^7���@B}ea���k l!��'��	�G}���Us�c�	&�� �#��AX�z���}���.a/�}��Y>�� t7$��޲���B���/^H~�U~��/��jI�Fg�C�}!9ܐ�^���R���$�G~o��ƕ�h��RS��eݶVѲ���E[1�J@��{5Ȇ��a�P�z@{�5�v`n68w}'�t�+(W ��3�#,Bʴ����LĔ$����Cx%*����+!0!0���y�C�0 ����o�9i\�Q ��ۡD�2��I"��A���>��}��<>��qY�"��(�P�ѿ������ݞ ;�C��1萂�}��pA {�9nȄ�{�u {�6Di�4Bml���aܦs��K��FR�4�뜜��(XޕЋR�G��<�dC�z
 T'��	;W�@�jE	k���7d�^��O��P �4�ZI�fA<$��HNw$:��7� �m� ���}�$�Nn}�ww��9$��D�(��$��r�0ū31̰��0��2a��s�3#j���'	,���,��ʃ��B�0"2	�K$�0�2�*�ξ��3rf�=��8�$��G�������@nlSL,� ɠզ�bm�2�W;Z�'��̣�;�t����<0���8l�0���ⱴ��2'�)��.��"H��8��L32���0�1�1�L֭��u�^9��������#ty4�8����WIw%��/c�5M�wQ���5�\��ۗ�+���J��S�{��z�����|��p�N2t(��!Β( ����ݜ�����l��y��'"{&�c�	�]~���?�@'����$���*� �g�뎓��䱨�xISa���5�c}�w�~���	����}<k��g���
��ސ���k2�mC�A=��Fټ�{�}9��� �C<G�ǜl1)�p��H	'wg��P �ǆ߾b}�(�x���x���;�f�{���D�P��r}��$��� |�HL�s��錠���y��9ܑ$������0��7�أ�r��Z'�Hvm.{98i������6�u����be������}0���<��Q% k����8I���	�#�S�'(��-y�6P�&�I>���c�	��zBO��a@�{�DB���G@Ś�w�'�� �= '�Ō�
Q�����/:�[�����}�n��ND�*s�S�М����?șUUUUT  6�:�:'M.O�M�7��~�[�m3GY^Bvl��(kj�&�����/=U+��ަ[�F��:c���X��e��<�8ۖ�.�qo7L�lö�t96,�FhM5JWq͂�X��-�Ӓ�d�Lƌ�Me���;RI'��M�v��;q�ў�WW�<d8��፣V�CuSm��v������:�������PD�E�`��>��'�-(�=����	'ç=�ˑ�Wr�^��<�p�U/�k<D���SVQO,�Lh#�߾���O�r��J#G{hy��D�M!#�I>�J�@�u���J,*���-t�y$�&E����ۮ�j�;t'9��h��J�iv�c�� ���9�!x�s= �/��80�i���dozޭo]����
n? �#�]"2"�P�>^T8I	߲~D��N�hq���&�P�U�Ӆ`��� 罳��ߌ$����6F7Γc΅
;�BN��Π� �\�-@����*tw����ۆ�=�=cg¾�Ug�ߟ�T����s�f9��C#qC�jC0�Ns��z������B��~��a'��8�3_y@P���	�-ā�C)���$߽^;�@���H��2��Nݡ�N��Eޒ|7�����u_�S%�ZB 6���@w�[�\��$$v��q�ʎD�>�=y!�-w��;�{+��DF�.>����;���{�
���{.��P+ I,���B@����\��V�9���>�6��y#���@�Mˉ�1��q�Ғ�zA��KGG���v�0���k�L(|�>�A�Z��ux��)/{����	9h���Pp���s��Uy8�|���O�쩕blI(�����	<�c׌~���@r�����m�ț�� ��eB�#�����ğ�����@?{�����6i���w)�B���Я���u$�8:��X=��}�O�}� u��� xM����$��1��r&����	�Vqa��=y'Ʃ����)Q�!�w�5|`6ow�Jo�n��z����Q���Q�"�W@>��w6}��<#���>0�3�}��D'΃��W�S_}�[�����W?~��)�`x?�	UJ��/�T D E��I�I$�@   �5ۭ;n�؃nM���씪��$�b2]o������2���z�Ly��<�<mUDn��O!�m�AqUv7&mǧ��^-��宄i�͵��ܬ��I��ǵ����������M�����3W��s���tuҪM�����s9^����8��`"(�!��H�Q5�Q�J����^A��=į$�w�f�C�BZ����s� >�p���x�
�yGp�ކT)C]����}�~=�ϱ�^-
#!3�o�$��ݶ�?�A���$/��Q�D�	'��O:�m/Y����F����]6mR6�G�n���f �6�jZd�M.�Ps�rYo�x���4�]�aP��^s��[�a�wַ���E��ۿm�o�,�.s�3?{��yf���� � � ���l�|W�g]�Ў��ا9"ם�h�@��	�����w"}�h P �#����{oy�6ٮ=H�H���oh	�	��f"�כ"�
=�-b����7R d�4��W��hA�
� ��'̼��k-پ �9(=��B�A�A�^�����k(������lE���HA?�͢=�o����y�Z���4�>y�g��9�p ���Pz�������=�%�׺Pw
��99�zko��\�6���E2d��ld�A����C�6;�s�|六s�v�fr�iiA��4�|�fH��8�'�Mb/1���>��Cp � ��0� � �#�~gֲ�v�-o�sJT�2E��L�q=`��a`G�}�p�� �޻�4(7�����Py �B�H�ߕ��\ݭf���Z� � Ѓ��iA�(4�=u�-� �	��v(	�Lh;����GX�[u�-��2@�u���44 �����ͻ�oV��=@�K𤪞���`�@�H���d[�b/X���8܋0P��w�*�&�� �r�*9!�}A���0��l] ����>��oU[�$7B!�*bZ�hڱ-+��LW�������;��^[��ϔ>�1�q+$(����>�W�ae��ف�TG;�/�hl��m�}��7�z|�|��|��Ѿ��wL�J�ej���x�/��G�FwЂ�$���أ��T`�z���f��Z��u^�b���}�� |}��z��|��Y^oⵆ��h0!]�%؄��5��wJWHl�u@nBө�l�]s��]���!8ˏ�mg��GI�}x��z��Tmb��d�ƣT�~�o�}U@���8{��;�<0D���צ�n��v���g���K!B���-p���6�<#@��}�I$�I$�InI$�I��9�$�I9������s��N?�>!����ѹ/����%`��i�j1�7x��A0��x�ē�,FǤx&�� ]?�vv�0L}�o�e���=��S6`I���L�b�&KDPo��������4qH��ʀѤ�[�||2c�z{|�1$�r�aMbD$�I�AV��@�6zI�u���є�	|��!�u�.%�9�myu��tPa�������5���N �\���զ�                        $��2��(�%0]�``�������#�wF���㜳vR��n�[c#;suW/M�ؑ��+�-m�2 ӶIq�铣��U��!T��[d���22��i���X%NM��q]Q��ղq�՝Y���*<i�#��y2A����yסr�n1�����[�0��^���g���D���"�4`�,h��q/n��I&JWV�)L0���MI]m�7f�VƶE�ڢ��m���3�Y�&�4b��KT�Ua����(Hnm���nu,j^�ջ!l�ٵqO�O ̯U`L	)����5s�.��1m3j�f0��M�TS:�T���6�b�I��͔	��#r/I�m�EH�m�&�4;tBl�
��y:��lsƐ@� 9[���IO	pb�K̩�hK]WTkɭ�U�1���PUA&nGp�.2m��:ү$�\��2�,XKU� �N[`)%9a���e�uT	p�-�
N,����jL����EV�t崅Ս�*�84;�т��5 �ݺ&��nWn\�kI�k;tl�;k��\skن�	���&�R� Y�Z��U�d�9@�����j[�8�jqk��[�K���m�[��7�j�4s_�/��U�j��IM�'��a����1f�ֵ�6�E�J��+�Q���5C�>
�0��-���ڌ��C�MIwG2�Zj�ӻt-�9H�G�\����zH���I�%�
W*����  �K�Μ�f�c��e.�R� �C�f��fƫ�_w�t����V�; ���ug��?��7],�ȳ�}?nS�o�$wc��&���0�9�y}jN#'�8���\��]�]wi��^�C$E�pR��(s�z�g�}��g���"���	4DK@�s\�6׊���Ntq�V��S`�JK�١l-S���:z��u#���\���y���c��� �Z���%ăz�_�M��a�loZ�P{��N�,I���]�u��"~7�1�%3��$*>�k���U}���zwb���8,�?��v����'��`K6��v�k"K��G�I�Q�R�R[��)6�˲��LqGƫ�~��:?_ߪ����ƫ>�_����&�Ȿ����к��"�v!��<<�+��@�w��5h+ �@����p���;���^��c]e&�,�8u�G/���Os~���8Z��`����9�vG��t�Us{od���r'���oGK�w�k�����51�ʥ&�J�,����zzm�����{�v�G��!D�qׇ����x���u���i��~ؤ �q���Ƴ��
D��W�g3�^�a�q��,�NG_{=o��<l���_g�{_���Ltf���[�wη��'�r���tV�kg��X�lg�&����;[^\�H�GDv8�[�띷[�	�w_=Ѯ�&�,%ʼ������S��Q�8��ʀ����"�o�8��u����:q�	F���3מ_o�����w��Mǯ�и���� 5@~<���cxJ?�2
C����;�f���ʪ�m�@ZMY��:·7���tɰ�S)@[n"�.E*'LG���S1dz�Ͷ.�Q�hj�Ԅ��`�f��UP�3$�R^��㘙�x�c�L@ёpfk�&�ʗ�S5��7	mF	)���싶�:u�U]�t����8�j2�\���1
�����u�ct�ɡ�Ku4SV���JJxNO�I��:��ʪ���� K�'����Bm-�z��)�;ۍ[2����ҜO��6�7nܥR�AG1�B�[�iH�����Хu�h��۞��Qs.�^�uj��h.M�Ӡ��u���\�n֜l�7$f�8�h��sev�����}]ڻq�;[��*�Z�k��'VHMY���Cu�7*�,N��{��T� ����t%$B���@&��w�4�-��^��YN3�a}���t����u���N�i�ް;�c��];z뤍�dHH0�zS�v���;�����<��e�r7���.��Ӄ�������X7�����"��a�>��H�n��������a��Sq���c�(Y1�(z}�@?^dg3~�����Y���+��D�11;��H��e&-&�2�B:�T =�1w����}`m�Ӭ�J4����n���b����>� Q��Aq2̆vLk'\8HS��Ƌ��G
h����k����}����1�뮊�kTQ��8&f��+�ů1�ׄ{���0�y����>�߶g}���M����l�y��9��`�t?��L��O��W�f�v��}�1��h5�6NY�1w��c��0��s$�N9�Hr�$���p6�;=��4cEB�Y��Wf�,]�zw��<�b�
��r�����u�6:Ɛʲ:u�ED
p��xGP������Β�)�cQ�v�i���l�,�A�A@5E
����$E#r�:��ע�:��OzM�$"��b.]�������v�d���68�ۚwN�����f��p]��;��Ǧ7"��7t:��]�;����a��9'(��������\�֍���A.�bȵ�w������Q��A{�c���i��T{�Ϋ���;�`}@B�!��>��2m�j��I�צ�    �w%l�b.9ə�bњ�8uWQJ���b�s��[X�Ĳd�v�$vP�[��v�"��̷*�c�T򢀎;rtYF3As[��m��aC���@�F��Epj�b��r����+�vaʲ��s���$y��;���Y0T�{��9.���� ~�W۲X�����TM&a�k��c��4�-�8;d�F21��u�܂�i=�c��]�ȥE#N>fl#�̃��e_u�H��\E��i���wu�ލ���_����4 i����]�c����M�$�3�'hG�Zw.�;�k���'m���\��'K=�ߍ�.큷��P������/��(��+�w� ������P��ޱ˶/�:���O�݆T*:�<��]�Æ��A�q�,���	B�N�g�#��m�1g}@�F/
VN2�f5_��~�U���`dt��I230�$l01t`�X����]-2c]�s��6���j�}��嫼c�����݃J$_����";�� 7x���T09�>ǦD��s�v��h
�9C���I$�I$�)$�I$�Ns��$�I$�ٿ}����9�$�� {y21
P�'�z`���K~��������8u+�A��gk�tm!zp4�Chp<�h�0��#6Ns��,�b��Nma���z��F���~v��믭������ь���c��m�U��8�>��x�=�Ke�y��$zA(B�IC��Kp{`�{m������0m�@ Ymƀ�ƒC��0hl8�a��0`��C���4>�#���p>��{��b|�͂��/�͑�}#��p�*g�KI>5�G�k��\P�}X}cւ��(��U�������`����r��r�-!�"�@�i�ly�]�:���W�HXq͝�����<	�q�r�W��l�*i�K(ͪ��t����~g���7��0H��P%��8����W��Wz��s<�G�
�)�1�w�s��h&��w]w�N�E�$q�����f��=�W3���O���l@���"��~��U�7��1��A��b�.CW{�Ne�7��c�I$�i��e��`5���Ͱ�0��Q�������t����;�_t������%"�^�c��	z�b���t-#f6�\���7��yf7G�����ь&�3Q���1w�a���>����+~Z[�J&�$NW3>�����^9��~(}D#'_]�    6�\.l�v*�yŉ�1�4��׻-��]����k���M�C!S�(�"�;\����#-\ݎ=F�m�x�j����3�/�	h�7m��v�q�烵���v��$�%�U�A��;V۩�FH7��&��\=��qAnW{}����>m�Zb��ҏ2K��u�D��x[�2������QN�3<���Pfu�/^�6H���!H���Lw�ǀ� �@
�z��s�C��1O�wwܫ���ݱ�������&շ)��j��(��=�1w�;�'�����Sb5�GA�8qZ��R��5�����%%�L(j6���J��b}��Ϫ�Q��	�Ƈ��4p�`g�l��r��L���T�ǃdG}��{U��ɧ3]p�>X[Д'o�w|���=�<=����NB�( }�g~[�t��7`�m��Y�P8�n>�u�h���u�����I(���=s�&�quq߷�v�л�p��L�"���L����w����kMt�w�cd��s�n�U��V�j^�Aͷ���q�zl\���	�B��q��s<�{~�Y��WD;��9��w-�w�h'��N�f0�5{�����Ӆbx�m�$ҍ���k��Zxk�}�5�mi��6u�f�2������u��f�8^.��Ӽ�퐐��S�&�;�d�ݡg��]�]��CTR�q�x�q-Ԉ�3'�3ν�h�9�dFb-����Aۼ����9C���GP� � 4� �;�Q&���#g�lF��~u��N�#K����Dt�ݒ&$�֍�#�{c��a��ZsM6m���Ŷ�����?i�uU�}
��M>;^�/��,��+�M�6�����71��C��ጆ�mw=����e��Ϋ>*�ih�Q	��7vWv�9�|}��S�_�����F:��,�C	��Ӗ�#�^��M�rbI}�{�@˲����� ��b��,�]���=�Ϲ&�덂x藙N��qsػhP�Kuׯ�����z�SI�y0��oOUЃ���1C:6��sև=s��DWY�)(�#��f�����C�s8ʣ�N{����J��p���i~��ˡ��s�+h��y���{P�'w��m�ifѱ�0�Q�oFs.�<#rޛ$��d����^���q>����H�Շ$a��N>���-���Yݸ7�"Ȓ�E��� �~�}�u����߮�����K��E.;���g!���{z�����.�If9�*NsC0�G�ScC�LϨp#/��	�;�ќ�u��:v�g:����p82���U �Ue`�R�0GmW~�����aw�j�s냖BZp&�q��ou���?(����w�W�1�P㈞W�5}�9���6�3�r�P/����$��"2`m�\�ȍ�Qތc�z��T�hy��e�r���5�����olQ�[�w2����}K�S�=���oq�<���w�d#׌2Zm�d7!�l��M�U���n���	E��)pa�	�|�O���
T,
�%
 T� i*�PI��*���_>c��lBGU�]�\&5�hU�>�7Y�c�x���3��Z�cJBT��-5���x=��H��]��v�5�IqT.4�,���j�Z���i4��pXPe�`M'!M:��f���v{n�7b���I�w�Y�7�<��s��IﲤaA�Þ���/s/������"֝�H		;��'ηq������>b�d�X���a��{���d�[X�[��꾪�m�{o;��ߕS��Ic�,Uo5�v��tr�l��ƙ�-`��+�NT��|��o��-b�e�cT�P�_�~���u��?u"3�CY�TFHT����:w�#�ۈ��Zp&�2�,}@��͜�^�d��V|�^a�P�q�>�����lX�������    o}���I$�����ww}�s�I9@Ug��H���,xT�e�wLFinSu9���ts�
�0c�h��bGk֕���R���麸t��ZT�l����S���
��AO��N�"��a͠�w10�m	���V���ps��!�<�S�^�h���|tE!|�]RB���KIz���K��K:�1�t�N��W+��m��զ�                        &����)����7E��ܙ���E᭤��=�$�9ɘv6x��^B�<�M۝P�l�+����<�Y�`Q�����l��D�A������d�-��dճ7.�6� eRü�ZTܽ;u�s��-�K��N��&��F���g]gS��[��#�!��ޝH��5�xs9�x�f^�]�kjw3ط��VC��H�.m%� �J�%���d�� ��m���[���
�Ʋ@f��Z��&ۅuDtf��FG4�,aj� �j�Iy�XxÎ�]���ڛ
z��U.��p,�[k���`�'��歨:蒬:��Ί��8��۲�-�<���:�i㝏E���k��<�!�8;u�m'))�ݑ���lM�HV`&0�
�h���.�s]�'���\v5�V҄t�d� ��[j�g����{u�v�a�zC�6��� s�1���� �j�ͥn�Q�Vd9a�U��浚�!����H��LT<��2�/[���:X�KU�l.�(��E�*��A��t�jZ�n�cF��ciKf��`P֤3jn����F�c��]�p�v�YݰUUrA�h�᪌���\Wl;qg�F,�	�g��$T������J9������B�*s�z.���d���R��#@������- ��������i�3>w�{ٽ�f     �"J�/6�.e�d����:&��8�A�=yvP��֋j��4�����n�(N�[��	���cK{B�Cp��˜�x�s����m�L'�r�[M>�$�;�HDiZ�y|b�]��t]>&40"�Ӄ���u����F�K��{������Z[ثM�[A:zw�Vܙ�$�g���P�$�$����Z��gm�#��?�P
~դr�"/H
����7dv�>���7�z�{vK]�:e�0�-b������g��Ȼ��X�1�J����Fe�f�]:�1���@�1�	�ien�2  �+یt��I��{?�򦖕q�sf�	�q�%����{m��KZ9�Q!O�}���bϺ�(��݃&i����n3
i���U׀�;޳��}��+c>W�G���#��x�#-��|#n��$�r�b���'�n1�یY�U^
����/H�PpG,{5��P��^�}�bܳpmPÇy$�mWK5�t�I��%��r\�C������]F���-����g-W�w�83��/�=f�)>�Y���^㭻}6	���ӄƂ;����c�������7���+�VY���*\�>ª�핷n�}�^��x;e-0&�aFSN���Z��OGw831�.�!D�l�� �!N	��v)�]�
�m �\�	M�m�c��x�;����]�u	۩���a����;�뾷�O���}j�l�P��Nto�үo ��(��ۃn��07-�[�}$ݪ����� �x�
@��}�w�}��Epս�	\}��e�཰�Fݺ��#�"�����c�L�ϐ��W��hWj�c��]Ͼ��{v�N��,��ON������n?N�1�؃;���7e[I�SN�w`���u%w��S�#r$�G>;����9�ǅP<�b���@$b	ZG|��ꡛ��z�A�U~� t5�}�'_�.�   Mh㦲���ǝ�Ya� ��!�[��������ְ��mV�5
������;Ҝ�\��2O���Zfq�Kr��,O��y�7WTPlm]��nV���]�"K����goZN�s�!�m�B��� ���w~{���I$���*��,�c0���	��h[��:�[b�S�thZ�$lG"��d�nkyk�C�y+؆���$a�ԯw]t�Q(�5\���
���k�f(�\}��eʿ[�۸4l^"2'�t�-o� �Ǧ��ў�b�g��TA�O�=��o-�ø�����V#ec����B��.���kR8�ݲ�tL��ɶ���g]=?}����*��0^�ydnA6�Q�`;�����4�bZ��F�M]t�^n뮶�gK����� ��]��/-���Ln%j�~��P�gc��P^���;z��f!���#�1�K�Y��M�W����9�vF!��$,3��1�D�t�yL���nv;r�10�&b����+N����ܕ�|�0"X�pF�4ͼ^c�^��qVt����R��9��;�>�P���:?�4&�D4)��p��2�";e|��n�����r��{ 9ۃh��@�nG��c|  oug{���z���d�IH8�F6.��7%p��������6ȳj(��P�"rBI�("q}�/-�wCy�K��!����RG,-���1��C�A��C8�#P�5��E�>7��bV��p^۬����{D�+���ث����z�(mP�)H��@P�:��}8	>�^�	qWv�i���=�1g�VG�EZX�$	��q���X汢�0	�ٴl�@�D��C����Jh��}��r���k�T�����E�PjӮss7�H�S�s�����oH���7#����Z�yy�ҷ͠G;�tu�A
Q( R!�P��{n�z��c���	�wPm��H�I�'�#���i�U;� _�
>(H,�"<�-Vk5����`   �m�,];,r�`Ƥƺ�N՛G1t��4q;L��������]l;7V��^�A�T\�]�
�[=���^�fx9�feG��Vi��wfݬIE�--�<a͢�>]n�g��k�ϝ��y��]-���Z�'�rNrI��C�����}��ȝb���͹)hsB�X?�1IN����y��B��F��#��Ჺ�Q������j�N�� �f"�\�uW7s89י�۷��9DX��Y��U�{`���+���>խW�G~	MEQ>?���/F����n��N�<������8EE�>�(RDn
����t�������f	BRu����P$P��H((C>�E7�I(�\��v�z�ذC�p���I��]����5t�s����3��(JNy�{NBP������9>��ȓ�''t�o-mcv��)9�m9���Rҁ��>���J����7	A�?\x��H�M�P����9��JL���vlJ�޽�n��5	��`�%'_u�̞BR{'�=�=��[�e��ġ� �:��&����3��(J��]�y	Bw��ؔ%%�B�ka�(�\��((jX��H��s����%	߾obP���ݤ��s����-�ߕnΪ2����]BȞSs�u�<��]`�٨�n�ֵ�%	I��{��'3��7�)JO��I�J�C�gy�P�Н#��.(����DP��
�������O3��)9�o9C���DP�;FY��i�@�@��~�.�'���)N����7�� �   _���ۻ��s��H�j&� �	UE�T�m���44��u�^����m���L[��a&R�dN��H셺S�e����R�CR��;�K���=�q@<O���caƉ'%�^S���Ґ����AJF=	 ���r�27�ti�q��Ne���:<g���'K��w6��yUʃ'���uĖ�<H�C��jSV����w��^v��댝u�[NJP���͉�f	Oqߤ���V�f����:��>��1w9)I����9	K���9��L����t���;�ǔdJi
�hs7%@�B����	I�~�7	Bu��`��']�궫Zq]m\K43���Ʒ�F��e�����}���S�r)�EHP�I��M��'y����w�$�%'��u���F	A|�'��$�P$P&�޺��γ�)7��9	Bw�ڔ%'}zg�zj�[��'P�'��f	BRo�;�r�a�O>�{���ϴ���&H��e�7ku�f	C�P\�����}����ﷱ(JN��I�J�6@}��H�o=�(*����p$�qE'(t��<���J���>y�I�%	�g��Q@�� ��H~V�I)&�eF`9�c��'���Υ�]�ڂ�V3h�b�˭��	��y�M�P��:���ߞ���%	�y �H�M`#wQ�9jr�H�H�S�g����c�JN��ݧ!(y�~�ġ)?wޓr~F}�Jy������ٽoy�P���߻NBP�w���M-'�{�ܥ	ε����߽�����V���'P����߹�(JO��I�J��f	I�2~���6�����@�hF��%4	����"�_�OZ�� �2����ǐ�'ݞobP��ةѬ?C�٭:��g�`    t��;��lN�:�!�5�L.��n84H9�:�X۞p�u�%������-۱�����4n���):�Ӎʖ��ɀ4�yq�`髳̦Q��=�Ӡ���1Z0�=��E++HC5��Q��$�ri�'FURM��Z^h�#�q�nY�YC����өl0P�w ��.p���e�����'y��	BRsud��BH���"��3Cٮ��)����37ku�f	BRs�|�r?�#!���{���d�'�i7$P�V��O� ��;��I��M>Q��.B{�w�)JOz�I��a�N�<���)h{�~�9	Bu���f�Y�lխlz�!��'�>�n��3���X��������:�!>���BEEw����S�:EEK	BQ�y�m:��>���J��܉9ry��J�g�Tr4X6ӊ�Bl6��xWCQ�k���V���9:��^N��yߛؔ%'�{��
!r���K@���e���1Ȥ�!(O=�{_�!�iJH����K��=BRy��I�J�ϳ����r�P$P�a��эFr
�I�^�7	Bs3��(JM��{NBP����%��;��=#=+yl��o���=�}�hL����=�r����JC�I���n� <�z2<��V�ֳ�(����=�w)Hr��y������4���:��0��EJ��W6H��M��Hb;�v�����+�u����D |F\Q>в((}�		Oz�I�<�$�k;�O�9	I��{(p���х(7򓂁�(#C����|$Bw��`���$��ǻN@�C�[���4/H��I(
{��eq:��=��1|�����c����1T�C�.�L	�}�ִd&}��|�%)?y�I�BEG��b$(+j���{��%	��bP��u�py.u��r�峐' r?{g�z�%-z�����w�(JOz��ys�!.�Z�"����Ӑ�'���U��6�@؎e5��3X �b9�p�Î2n���y���k{��2O��\�����:���P��}�{NBk0O{�{���L�/M[�fY�����4b�9)I�}�i�uB}�ؕ�!�~��I�?&JQ]�j�rݭ٫X���?K�y����!(O;�{�V\��<�nH�{�"		���a�	G�D�GP��!�sjP��w��p�%��X�!�/�z)����Ӑ������E��e�C�A\ ")���%�w�O��JNk�6���=;�g s�9<��ߕ�,fjk� �;@3�p6�n��v���L�̣-�]��윁9/��' '|�$�2��7�(JOz�I�t�DP�q�EH�d�B�#H����Byߛؔ%'�^i7	B.�(bB�"�;�C�쑓�v��B��߷�(Jz�A���2�<�
����A\"�"����n@[��J��4���.gZ�(JO�u��N�(?#����^�$����}V\����fq:��.��b�%�~��v��P���{���ךM�P�Ҁ�ȡ��A]K���}b|w���`    �J����Β�դ�#P%铷u�S�2¹�z�s�v:wV"�\g-*���!��B�	�)p�Y���Z��p������E��@��#Ue�pG]���ʸ9�r��g�'%6��:��!���/V�x"�_������+9d�r䉈Cq��B���'�?�;]��T�=.D�2���f�3v��k��JN���NJR��I��y�(JO������.gZ����z�OQ�di�P�	76mz�Hwd���I�J�<�	BF�s.P�uB�EgT0"Xj[�P����p�%ε�J|��2��w�n������{&IIH�a،	6d2r�H�H�x�"�"�'�뽧!.�Os��J�޼�n�C�ۺ2#���@�s%(O;�{������rR��3���9����=��T���m#,��&JcX,�Kf1-�fʙZ4����9r}������rO{�I�J�����I��	C�P$P;x�%ģ� �H�L��[�#�j��d�=���2w��(Jy�^�9	Byߛِ�`�����/�}Yo38�y�d&^� ���ߞw��J�=�ġ(�z��'!)J.��ּխef��	BRs�|�r���7�(JOz�I�J�u���<Й	C�g�k���ټ޵���	��bP����p�'wZ�(JNs�m�%(O��ۜ����f��ԃ+�J�I��R�h�lX��MQ�4՗]lJ���i�J˽`�%\��:��4&�
�#wQ�$቎ԯ���Ru�~m9	C�w�6%)I�}�v���:��^e�oyl�k7�P����NJP�y��%?�A7z�(��XMb���|�8��j� �O>�I�J��]��	��#V쑒�RNP�5H�f��9%'����%	�γ�?d�u��Ӑ�%��e{[�ދ5f�%	I���=�	K�3޳��(JN��ͣ�Wh3Cל�,�DP&�}�l���Tm#���6��JKX�قP�H*YM���Gw9=�Wrg��P����vӐ�'����	I���9	JQy�exҍ�B�"�@F���J"�"�^H%	I��7	Bs3��+��:�e<EDۈ&�(t��� �H�H�}�p��:�;3�5���^����߹�[5o-��Z�ԡ)=�t����u��`��!�I�si�uA��ҽ��	����N���slJ���3��`�ۊ'�"�"����R���~m9	B{ߛؔ%'���r������n�6ї�f�:�`Ю�8�b�Z?ӡ��-��[g N@���ߞN��'����BR}���r��3��(JN}{U�3{��JL��=����JO��I�J����2����Ӑ�%���6j�V��(JO}�C��!:��0JS���y��%	�~obP�={�G��0�y������1J���<�r���7��L�Ւ{�t���c���
5m!@�@����((e䂊��}�n��Z�'�d%'��� �m�` ��3}���s��CBɪ,%�@=T��]��9�ڇ[�!_��v��I���D	�g�&��A�1h�X Ԇ�e�FT��fL0��; �C�5�}Ff	�O.������pkj�-V��3:��������0#���u�I��(�|l�*��<=��}=8G
�=�:{8��sd������"ĸK2�0L0�cc�̃]}ν#{.���q�z��5����n��z��6%�0R@!	�Jy�ޗ��XNٿ�w^�p	6��dkh                         m���!�k�L�/sms��/\V�м��sv���,MH�&]�l���VЕ=�u\��� ���\�K����ml ��::�j�n:��$�5��e��v x�:�;�2Ԇ鍶u�s�������	��.��s��)�z�.T6�+4���P�$1��ٍ=tbFI3�p ֵՒ0�A��n H��#�������UU:*���V-ϓ1�Ē�n���Cg,��@�G+h'�s�`۳��m�����n�
��^��ζ���j捘{:,�@�S�>�~�+v�۱$<ґS2"�k����Tn����sɘ��F�r��k��B�&���(��R���m�e|X(;n�"[{^Mu�p��ss�S���sd��7Pv���thv{D �wV�X�n=�ˇ�+j~��}��nq;�U%�N5�^nE�K�`]ͻzB�g#Q+uí�Fږ�m)9��LQ���6���6��n�+e�W�*��ܰb���8uK� �U����'���vh!�-gb�.�v�NM���7fҀ5��ln4�;Q!m ���TB�t�듶!$w ��0Rͣ�icV�ew`eWn8��S�U�խֲݽ捛T4ǡҜ �'�C�u[V���Ӫ�yK����ܢ�o��v�(v$��vX�K����P��H��$�I$   v�kdע$����`#��1V.����8%{�o���l��3�� ����ɇ;=�fwNd���?X>�v�G�?H��%���4A(!�d�;ޔ���
�k�ڤ��tu:���_s�zƖ�kl��ѓS�tA��	�a���a$���s��W�W�wz�$��{�eu��Һe�6�D�T�kb˫7�_����n�N�"e8�0F|�dP$
��(p�F�o Ԟ��&�(N�֨J�ˮ�ޞN����>���������L��&�(Nu��BP����Ӑ�(nd���U�h^�󌤛�'���<�Z�(J���������N�H(H�hn�t!	-x )L�f��Д%'^��Ӑ��Ϟk{����4���9ֵBP���G���m
˖^����������@�����p�':֨J����Ӑ�9;)~�Y�TH�4l2M[P��x��ࣳ�9ɗ̖�5a ԃ� ��M�t!	2�IP�L��=�'��*���9�(JO{�#�^�f�3��%	��'Q�:~A4�3}�:1>@�&�<��2L�|�r����7�(JO��I�?�I2=�Ƚ��0��7���(JO>���rMI��w��%	I���7	Bs�j��)<������a��ָ�BW�{�6%	I���7	Bs�j��<�N����r��Ϸ�Zٻ7�����BR}�M�P��Z�(JNy׻NBP����&����̼_Ҫq�-��y��xc��G�x�ۂƗ�sӹ��rnG��@�C=hP$P&�r�P����x"0�%'�{��%	h��
QR$(+Hпg%	�<�	��bP��w�p�'3:���X��I� ~�~����Vl�o7���"J߿obPu���~i7��BP�b��:��P���0J	�߯�C�P$ �XF$r%)��b�"�#�Ʉ�v�wn���N��"#:
Q$9�.��P
�U}��o2�w��{�Uv��/.[]�_5k@��۞qrdܑ�����2�{����V�\�f�8���#|�����u_�$��p]��a�!B8��1��-Wv��8E���RnG����i����}ʪ`]Q�4	�B����3y)EQ��^�A��2�q���U��+rH���'S����go<�t�oe�fԥ�]����t��%��r������-�}Ԉ��f�HĎ2[Q��������Y�X �L��Im�%&�೺WH�^OP��wηq�8�+@Ƣ-��,�y��P�e���*�ON�qb7875���8z�s���~� 0TC��~����5	U��k��{    �Kn�N�ۍSZ�۱ŸV7c`[�.��G]�m���Mz�ʑ$B��\]�l��v:����g��F!˕-�#���9U(�:)��7�Ŝ�&�i��W���-�&.� �ͬ�uV3;UvèT'9��rrN��UWbtl�b%Y��������;�;��l����l���lC�U�g�0�k��;�I�q����#M�����^�bUP�=������U��v�WwtA���_��j^rLjG�{�Y�ه�C�n��	����-������*�}�=x�z�d�[�z/c�=5�r�9籇��g2Gcnx�T$by1!��z���$�_ܼ�Ip�@Ƣ)�W����}�  ������ƈ�f��IF$%��ŗ��c�ζ9�	���x!Q��u�[�HI�\�޽0�K�!&썏��#��q#�w<K�2 }ߪ���O<<~Vؖ���Ѥ�CbS���͈Lj���J���k[�V��o�td�H�d�)n=T( �_�j^q������R���uyP>��I�1#i!��ڜ$�섞e���� �X���i�~q惇�S{X ���ل�ܐ�,��V&N��^{����a';��+_���I�#q���cQ6�	7y<xI���:��� ��X�I<����]�3g]L��m�8A1�� =B��l��
3l"�>���}Q�����+��������0��\��O�d�H�7x8I��><<M��#H��#�7!j9m�~�!'�xa'ޱ��R>ݐ��g=%"JG	��R̞0��~�qs>��n��������0Z* "!�_*�<����e^�!��(�܌���	9�!'�mMT�̈y>MҪp.�V[lb�N��3g�H���98��m3l�)�v�}���ځ�{���P���J&�h�������i�'��D����#�F`kX1��c����	9ܐ����/��_���O��
`IDK��xO�T��BO��s����Bv��񄜿Fz	Q��|'���I�]{�p�v�a'��	=�@h��Og<'$��9I9d��1�UUUP  )���6�n#P��N����_���O������2�RGn��Vu��e�t�sl�9Mp���)���b̝���j��n�	�p0j�e�IꦗE�����Vɴt]W*�%��z�`��L�khf�`���.�O$�?�$�hw��35��-4�.
�(���f5YZ��--3o�H���Mۆt��W>�{��1��0�$�p�v�g���}�/��� ������F���ߥ�VHI��]��!%[�\$�#W���%�8Oԇ��B��܂x��	7�;�p��2�s����z��o�''���Y�=~�]U�MYRfPS�GdNwn�ʝ`�����7V�d/���P/�0�ܸ&�v�
b(��)���/��(U*���U�+�wNO�'���I�v���fO0���Ԝ$�ސ�}���{���(y����v�=P݂�2a���=��?y�m�A�(b288IWs��M���nd��פ y��Um�f�K��f��>z&�P��lf).^���q��1��'s�y#��Nw ��\Dݿix�Abl�	>ݓ�l��P�v�a'�pBO��R����.p�+ׄBM۴����6��$�F�o` ��������|||}@?:��15d Z��J��,�� ;RE ���������n'z����8Uv���H��8BM�]�&�\�zM��`��i	6�t�,X�.
u�u��^�� �(�]kg�a�o[q�^�`C��4`pC�B{=r�%�����$�z�"P��Y`&H"H»�ؗ���z`�h�Љ��$ ���8�yu�|ߟ~�.$�G�UZ�E�6!ع��ۧ4�EFҼ�=v-���68����{y�=g��뱵����_�~\�G�I��1��&�m���y��nHx��$$߲I��
�\�⋤�݂w2g7��~d@��+���3[�Q!���K��s�=;��qۗv�8�a�!B8O��͐�R�88I��>����'ۓ�D��M�!o���A8��nR��8����"R9x	�R�##��꼐�M������"{�	�����J8��=X�$H���5�ϯ7o����z��6����o�bH��~~l()�չ�����~��'���M��v�EK^�#�]"��#����\7i3X�
RZĖ���f�з���#ģRZ'��
{�ڄ�e�H6��'�AgY�D[\$޼��P���HI���	k�ا�Z���0#p��	>�HI�d��/Z��[�	7݌7�"�2�Q�R�{�R8��	=��	��÷�N���$�PF�I���I�SZײo�3��ŉt	�*��TMt^��|N�_.�    UU0�+9���*�s�+�Itd]��F�����&��C0��F�e�6[�4,T�:���̝�:��l��I=�Iϥ?���{�~kvz���]5�3u���(l������\1�I��ݝ�N�t�:gH%��k�u�Z}� �P��"����\�I"M�Pr�q���ū���n�콴�x�b�^�l�qs�Q��� ���T^HI��?�6��z�����)G=$�߹É[�	7o�G-�3�B���}���CZe�0BNp���	7o=K���$�l���b%-:�q��I�P�����b�M0��rW}��'6�[MB�=$޼0�w�Ow$ݽ(O��t�M)�j[U��$.EP��pdn�MjbdJf`2�'wgy֏�w�$�?J\��{~�7�D\Q��	7�'� 
U
\�C��~�W��V���wn��y���q�RM�ڒp�w�BO-ᄑ��uv��ސ:���KQ�����[	7y$H�uHI��psR?��?!��&��rv��/V���￫:�z ~��'�����®�L��b�����icN���#�ӭ�Ѥ$$�I9�HI�f�p�}���DNX�':�)Y�C�'8A3T�yo����b'l䜡B�+Ic�B�$���'l�~�Pg�"��B궟�D����������W�y��eK�bgd�g��f~�$�섛��yoL$��0��q���&�d'W«w�$޼0���	'���FQ.(T�ѷ9#�1É<P���-�5-�+����e÷@{�@����i����ޣC�y��m��T:�za'1ᄞ�����I�Y��-�q��O��	=̘7~�{�� ��Z�Dd6�	7�%��3x=�O^}�[�?�N�? ^����=�zpg�0�8D��	9���� ��G@{���ި�}�oUZ�t��ۏ,Zqh�e݌��6���%q5&��`:���<�IWy�{�!&�`�R+�
g��B�𓙲{�!&�鄞+�<(W[7��7��b����{��â|Q=�N��g8�����a��Q�� �fOI=�q$}� <K��	=�s`3��AY�~��=�{��@￶��e�߁���#F������淰    my�K۲�4��lb�u�H l^�`q�\JK�E�3��<Λf�U���:�m��י��.��<�����/����4s9�Y�z.����4��Z��Ͳ��/n�9�]��}l��\�I���U�F�7����rz�B�]P��J��-|����Rgк8�����8n�(�ͦ��<���:!�M�i�p���2{�! �� ����	�Ix�CZCXM��������_?T��A���A,�X�t���BO�%w�qq���	<�"!���68H=Y�n�BOw$'5�I<���Y2��:�\��vBNg���;��$��P�~����nP��糷1��̴D��=��k��ayn	B9H7�IϽ!&�d��~P�w�n����j(�	9�`���EX��@����l,J������L�|%
J�PP�|� �%w�{�!&���!I�)) �'��B	���wroK3�BM�CV9%G�����p�������ܐBRZj��Q��M�	=�A	=��<$��#�wx~�U$�2Me�S�4����������Wa.3b��r�'q�	>̐���!'��D1�j��+��ĊYj{�!'/7����푩�	�d	A�No�$�2o���u�KT�)[-IZ(� 9�9�}ߠ��v|G��m#�R7�!&�`��^A	=���vFư$�Q�8������a'��{� Ԝ���{��m�[���k����ͻs��B�^�ĀĔ�(��I������"{��Y�I�hb�!d�pgSK&ɔ)#o$$��u)��	'H�-��B
.p�{�jF�`��K.I]��	;vc�}�sv�=��y��~|�뺦��W�R��dTu�>o�����R5lp���>J�d=J���P�賮��5�Uڻhf�ٞ3v����q�`�z�����Z�e��=�C�߾��1DO/ �"�x��`�#�:�l��T l�l�{�!'�['*�q�)"�Q(�	7��[�%�������s���lD���!<' �}�	6�T$��/��~PBu|6jZ�Q2cqA�J��8I���H'w�!'��$H��Q����DS�eTS*��G�P"~�����Q��[A(Ŝk�m�����o�<Ҫ��h� ��P�kT���I�BF��0�T�p�%AJUC&$ʹ�Y*͚�A�)H���,E2���BE3 J�(P�#�1�H�&aX�ĳ�� ́�U�"�P�xD&��D�D-� �B�)*�-4� b�%
�IB	B@#@1
R�BV`�d&a�:m�
2�R�P-!IJ� ��д�
4+H- �( fD������TfT��o��f ����e2BB �
P;�z7`��Ph}�qj �E1�E0���!@ܸ*B�6�P(��kH�&���!b h	�)�E���Z�y��+co����?
f/Ys����z�,��;��Щ>om��me�ʪ� ���R��%��"��MU_�T�u��'�,������Y���Ro_��s���/�D\vn��~�"��x���*M��
������_�_����
��;>�����4X����9�/���ۿ���Z��K��%O���_v�W�}��9��1d��
y������?��Mr��믺�>��̬f}�s_��kO���j�㎺��*�>���\}˜�����f?��������!(�ʁ&2���2(
�@ �F�b  �b�VfFH�T�R!d�d%��BYFa��BQ`�HBRa$e���	��f (�V)��2�K&!a�*A �,2�@P#+,�B��HH0Je��U�2J�C��`�����)%�B�$,b�>�+L��o��H	�s��ƭg>ٮ��o��~�'m�1�����H��'YmT���q���/k�~b���|��cc�>���~�����>���P�_-_�m7��~n?ʿ�|�%�?��o���¾?/��n�_������ϕ���������]T�=}8��Y�����f~���}?_�s�~_s���P��}��O�~��>\?E���j};8���s�#��~y�h�ݟ6Y�l���?؊�51��>}K}�t�"�3|���2%O��w[\���k���?.:sU!M���U�>5R��C�G�~_�� ���o�����z��d~�Zϯ����&~w�*�Z���}�UHS���#��'�U!O��R�Ǉ��������?G��
����n��d��>�51���<�2�V��>�9�W������qu�uU!M�i�7��4��=��kٯ������柟��D��|�u��	��8��_���>��?���m~�Ew���*o���AB�K�kc��4q���S��X��X���[�bW�|=��.�p� p��"