BZh91AY&SYL��m��߀pp��b� ����av�   ED U*��� II( (��� /`� � Q@ $R@�x   �IJP�U*R@ �(��HIPI%R( RUJ�R  
�T�QIE�      .     `�
     �=��+=�{j�o�{o>�R�� n*�;�93��Z]n,� �{�V-�8��  >�5J*��� MR������
�-T@ /��b*�ۧ�5yj��(      �@�4N� ɥ�\�:�����qV �&{����n���+�K  �[��r�� ��J���t�� �A���1�,��v��u#� �*����n�ra�s�t�� p�
@  � � �P��a�NF:�-B��x���&>����� ;���p ��h��r�x�=�#-�4�:���H�� g	��ɮ6W�O�p  �  @ =*��ͧc9e]9s�Ox ��.-��g��v�Y�N �N�oyc�ۯ>Χ�xث�  �w���i�6m�5W� 9Vl*��OZ^O����w(�   (    (14 8zVOsS��'B���s�9϶�p�g���x̕�Ү� �2��r��<  ����ت� ���S��aqe�8����U����������O^�>����|M
         =@��U*D�i � �M=M��S�R�@ 2   i�S��Q#ԠF�M2 Ob�R6�� @   ?�2)���*  � dd  !H@�DɑOL*~��Cz������z�"~?�������z���o}�u����@UU����b
���UU?�����U\H� *�����UWW�%�YUU���- *������_��^�!)�r
��0�r���m	u��8�>_��9	ܛ�,{��%o0v����8�K��9h��� 20���Hk�Ѡ����i�����Hy.9	A�ܺz֍=GT���Ե�7k (���jd�X�F.�G;�y߾�r������<KV�3BY�2�kZ�H�^�Ύu�5��8�٠�厹c�7�OVkoO.��0�c�5�<J\r#@d%I0`�!�r�x���r�83�o�s�L��r\u;usz#p����:G7NTjՄ�޻��3��7�aӽ�f�{�l������'z�6��%f.��zӪ',a�Lc��w�zZ�mu==��؜�3J�
r�,i=5��2M�r���n�O'4�+3�X3��NÜ�p=�I:�ܚL̖�6��t�u�o����J:�Fs�7�Nt��I�%�9F��ݠ�o')<�0m��6f����4y�n��	f��<��o���t���}��|�m�����y�zj,t�y��
4sQ���DK%�����֝�?j~��Z�3Zp���o�Ǿ�[3�i���Fo��ތ<#7�:��5�z_/�㌜�y�u��1�V�"NF�����H���1�O�#�����E�����I��Hݛ �Y�������٢#<�z+�<O�T�8��w5�(X�JP)��/&"��X����ܮ�$�-o�&�EN:��~Pb���`:uz����S&��N$���<�P�	BR�%	BP�'!(J��(J��M�������&@e��ԥ��N>�ҍ��7è�%��4δbG5�9�޳�Ύ�a��{'�l�ݲ:ٖT������s9��Y�5�{N'��ь����Nkf�h ���hd&���0�-����z֤��� ���C#ӧ�|�شe֢�22�4�k��!e�����~�-m֯�sӠ2����=%(�u�E~\�B|���oԞLE�Qi5.�uη�Xvp�9zP�a0k$�5&%m�]wΎ��^��78��������CQW����Z��o֯�@��%�-;3EG39�yN��;�)-��Q�j��Ы�;ykV�&|&�MBRx��p��|r4�3�4n�y�h�1ǝN|��
z��y᡻����<߆��3 �q�w�x�=�5�w�]�0cL��Fl�J �%���맮c���A����Ӗf��wD" �l���o���bQ�ہ�a���`3����^�ɯ;3x�$3!)d�.���o�޽�߇s�F��`M0�	��֬��D���0�	BPd�d<��q)w���:<O7�z��L���%퉹�0rPi��$!�0J��5&�"��x�Å����3NKGfd�4�&JcBP�DI	^O7�O=�p�
D�܉L7X��v�G,�2�PvB�:��(�5	�J�CP����9��8kn��f�=޽����
x���gY�.s���cphْ`Y'zN���^s{���Od�h�X6p3V:�)��sxټ5`h�7��yMv���%J2y.P%�ԅ�5@���LV�9�W���*g�#��:1Fŀ��ܚ�]�Q	�Z������[8;q�E@BM0UE�\��CRd�Փ��ֳA�>�5םpΛ��r��1�oDʻаL�*b�`�4�&�<�����J��ĨYSx���~���)�M�a�	�k{�6F���&�a�7�Ӯ͎wC޺�ᇯ7�ӷ�s]��%	Bw)B{&p߃���0kEzz��<��F���`�1��(�_r�$�p��1�u��s���jN��OZq�jĈ�Z��d��#&�v�q-o[���fY��=�u��ގ��7��p4��i�Z�Z�y�5�Y�zf��2*Mյ(r�Ñ?kK�D����Х�_YW@�M+m!yz3]�&&`hwi8�����Pu���;��kI��XoM����j�Й8�"AL�V5M5V�UC�V����]�|��VZ�u��XF��r-녚�xճ��rB	�����8r�)��!�%��S�sږ`�<�HS(�zZ�*$NH��G��RlFOT��3��T��a�X�-�1�*ua$rF��Z�;���\�Y�M���I��n=��V��H���7h77[���a��N���p�c'G��y�]\Ú����l�[�3����a�Awh��B�c�BZqjth<����u3�A��(MK��!�����F������n� �l�Z�l6����ӳLj�q5	`�ދ8��24o#d�q���c����=jv�.=�Á�`�����]��5��kF���&��Fiu	�	[H<��}���N�����r�:ߎf�2,��z��lԙ-�:��o,I�o��v���|;���^�o�u\��}0�z|6(% �P��F�w&&C�����ù�6t��M��w��1��3F����ٱ��U���7�z�n���4Ƶ��#kҔR���ը՞�]
fi8��^�Z����N:�K����B;íu��#L�4F�:;��\�.�f*\�H���'���$\I���(PѦVͬ��4%^�<MUQ�ǽLg��u%繠��N��fV9���gON����pȉ�	r1'��\�̭��٭�h���革l��m��?LJ���ymJ�G�p�fG<#�z���n���N�Z�N�O�e�aI�fa#5	�:��k18NF���,��b�f��zu��Jt�;�A����8[�sU���i�i��oc�4p�ӑ�x�2xka����(J�<7۸3Df��F�1������(����د���in_�9ݭ������Y�3]�uެ:=��8�4����5t󚻳��zEf��噠p�n%	t0P���[�JK��y��)���@����P�a��фn���>����ʳ�!"x�(O�����Hk,C!+Hde&��6��h�8N�2��5ѫ�g+��%@h��(�py�;����n�2�ixuF��9��5A��;X�c���Оɉ���=̈r�m=�b�������Z�u��rK��=���j'X:�c�n+�f�sk4�O(3q���4鷹ٛ
B+FA��7!��m��ya����	��g0K���:�M��n4�g=��&A���I�%.9�P�u�� 0̘hǏF��]9.rrl��0:�|ν��ri2M��c=�%P�c�_���ꢧU�N&�����ߙٻ'^�s8Y���w�iM����7F���P�6�����-F�#f���d�k�����wa�F�כ�]��u�
��th����&�m'!²TPE����Fxo�y�m��̌1c01h��,�sR��^ζ��;�37����y��q��[3���lr��cQ�S;���2q#��e�p�@Y�����u�m�(M�1g�)Z"R�Rȑ�T%�O��ʨ|��h,u''K��'��Z�;3�}:/H�:X��ċ"�3!,�ʰn��Ì�h�,L� �Ic�
�5k/tw��[�h�������N=�c۹�<��]�ۚ5�4�.�փG����;�[��[i?!2ܢS'�<���_*®wȨy[H<�vr*����Ա&�����0�4�D՘cNK[�q�����r�Bu���(N�(}Xm�)��[F�JI���YcI��� ��ʌ��!;�P�%;\�ˮg2M͐�99#"N�� �jt�r��,��@p�b�&�jѷ��Q�Rp5�z���l��
�9&�-�P�Y����̌8u�~q-��&��n�udx�y�c�9��X,�bit���� ���Lzb<)��X�5:u.h�zakI98��wo����I��8��N�;����V[+N�<�AֵGAy�V,d���`iMl����5���BRǝ�� �KDzDP�c���C�~jM=�S����i���=�BR�Lc0ĝBl�������":���n^��\�NjY�xN<��sP�o5�[���3GDOA����#�ᢓ�2�S��]��s�j0ѣ}����9��h��)J��ں�G�ќ7!�h�c�#Z!)G���Ԅ��Mnoa+*��2=܆y��i����2p5�}�Xh#"
��I�My�8nO`�J�֓3�`����l�{�39�|õ���\�~hHmT�C�^��0�����[�kvA��k��î�Qs9ے�'p�	BP�%	BP��	BP�%	BP��r���޳��VlBj��(J��L#@o8k�;�;ֻ���4���떂�!(7A�p���`�h� Ɍ� ���Y':���ގ���!��q��jX�FX�Hf`I�$���Bo1���Ә[7�zS8�8Օ,`X�A��Aw�.��ޱ��V!��&^��Z���s9��4a��LkO��k6�Hw�����20�EN����V(:�����֡���k��ɬ#xg}��(��rNI[�Z����F��)"�{NA)%�ZJ^�,����O:IA>�+����h�mJ���q[<е�(w�{����ks\�8A�y6n0c9�dkk�0��mq��hf{���t�����K
��*j��B�<�����I���!.�lg6jhָc]^o۪�6Db��s��3̺���o��J��G+&�_�d"ZS=����������(2mL��Q1N�dUb�Do]{5��h�s��=N�f�0*3x�4�h0�X��N��c'y��=�ё��2.xp沤��9��j��j�Gz�d00#1�rt�&&f:q��̓I�bq2�g	ލ�E�a�{�BVR�v�B��CQ�͊<q���J�C
c02_;5/nC��I��S;z!�X�h�u����̷�����UUSU5UU P�`m  ]�   �            �      �2˶� �� [E)� ��      � �  ��`�C��#�Y@     7m�
�i5P`9���  �s �6�m   [E��  ��  ` �           0        �          -�  i�� R�������a��l�5�6�{]���Pm��k�y�m��������fj���+�僶:�P���=��9Ǯ���SP渕�iZ����ݮR�8���FM���ڸ�]�vJ.Z�{,ʋŃS�[F��G ;�E����USn���.}/N��������bf�v��۶����6�^�SĖ�e�^�xٻ^�kU��Т�xy5i{n�'F6��g�e��%�=�+��p X����^À���*�` *�mù���;:�Y�
�Ke�$5T 8l��]m`��m� մ,ç6�ʇ��
����]��ՉI9�ϥs�  �M�M�+vi6�knZ 6�T�R�6�Gv���@A&p�Bn��ŲPH���$h�l�P�R� �Q��U[T"ZI�[F��F�i; o��gIzk�mqm �[�.�m��M��Ӂ'-�M-�mt�w  6�Zl��h p�A����  �m�����6�;:λlN�#m��[x p�,;kz�8jt�ie��fZV�m��� N�H���k5+P�uC����i$&�v�ݱ�@�G�pe�z>�����h���A9�Q�E�����6s���3�v� C�"=�n� *�<�@�UU�m����zY[vI��[B���j��PG�2|�i'z���N�d�l�]Vԫ۲�.Z�L�n��n�M�R��m��^����HJ���U]n��7�W�g�e�FdS���&tU�$�*�����uJ��ĽP��GiV�s�����o_Wű�	�mcIYim�Az���P�y�X*�^�j|�UJd��kV�@�݅�E���X�m��/^��h��%����B��E���6��gm%l7�r8#��@�j�j�����P�h-��I�(���+�uڏ��m�ێ�*�U���eC��`��5E���F�QX��V��v�� q�T�
َ�<����j<;ڲ�[��w9�C����cV;\/=[����K�dշ#�-'&��{[(�T��À�,�4��@P J�T�`.�	������!*���'kW5���H�lٶm�l�kuu�m���W �J[@�v�tćKKL�[m㦶0�[n�Ҁ�l�)�Jܠl�[BOKT��pl�$==���6� �@:@8j����I�z��U�t�WJ���m�`n�[�E� �i	����u��Y�"^Z�t�Z�ݞ�vIҶm���kXH��m[%�ש���l�`  ��m&��Z���[J�Z�8��g- 4���P�!����Uaù��V��;��	@�����Hmݰ�&ٛ�v� $!�sk��ɭ�Z��� $n�m"�V)�m��UUR�d^��s�lb��Wrmˬz�3�\�5�㍵h�J�9�l�[y	�GTڕ��\�J˻*���xVTL #�i 3B�.�P�`�cix>Yq��ʖ����턝������ ���:�U�4(UT��k���Vݵ�O���MW�v%�`)@y�����.�EZ�P6ʧi.�Zl[[-6ۖ���H�Π  ��6�*�%�ڗ���<����iƚ�m���j�sl� 6]Qsv��f�e��
���qt��z`M�p[rm��/]n | ���������m&��p� (0` ��8�/^;P�6@b�y22���i�f����i�Pp6Գ��m�G�;ͥu��M�NQm[�Y㮒v�t�Ͷ U��*���	���-$�UU*� �Hm6ͱ���� ݵ��� ��-�'Y�`Gf8�gp��]]u��l	 �l 	N���s�]۪��	I7[��E�I����4�̘ �a��V��F̭Xh�fݝ[Mj�^�*��Ӭ�UKмd�[E�WS����d��P厵.�'{����һGS�7
�\ZÁ0P:�ɻn+��R�em�^����v��z�n���ݎ�に�umf��2�=�6Vګn���*��[����mU�<�5�@^[���.y#g8v�x�VK��n�L��K�v�&�����~���*tK�u0���m�j]�Mm�m�UK9���AX��28��7#�{�V�X�Nݕz[�vp[���(7l9'^�:۪z˶�r�[@S�fjWa��v����g���;I������[l���Y@&���%�ťUz�eZ��ѫil���8�-�[�(Е�֚kv�v]��ev�kl����մ�uHh�*��=U�+vn�U+���(8�2I�M���n�,�� t�M��*��^ڀ�`���H��sknJl���H�ک[9nlm�p)E�lXa �kl�&�l��Vܴm����s���n[ls7!�Hɶ�j�[�I�Ͷ�kn	��  �����H$Ѷ;ͱ�}Amkm���Ē �u۶f�[m���n�i6	�[n$�a ��o;<�:�4 ��q��)# 7m�m��s����=��h�uV�܍�I� V��\�n�큲д�8HݖLHH+���ۤ ��d�� u��a����mDu��z
c��j���R��]]mlKX����  [{I�E���*Ģ�������`)V��Z�e��Vղ�j�[@��m�`���M� m�p�lknZ���ڶ ��l�5l�l���W���>	-����m!! .���$ �� ^m[-�lHm   6�-ɝ� #]����5L�ì�[m�	 $����n�a��$ �ppm�kn�8�m�f�	����m� 6�l�ām[@�$$^�m� h �ݤ�6�q��$���  [ӎ�[A��km�����m�i�(�dT�&��n����  ���i$� �5�Mvݵ�m@*ƅn\�UT9�Ԇٮ5�lT�p!�M�:U���x�����2)*tִ�:KjA�ƶC���l ^�p8��	� %� �t�iV�[q�*�
S����>_ҹ�a���U��s��@  �mٮ�(	z��!�+q���eaI	6i6�n����Ӭ�մ -��.�j�U`%@i�6��8 �E:�88   �Uc��)v���N6Z�m�� A�V�`6����R�T� �S��V��n�  stRۦ�J� 
(��P�R]���f�S��k��M i��I�g3�2��عt�I$2����i�I^�U<�JKp E�%���^%�V�j�@vvwl��A���[BF��m� ��9]�����(6��p���  �m�$Yvۖ�@ �	 8[{m�m5�<���UUm�U<��mٶYLm� �m[JP 	 I� [N�'�ml�d�m�   �� �k�m�i����` �vֺ�91URe8^�Uj�	�F��Lb˱�Rݹ�&����;���`������� ��AJ�WVmZ*���e[.��+P&�]��a��d��� -�gX Imm��p9��$ӡ�fT�[`  �m�-��m[�� �B۲�6��i6k�  ���(M�-�-�m� m&ćm&�6ؑm9 m��]6�H�#j�Hp h-��� ]7amրlӧg���:����m'@�n�Y
 �PM�   z�$ֻ�:���I���  ��M� �    �{e� -����@l�m�� l�m�p�p 	 h�i.�zж� 8��H�`H�m 8	�  �jM�[p �`8[wlH�&�  m�����h� [@ �H[vͳ� [Fٶ� m�h��ٶ����i�{���]� 	nݰk�'@N�h�`i�   V0�`�.�`6�� m[9����mz��I�ݶ���� ڤ��h	��� $X����j��[� p�`�[ZM�.�(��J>үO<�(2t3:�ۈ)����Z�gr��.�.�K\�R�k�~>��xX1ٕ���^jvT.��&�vj��Y25�id�r�۶� �b��0H��m�� [v�-�Kh6� � �m� [@�kn ��v I E��n6�     �h��.�ۦ��һ 5�km�l��Y^��ݽ���-� 	 �`۶�`	 -��a�� ���[pG��m�E��^���,0��� Hm��6͛e�`v�d�6�H�հ `K�$����\lڵַ��{ս�����_㈊������������?�����_�o����"���O誟�?�΍����I@$�(�&���3`�@A��!R� �/��A��)�t  #�4�$��F�A��{�{D�B��)��� :�@A��#0px�
��JtiU�}�d��OU�E �v��׈�tá:'�!�8�G�^ �����҈�����pO"���O4*�}D��p�S��D�T�Dn��@�tT�T�S���4+�z
qP��1�c� R�0XA�!r�z!H!I�<P�T�!B J$!D�P�hM q|T=P�'B������������!��*�q�88���=��D����T�IId <U��=@��� ��$UL���$}�����P<D�A�C��P��v gzT=E�P '���zAm�"hH�����DS�$!E��6Ӏ�O!G�\%�A	5���'`��(y���d�h%`���	d
R����(b:T�a�`x�������H���T2 ��;T^Ƿ��M�P�bv�OW���⾩�
�B	�zx+ő���!��<҈=��oO������'��������k�����"!�8e!)E��3R�C��P�H �(�Pt���b$���:���   m�7�[d��` �l̘��ն��^�8;m��    -� �����~˶�C��b'��1ˎ�\g��1Ȉ8�L㵴�b��A��S�d��t�kj
�K�K�u�����h�J5��]��`q��ckb+w�`�p�3����p.����kk�����P��m�x&�)3U�ֺ;]�Ad�Ŷ��'gU�3���>�vݑ��,i���ʠ$PS���v��,���b]D�d��ٜ7#Ŷ����iM�	@n�$q7e�muµ9-[nc Gps�E<+����l��Z�f���u4��2N�Q��䞴��su�9��]�9���]�|�5��mt�ٴ� �;ume� ���2E�(�^n�W�_`ݚ�;۰8��R��5H��-)g�����Vˬ������������\�y�g�l.���A�μV�ڎ<Xɇ��˻:�zv7c���1�m��q�}ݸ���;������/V��0��P��˴j���<���uЦ���ܲY�nN��rI��A<���zy-��cј ���H���6䐦���ܦ�V��gt<�m�`�pf��{c��VKP�^R�ь���:)[eZU��J���q�<r����U�+�{=6'��1�Wც
U��7.��F�{�ݺ��À���|ܞS�q�I6��X�C��N3�zFWk����2�k# 1ϢR
y�g�d5t�]q˧�]�v�w[��N�	2�Vʣ�m\�v��PJ�<�s�y�����U@PY6�b�Ҹ��y�Rݧ;,�:�v��[�:N�\��v�S�=��v�,����h\;���NK�VPs�-uR�Sɒ^ZCKB�/\=VĽ��ʰv³�-V�sl��9��.Z�� g��m[nvc�ݹ	�#����v]p\:�]��Fy����UV�j�哏
��UT�ck=���^�j_!dM��{N�h+�ݨ'��C�����D;���Ux�Ap���p�S��I�0( ���ꏮ����@ڌ��w�g�j8�.����r1.R3��F�[�n=�3[p��s��X��\�y�On��׀+{vKp�Ěr�{cOnɱV�i9����6���]�.�N���[��o'c7��p/v�ڃm����7j�}vm��d@&����&t��ӻ-�����Mc�;����rtn��u�ی��n�a8���ē�Z��ls����(8��Z7�ЇH��t��7�3XDfwld��sˀ��q�*�xplxy����]�<[��Iϻ��/6$
��T�w:�+��lM ����s�����ϻ�P��:�E��0�L��34�u*67��w��/{���wGx"e9���&F�U�΀ǻ�@��@^�R�5��>��Q娈��@c����/{�P����~q߿��~v6F+��A�<-�t���l����ݩl��vۛͮ��ݦY�[jիm�5�t� �we`y{� ���X�.�ʛ����4�m��o��TbԼ��%�����1��}�{�4�˥Js2C!ˆ���Tlo:�E ^�M{�J���9L62bZ�0&�]�w��/{����@}���+�IM ����t��t�67��w��׆���P+�kv���q�;u�]���ϳ��U��x�^�!�E8a4�d��N������@f��1��P�t����Mմ���v�`_�� ���X��x�vVJ���ξ�Dt�I;v��>/{���iy'���a(1`A�1z;CW��e`_�� 7�yrVĚjդ�k /{����@c��1��P��92�T�lj�M���vV��ܰ��E ^�M�K����|�}�!	�j�RMl�Ӎ�:u��*��X�q�8W�+�����t���I]���@��E�c����/{�P��)��LKS5#56��l�wwv��*�>ԭ����zϊ�V��m�����h��T|�z���_w�@f�qb=0H1�D��{�J�ǻ�@c��u��)��"`B�N+�UU}ilxՒ.�	�i+�ۻ�� ǻ�@c����/{�P5��>��a�Oi�@����
茰�W�j�r�mZ��$��h����V�t�7l��L������/{�|���>�9D����jնƚ��s�7�ب{�=ފ29GD�f��p�m�}ݕ�}~�,%߯�, ��x�˦Bf	dTCr%P}���;��_w�@��@^�R�5��&ӷt�&�-5�}~�,UU��=*�<��r���q$��$����������Kv�k����ݲ6$�m��82��&^a��sZ|ܽn�u�7:�yG�kb��O[�	�m�B�K�0�)^�9��Q+��Nv���r���Nm6����.�gsȏ�YONܼ�՜<F��v�mH	�N�m��p-j�v�d�m3v�͖O>iQ�r��Xן�K��6~���D�;]4;vܠv���Ϋe�]��-�^����=�������9L냏WR��θ��5��\�?�v�o�����+GE,nl� ;m��������^��߀ǻ�@gGq`
`�c��������΀ǻ�@��@g���!��
&e�2���t=ފ ��}ݕ�z�y���v퍴��_�w�@�}4�u*y,��t��<�J�WJնƚ��s�7��X����ǻ�@}�䗱j���"ff ���+�牻b��8��r]�ޱϋ����ύٱ7jt�I7��Lvƭ$�o@������x��r��V�t� '�F��;WW�����Uw��?��;@��SI{ދ-�TPw�M{�J���j\�"`4=ފ ����� >����⻑C-��lM���I$�w�M��Ԩ3zh{��w6�&)�Z&fh��T��4=ފ ������[�h-�^۞�s��Cv��g�+�f{=��u<��@y�O�DL�D(���ʠ��1��P�t��Ԩf���B��-�i��}~�,�_���>� ������<}^�֮�M]ӵt�k 7��|��=�� �����3����˼��^�E�����+CV�m��o����� ��z(�h��L���,P�J���1��P�t��Ԩ�G���Ff�O���<72gGe�xy�vt��#��=;rN��|��������;f&h{�{�4�u* �ޚY�]ȡ���&���s�7��Xlo:�E���	�O��D��{�J�͍�@c����3��ߊmR�I�wm����~���_���Uu��� ��PL���r������ҷn��M���ܰ	UO;�����Tlo: �s���,Q
v������[��6{h�v�t��ɣ�s�t��ٳ�C��t'S?m��������΀ǻ�@fG(��b�4�M6��vVJ�v{�K�=}�`~�X�us`����$� ͍�@c��-�tP�Ԩzo)��e�dP�]o7�����@^oR�3cy�ŧt�����3���z��΀���@bߩ���򣶺l��k��j�S������^W�n���(=dۤ�l��ܶ��q=n8捸�ё�6DwQj������Ѥ{g�ⱶ��>s�����m�y6u�.�WZmG0�^*��9�݉���lB��2fZ��:�X^ѵ��L�N�t�g'��qk71�Fܺ$b��y�'[GF�X�۳��֦K'���l���I�Ε4�N�q���4q?*� t��+����fDdo0��v؊�i.v]'[F5�u:�0[�Իb���K�r���t]�$�
�hk��{�+ ��y��z({�{�{�L�"LK��Tlo:�oEo{���ޥ@z�~��M
ݻcm7x���m��(�y/$�o}J�ގ���=*���Ըjf%���-�tP�Ԩ��t���}��\�'j�v��M���{�PoO|�{�Eo�����M�j ����.���̮�[nm���f��Lqۓn�Z�m����պ�d�N/.�7|�o:�oEo���^^���*��JcAt7B��JӼo�r�����!�u&�� C��y�u�f�*v7����С�G03*"&(}���Ԩ��t�ފ7y��	�L��D�P�Ԩ��t�ފ�wE�����A-Ī����G����ot����߂~,E)Fݠ��aNxu���t��[\g؎܎��ۛ٘��'-����Z�&mi�}���Y�җgoR�}қ�"Ijb��n&=۝Գ{�.�ޥ��G�Y���t��e�I&���H���ؿ������N-{���d'_�?o�<^�k�C.m]�<ڟ�H�С�U�tB�?��;�<>Ok�>�{�A�)����o��zZ���Ɵf��/�SA�x�����"T�1
z�P���ި.�8�ؙگc�[���D�C�Rx9��gE���BE&'Z��;#^�$�,\4���2�"l��=����!x�fà��G��$PI⋣Z��e�M�H
��6p�Bi�����GNפ!q&äG���y�v�n�1�������MG���~��OQ;Sb�����b��� �� h�G�5��mҩ�/��><��:��qJR��<��R����oe�y�kۭ[�Z��)J<�߸=JR�g�}�JRy��}��������G�(|����{�f�[��wz�8=JR�g�}�)JRy��}����߾��)J<�߸'R��3�3"���n���*j
��&*������-fL���f�c����y'�=�j��kZ޺@�);�����(߾���(}��~��J{�}���)I��C�(�*Bj��vvԕ� �����>��߸=JR�g�ߵ�݁��l�;�;��*N1PT���o-�g�(}��~��)J{�}���)I�����JS߾���);��uL�)�B��(����g�݁ݶSn�JRu��}��R�����(I��2�FL��䄦���0�V��t
����{��>]��>��ԩ�(����f�l���)I�����JC��c���fwZ�[3��v���A�0Ll�X��X�v�y3�
y\JeGІ4YV�n�\t�m�\��J�k���{ݷ�߿Ͼ��)J<�߸=JR����┤;{䕳������eT3�%4ζqJR��>��R���}�8�)N��%l�;�;����݁݁�{MMU3E��o7�|��|��)J{��s�R�����pz��=��qJR��>��R�����ϴF�[���fo|R�����ԥ)��}ÊR�>y��pz��=���)JN���3�5}��o[��|�)O~��R���$�����)O�~��)JRy��}��R����m��?��j�"�D��UP3��ԑ譬=�OF�J����v	����Y÷�ٞ-���0�y���ųR�d��&�����*x8.������=�u��K�1ѳ���8��g����>�9:2=.����&b,�3�{��>w]>��uf����v
�n;b���*`��/-����,=�㶑Y�춲+�;���ml���+��m�eK{���{��߻����#U/k�!x��nx��2������`QOSG�q�cq�:ֵ�,���3y��l�JR���}��ԥ)�}��┥'����O�*�R���u���;�;v�$�0ST�STQWswv=JR���}�)JRy��}��R��%mn���[���w`wo%J�b�����Xoz�f��)JR{��}��R�����)J>�߸=JR���}�)J��y4ʦ��j"$�������w`wm_}ÊR�>y��pz��=Ͼ�\R�o|��|��^L��������d��kg�(|��~��)@U'�~��\R����߿pz��=��qJR������?��ob<l-�6�=[`�)�����@�el��s��p��o��]��ESU�U]������	)�vvo|���)J{��p┥�{���)E�������
�i���vvm�%c�m~bz1N��a�:������)J>��=JR���}�)�Us����a�e��Q��o7��z�v]�mn���[���vnvQ˵�)JO�����JS�+�~�kya�o{սl┥�{���)Os�~��)=����)J{��p┥,��$�b��`�j�*�����w`wm��k�R�����pz��=�߸qJR�Ͻ��R�������j�XZ����]<��N��c�G�f���y�z7fE��6��f�\j�M\�^oJu0S���o{��}��߸=JR����8�)C�����@wmS�-݁݁�：eSME5T�ͽo|�)O~��R����}��ԥ)����┥'�����)K�~>������xf�ѳZ��)JP������R���{�qJ|��c��	��&�Q&T����rs����ԥ)߾�ÊR�?y�����M��TU5\T��>���w`w`vߒV=JR�}��8�#C�����JS흖��,M T�D�E��;�;o�+g�J���}���R�>�����)vJuE��;�;s��%�i�"��&"*��]�x�on����<Zގ}�ndUColq�k�8�P��=��D@�ė<EMEM[?û�w.��R�>}�pz��>�^��V���䕳�����4z6U44D�LUT�4qJR�Ͻ��Q�S%?~�߳�R����σ��%��ݜ���d�E��k-��n�9���)O~׿g�)=����J{��p┥�{���)O>��lַkF��Z�{����R4����pz��=�߸qJR�Ͻ��R�">���@�+��>@ ��>����3�R��}料���4n�ݽkZ�o{��)J{��p┥!߿{��JSߵ���)JO=��=^�m�v������^xư���+6(�vI�:|uB؏p��%��S�@�:�����]�2k[��͹�f���R���߽��ԥ)����┥'�����JS߽��v}Zjj�ir*�*��.j�v=�^���JR{���pz��>���R���߽���!J}����F���o[�[�qJR��|��R���k߳�P	C߿{��JS����)JN����2��}Nf������R�>�^��R����=��ԥ)�����'�IL��?}��ԥ)��߷���l�Yk{ս�┥�y���(�	�����R�����~��)J}���┥'��4~}���{�;���j͛�T��Ö�=��-+Om�C�W�mpV�ۓ�[k���{n��nyq^6��st��P��ێE�6��v
�
�����`K-����>d�n:4V��1�{P\�i�݇��pd�f5���8(��v����{jmC�w7^�'��m-���;�w�V�-N�f����ZMͱ��8x�q�;L�;r�y�V2r6�%�׌�m�b�*|"��Ѽ���k,��̎��{h��H���s�'X���-2veٵg��Vu1׏�%��h���kﾾ������o{���~�)JR{�����R���w����)C��~���R������oZ3n�j7�n��8�)I�{��JS߽���(|��~��)J{���8�)I��M*�ʨ�����*f��vvZ�[qJR�ϼ��R����ﳊR����l�;�;��2������h��j���8�/��!���~��)J{��~�)JR{�����R��߾��)J����{Ѧ���f�k��o��)O}��g�)N��߸=JR�}����)C�~{�;߭�v��~��p~3=:g�pu1���\	�N;���\�"m㧶��r�ס���y���֭�������8�)I��{��JSϾ���(}��~�=JR�����)JRw���S����ޭk[��)Jy������i�����=N��R�}����)O=׿g�)��[>����G�UST�TNkw�(}��~��)J{��8�"4�}�pz��<��qJR����M*b��b��������|���vR�wjR�����R���}�)H P���l�;�;��j�����z�F�����R����=��ԥ"�}��8�)C�~{��JS�u���)JN�#���1k9�v6JKs��W�p�8�&n�n����\ls�l�d����{��>�EF�5<=JR�}��8�)C�~{��JSݔ�ݝ���{U�������eU1F��oۚ7Z��)JP�ߞ���?
�(d��k��┥'����JS�&VUU���~�6�~-�wm��i��JS�u���)JN��߸=Ht҉ $��q�A ��"A#!	,AT�R�0� ����;����ˊR�>}��=JR����}բ�u[��5���
N��߸=JR�}����)C�~{��J�u���)JO��"�RL�[>����JP��pz��=�_}�R���{U��������$i��j	n�Gs`��x�/�i�Z�73ɉ�B�.�9�}�su,DESMQ14[��>��V�ԥ)���┥'_y��^�)O>��n����ƴ�b��b��������z��=�_}�R����=��ԥ)�ʑn�����[>�����fje����oz7��qJR�����R���}��)O�X\��=���JS��~��Vvo��ULLIS351Ul�;�(}���┥�����)O���g�13�R<��a�4m��x>I�7�\�)K�>>������xf�j٬��)JP�ߞ���R��?uwE��;�;}ں��w`wd�"��=������}���!��̖;1��XK�܃��g/Kֱ��\m���)o^��������Oi�{w�ٜ�k|��)J}���8�)I��{��JS������JP��u�������=<Q1,@U5Qn�JRu����� �>���qJR�����R���kﳀ(Ҕ���م��j��3z��o�ԥ)��o�R�>��pz� )O~��g�):��~��)Jvg���³5��e���kw���(�d?y�߸=JR�~����)JN��߸=JP~�߹�������&������Zj�����|ؔ��}�qJR��
�����)O�~��R�>��pz��6z"y�����	#A&���N^�� pt�K3��%���h0�������fS�8���x��a�^��}���u,,-�:���q��D�m��I�|$Il5��o̜����`r"h
�I(I$� )i�ǧXP=oQ�'p�URF[8�;u�s��tP��`�݌,2E(˽H�A,��0�p�@]2C	�;9����M��j�i����bg}��� �E�k��gB���ǃ�]�x t=�^\÷k�8�4G}	�J��	*�� Xt��pZv@�g��i�����4���,�u��b�]�1�+͠�:;z�0�%V؜4r�3�ߎ �s@�.�>׷���ofjַ��   ���1n�  �m�9@m�6`ӭc����    -� �o��_��u�����#��Aa��X.��a�#d�l���\�l��9Xg�u�,���Uw4�;v�S�:�H��qv��ݵ�l���F��Kq����=�$7g;6�����.�f��-���t�U�����8�Ɵ緱���\�¯DuXx����;�O/)uj^�ոKWL�pk���H��8Qe��vs4�1r	�N��@ݹ�k9���n^�mCX6�z�� �[.Ζ{�0.�;!'�#
�n"���M2N͐N��q�c]<JHN����i���Y�;�5��;6�����?;��Z]ݷg���Ǩz�m�0D�(-�'Z�NwRҽU�O�Ҷ����.-�!��,Y��`�&�fG���||�8��Gl4��+Ս���5�j�6:8gm��,]'8LY�>��k vlq�Hqn�u�]�6a粟.����=�L�/3a��Y�Ǜ��p�r���dpLM�u��뵭����2�"�3�L�[�'Es���6��Hˤ&6�����s�;�AR������z�N�\#����@�d��*���k�� �n�Ph`\l���fպ�Z
ZU�lb��vX�U��At+9{�X:(�S�W)X�*V��h�Dt=��5<r�� b ik �uq��k����w8)-v��=�]�́��K�����uZ*D�uٴͫ�X�C��z��d�P��ݍ
jR����M�kuL崻D�a�A��]��l���v*�$Y�֑��R�pP��콝�bY4v� e����M�,F1S�=���7l�\7+]W�'\�r\sR�V�V�t��	$�E���nі�ݸ�H�\�pjڝ��4N�:9��&
-�(���Юm�;n�Zyz2b7D�@���iѻ5"���ԥ�r�T������oh
�c�2Nv+]&��f[4�f���� ��-�(|2?>�C�<V^�j��Q'�(��z�a�@����Tz�cp���U<mV����ͮ������(����g���hհml&�z��[Px�+�O��Pę�J�&��KI��n�<�/q;pc1�\����..�Ro"f ��Lȝ=�^���i��NY1ڐ5K.y���]�8� ۃV�GGGt+uW��u��&���R�\=��ڌ�Z�7d�bE��j���c<n��Rj��;5��{��J ~@z蹝kZ��6a�7՛ћm����P,=;�Y�ɶ�t��v���d����{�[빙��������*������z��R�����)J{�߸�R���i(�vvo��iULQSEL��SV�ԥ)��o�%({�߿pz��>��߳�R��w�pz�iK�~>��[ַ��u�z�{��)C�~{��JSߵ���)�����R���}��)JP�痿ލ6��z���s[��J��}�qJR�����R���}��)@]����)OO����k5�-+{�f��┥']����)~�\R���=��ԥ)����┥'�uy_fDd}�Fl¬���F�x�g�j\��n ��-�	Ҏ�]e�u�g=�����⏃9��9�-o|�)O~�\R���=��ԥ)�����~2R��>]l�;�3y�GuD�MSLMמ{�:��L=` b�F�:%�ȘJ���vb���JVŁ��Y�jT�vg��kL�k��b���1�f��Ix��7J��:G ���{�)6�+��Sb��E�;��՘�H�}�W���������^�t�����[J�m��4X�{�j�T�|�f �����R�B.w]M��2�չ*=lZ�zN���nM�囉$��,ڬ��t�w�٫�_m�� ���E%����@�0��қT�?ͷFbO3@褼�U@g�V`�"�=��^s3C�@�uD��i�%@ӱ7x���۠t�}^����vkwf��z� ^�Q`|�aD@�DTU�����˺��v�����=G��t�꾹Av���t�3 7�� ��]׀{�t��s}��}�����L�v�1��V	�v�M�6.q�Fۑ�b��]l��8���h&ǯfh��wޓt�� >��{�)6�+��Sb�����Y���H���^�R�wfｭ*:�'m1���Ot�� >��~���K�;�I��*6R�n���*H�,9�gvh;uu���,���ǊJ�2?H Ă�`�A����o��Uy���i�iz��*������5JQ`s<33�����wW ��W�|̉4�Y�4����;c��2��	h���ȩ����dg;�w��z�������>�b�Y�jT� �{U�����(�>��D8�T0��Y�$������L�$R^��n����>��Q���tZ��� �{�h)/�~�6{��G~��J��ة6=�y��33�)E��ڳ IR,�~���'�r�J�T؊lT�w�l�M�?�~���� ^�׀%)E��3]C�p������"�pLgтf����4��q������5�0�89�n�ex:��i��"�UI��d�Kné��5���30hMY7�����NOcZ�X����R�Ccg�L��Yn|Ks��gn^� ��WS�Ԑ3ٮ:8�s80��nm��0�]�]����c�{s���#���\������P���q#;��YWg8�vF��N�u�m������{���{�{]��(�+ێMGn�0����w1v���}r����Zas�is&z��-���m2�Vշ��}���� ;�t�)J?1���ـ	suP��1�%4�Q`��胺{���w�0�"ݘ��Jؿ;o���̵���K�7���� 7�����Gj�,J��v���o��t	#� o��4
d�(�>Ka��PP<E4EV`	*E�����uu�t�E���f�!JH�KڳN3��za�DX�n'iݞ^��-�v�9��rIx�v�=�t��K�vZf }���K�7�&��H�}�_RP���b������E%�figww���n,�T� �wU�3���4��i�����(j�Z��,���H�UA�wL�$R^�u_G`;N�e���Ot�RG ���4	�a���;�|��0.n������������,����9����0��f ��`W�\�nJM�ؙN�@�p7k`�h�5����9[]$Ź�%U�-����}�j�����<ĳ3@�Ix��t	#�W���J�*�զX�m���ĵfs�;�3C334�\X�]xR�[��8$j�qᨨa�)�f�*���ʯ{�߹���%ܠ
��*@�2�K@�JB@z+�@��kﳕ{��}�Uw���HĈ�p�X�J$�����JR�<�f;�;�37w_�Bd���n�!&ǭffh)/ +�ꪭ��xJ�`�u^���	�a�{Z�7n�c�y�[	�]9�%�84�.ӈ�gFmce�>�B̙�V�'s�$������T� �n�wvf�����kF��;nݱ��I=�$���U o���	JQ`g�Vg;3C34\�MT�MT�K�SLU��׀%)E����Y�I0�Wt��_�O�i�����)J,���%H���wggl}aS���9o}{�:���}���[��M�i�����I0ﻦh	JQ`s�h����fb�y
�j`%�.� Z���w[X|g�^D�8���j��7��_o�g���x�h����,>�W�%)F~�7����Q0.�)]��-3 >�u^���{�f�R/�ٙ�xyBi�h���`��+*n����{�f������^��S0�62�v��w����M�:G ߻�h��}:���wmڶ[J�IR,�=�� �)E���Y�]=�o_����͂.:4�3P�	v��>�6�9��x9�etf�<�v�\.n�E�A����u>����I�NTrs��<e����\[٨��s�ۄJ]J���qv��o\��n�哜ܻN�u��dMOM����:��5ŵ�S9u�����=X{�c�5=���شa�-�m�<�N�ܥ�ζ����l�kc� ��(�c jv}_�{���wwso���W88��֘z��o]qg]b8ی��On�S�v"-Oj�{����ԝ&�����i� �����tR^ﻦ��	$x�t��_�O�i���������۫0$��3�U��<A����Q14AUTEME��K� J��3�U�	JQ`}����PP<EASY�;�%V���Ù�v��.�Ѫzh""hj�"b��,�-W�;:R�X�j�%H�9���e������1ڑ���]ѻh�]�R�7�.�1�+6�vmt�m�6�۰�t�Ӳ�_T���t�E��T�gg �Ӧh�/-4��C(mګM��M�P����f;���d�E�gf�;����]xR�[;�3��GA��+e���Ot	#� {��4�vvaٝٚ��}˳ ���`���ڻ_��Vـ�t�E%��t�ٙ��%H�|�S1/S4�SMq5w�%)E�;�������"�=���u"�+cN�$�˻c��j�vW�/i"���ٻu����������`^���s��*�jӻ�@[n�x{�n�$p�|�_�3;;����=�`{�G��1��ݍ=�$��L�$R^�f�fwh=�����i�"f*�"���.�T�Ky����0� ΐI!Fzq9�z��vtg�p-fTŅ�ŔfBx�x]�·���ͦζE><ѶS8��Qk�<�uR�؜Y$&5��;eX��)�Q�bh��̃.�� ��y�o};���p���;�0�h���C�ON]�O�xl��H�j�����!{@�F$�p�WQ�K�q�����D|D8)�X�{��A� D�#��:�N�W�W�� z�:�h�{
��oЪ�t���N���������`�����hlz�ff�UU����}:n��8`��3@��&��he�Ui��6zM�+�ꮑ� >�j�T��?��tptI�4Q(J��-s�8{�V��[�|v�k�����1�1���7W�йmF�-=��~����� �{U��(�|vwx�{� P�����t�n��N��`{�f�"��Z�`	*E��; o�ژ��z����h����)J,Z�a�;��A��ŀzI�����4&Yhmݴ��U;1�۫0�"�3�J���wfdX�t�����}��߽��&pݸa�*
��R�X���g����'@fw}v��g͈P@���- 7m��c��G�/��4v��J���#�W���x�w{���y�0Wm���+n��0}�3@褋�V3�;3`�"���֕-T�&Ƕ�fh��}�t��p����+�UUPwu9I���j�7�n��5*E��;��}� �)E�Ӫ�Ci2�$���@���~��� 7�I�E%�}u�J��Mն�_�4[f oޓ4
�U�������u�^����W¼ 	�Q�"d0��@��v���'���Kv�.�CU+�!2׎����qn�;:u��a�n�Hl��&�ql.�	<�-u��m��CR3n�B�y�n��3̝������N�����8��\����o]nTy�n�1�u��'5��=�h��B�x2tl:�V�v�;p;����m�\s�E�U�^��XMk�Y�1���N�!Ìcs�N��]�n[Vz\r���-�����n�w�{ﾹ�����W\�-X佶5�\#�=c�U��=Z�R�we�;��_}����U4�d�]�7�X}�Y�jT� Ͻ&hQEQڴ�-Qm��N�{�3J�`�J�R�[ ��({��]��=�:G ߤ��tR^�{��_�6�Wm�.Ҷ�� 7�&h��}�I�H�o��EH�c@�c�O34�K�>����p���3@%�6���];bE�Mn�=�:����;Y�̛8��:ͻr�X�=,�ԎnM7t�e�Ui��>����p���3@褼�p�t6�.��Jݽ��^�����["P��D|E�����4�p�>����.T�n��-��n�0�zL�=�� ��ttp��H+n���6������_G�t��{�~��4�R�;V�jՖ�t�f��&���{�f��{ ���<|)b~Lʅ���Lu�㬤V6�iҎ�]�ܗ!x9�`�Q��u�^�vZ{�{�� }�I��8`}�n��΍�]�;���t[f }�I��8`}�n�����ƭ�d�QYWw�{U"���K0��fc��*Sbp�%T�qr10RS1!��ٙ�=���^J����jj���P۴�ـ}�I��8`����{��ӸQ�vۥli%n��ܩ�����H�>�R�wS�[C�s����kP��k�u�Ĺ�<kG&���[-����r��W������`>����0��7@�G ߤ���Վ���w�Ǚ�{��~�>����0�zL�$�.�J�,h-��fh�>�R�ک�������H����q�(�"����ݽ��e]���s�����r�t��� �9����t+�N�v�N�l���}VI-���ﾻ{���/5�?��L�l�4o6͎�`��n�5�'�6ܯs��\Ύ�8�׸��o�4��kWWw�{U"���K0j�~;3������'T�m't��v��0��7y�����ŀ{w��j�_39 �"�i�I�$��{�t�� }�I��8`}�7@�ʹQ�I�wj�����`�y+�=��`}���fvx��ŀ{��4�UQ4�SQd�]��"���՘�H����;�34�3C;1�$�"F*Ɉ�&������������h�(SV��4�J�l��=W����rVȸlp�]��1�Kf��n9�k�|<���0Ht�T�V�Y��Y�p��kli^ss��m�z�˶�u��C�;fRˑk���������jg�e��d�=t�H}�]��mm�rX�"�'��49��֞
k�9��`��e��P����nڷ���Q�l<���m�F�֒˻\���wn�:ܽ�v���Wm[�ݣuԼS�.`������:�������#���ݫ-�Ҵ���M�:G �z+�5*E��D%�@��Uf�R/�����uq`}��������N�v�N�l�����p�>��n��8`T��ƭ�bM�m;��5*E��۫0J�a�����n�f�:���i;��P۵V�0�jT� �y+�5*E���bb8{��^�&��6h+���k:ֹ�؜�r���ݫOBm�Ұg�r步�J�7�� ��� �y+�5*G3;3���f �SO5<��QO35E�g��徻�ʐ��x��\���r�}����� >�HRm��'����3@��n�Ù�uq`n�^ �����Ln��bf���tH��t��8`�ܗ�(aN�i]���p�{�f��0��7@����F�^e,A�7=���që�������z�(��l�ۈB̀(��d.���qm���4��oӦ��� ��WU­��]���&�4��oӦ��� =��f���*�N����%�j�>Z� IR,�n݆a��b	%`�'���/u��s�����'�Q:Mզ4��i�$p�}�W�$�{���654�S��V�䝦� �ӦhG�t��I0�8�JNZ�&�Hl�����`�X�v|Z^(�DA��:f�-�}}��ű?ͧx%���� ��&�I��zt��T��+I��lBL�=���I[X�Z� IR,�(� b�����&� ԕ��}���gh��\X�ݘѺ�h	�ji	�����kp��U��"��ږ`&gka؅�C�����CΑW�S�?g���=]���[�v�c�Y���H�:�˺� ]�V������xߘ���e���'��k��&���<�� �b^Ә�nm�F�e��}N�:�Y'Aj�l�=�I�E%�ޝ3@�0��q�I5V��Jݷ�E%��~�����׀.����ږg<A��C�����i�Cm� {���h#�Q�M�:)/ 7���m��'���-f^;;B�,���T�yj�ܪ_�����j�f�M�:$��>��x�H�<�p0�;3��f�R���g���EFXoݵ�GJ��h�xh���|�Rvl��N.�ɟ �(�3�)�"H���ғ�D����{��e�D�s�<|2����z|�z���{6�I�fx�yз�j�������Z@i�Y�S�BHf*�پ��]�n�0"}C�뷁�v)Xh�Yn���N��t���'ΐ�\��A�%�	9ۮ0ɹp4�i[�X!+=��Ҟ��H�$;�A�g0:�S�����*0M���$�� ՅE7�)��:�:����S`   m�m&�i7
P ��6��( �t� �6��m�l    m� ;+T�i�m�l�ZU{$��U��ж��St��AѴtc��Q��j;Nۨ.�%1sr��3+��D��Ve3���9k���+��ԗg�NΜ�v]�<�l݇�Sm]t�1��];��D�	W��v�")�f��^���҉���u�'\c�C��:��T�mּ֭��8[z��L��i���V\�;A����q���/!Wd:`�ye�`�5����<����t�¨���4W;Ur�v��6�S���+;�R]��(�s:6��VA���:B�ʒ�:�rv2kѺ������;��<��N$�m'����dxF�����Jgn�҅#6惇t�����P	ej�4pJ�F�����68;1�ױ�KդͣX^C"��B���MX�� �ϭ�n�>�w'��c��y܊t��/gN�ܳ��FNr��;8�D�w��GIog�&nU�ZnJ�)]��vD���<��67/����u�^ۍ�.xf�uq��Cl.$�X�5ЗMFP��m��m&pv���3u�٠)ݔ�]m.�7VO5�F۬�b�1�st����E53��T�t��s^,�����i�I�Z�����9� 
���KaG+��b�jWv� �6nЮ����P%��5c�՚$6x'u�N4�n�;�������v�ء���Z��\�!�
G��Hnze���72�N�g��.c��)�e��0Ԫ�	Y�[ԖQ%������@�4�8���D�EP�#�q����/1�MB�7*/kX�v\`���iy�V�5:�B���\��J���6%YYX�:xMY�v�(��@<�]R�Q*�F�N$)JA�[h!�H�:4Y@�-��u;*�̭i�.�ch��[k��p䭦���V��$Q[(���j����e���%v*Vz�)E^V +X�5ix�Bu�N�y-��x���7�D:S}���������Ҡz�@���x!�W���^�v[ֵ�dj�$q	�(Ty^qm�8`5ǵ��f��#Ѹl��`]�'[�f{nn��=8l�	���3X�<�ɳv��!�I��p�ݎj�m�β��i�v�U���E������˺�F|7Yi8�n{nc���m�iH:��)9)[ ^�v�wBn�Ѹ'i{U��I�h,=�;i�Ś�+��*��lVq��Lg��t1�����{ƴ���7;�y��N�u0z�Щ��y\�6���^����n�;���U�
vU�Zs@�Ix��K�5*G6@o�v`�����j�B"[����ޝ3@�0}�n��Iw��ͼ&� ������+"n���\`�������N��w��m'`ӿ�N�6ـ{�t�K��:f��8`'
�i;�Li%cot�K��t��p�=ޓt	gD��ma�mi���O[��=�[�:�VƱ���c��C�vⵙ�\��� �ܺ���Z� ԩ��g7��6�oW95T�OU4�d���	*E����ɞ]6a�3 �S`j�y�����C�I3D�IUTI3E��{� P�� ��L�$��Ig��SJ�5w5���=�6�˯ IR,o���;�&�tՖ��$� }Ӧh$p�=ޓt	rE�}^�d,�]"Ψlzy^��\B�WNw�v���V�9�f�oo30�eeګe�[Jě����$���f �%<͌� yr��;z���j��⪢Z���=�K3�ݙ���� ��׀$��jZ4ª��Zb�`���$��>ժ�vv�|�pЂɋ6(�&p����o��w��7@���JuiZj�ݦ�i���U_��#˗^��Ł��Y�(IM�g� �ڤ��6�^	ff�$p�=ޓt	rE�t�\�Aq&4[��
��c������<Z;���f�^�t<��{n{��nq��m�͢�;��t����$��n�.H��3@�8`�YC��J�Wi�.H��3@�8`�I��z����j�����fjl˗^ ��Y���0��4Q��*b�b&j�ț��vx����սـ(Ik��?#�O%�.��ΰGR�̙���ɾ}����oRj���&��v�����n�.H��:f�$�X�����:�L�=D4C1- =m�m��x��ڽݹ�;qٓF�u���UO$v���������"�*������j�H�{�&��r	N��M]۴�mUM�o���fgf�;���7���$� {�%MP�?�&%���� �wM�%� w�L�=K�t����$�Ӻn�.H�zI��� ��(
���T�����`�+�T�ۺ� �xg�a��	H%X�hi��Z����w��vqt��P�ƛ����`[�8�H$scd`y�ܘ�rl��K��'V�;^Ec���n:B�N��]=��]��tƹƎYOi���8܊������;Z��c�3�!�[n�m��R���(�� �=:t�ru*�"lΒ��'M��^s���4Q�L��nY��[d:\������v(��K��Mv�\F�v��,���{��ζ�7o	'b-�`-�^�U0=��gqV�7R)��&��C�rXwm�[��-&��k�N��� �zM��K�,x��rݦ��D��7wxR�_;�3�A�{� ����j��wwh�����j�i�����j���5ov`
Sbw�=��JR�3��jP�}�o�f�"����n��.�MP��j�ݫ��M`�I��K�;���"�>��B��i�-�n�1�I]�à��gs�as������l�G6�/O�滙߇��tv|�E�� ���ڳ P��wv�����7���I�i�����&���{Ve��<����-�xR�_;D�ssD1AD̴��Uf���`���)/ �{��Y�v��l1ZjĦ�Ù�>���{���{V`
S`}�r�ݵvұ4=����$R^��M�%� l�����F�+wN��å���o-�
�y絪'��ry^y�{pִ�E2um�Iմ�tӿ�N�4���t�\�`�I��K�>�J7v��bb�*k0�(�gh�������}�Y�������bfj`�&"�jj,�������glfg�fhv(��X��Ru&S����vf�d�۝j�0zyE�}��1ST�2�n�/f����R^��M�$R^ l���z*�Ph��;Jۧwm�����Ҕ��1y+����������q��7F��3ǋȼu����������aWu.�n	ƀ�'��7ckk+̅Y�%)E�b�W�%)E�;����>�v"TATLML3Q`���;�3<A�=�`-�ـ%)E�3���Q��SS0MIYww�wOtX�j�E%��I��r��˦��v���,ݍ��f ����^�?����I$���y���w���?�r����\%��n��@��E%�ߪ��Wݽ�����ڳ [��-��(�I��r��EY�<�k���F�p�q��rv��������Qug�9�Y
�c��~���(�7�Վ�R�X�V1T�4���:���h)/ �{��)"�1y+�wggxh7���&"���&*�b"�,��0�(��� ��������'��]�U�+Bj��*E%�/%xR�Xs333�-��`�(��i�&&����/%x;wWt`yv`	JQ`f������3�P?��"D$`�ITIBZ�p$XX�H��O7�?�G�V0��n�iIݶk��u=��Ƌ.txgux���ۍ��<浸��w�k��|�k�e����/fy-�:5�c����k��+�s��r��xK��ћn�:��S��:J�;Q��v����S6�W$���ιV�b�ɓ��ͣ��WG#��p�L�����vd�U]f���$�n�������@v�J�5���/�m�`'s����w�ڶ�W�ؕ+t�]�R	��̘뭼��`y|��w1^ۮ5�gq���a		M5%l]���<���-Y�%)E�yzL�'��v�t�����SM�ޝ7@�Ix��3@�Ix�P���v��t+v	��$R^ zzL�$R^ޝ7@��Tb�E$˶+��4� ==&h)/ �N��H������Bm���lu����$R^ޝ7@�Ix��3@���qI~%�N�J���}�H1�f��k�`��R&���
�d'������v�'hm�Wi�ޝ7@�Ix��3@�Ix�](�`ĕ&�'�U������C/r��p��'���#>�X�)E��fs�4A���!��:v�i��\���@�IxzN��H��x�m'v��hw�3�"��I�t	��u���	�%3�EC�MD�MTXKV`�����]р(\���(�9���11L�����s�6G�.n8�r��y(��Ӳm-�v�'�]n[�/z�S{]�6k��������65j�)J; 7�v`�����y�"(������cV��ghh;��,�]�������������"Jh��������Z���eN������4��$�bXLa	6�z4PA�	����)g7*f4N5DA	D�r8������I$QLE<��l1��` �I	�''���36 ��5i^lv�m�#P�&8��,@bXX��h�Ji��z����A1&���7��/�K�9��"��j�"\��b�%,�&!�jW&`�1Bp�	�%�w��G�1{w�]�f�Z�1���ʱ��2.��#����7�kDwMUZ�v1��@�6 �&�G���qB�UЩ���"Gh���� 9�@��x����:�*�:H�ER�KJۤ��"Ӽ��n�.H�r��"���.�QmAS-3Y�(IM�����9t�t�E��� ��3
�����b&�(9�gn};ykm���ջ=���)�[c�m؝�X�CBwi�WJ�m�$��;�tZ�K�==&ց.H���#-�I��մQws�%)E���ݘGwM����iA<��%wM��[N�4����t	rE�w��	��wT/�:e:t+v&��.H���"���a=� F\ȅB��:� �e!��v����z�ު��z}�T�$˶+���xyN�@�Ix��� I*�9�پi4m�jbG�$���7sp�q7<���K���%�F�&��6{�姞�1u�%�:�=�2O��~�W�zzM�	$xyN�@�U.��V�7v��Ym���7J�I�S��	JQ|�{��\45LD�S15�wW�V���������Y�}tw]�v]*acii�yN�@�%���xfv~�,�c�H�����Z*J#*�p�(�9ٽ����wuuʽ�^}�������@�#P�� SA��L�\������g�G[	��n	��6a�l�87C4�&z���U������)��Z�� ۡ�9y]lu�V���`|�KC7�k�����N����p0;1v�|��krk'P�;N�v�{ml��6c�9�:�`R�G4��,��m�D��s�a��77k6MY�j�죺|/YR�v̎�9�2R�.pc�����l�r��ۗ�`���Fӵ���w=�׹�v��n_��`�:ڵ���Ս���`�5/hg�Z�4n.ݳ�u��߽���yCM�6���n�6����7@�R,��)�v�B]6��u1SCU:���H�{��Z_tXڵfs;��3��<	O7Q-2�4DQ1M1TX�{� ��SgDyr��=�\X�����������h"�pww}�԰�t��0��G�z*�J]�n����&��t��U~��p�:�������.�J�I�W��)6�R�cS���P�8��<���-��s�V�EI���(�c�Z-�I��_�#�67T�d�.�a���Z�-�Z�5��{������Z�*R�&�ڰ���<zj�w�E�{���8`�E�nݻHM��fc�:���='Mҿ~��G�N�@�RP�wM��n���m`~�ܻ���Ł�����7T�	2#Z:e:t+v	��>�� 듣�:���:N��}gDwm]�;�E�C��g1h�;�^`��>4[v�HxD��=����IRL�b�n��`rtz_tXI�hH�w��<��ݖ�-�/-f= �tx���0����]K�
J����C��o ��7@�߷��`K� cb���ԯ�N�@;��B�]�E���EDL�`j�X�ԧ =��Ý��ܻ��6]=CMAU2DM�u)�9�5.�ܻ� �U"��fv}m���n�Þ��f�����ld�պ�p[Vݎ�q�R��w���;�+9q��sZ��x� �?���n��G���@�RP�e:j须I6���n�tp�;�H��������ӧB�`���yI����=:M�%��*J��]�]�J�0�N {uU��f���@vf��acaڻ?:6r<Bv�����.A<�?� vZ(�쵍��� �Գ �*E���������<�:H�b��h������Zŷb[�Y�{?��s�;w�8�qgњ���v�rۥ��$�������ک�u)�gwc�K���xk�?��.��	[V���yt�@=���^Գ<���2���!��fd"Z��r� ��h}���>��}"�J�wb���R�z����I��8`Q�Α�˥�~v��v�m��t�p�>��= ���,S����JPR�}������� 8�&���]�G����s���(ųlf�:Ź�%-s�����r��R�6�[�7�7<�93fd���\�Ԏ3Ct'r�=-X�����"B�;t�Լ9�vCٌ��m��������=��h�vB�:n4]6�z��<�zywJd��vx��ix��v�L�â�6�8����� ^q���YA
Q���j6X���w��w���?X���A��s��pgGG$���n�&�$c�;��n�#��X���)����hz8`\��wtx{��\���]%(�b�n�ـ}s�z�������R/�����`TDL�PM�U� $���K0�gg��uq`˺���D4�SQU5U15V����˻���ŀ%�^ �$��ʥ���c�Z�ZOt	#� I�f�.H�	:M�=P�.�*�bv5�1q��6ª���d�Cӌu�#�}��5��͔�Vb���n�Qc��Zf I�f�.H�	:M�$��"�J�ڤ��by��"ϿW�j��L�t	9� $�3@�](i���e;SU6Z�`	*E��r�����Z�"�*������&�09���� ����$��[�f���Za�SL�Ա5E�/$� �q������?��@�8`�u$���T�M6۫��*���������ʤ�b4.M�g�]*z����?��3
)6]�E�f&�f�.H�	�&�G ��f�.��K�[t�i6����n��;�J�`�+�$� ߡQT��v;v�V�I�$p����աN�b8��tU~e](h��� �t�����WS�	X� �Azcm	(s���㻳4��?C2w�z����Y�(���	����M �� ��f�.H�	�&�G~�D$Xۻ&Ǫ.��	)�9�ߒ�������Gr��V�ղ���������nH�r,ܺ�t���鴳�:u��֘3��:s�e;t�k ��n�$p�	�&W����	rE�I*���n�n�7�J�|� �w^���`|�,�fg�.�i��戊b&&���,ow^ �R�wvv<�,��E���j�i���۳o3@��,Ӥ�tp��W$}��;��
��}3@�Ժ��[t�i7J�m`�&��� w�L�%� ���Ŋ��nq��<{s�Y�Ռ�>��h��i�T�]��.���î<!�H�������_��o�+�jSn����R�G����(��L��t�_H��&���UW�߀ߺ(���v*M�U���K���n�:8`zt�yt��n���E�m���n�5R,}����ٺ{�l�ȉ��4�7B�`��H��I��&�Wy��uW����J<H�|�0|y
b&��C>����R�i$�-�,g2z�5��3�8!$äwD���C�|�1���������bgM%k0��M$�Ѩ��;ᙛSp��p.sZh�w���8M1؇`�� �׉8��=.haâ$�3�4j0w�\̵AAE-%�N�� U[#:҇�q��N��A�D�eL�Ah��v<����*�a�ү0WbkLh��yߜ���t	�ӉD�16���ѐX��Y��Rc��X��w$����tv$�OX+։�)"d��K�JR�/���D�8偖e�@a�c���d�9�IT�E�F�'���n�JO;,q��O���H<�yÂtH��8�g�Lm<�Ӡ�����@q|�Q��JZZh�
�����$M�:�*H�<�~���Xg;	 �0�/l���߷~��,�~˦�   �n���	n� ��  [�6�c��3m��   m [V���7�%�]V�P����`�����ѡ�d��Zx�,'a��� ��kT��E�Fv��!�E�5]vQ4����=�鶪g�"a\cU��]�r��Ό6�l�m']�n3��S�9u9�Kd�]�ъ�p��S�6�E�t�cc�(�;Z�����yz�r�'HG:*����q[�V8��.�j���7�v�h�`;wWk%\��t��7S�L�G[s�m¢��0늝�&ֲ�y�������6t��m���Smg=��5��e ����8�n�OK�C��1�r���9�퓌SDuܦ�ơ
g�]�ࢺ��4�O2�vd�m]Ie7����n�=�5]�b47e�uÊ��keg���_B޳8�*��\�K����$ ���ʉ�"c��Z�;v7���q&x����:��K�k,q���:�n��65O��F-��kA
�r���ʪDmۋ��am�W�u<�c=S��u;�l �`�ݱq<�9Â���]8��if��k�WWQ��`%i���T��smF���wiݞ�v:�j��{K�d�e���M�-׷)z�4�Ԁ��Ҡ+�S�V��3�̏Q��e�t����(r�z�.l�kh&�t �)�^��c�`�,��Gv�ΓK�cDh1�U㇂g]�Qǣ�<��qȁvA��+����9j:�� ]T��;A�Q���D�P]��Q���t�(�Vؤ++N�2���v#@A<9�FFvU溺��*��(�!�6�n��c�b�m��f�vfܼ�l�5݂��`��m�ghs�tv`gf1��j�1,��J�*��@��S"�V�Xm\�R�f�J�f�yZ��R�]�*fWf�����;+l\K'-\6�8 �i��<��m�Vx� ����F��E]N�d٪�CF��m����Vcnv6��v��`ņ�����(���)�TP�"m��S8�Q(�%TE $(R+$"�4̍PR���BT0�� h;>���M�'~�]�����?���e-�����J��&��{5cC��Ъv�Bs�$z[v(sNWc��a��9ļu�γ�On�n�G��Ob��7;.��F�^�8�4������l�n�lJ�;����ܤ*㌁���ڞY�D+RZ�2���'G���\\Bv�t�VF���R���՜�uq1�o1��s��n\v�9�Xݺ��i{l��(�-��ݮ��׻��������=<�Ż<�r����kI��]�xΗ�8��׶�sr��ʼ�]�!&�M��t�\�`=&���U�I0��LN�����Ř�4	)�1y,�T� �n��ٙ��]t��!�Mұ���&�G �t��K�,}
��]4�	ELL�`	*E�o�+�$��ݝ��I��q-��(��L���	)�>I,�T��:�:���<N�6�>v�� n��Ov9��vm�_U[�ϧ:ۜW��x����N�3�k�~�����>I,�T�wgl�]׀v�������	!�j���$��;�@	|���g+|�\ _-W�(IM�; �]D�r���ba�&�@�8`wt�\�`$��u�J���wn����6`wt�\�`$��~��8`��?��b*�����BJlo�����,wu^���tP��`n�%�������\�U'i͛��s�v��Z]������߮�7N�制��n��5�}��������7}��پ����5p�<�5Jڴ��G ��L�%��t�+�U�t�EZw@[
i�`{�s��Ͼ�\��	�O!I`X!�����ݙ�ww��Y�|��`g�	I�UKMQY3Uw��=�6�˳ IR,8fgh�׀v��*�^����]4��6N��I0��3@�$X��J.��&���U�j��;9��^]�gţ�r��j�X�Z�O�m�]����?>�e7B�`��H����"�fl���v`
t��G5DS$�KTX�^s;3��A���`}ܻ0�"�W�ߨ��G�ScjӢ۳���%Ħ�ĵf���ŀ%�� P��[t�i6����6N��I0�Ͼ�U�OM��U�[��r�{�>�J�.Ɲ�ջ���G ����K�,�:n���RW��j�v��ݝ���l�t��@�-�<
=k�S�rm�m�E.F�'v���L��I��$�%�������3�R�	���	i�+&j��	)�wvf�=ܻ0�(�{���x���	��)r�>��*��ĵf ��Y����Iu��� ��*&��Sb�`��H����	)�ggcK0��-2К����&���,wR��{�pwwu�_}���W�xlH��:�
A�q����?��sa����MT�x1�!��Έ��m�Z�M�͹�	�����<@u�=��6��]��u�Ǘ�V`9�Z!���筰iq�3Q]�Qȗ��5�r»��4W�t�Nʋ��ۣ�����U=���-I�箻9��X��{Q��'[[�q�mkI��Q�α�5�8�ԗ:ݭ���۳�ܖ�4���n99'��qj$�U�%-c����l!�n'�P>�p���s��{k���ώ����ѥ�!�3&�i��t�b]LET17v�����<�Y�$���t�k@�]u��[t�i6����<�Y�$��K P���w�>\2�憈����&*"f� �����n�l��"�6t��K��t�E]�)ڢ�0�t��%�����T�� ߎ����
�c����	rE�w����;���>�K �ffvhnѠX����G\Oq�[�dcۇ�zs�b��C�1l�5��Î�uvz���g�:�=SU8���%H�3�Ռ�(IM���*�w�m�ح�&�@�8e��ߨ�ZA{�\��� ��Eٚ��ٌ}���tw)�3}�0���*�N�E��M���mh��f�������}>�V�SMQLE;i�h� ��M�$�����%�]t����v�hV�X�~�RG{�mh� �t��i+���Ϸg�u
��E��
����O.|l.�wA�Z�*H��Wn8",$~�[o��H�3}� P��7ڳ Q�L�<���vS�E�`�鵧��.H��t�tp�7㤲�t6��Г�ھ�~�\��<��P�@H��IФU ,��h$�H@��z?� a�����Uן�6�z�JwI��ںt�;m`�t�tp�7�鵠K���*&��cb`[{�N���6�	}"�>��7@�WW�-����wWJʶ�[W��|��� �9/u�l�ݯ���Z���������T�� ߽&ց/�X�{������#�SCt�:v&���jSi������`}������� WR�K�V�1�m�[M`zO��'G}�Z����%]�lv�WS35����]��۽����V�|L����Wc�B���u�}�b�t�wWn�bB�� �zM� ���V`jV�;3�3�n�qo��bv���	��^���ܯm�9㜒q���{u�Kק�,1���vy�9o� Ժ�����>ԭ�����j�l ����wI��h�I;m�~�M�>�2���6������Tm��T��rṛ�3���y��� �呂���t	s��U�E�E��T�:�7�t����h���^��P��T�	�t�7cm�� ��<~�M�=�X��Z�~�,mZ��~v]�6���J�r�pg0�rl��Јu�9 �ָ�7g���!\�r��ud���v������[�ɻmmI�<�rU��3p�<o<y����[/Wm�jHێ[C�Z��=-G�m���n��4f͆5�vۙT�6�ݝ�М���O��ͨ/ݻi���U3;�@sWW2��.�n)��EՔZ����j�t>.N2�ˬ:�z���{{���mX�;x+cdn�JF�ׁݺ�ٚ���;?��]��w�Gu�������m����i��O����+ Ͻ��3��� {{���!��h�(��մ�{�}$��7�t��� ߽�3�.뗊*!��i(�	�k�j�l ��Vt;<}ڻ0wu����ɢ�(I��{Z���=�t��X}�Z=Wҝ�i�)�N�o ����%����@vo}j�;{�7����θ�g����S��N����>�ݵ��O<��h�u�w$�Gj�wU>�֬��{�w���;�t��zG�l�M�%��8N>C�C���c�Tf�֮W�+� v	`N�4�SN�$��2� 5YX�&#�8+�����O+�~�|��<�f�%m|��л���J�*i���
������1{Va������^����l!�T�T�UPT�U�;���v��ou���{V6 -�V�F�*���ݡ���zL���M� ���^՘3���: a�&	�F�X��{M�ɞv��;'4F�Ǯ�u���lj7H�w<oםٝ��^*���*F�f�*��^���;��6{���e`��*���Rb���րN������X}�6����_��gJwN�T��:I��ʻ��~몾��r���_�]}8���A$ȇ�q�#[�e����\��a03�}�b��v9��0�E/p��e	m�ԐDCk��A=PC�N��a��k[��[#��8�C
\�K�f����|6� �rz�s��a!����Z�"�)�@�$�AVC�I���u��!��郦#�`�%::�Q�=W�ڽ0x�=}T �4>��v��}�<��C�d�Sa�=\yb�^P����K�����`�}4��Tn�T��n�I�ޓ+ �&րyj�gfs��Y�(݆�h��T�I�e�X}�6�ӣ�>��zL�߿�����a�]��M�P4����'��iq$��v�XL��e�ҧ^ɉ���4��n��yZ���Ot��&V~����zM���p��n��m�I7`|��3�� [�m`/ov6 yj�{��]�lun�����2�	�鍃�0�U`/�,�>Ԯ^*�x"�j&j"��9�;R� 7{��_jY���Pd�A8D� ]����t�T���
�44&��ޑ����ݫ��w���^Ա��yJ�WGS�l�ݱ��q��Ka�ZN��m��r�uN㓯HZ�7!������*x�I��&V=�mh�#�=�UP�-EQ1QY�{�[_;���� 7{��^Գ9�ݙ��P���D�55SM5�ڗc`��Y������w��V��IYM;lmӤݍ4�c�J��K0y+kn���6+���6�:V��'�M�=�2�W����Uy��o�|(�}U%BaOpQ��;a6B��=�˦����CU*X�6�<��d�q�4קv���T8#�h��k�5[r�{mk��u���Qc��ҳ9����L�=�kq9�����6a��u*Pm@;��9�H�Ԭ���3��c��uF۰��vHs��되�n�"
��o<�.��JMv<��s�t&��1��u���pp�W;��`�p��ⱈ�l�u�J6�n�$%���ɲu�1��礻���{�=�w}�o�A����܏>���m���W.ۡ,$��L���fu�'a8MW`�[X�$�����V;�mh�#���I��&/֝_�-����n�	��k@=�>�n��I��}$�V;`�
���Ok@=�>�n���X�鵠,�N��iۺlm[m��&���X�鵠� ��*7t��cb�wv����X�wt��zG�O���N�X��
�E�V�vyY;n�����t��$��yN$ǓF���P벣�]+�	0Ҷ�B�� ��6��J�������u�������5EV͚��޷����>�|ք~ �D,]��Z^^��L./�7�Powִ���+n��mҥi�}�n��%mg3;�4Gj]����`/!J"�*)����bk09��7z��;R�l ��x�����N�e1�v��OwM� ��x���ގ{�~~f��r� ��h�:`-q�%�6�"��;j7�ݝ�ܷ\rN��2X��%V�R��T�wf|���k@'����Ӷ��M��m�}�fs;�4A��Ł۫���J�������uT5MTLTDT�`�\X��?�g�F� �b�"=�w�`r�Y�(M����&&jjj���Ý�;R� 7{��_jY�{ʑ`z礬�llm�v%m�h�#�_y+�=�H��� O��I0:cFy���&�����Ksسc�uHt�[��kѻ9�1�m�]EM�#_m�?���n��G{�6�ޑ��.ʸ*)�&b�bk0yR/�����]����`/��g334A��4MCP55T�n���y*��K0y+kjL�j
�%��"�fk�7{���ov`�V����0;4�CK�U$$J0%� IIFV��C������gU^��#�6Scj�o �zM�?�~�U�ݍ�v��l ���Yy��*����&�;]J���8wW:����y:[��c�ٻ�����i�W��N�*ح��O4zL�{�6�ޑ��I��]t�J�
�4�b�� ��M� ��x��n��I��z������Cc�;o+@=��_y,Ý���x7{���]��u׮)[t��n�+M��I��+k{ڱ�9��#R�9q��@�[���i��I��_���+@=�*�_y,�>�v�Jɕ5UM35LX�Ip6Ӥ�':ΜYף��r�ۧu]7gN�������N_�7��ΧqLD��y���3�h�*�m��pj���Q�.��`�\g)��I[��͞��k\<N1��)���8�9�.M���n�.���W��b���<� r;i�aRѺ��1��$���	c��v�u������'�Qw[�T�k
Ǳ,������{�w��{��;�'"b��X�g�zŻ.5�{S�Wnxz����u�lGP��7e-��qv֜������wUX�%������@{�����bZ&��bZjb*&f��wU_;3;�������m`/{V6 yl������o �zM�>�e`�鵠� ��F�;l�`ݗU�ڕ����c`�UX;��{V`�u�T�J�i�Г�Ot���U`%�Y�|�����C' ����E*u�Y]�@ݽp�b��S����m��	�j�I�ĳ0)'N�$ؚ-�yZ���	{V`$������ P� i��������&��Kڳ>a��wjg�)%m`%䱰wU_;�3D��� ���������=���^Ս�3;���{��%�'wEl�N�9��;�ẁ�U���f34yWt`�P�NƨT��v�{Z�����0�R�/j��9���F���%r���Зd��F=p�l^v=�&���h��mӗ>u�}�}�=�tL�"���;�v`F�6^Ռ��uM�=
��:i;�`ݖ���Ɂ���k@=�U`%�Y���3��0����i���������l ��U��㳳���Ad�`	",�"����Ν����x� �jS`|�Q�±:v
���yZ�tx����Ùٝ�gvfv��]��t2�p4�SQUUT���U���f�ޕ�8v�� �tx�r.�J�'i�)~_���u��猛���Bǩ�]��y\v� ]���6Z�*H�N��.���L���_H�Ot��� �M�:Ke�]U�`[����>��X���}�E�o}v?���g�=�����*%�Zjb*b&���tw~M���ـ}	)��,l ^�SKMv؛k�W��_���t�I�U�}�GU��
A�i?
�J��xm�!��f��������^>�mh~�	��t���Gl�trn[,��su���r���7v�>�Q�^n����/n�s������%��o�TXwV33;>�Q`{�}%'N�]�c�6���x���t�}$��%�_i�m������n���:��ٝ�_$����x��e�.���L���E��	��k@�� ��7@�r��m�v�� �I6���	��z��>��*�O�lC��WC��t�-)�����`�Bql1Ij'9��1Y�	,�L������@�q����:��a/|7�a�Ƈ4@;3hf�7�XM�da�$0#bj�؆�C�Pl�`�i�N����6u�_C�Q����̅z�*#�f�g����N��9�qM[�ovkq����l\�a���Rz�jdN���X9�Ă	�f ��#�)��^��g3j���Έ"�ptD[�(GY�;y���&S@F'f�)S��?��AxFB|�n��&�&���۱�M%AZ�*��#���"< �h6T��#�{/M4�ʣpAAHw�BiE�f@`A���dY'52՘f"� atmV��	��@d�	�UALl��vhu��[�ӏV��{S��w�_������=�����F�   p6�����Jk�� $m� ��e�3m�8�ݶ[r  ���-� �jغ�򎵓�L]lM���Z휻�:��5@t�u�$�S����{|�ݛu=��@]]�s���Q�	��=��_}b��`Z���T�*
��!���]�q4�DwEm�Xf��!���GV��$tZ9Ǧ�[��;��[�9��7Yڹ6�b��w�ѥ��I�u�6#�$�'B�-�uI�sr@n1n�wX[��\�9y�����vl�ev���+��;1�m��M�I��*�4-i{��4 dz�rjr�zM�Q�u����]��,��We;!.��t�vk��Z×�]�g���[�m��	�{;B�����B��t�z�d��LpC�U�/tJ���]�j�ǭf�Qm�*+%�W�z
tY�CUe@>Ŭ�M��uڕveD�l�,Z^��t�>y�c]3�N+�Hk�
8��mz:��Yz�m������/i�cr��V�Ό����]�Ͷ):�(��g�0�h��&ٛ����2Ô�ع�#Eȳlkgm/,n�s-k�ɫ�{sF�j������[�3-��n���[WJ�ʹ���uXzwC���u%���M+e���Uv1N�dZ��b�}ϕ�^�AM,V�4��N���r�]�傕h
�ۖ��Ǎ�Ƥ��ʌE�@��R��2H��Wo6T�d�.���]+�ź}7[rx�7I��HShD��yܤj��2�ۧ�7GkƗZ˶�T�f���T���=�9M/9WiWi�;�.ڤ8S��������b��TspLuٖ�W$Ryz��2f��̭d�ZI�q-^�"N��ڞ`�f8Nc�z
�U�> �ڗ�����qZ!(�Uca���;5[mUvQ�հR��PNl���kK�l�*��8��4�`��mҫ�	��_B	��jC��1�pja���Cu+|Ѻf��&�[n�5���`�g��gm�:�
M��[F+�����}��~��$v�="h}U"	��UM"�C�h�	�z�� y����i^���39淼5���3z�hِ5 v��!��Y�0'u'*����+nՆ��*�I�=}6���2��Y']ә�O/';�����cy����s�l��NƔ���F囨�=���RgE+�Qշ�M�ݼ�3Э�,z0�=I��Fy	{�\�3��...zb��u�zۆ�ڡ@ۋ�ֲ���Tk��4f�'*pc������1��rݷ\�ظ(R\hm������{۫�nߢ�نݻQ]�^ێV�s�l�v�X�s.6�]�j;lF`�����U6�
ձ�Z�cj�y_�;�`����%��&րw��j��ӱݻ���'wM�;�K�'�M��:,�ߨ	]�H˧M7t0n�ot���%���vwv����`rK� P���	T�]&�lM;�'�M��:,wt��~�)/ ���JN���uE5Um�z��;�]��-���M��v���7lmU��i؋I�o�.<�nNz���Eێ�'��������p�y�E]6��dm��"�Z���t��	��k@�΋ �����n���-'�yI�� ���2*N�v=}��lr���fh��Q�4UD@RL�X����=T�wV`�%����V�vҵWcj�{Z��<�lIv`�J,9�٣���6 N���jݻh�C�n�	��t��	��k@�΋ �Q/�.S��c��+8p���v�Ob�1�[�m�q��{S�n:�;��mH�"�eӦ��`����%��&ց�W�'wM�%��BU(�i���*���_jX�������.��.�})E��F��k�j����������69t�۫0���S<3�����m�`�&s��>�U�~��GU{
�V���n�-5������t��	�I��z�E�w�J���]	&ZOt��	�I��z�E�OwM�;��좬
���P�V;����x��lvO�t���֓l6*�79�}�{��~����U�w`4�'x����=s��'���r���tt+V�IU�ڴ�ց��S}v�ـyOtX�K �CCt�hHmۻm�{�n��)/��W�}�mh��	^�;�;He�n�ot�Ix����=}�`/ߗ���ʿ~��l�h�D��B�M�۶�,����3����uM���� �e(�=�껖L`��@�Z�ڻN��q�Nl�v#�0�&���9���_���w��M�t�LM�h��	��ܤ�}�mh�E
�V���n�-5�Ow,�fvfv�<��,����=�m�����'*�t���$�I��)/ ��M���>���I�e�~�˻���}�Z��,}}�K�7��ЭXݤ"�m]���z���gwu��^��Q`/�� �g�����Ƿ{�{���]�B�K�� rF�B�>&t;�]V/A-MmG]
u�ӷκ�<h��;L�����X.n�e"�	X��z2�8ܝug�$�}�����n�1�ď'A
�F��pc�wFL��X�p�"��Үy�:���q�.�A�3ue]5��`��<q����}����T�i��`6W*v��N�k!Ҽ�����m�ɳ�s�F�"M��]��ۻ�Ώo��4���+,Cd�#p�(O��.��9q����׌���U�V���l�Hmۻm�����r��	��mh�tX��Etwtؐ�CtMV`zR��wv������]6�ڳ9� �L�X&x&!���������wߋV��7��:>�����P��$��Ιi�h�tX��n���Qa�ܻ��9Kt��MD�UUM2L�P���`f��:���Ձ�{�--ߛ�~���<Z�b�#a��2U�q�EC��3;�����e��6�-�en-=�>����mh�tX��7@�\�����e�Гw�}ޓkUS���_��&��`wI��R^��bcv7i'��z��`w��?����=�`yov6 }퉑S�Q2UTTD�X�I7@��K�=�I��z��`_&UD5T��%UEMf��(�9ݝ�w{�o����`}�K0�SC"ZBӎ�+'랤/l�	hªq n9����P�M�ڛ�:�;^�+/�����I��z��`}$� ��>]%ebt�Ce:M'��}~�}$� ���N�Z�U������$$��}�]Uw��o��!I�X�H�r�;��C;v���侾��6)�>BR���i�hbfi�f� >Ԫ����lѺ�Ù��}��`�S�Q �TAEASU`{�V6�� ��M��� �qV�m�T\rN���h��W
��xR�]�r������8u��a���ٴp�B7�[o�����=�K0�sd�+� 5(�'�*�"d�������$�9�����Vwg�u�E�u}(���I[v�� �H�};!�u�E�{ޓt	�*�**��i��������gwv�{��lB]6����fha���f%���յ_�d��	�����ӰI6��]۫lcuM���Y�$���y,l���{�ߚ�����v]����Y�H���Ƃ97T�t�Oc5��k��)��u{\uf��t��Z���� �H���ڟ���&,��vQt��ВtZ{�D���y,lcuM���Y��wOt�C�����m���mh}�`�I�����%��vR���v�=�cuM���Y�$�Þ<�ẁjVп�;��v�X�t��,~U�0��6���;3����+��:�I�H��p����O�Q�)vqt��P���Y���g-ݴevO1�g%���=�������֬����מwI�ާ���1Ԃ<�I�G]7m9�ώ=`�{8 #���9�s�<H�jnUMۖ�6v��[X��˂�'6�m&;y��W��z��h��z��.�`y��b����1G��4�sJ���byx��,�k<u�O���-���V�]�%�w���~��Wc}��ߪu�ɠ��r`v�e�u���ݒZ��d�sw4G\<ݺ���a�4����7嶌cuM���Y�K��X�hm�Ӷ��N�h}�`���$X�ut����+M��;Y������M�>�"�7�d4�](u���t��X��t��@�wt��m�Х.��twD@�ҷ`$�	=�>�"�7�d4��w�n���ĥ�@�e���˧Gg�m�ms�f��:�܂�j�۬d��m����<�R]�����[k@�t��=~�,ٽT��;�8i��q2C���^���z
�H�C(C )L�0�BH��� �>;C��`����m��$����.ջ�v�XN�۠}}"�7�d4_tXW�Etwlj�j��*k0�R�5m� �n���ի��?�TK��n�ݡ��M�������(���ǿ}��o#Ø�Bd��βk+��V�t:�.���D��Ѷ��\3W4��fVV'N�Zt����4_�,�}~�`Ӳ�WJ_���$Zk �{��_�X�솀}�>%�weJ݀�t$�@����]{�����\{��KXh ��RP��D9]0�C0:
H�t$��>J|'a	��8�*�I�F��аA���v��J<�A���{�a���1�g���g�Yp �]�O���a����̢}^��G�q��{�"�i��gS2��I��O3������ކ;�=��{��5��+�LV' %�(����ĂZ΂�x
v@RoN��@d�.[O;y< �z�;S��2�ל6
xo`q�[o�x����'���}).	���!��H���OS�����:�$�p�֥��
��LOQC�t��6"f���gvfr�X�%��R�!�����������q�K�������wff�J]6�GsT�EM@�35A56�;���{�1�}��}j���7�o��%���m�#�+�6,��SۋqH�T�m�Dm�nhָ \۵`H��m������vC���<������5I5hm�=�>�����txw�n���Bݺwv��m6��6I6������t�tX�ut��N��I���7���U`n��>��l���f�a�ޡ��'6�����
��<��~���ًbv�N�]���t���vC 7ڪ���H���i����J���uy��ɟa\[HG)��ۮG��ll[ko',�etN���I�
ӫI����������\�� ���.��h���"�"�lKm������v`G���ˣ���*j��&�&��cWM��}~�a�F�K@�u�G�n�&j
�����vx^K��=�6%���~�W�G
!�U���������Ķрz=�l�j��A�#�B`@c}ϳ��oxj��� \��J��f�.�M����]�O<f_Pc@���<X�8Nul,sj=;`���r�"��Wv��f�us�زm�]�cr���ҁ;p��s�WeLr��/c�KF�
�eѰb۫��)�n����F:�ݰnY�5���;���x���ݱ6ӳ��)t&�Mȭ�����ג8���۲q��+�S�<�ذ���,U8�h�	�cww�?�w{������$�{on|�:˘�e�%�)�܏#wF7n���kc'Y��"f�v��Ur۠�ET�3��o��=�6�f�y)�G.�R��,"&%���iX�����wuf�y)�1*J3�ݢ��1MTMEUM4�S`$�f�y)��#��|`}?�>:仰.�v���{�}Jl�IF����ww=��0)HWWvS���uv��7��z����M�>�"�6�qe
*�ZwA�'iN����xN�2.$�(v�8z�9��f����v�1Ӳĕ��z����wt��,z9/@�sJ:e�]�v=�����ʼ��~��3ڨ8���fwgjvvi*))�>�IF��������D1��ұ�4�@�� ޏ��}�`�t���%V���i��k �K�:���;��t�H�	��遉ӰI�t��/@�� *��~�W�}	)�1mj����Ҧ:H���y۬:��WuDq��1�5v�s�i�On�|���8Sϒ����6��T܀������0�%6-�Q�nΨ�ƩE�Eҷ`+N�Ot�H����t���7J����Wue���vYm����ϖ�0��S~;�㻎;h`��*H���U? ��5���0�ޛ��I����h�������4���}}rE�o�M���(�ݶ��7m4����n������ ߤ�Zr�x��}wW)ա����y���4��������n��.�fM���:\Z��=���5
�C~�[o�� ߤ�Zr�x�z��('j�v��m���7�&ցܺ^�{���G�U@O���N��N����yZr�x��M��� ߧM��U҇aM��m:Wv����n�}'��]w��tu\�T�!\���2�DGh����\�_g*�ϱJ* ���bi�f� >IU�������S`��,�ڳ �vgd�2�q��Fݶ���z�=��z�\�nh�87](�I�v�rnS
��V��U��_�+kޟlXw�g;� {����r�`wm:����Ɩց�]/ �rU`g�m���ݠ�݉�L�-0SUEUMTX�]�ѩM����{�����K ��Q��wHLbJ�cOt��X|����=�gw�v�� �掞&�Y�hi��m�~���W��r�>��ѩM���v�`�!�Q$̪��I��`Y��1�5&R�[��-�7�}�V�eMu�V#90�a�rmk <uS�}�7Q��N�L��~��F��N�I�g.�f僦�A����;�����'g�c�*k�x��';de������x�����[�eSۉT4xA�$ۊf�FB��՛�h;mQ��9��Nr�e�����b����X�l�Sr�HOfwI7��
5�oU��3-۳F��T�����߯ww{����F�E���.B�2���^��: ��٤��Z�գ�w�}��MPT5<D�`Gr���Y�}���m����Xܫ�V��t��T~7��}�P�u*�Ex���[�4�iդ�@��E�oӲ��vx�F�ݫ� ��e#A�EDE'31@^}Ԩ{�}������~c�V�V�aok@��E�zwM�>��`;������Q���2���+�ܾEC0�Q�������+۳�^VV��[t
�I�n�k@��?�@��E�l���>�{�>�(�����o[못�~�\��X gi(8��NiA0��*�G@6�3�0���a����7T��՘�U��S.��M��X�����`��t��X�ut����+m�?�YZ��,Ӻn��� �N��7��SWe;vƚt��XӺn�}�}4��J�ǻ�@ZX|!��D|�o%�n{�).C��Z���i�P�y���N�uv����,Ulv���y�t� ���P�z(���7���6�)&��e�o �N��>�{��t� �E?1[���I���h��W{��uz~	����Jb)J��?������Z�t
�I;v�QUS`}۫0�J���kfvh��ŀzQ���I&��� ��xym���{�6�uf��˘��6�r`��6��ی��Jʏ�h�<T]nҒ�ݒ&��\�j3 ~$�ߏ�P�z(�w}v���@}�˾T�i�b����&� �n��f�=�v`����7Ӳ������Nݱ��"�7@g��]�g}���u*67����*$��j@��h����gvf����}Õw��9Z�Ia�J���B]ݝ��ٙ㢺��yOq$4�A���7�e`y{� �Ӧ��#�����ߏ�F�^�F8�x��v�
Pܞ�F��<�V*��8�mӎ�7�(�����U[.�ց�]/ �Ӧ��#�7�e`�y+�@�T��t�M���M��*�3V�Xz}�|��y0��j&����ݧ�������X�^��>����(���;�M��x����X�t��t� ��x>�ҝ4��LTL5K6��uE�<��]� j骹�p�_����� *���h�����������sn"�:!Eܠ� �(� �o�_��������*������������������?���?�������q�W�j���[�?_�����������������A�~����������� B�/g��c����������g�������
�����7��������ӝ�������������W�����a������u� ��JT	�H!D� R�T�Q"TH�`�TH�%D�D�Q!�eD��R!HQ%�E�THIQ%��R!Q"EaD�HeD�IaD��@eD�IQ FHQeD�Q$H!Q!!D�H�HQ&H� �Q&HeD��IQ!$D�d�eD�U�ETIXQ%@Q%%D�BTH ��BIYQ!`�!D�%D��QH$�Q��d$d$` `!$%$$�� ! !		d&B$	BB  $P��Bd$Q��@	�� !��	d&@�� ��$ ��B`(	d $%$XIBUd A��    H	B� %d!����� ��B`&BI`$$��I 	d$���$D$$@$$ ��Dd$	`	Q$$RBU$	��I�!D��RB B �T��$$D	@ ��U���de��`�$I	�e��
@�D	$%a��	B�T�"QC � 	IP�%B� 	��
�Q(B�)�`%	a	R �BQA�A�!U�$�ad	@��B V�(��(F�J����A��$D�aQ!F@��B���HVQ�$	BA�F$�`T�aU�a� A�dQ�%HQ��`%HFA�
E
A���`aR�Q�D�eAaPFF%A��a�`�!A�$P�!� BQ�a�aIFT!QIQ�%Q@!%Paa�dIF !!@��e@�	PeI@��	aX�!@�a R!U%�	Y@�P!%�����6~������ UUc����?�G��X��<��3�UW�?�gw������������o_�����UU�?>������u��0���0�����U_�?�g�b������3���g6 ����s��������6|�����\<��UU��/�����j����ّ�����㣑�?��U_��Ͽ�UU��?����?���Y��x��ӫ����O�w����\ßӀ
��΋?���sF����v��=����}������������o��t ���������h������d�MfVED�3f�A@��̟\���1 Q%H�
�UA*�
T�PA �Q"B!J� 
� $*�  <(* ��!E@J� H(%EE
B �(�D�B�J�� �(  	@),     ;�    P� .0�}��z��g{��{��zX }:{��,���sۓA�����A��7  ��E��}�P��F{�\cs3�kgM���kװh⨏w��M�n��x�u^��5z�����   
� Ib���}�7�� ��R��R�g� t� \���Y@������M��JR�Ҕ�,�� P g`t̀)F ���(,�)c4�.YJ
=Pv�t 1@��:P;:P�R���      %\lN�)JR�)@�խ��I�{�s�[�(9�e�0��\����MҼ��(z}�:��{�^Mp  e�nG��2��x }>��5r���}��ϼ��=�F�� �Ϭ��,��es۪�����  
P  
� P}���N��=3�p�O�pN�U�;�Z��ϼÕ�
aР�Ic}�Ϋůx ���w��c}�
<�g�#��Ѯ��K���=N��)W�Jre��c��e���K� ��   @E,������e8����j��ެ��
�y�L��+�_Zriw���=+� z}=�S{��O��  k�v����J�������9����^�}��;���`���2q�����    OPT�ҕ* �OB�%J�41Ǫ�Dʙ �Ob�Pi*��db41?�%�)*��db40���ʔ���"t�����l��s��Rw�gG��w��e@EW�w���O�TU����"�QT����$h��B�6[;��������fS�(5����`�!�W�|�j2j�PF�ҚO��\�6�E�=l�W��s�ml��z��Bqf���D޺'7�h���KHSD��b.�5�'�������@��P2k�>��9�l�SbDd�K���$)Ϋ������e��$RB��5��Aˤ� ���qi\�h|�Zƽ��Z�'S��5���U�s�Q%pU�B ����[�kTƔ֐�9t]-��|��k�}�b��/u�O:$U��޵�y��pFD&��}��w��C�K����$��04c+�T�B�`A�D
,�����@�A��(j�����5�,a6�@�
�	�(E��# �f$k b�E D��&dD�	f�uXf�����ھ�q�gU��z�D�9@#$�)�I��-+�.�'�s�#D�P��B$��%��E"H�eH{���sk�[L�;΢���`�kxc���SW�Bi�	�߱<��x���! ��*��_��٤�����#_ЬHA#�`Ŭԛ��8�oZ9� jF��t�[��3T�1e1��$~�B�F����d�C	߈L�2�!C��.�aR0�l���`�D�
bQ�I	b`�c)\$�ԍi!�
o\��tޱ	����Y�Xd�;p�k;��B��$���oz\�ή���C�bN$&$dX�-l2�kBk)�ѻ��ZE�XV6%D��v���� ���2sn\5�Ulj(��KHy�n�	�[hv���f'�,\ڏL�f4$7� �q��5�H$������ɉB���s ��?@�;d$7�k�Ƹ�.`���ME������wf�¬HL�R%1`a�$rR1�����ф��$.��F-U���ԭV�V�P�{�^�����mn�hE�[\ZH�w���=N�ݨ�c��p��Z4��i (�O&#3C�i	\ѫ�Zd"[��k��c'C����}���D9k�Sr��nNʌ�p�o0޻����IdJB��a�n�Ei#JU���+k������oW��I�ɮ!��	 1D�� `Y�X�0�%�e�=��P{���[aL"HF%��j�ą"O��4,0\�`�Y&��zLH57�ͫ�����L�	��l����Q�hMEE��HM(��0Ȫi"���"$X�tc�!.T�H3�)�g�������5�2�H\֩��ū�Wg�)�a�����A�����$�2&Cl)��c:��~#�-H�"}���G��Ǵ�����>���w(��O��E�Ü��=�W�H;v��F0H�9[HZ����iJj@$`�`��4�Ќb2�%�w�Ǝ:x�X%1t�^����$P�����{�WZ����M%*B�#K�fE��rMo!X�2%�ʙq������x&ڟF�]l���5˲�,q
hf9�eM!<iJ�E��SN��;�2$�]�����e�F�q��$f
��CR�����9��<�@�hci�a���!�l��%�\��dN5��I@�X7�xj��@�i&�æ�3@B�HT�jv$k��d$� ��������	@���$
+���4��h����$��%d�B	�CE۾M]��ީa�ۄ$�ֆB�?��MH1����DL`H��_���?���+.�o� ���äB�F�+���#$
�D�H�V-bK1+w��{涮�U��t�"�H�cE��	 H�9����\IR�GH�m���#��Zp�̐�r�k0��h�)�!sW��ݑ]ɣSF��Hoj��0[���t~1�_���$�t�������iIMnHQ�V����BhUy+�WE�4����#�t��������A�$�D�1��͘��C1�}ٗ9��1iqoWHMSJt���-(�p����Ŵ��{�)� &��B @8���IƤ7��t��4L Q0�0�:�k�su�P�Z�YĞ �x-�i�	ˮ$�3um`����.����yŬ\1Ŷ=խ$5�ĸ�6��D$�<��-�UpǊ!!i�\՜���E�k2N�a�4��zK�Mbj�Q�w�%0b@�\k��/D�ߴ<��ܽ�4���ے�$���A�,�=i��kJ�a�\�"s`�1Y��4If��<um*�]Hjbp�,��4[�!FU"�M��ik-�ц	�1�R|'Bdޮ~�����;�p�;6&�U�Ѡ�6� ILP�dX3�~.���ɻ�5�G�y��}�[�!e]a����a	n����%�h���A�*��:�qmo�޼4{o�S���M��{�����4&�)&�:���9�p��K�h�v郔��%A��54��n`���ר�R-�j"lpJ#��'I74��#��kz��ښ�Y���ں�H�J5a�V�M���ܢ\0���D�)�G�$"���`�=���u�9�	%�:���э$���"��\�	e
d�	M�jM5���!�HU��2L�$��G2�vB0��!��3F���s���k����L�'��9�$��Ч2O��'�G��r"\ωM
�B�@�F)�D� D�) �T�B2$�%�''V�.$kk.����U�8E"?�ȑ"A�aJ2)$�bV6�d�r�+HN�F��X���M��� �R�kB�TЛ��4��ŵ�����o|�q8��&�1�T�4Yٮ-'�����2I���h`��bK��Jn0�G��1Lap~L��������d9)rC9լ��pB�V���C"�9�ou�0/Q��P]ޞ�W�:����g�o6�"GQ�h�`D��;.�{���647##Ё��D,(1#�$�Xa.i���
`aRl�5��F;��5��<��%�ILEƂk|&�!sT淇,S����f�F�����X�\��Z�9n�{ιX��$��7pL������?B�˅�]�\K���o�OX��@�m)Ŀ��6��(F4ҰHB��3��g��C�~aHэ�\����5w���H���cH�X(�\�=w�Ӭ�yu�Ť@�!tS����q>�s��ĉ����^k�3��3|�ʻaĆ����LF"�4	��z��r$&�wZ���tWt��l��P�����K��R�	��re5t��`�w�	�	�|��G0�XR����B.�":�`��C�Ё��5�7{'ow��߶���]is}�~5�2���C#�B,$9rѣ�
�i&�֍���4M8Ĺ���P�0���?b�~9X1" ��&��g���e>�+A�i68��6 @�pm�|t~����aQ��SUx����$O�T4�j EH�\5�K���a�3�3�l�d7C`B���2F�(XKY$K�"`0�A��?,��������/YpH5�
�ܡ.O�M��Ȑ�l�V[yv�T��?0�c0M-f��I��hbokZV���:�ѷ�("F�"��߁!���r�i	�1	����.w�����4����~ IĻUM.$�7U�A�J��G�b��E�U!#.Y�=��$?BU;ϙ�I.o�?l!O�ff�I�.�Pɽ��K{{ˋK���.���h��=��-�S��X�)��Zo�3��!���Z�Wm�Ux�ߧ���}�|O���fs�6���wL��B�{�ev��H�07R�*��4b;7AoʏJku�jdJ$XcX1��fSC�F�����0	a��5���}?��(Kp�G.ȓT�lcr���a��,�a��ޡ+��q��:?Hq�L��P�G�`��`SPB�&�����s�J�F�$�~��aC4
nF#chޭ8f�Ɯb�&��(ƛѲ%�BH�4m2M������Gm0t$a���[�s�~f�?Dє$H�I��Ĺ�fčt� �ʴ��2��1EV�7��$0�TÝ�<[�*\mS�`�.�~�)S�-����e�!$8���� �MԠ`�(���"Q��%��\t� D�V�8��$!�hKR$�B�0�K�w����3\�1�<=2�S.��	!		h��3C]�C�T$�L�؇����%U��h�I�5�!]$(D�@�F	��@���A(��	�N��Oz���zz�^~�  ր                  �m����� ��                                      m�          �C�          �M�  6�   � ��� �      �   ˶q�KZ�Z�3s��k�EgK�������s�v���h켨r���e��u��@]x@V��8�C`�uW:-�_��D�����H0�M��U*�uxX^����û@U�ݯ>^F�[�ҫV�MK��Wh�s������ Aڠ��!��l�F�C3J��km�4��%�ت�J�V�wY���u�`�m��n� ��zߵ�l��5J�*�bdAV�D�2�������s��s��vjsէ�3\�--gf�\�q��UmH�Nݫ�� VRڲ���J�>����t�����8�$�ݶ X[m��S`� p9�plI��[@&�m��l.v���L����[���nWx�@E��ٖI٪^2UT�l -���mf��Hm� rKM�&݀�m��k�  q�Yƭ�ۺ��m��h6�`���R�  �����iV�g3p�o���-�l�dʴD�ɜJ1#�m!��$�dͶm���9�h $4���ݶ $�`�p 6݁m� �c��$�褊PX��V� $  l ��F���@h[F���K[��Uj��XP�/ۭ��Ē[@ ��:�e3О)O$��i�j�u���u�� ��Ad�'��H12ir�PR���]�jU��  ��H>��]���H6�Ni�� �  m[mn��� m�X�luPӪ@�l�R�آ��h���KWVAg#6�X6��c�h��6���@:�~}��nq@q�� �J`Եsɝ�VVΉ�꧖Ie��,�_K� [% ��m�`l8�`�#I�v�	{4�v�I�.n��Zt5u� ����\�[d�  ��t��Lv2�V�<?|�y�fQ��uc�@<��C���6;]���L�ӻu���Š1��sеZY��i+��ҝ�����X�h�ٗv()U6̥�n�U�w`�Yc;�P@�l�C�n�d�mj�u�t���7m&�b"nڕ�^�� m���\R�>��[)�@]���vݳe�X�$�l�A�
u+Bf&X*��]J]GG
�mJ�瞞*�v�l������5UH'�}j����`Zꀬ���Q��<���#]5o.�M�^��:j��<���UV��8ƅ�lt�ҫv�W&�v���M��.�J7nݳ�v�'������}F�2�7��*Wu���[���;�U�<�[��ڸ6���R�m�AX�^�U���XBWdy���B[�gG#�V�������;����!�ds�B�v�RI$3{\J ���+ڭv�ذ�mZN����B�J�9vd6B����9�1E�qڔ��@�.@l�M�ml��<��i(���#����1��*�Tjbzv9�u�6�5U)�m��-��ɵ���|&.��z�=��R����b�r�Sʈ1��rŉ	6����&��aV��X8�Ht�@uBB X��)"��:�6$�m2�l��K��U*�����j��;�)3�=\���Bmc�����M����D����*�&���� )+���a� J�6�7)[����UT��3��=* �g�G�#��J��m�tl��ݔNuֺ�eL⓪�;��%�r�<�p�i��@�n�N���	&�%�.��C�^�&-�g0u5�B\<��z�T	6:�[��Yv^�a^B�T�]E�$�$ pM�7m����f��+=�eu��kh	��`� [kcJ�6ݜ2	�� i6�$�II��9R��*�U��j���Ӂ��Y}X��5�M�d���
����U]YV��z����P T�Wm�J�G����ն  ��knگ6UmU��n`��P6�UV���)��Dڪ��2��}/��(lR�Um�mUT �qKK�*�Sm��jj-se��� Æ����	Vwg�]�(#g���kH9��շ;9x��/xV]�yUx��L�g�7`r�.�������[���"�7[n����mv���^:6�K6����!ʹv噷2N콨�9=[;�2nkb����g�+3��sM��WfRT��Uj���)�r�8|@Mt���P|���$I   k�8�I�[@K4���u���	�׭�"��kd� $h�im�kF����j��'=�vy�8�8��f���#�hH�I��c4�Q$[R� l m�� ��m��- ��i%�4���X�T�|Kimp2Hl�6��m�l��i5�p[D�[�� rpă�Zƽlڛm&�P�n�$[@ Ͷx�ڦ�]K����0�PU�eX78�U�Z� ʦ*	6� I$�D����Fmg�m�$�)R$q��[%!��$���m�  s�m�`-��kM��Em���  6ہ�l� ���6vշ0�\�U\lUuS���i=i$�M������6���kՆ�ٶ l��� $Hpx5��5��V��%K��$�U��FL�_��u�/}YF��� mns���:����-�@j��+u*�( ���I��� m�$l k[M���['WM���JH�ԃm�%��,�۶��`��6� -�ɢ��X>�����m:m�d䪉w,�u��*�tja��W!8�[J�s*h-���4P������5v�	�6�  �k	6���u�m��m����(�dz��x � )j����ʵ� �I��i�� K�i�ntW�n�v���m&�]qͻl\:l�B����lH����2`�[2t�	���6�U�͍.Ϋm�n�{t�w/S]�����x�%S�b@bSh4Z'c0����G�j��Z��m��@+.� T����]��%���ͦ$�7�Yea��������k�����a��%ꮠ�f�y��jS��1l�.ڠ�HG/%�^֚X��m��� m$M+�U��Ɨ/T�� j�x�8�k��,[Ѻ�6�<�ԑ.�����L�Mv ����el$��۶�9��V7gAUTM��y��g��&F #�9�r����K@�i-�ѥI�Ax���% �l]nm����n�7 �v�]3m��V�i�8�n�"��m�;m�[I�%7j��5ָ�U�a���dd����oVS�̮�%�^�cl�E*�� ���9�P�jU�vUj���mw[E���-i2͗l�pqěi4����*�b�
��S�'lr�*ඃ�R���Nu��n�Hc�-��oIjٸ�T��T�r�<�:�[S�m�� �o�_,��l@RZQ�ݹ�X,�h,��peÙd��]��эJ�c�Ӣ�86XۉVw))�ܻu[U܇&�U�fVW^�-��`XiF\6C`6�$���nۤ���}��1�gl6ۛkn -�psm�-6�#�[x$H 6Z$6طT� ��J 	 ���i�$  ��m�� gK]$�i-��6�`rG 9���m��`Cm��T�=��۴i��VTᖫ�q���]$�����u�$�ΐ�@6�'l �+[װ,k��vٴ�UR�*�� �S��t��՛am����H��l$��2��A#��H   -�㜓Z���h�DK���%,��E�h���Kn�u:��p5T�8-�T�����m��zkp`�ۖ�m�H	8D�� p��i!�l��I6  �U�����H���m $	 �kh���` v�C[\  [x A!!m�[	&0m��v�`m�۰;mmÀ�P  -��`Y����� ���D�a�  m���BCm�h ��h]0l[���o��u�@]9�mJ�{9�3L�^sm�5Mq8�h $n� �m�%�"� 8A� ��f��fض�@��m��hl���mh$['Pm��Rf�ZX6��F��e{=���ҵU+�\�j�UʷP�m�iؑ��8 �#�D�I�l�8�  \���Hֻm��V�m�-�Jm� z�$ �l m�e���m�[@ .���J8���T퀪�*�9��Z���� ��iX-�m#A���6�I�m��   �oP�`KI6  �!V�M�[6�	���@�`H �Ŵm�m��m�ph%#���l@mZM�d�l��FB�����UL��6I��X�̭&�cm�I�����[и�f��`�򭩬�h:�CH�/(/+@UuR���lF��P6s�̫m�T�Y^�X:�M����H-���� 6�m�m��lm� I m�m� ��  H�ְ$t�hI۶��h�uU�7\�ݞꍠ�k�ADTU*�O�q@���M�H��ҿ��(����*5Ї������8ϒ)� @u���0m�"��E@���� `$	>�"�6���ƕh]&��L8��� �(�]��І�Q#��*A�!��)"�)����L@*D�Q5�b)�CC��~~W��Mh��a���� �?'��]��!��8/ tG��z��� ,��˰>������;^������U� ?�����q4�|����@�u4*BvJ��@#���
` ��S��"�B+ ����Q4�?&T� :��|*���W���M�@]aЀ������hR�x6~D�>A1^�~ �E��R�/V 0��"��tN"'��DG�`��X ub�QM!�~��.�I��!�PG.(�U>P���jQ� �AX��^)��'������!��~^�%�����#F0�H�&�4c�"�#2$#$`�,! �����D�@���� b�C�Aq�	?u$P�?�O�� :³`�"d D� �B)����,�#H�Y$h�����t �����@$P��!H؊X��Y$�K%U�U!�|�Ţ?T��$�$D����H;�G�h8!��! mN�Q�Dv ]��8D�1D'�#��T!H�O��*�Q�t��E	�(1AX,Y��$�y�1|i��m��m�� m��      $� �	 :[Gm�-�  n�Y;F����,�u��B�8zݹ��3:۶}u�cg��
�^�=���r�]p��fp��(=;�#n�65i�NI�k���U.G�gwgm-��nweSd�0��]���L�)bgTu�<���XCT�y6p,fç��5�q؍-mҭ�z%+t��̫9���VKɀg��9�٥�e�6=C��Z�Q� m͏����͓�l�pL6�$����'�k�; �ںGq�n.+Zy�1��1.�%�����3��e��U.qFZqC�����]/1�`�S���:�ۮ�܁mΐ,0�'�.�8��cg��;�� sJ���=9�ͫ�����cmca�睋��Զ���Gn�\f��"e���Iƹx�2��P�h�m1GQ�v��m��U��<nJ+�v�zP^ݷ<�礎��O-k�;���7R\�gs�i���9e!�.csQςB{q�v���E$�sY��l��s!6�GU��.��K�;��'+wj�8�2�ki^�WLP9�5ԼuA��r�<oU����k���9��P�1g,�D���u��Q�{e�l�@��d�^]���6��X�U�VNs�hom��n�d���\�S�q�rݭ�W(0;�0�n��o�`���z�m�͝��6v��l�����i��"ݮ�����ĥxL���J���q�۲{;:�ɴ��Sh�@Ӳ��p�a�����̹9�a��g�8��P:%%۪�����ζ�Z�v��혇���X�Ѷ��5S<�;\���-niC�:R��*=�(Y*5� ����L<r\Z�;l����+\%�8�ݒ �C��'l��� ��v�>�X �s�`���qX�I�P@�++!5UR�nFM��m�\�<M<���VCt��g\�(Kóe�f:SguK���z�'<�;(8I��6�`�Ĺ�������*���;܈� 0P8����<C��T�U���u1E���(�C��~ڐ���Xu���]�:�\���pn�w:����S��U���q�T9��b���7Lrfx|�׎��caʣ�qũnl��x�� �7��6�4
X��s�l�ۂ��t���ĉڒ��9�m�2is��xq��	׏G	֞���m'y[m�lۂ�*����v�tu�X����ۘ.�ɡ�jUa)2�Xv+g[j��n�m�.υ@�Q�2��9L�3.LG�ls�;9��ex���q���C���]�;s��y���y�ՠx�����?��A�gƁ���*l�Fݵ���=篖cg���`���5ֹ�?z�	��T���n-�ί@�ޔ�9{k�<�ڴ��C�bWH�5�=�zS@��@��j�=W:����,.&��A9 �m���V�����ҟm������f�u���RI��D݉�9�����ӓvyoPݞQ4�5������$�<�ڴUί@�wW��@�,�&���������7H)�:�z��@Է��nI>�����V�����G��I�&I4O�� o��:ϧ{� 7���<�[0�26�0�8���oؑ�?�Z�e�h�z��x��1b�JdRM�]�@=��h��� �m�����o�lݘ;N�q���f�<�K�6�VK���뎮���`��XM>�sm�/m��7�{s��=��Z��4=v��������� ŒM�_U��� ��np�k�脔�ѥ2����R�l��� {�x�Ss��$D$"��Pr"0�J�\Y��4�ˠ7��=�y�k֫8%�iI4=v� ��Y�z���
�W�{�e�	c��m�7"�s��=^�zW��<�ڴ��@�H���ݩ�ͷs�]�b����#��W'��GU�n��9��hv^�nuvu�}�����zW��<�ڴ��4od�7S*,�r����k��X�g;>����4W�^�W<W�I�%*� ��np�����o� ��Հy��2�`��F��s��=]���;{�sr{�&��� x��HZ�s[z|���V���pt�VM��^�U��9ڴ��4{���G7F5�:���7�W9��U[��v/�=/�ٺ�V�틚��0� k����@��z��Znu�~�W~Z�� ��p��H�z��Znu���������d�X�bdMȴ
�uz���>K������� �)�4J�E�Z��Q�i�z����<]k�*�����L2Q��G�zW��>������>_e��=;��I+JR &�wr�]UN�ãnՌ�lhy(�����7g�n9�my׍�2��$'ru�R�;r�^�n�6��W6�-��6�;m�6g�튷lS1�V�����M���`�c��R�>n����ⴁh�\�'�����A�d0}ŀ�7}�l���FR�<��I�.���\̷]]�4�ݶ�s�Ѹcl��ʹ݂��e6��k���R��7�ޞ��wt��~��u�u�8��э]���`9ז���nڭ�z�#vQ�-������'L�6����@��W�w>�@��z/j0�2�@�0�@��W�ؑk�-����+k�;���l��'���H���h^�@�u�@��W�\�[j�fYR��S6U��DD�s��=/�zW:��}V��Yq��İ�7���^�Uί@��U�Uz��ı/�щ���$�1g�ŷ���m�ħO\!��%�ۙ6�Ŧ���%�'�Fȓ����=��^�U�]��OwV�]�4J�E�Z��gu�rp����D ��$"���, �B)D'�]�� �TM���J��*k�V �ϫ rֺΉ��S��Ɣ�8F��>__��ⶽ��^�˺��¿�ĉ1��.��9BQ����:y>�gu� ��zW�\�M�$@R-��^�˺��k�<�ՠU�;�!��{��N�g�퇭�5q��λ�),�����nط0��<]�E��x0��ܝO�o���^�WZ�+�hvZ���f4��X�x�$����~�����h+�|�]��{Q�8�ؖ9"�Nw;۹'o�{��t)�lC�y�K:��sOW�@w��z��w�T�"1�(�Z]���uz�j�<Vנr�jǍ�_�d�c�#�9wW�^v��mz]����6���#va1�vy�ڍ����Q�m%���]�upm=B�����KW7�Y��M���h+k�*�����*�Y��S$ƒ��=�mzW-z.��
�W�~H�00�|	�"	H���~zs�
�W�x��@�_?��$'���H�>��V��О�{ٹ'/{�ܟ�`�o
��Tڢ_�`����7$��}�-���dʙ���p��8(�_t��S��;�U�g�б�c�$�Ĝ��@o7�p�y�!�wn��9��ng����5:�q̃bXHI�岚^�W�w>�@���@��R�P'�FȤ��*�9�rJdn�N���v�Ҟ�)L�"�2C������Қ�e4
�ί@��Ja�i)��Q�G�}�M�e4
�ί@��^�W�W�SJ6�4:�hgϳr��^�M����d�$�I$`��t綕�7nî���aHҘ��v���Q۱B]	牎�p[���w\�����[{��a5��=5���[��2�6�8�q��9�]
�Y鋰�ru����[����{L'k�-#J�W��xV��(׭ē��Z�h�{OY��#��[�ؐ�xz+��. x95M�籣$�]"�;��N�Cdz���
��331*�I-f-�X�eGQ��>�?r�o>z�g]��Y }<��sẲ�[`��۱N	�m�\���ֆ�ͷ�v=��^�{�49ڴ9���X�4(cY#�=]���S@󬦁W�k�/���B���%	$z��Z�e4�~ľ]��r��y�FE�8�ؖE�yl��W������/���=�#�D�FO�H��ـ9��XD'M�~����v��~�����u�z�ͧ.���}�ۃmY6ѹ��*�蘶뤻���k1B��79�}4X���`;����p��9%	$� �v}������&���p�ǠU��͝�D�%�+W�l]����ç���wY�r�@������SJ6�Z��h�m�.��]�������,m�� ӆ�y�٠z���]k�<��h���c�cBxؠ�)&�����9[]�	{�xzm����]���c�}������U9[9����v,�x�ٳy�!�Z2Nۧ�a��kT�m��6,���� _�����I{�T�$%�m�x�B����K�y�.7���,$�G�%�9E�$�e�o�$��dԐ��_�}���__�^����:�zm����뽶���K�����^�@����3�����~��h����*hB������N;4�O�yٽ�~0�[�{�챫����ׁ��۔*��wVQ��no��DJ� @�H�!�@�/��h>�"]���S:(@�bɠ*5�!��B Ї�8�{��0��w��}��˯�a��A>_l�P��������~����0N~�n��>H�,`� $I�LJBw��c��q��}���tC?) F,� �F1! �$�t�>����t|��^/��W`�^ J��h*z�J����!���1�7&�}���o�K���o��~�QX���ry�IޮjI/zu^x�^�Z���RNy}���m����Wv��e+�]6��o|��������&�m�y}����?�����??���(��:�B5D\��2��LM�����t`��v�Kn�4��w{�|}�BK�&� ?���g�m��{�{m�����%��1r�߾�~{�m�pB?)�5drH:�)4�m�޻��춱����߾��=���|M~�K�Z������ݓ<��<��������I%�KW�/���χ�$�\���%x� <X��6�(G#����}w$�+�Lݶ����9m������5@(@?A�h*�� �ӊ�L���߾���H�l��k��o����m��ً/��s��>��t6�'��}���;�c��x�Bw��x�y�ǩ�3��c���gq�q˗������N��NH։$��-�x������KޝW�$�������N�Ɖ�� ��'�$�����K�u^x�^�(�$����I+���7�HcQ�H㚒K�o��RK����K˖�<I$����K�Ag+���$N/<I/]��I$��l�ĒK�ɩ$��U�%[0�㸲&�lQ	Ƶ$����K����{�v�o޾��m������ox���-u��OK�o�$ ��)�a���kDjz^�wl�H���������\��$p�]���c]<��Ͳ��u��t�oP=u��y���d��Lػk��ݷpiGt��FU��t��Od�ԗ���m�\���7H���wo��~�K$�]�D�]�"C���kl�`�;6^�I��f�53i�n�jG��-�V9�.� s�(�t� �)��v��`�Gsgi����\�Y�Y��Ն�'5�*	�AH;5��-Әز��N��[��V�g�Y���_84�r�-�m����6��o|�����ZԒK˖�<I+�2!�*%�,JI&����U�%�v��$����<I$����K���YY&&&%��8��$�N��$����$�u�RI{ө�� ?��{axL@�� ��[<�$��jI/zu^x�^�jz�Kο?�d�|: nk�� ���_ ��g}��|�m�ϾsM��:�뽶�;�A�D��]N�I���ls��&=-�y�Ī�1v��Rr�3Y۳�h��7��-�a�55$�t�y�Iz���I%��g߳�f{�I
ߜԒ\�E�@�"�$��E���3���������u{w{m����M����=��Y�I�G��ő46ڃN7�$�}�}<�$��\Ծ�$�}��Ē���oRI^��/����(�x��ĒusRIwKW�$���ޤ�^ܶy�I^2ʌmbP�G5$�t�y�Izݭ�I%��g�$���K��b�Y�k�(۲[UNU-�}��%�6���E��ݵ�Յ�g��-���5A�v������G���_��� ?޶y�I���$�w��Ē�����	FF�4�r7�I%{>�y�I���$�w��Ē��[Ԓ]��X5#o�dQ)T�{m����M��=�M��9�`�bN&�`C+rT$B	@ˉ�P�|!��?������f�߼w��-���vF�'1�'	sRI{gU�%�v��$�{��<I|ӷ�5$�?��_d��#vG+��o�{�i���������޶�����m��{^7����f}>�|K÷f��\�p2�̘��5��v;r�;WA[h�j�Ň����n�s���F_RI+s���$.�椒�۴�3=���������_��_Äyx!�k�� Ͻ�����%������om��?~�M��8���_��{����ޭ����;��M���ߏ<I/[��K���k�/��H]~wM���4�+���h��M��Jv�}&�m��{뽶���K��^��fb�Q�DXU) ��N}���k=���-�V�P�c��d�m��.��m��9�}.�m����|s�z�K�	Z�)k�(���1�s�]�b��gh�7�Mo���A:K�M1s���_�k�H���I�r{�I��jI/=�O6�|����nF��W���m����i�붻e�m�������I[_�零ffe��_��3$��D]�ˮ���WGQ����m�ϾsM��8�뽿��$�������}�_����� �4�Sr=I}������ĒK��]6��=��o�X��Jߵ��4�o�}��G,p�/�U�� ���o���������o�{�4�os����m�k#���@ �)�d�R��yg6�\)dXŭ�	�<�m����P�h��u�2<�Ԣ9&�C���`�=�m��,.0n�v@[��'L�-����7n������};�����7Ka�:g���]��NN�C�.9q3�C%�mO7�n�t����D��f��hf�e�\�Tg\��=/S)�M�r��"s�Y��`�n��K�x�X�yk���*Y�,��%�(�w�rV[n���.�N0�Fu����n��6p�}��lMj틚���;Ր�� ����I}����K��=I%��u�~�֒��5$��T���1�5���<�$�;S��6���O<I!_�sRIy�~�_�T�������? ��_��$���5$���W�$�'jz�K�g����J�tD�_���{���tߟ��jI.���y�Irv��$�~���I/{,5��b�H�sRIy�y�Irv��$�~���H]k��K�b�,I�U�%m�^C�cV���]l`=z鬔��m����Y�7e����o�>�jx�!dc�� λ��fO���x�[�J?H{k�p�0_)��F�r۠6��맚�b��N��A��,]Q�����(lqFBIG%�_�ΟN y�y����c���&�7�LqI4߾������T}�}x˞���"���e�܍7K%��,|������@m�����y���0/��T�5H�Ww8 ���(��-�=���� ��j�Z1c�Ly&!�b��X��:�H0Xx}�.n6��ܛ-/V�ɱb�E~w���>��̮����-��v{����{�7�j�������r�~G�"�8�� ��B�DU��Ӏ?���������.��5�#��H�����rI���06��@?$*�Q�� "�T�V(��%ѕ�n������JZ���-ML�SW83��x�]u��w�ؽ��σ� I�m�1��h/m;�:!D�}������ �n�!�S�2k����/[�ֻq	b狒pW�\��s.݇��������Oۇ3�<���v݀}�}t�=�s޿b�[a��~��c>�<I}�6�(F��<��9�2�׀zv_^ =�yВ�=��r0Ƙ��c�-ߟ�-���0�(��UGw}x����7Ȧ��f���4�q�}��/_+��o�@��j�?o@P �>*l�S�bs|ZE� �F?͑ENM ��xЗ�^}�����p���x�^\X���s�\sՌ�ݗu]��I^x3��@0������������I�HuӶ�n��g�=��zh�]����Y���������B�ʜn����n��B�2���o� ����Q	b��}0_)�q9#u2[4ޯ�� ��xtD(I)�����Հ~{t���Xf\3u��������*g��^ �}����X$�|�(��m}��Lg�����O�nM�]�@��I}
!F��}^ m}����0���������.Wf�ؐ��RF:�ī
F/M�8�&�v��~w�$;��'��T����ȁ�)�HŁ ��!�dػ��XE�(����j9Dvk�>��.ͼ!T�~9a4��$���- P�Q!E�@�ĳ}��$%�F!� 	��?�b;�����@�+	�j�Hs�4�LeR�
�O��X�@1�O��!	 8?��B@ LD�!��i����P����5 ��2�B��]��jn M�?I~��2��G���x1�(``�`����{��w�=��?�H   �:�       K)�� � [G�M� U\qu;;��vy�7^ʮ�!��v�u�l�,�-5�%#:��讬nX��cvh ��R�A��n؀NȤ���櫶��tqm��[-r��m�a�g,d�.��9���S���;c�#C+F�"��6 �����l�V��k�`�Vd ��RLh�;,���D�0��yN��/a;N�s#d�B�\��u9���k�N4ƃt;�N
���=��ہ^}�u��^.lqO8�F�d��W�%��"�\T���qt���n��Lhcgm�2��I�z�.�.�fU;�\���kz�lq�9�m�������
�u��`c0��Sl;m�8yy��M�O-���A��n��v�[���;<s��2aN��vئ��}H}o8U�GHt�5 ��%Dpjق�u��
�֑�A.�	��g����k-ۮ����e^Վ|�5[���*p/Z��#a'.YT�ゝ��l�l��:�J��.�I�ۧ�� �=�֖㫖!�X��3n�D�5�dZL��&8�v�)8�3&�(��j��YM��n�;KΩ�IS�϶����n��~nɵ��ztq-��d�cu;�Ne��c�M��v�v�s��(� y��[���/�n������m�m�/�'O:Y�g���@jQPw���}���`5�1��<�����lu���땣t�U�zf�Yq�Q��WV��Iny���e�n<j�vD|�s�9ےN�2렫�k>Ɍ��8�t��tU*���VV*��Ůݦ`�!Bv�me�#ՉTf�T�6i:��,��[oJN�����*�M���qt�2�I����N�՛�i^ӆ�c�R�&��`:�R&	^}n�hWY`ڨ�i2pTۆ؂��:��$ +am�8q��j��m X��bY����&�K�h˳�)'9cm�\�sn-��^Ǵ��6ؐ,�F�s3YkWQ�I��(�p8�ȁ@�	O"�/�|�@L� >G�@�W��?+$0�l�,����K�[����!��.7m���v�2M[u��7d�؋i��n9 ���/�����{˵n�B�����ް�;~i��ݞ�>�`T�;yy��8+;9��Pۨ�Ty8�͹��6��c6�A�n��S����/jn���Z+<p�J��JBb���C]ud��Nv��.T���m��@�]�	9��9�a)���Vh��I5��̢�]�+����s�x�?�)(�޷�㋶�<^�gu���3�n{�)�N�תz�0��w�e��~��4ư��/ �?���{�[4���������=�O���Zl��^�=����B��DUw}x_���s�fg�G�����I�rh��{�ه(Q3������xϵS�5cj��k��>�X�{��4�>���M�%
&w�^��,�V\�Qjjf�j��7����DN���ϯ@��)�u��I�H�S�(�;n_k�5��m�Eu\��8��DN^Klc�b��wwwMᛏP�sm)�xݟ}4���y�>K�
"=A��������vT}5:�2�3u�����"X�%�~�}��!�4D�
�~.&1�����,N���m9ı,O���m9ı,K�ǽ��"$P��,O����0�2ᅺ��ֶ��bX�'{����Kı;����KĿ|{��r%�bX��w��r%�bX���������2�Z��M�"X� �'~��6��bX�%����ӑ,KĿ{��ӑ,K�H��;��M�"X�%����k*�U��ų131>�����KıF���[ND�,K��ND�,K�{~�ND�,K����w�[@�{yv�����p�q��ƍp�����l=Cb燚)���	��Ґ�`�\њ�ӑ,KĿ{��ӑ,K�����ӑ,K���ߦ��B~��,K����[ND�,K����X�UFꬶ�n�l��L��]���-�Kı?g���r%�bX��ǽ��"X�%�{��[ND�H!�2%���|�*K$*u��k�L��LO����6��bX�%���kiȖ58��ș��涜�bX�'���Zų131s���&�*���ֵ��K��@��>�����"X�%�}�kiȖ%�b}�}�iȖ%��X���i7�O��c�Y�Gi�+V�,@�.����,A�.s�ٴ�Kı?{��ӑ,KĿ�>���L��L��r��Up�us��+i���6oGN�b�^��.'um�ZO6�I�alw�)K��0�SY��ӑ,K�����ӑ,K���{�ND�,K�����9ı,K����r%�bS;�և�]Q��h�Zų13����6��ؖ%�|{��r%�bX��ﵴ�Kı>����ĳ1{���D�)�����-����X��ǽ��"X�%�{��[ND�Fı>����Kı?{��ӑ,Jbf.O?�!du�r�c�Ku�f&bs�"#�3����ӑ,K��}��iȖ%�b}�{�ND�,��!8�*0F
F�x�Q $U��1 '��QN���ȗ<}��"X�%��=��YJjC4k&kW5��"X�%�����"X�%��EW����ͧ�%�b_�kiȖ%�b^���ӑ,K��޾�ə���X���c��Kw@�n�Ÿ����lay.�:���h������_���۳�љ���Kı>�{ٴ�Kı/�����bX�%�}�lyı,N����Kı>���3ͳY�5fj�֮ӑ,KĿ�{��r"%�bX������Kı;���ӑ,K��=�fӑD,K����}r�1�����SZ�ӑ,KĿw��ӑ,K��{�ND��,O���m9ı,K�ǽ��"X�%����R�XLɅ��Zֶ��bX�X��w��Kı>��ٴ�Kı/�����bXb^���ӑ,K����Z�v4��+��-��������{6��bX���P3����[O�,Kľ������bX�'{��m9�31�ŕ$��������m��[�t��.�-���uҥ�I�́��ݝA�LY��#� S	��W ��,/:�g���}�v:甛H'\��Wf0�\Ǡ�����%�=�X����^��%��KgY��e�]˭9k*롺�a�{B��5�ٸ⭃��r���
�]�f5�qVnK��U22�H��Ɍ&0���^���t\n�<,8]q[5�.7Y�h[_�X�\Z�����NR�G���v[i}��öz��\����㝝��N��zZW>�Y�ZviE �PF�e�k�N%�b^���ӑ,KĽｭ�"X�%���~�
�A�L�bX�g���-���������F���'+v9dֶ��bX�%��������ș�ｿ��Kı;���ͧ"X�%�{���r(-�bX�Ϻa�YJjBUa)e�ų131w��Ʊl��N%��w�ͧ"X*ؖ%��OkiȖ%�b_��kiȖ%�bw=%;|jf�L�5n���M�"X����w�ͧ"X�%�{���r%�bX�����r%�`�X�w���r%�bX�wP>S�lv�Yk%�X�bf&bf'�|���"X�%�� @@����[O�,K�ｿ��Kı>��ٴ�K�L�Ͼ�>p�ƴn�NX�Dd�=��b�6[N���wV�Ӻ{Em�=��.����q?>��Ʉ�i�-��bቘ��������D�,K��~�ND�,K��޻T9ı,K��=��"X�%����(�c�q7Gm�ų131w��fӐ�N(�8 ݨ�%�bsz��ӑ,KĿ���m9ı,K�}�m9� F.DȖ'���ܿ�kY��m�SW4m9ı,N�_��iȖ%�b_���m9�Ŀw��ӑ,K�����"X�%��0�"T��ezų13�(b����t��bX�%￿���Kı>����K���N���iȖ%�g���~?��Iw�}��oq���/�����Kı>����Kı>���Kı?}�~�ND�,C{���ߜvDߋ�K���|��&8ӵ��Zw&��[yƤ��7g9������:�8�
Ude,�X�bf&bf.��mk�V%�b}�{�iȖ%�b_�x�� �%�bX�����r%�bX��I{/ʖ�%EnWmZų131w��?�H"X�����r%�bX�����ӑ,K�����ӑT131w���n��-q���f&abX���=��"X�%�~ｭ�"X�B�
��H(@�F�$D!`*F*0Cf���@��>����Kı;����Kı=��]k2��)n�Z�Z�r%�`���~ｭ�"X�%�����"X�%��u�]�"X���AG"g��?���Kı>�u�o�RD����L��L����aȖ%�b�����iȖ%�b_�x����bX�%������bX�'��>��s��U:e4�km���g�!wVk<V�����<<��n�X���ړY���%�bX��fӑ,KĿ���m9ı,K�}�m9ı,O��m9ı,Otվ��L�&[5��k6��bX�%���kiȈX�%�~ｭ�"X�%�����"X�%��w�ͧ"(�"dK�x���K�`��_{�[�oq����kiȖ%�b}�}�iȖ
X�'��{6��bX�'��絴�Kı^��mF���VFR�u�f&bg�r'{���ӑ,K��{��6��bX�'��絴�K���!?S�N.�'����m9ı,WgC�ʖ��N�+��bى�����｛ND�,K����m9ı,K���m9ı,O��m9ı.�������0J3e�k���m�+�����G%�\댃��WA[X�����{}m��� �N��Kf�p��L��_��[�[18�%�~����"X�%���~�C�,K��w�ͧ"X�%����>���ۄ��2�Z�ӑ,KĿ{��Ӑı=�o�iȖ%�bw;�fӑ,K���ﵭ�"+"dK�2��c���ƣ���bى����������Kı;���iȖ?°��>��k[ND�,K����[ND�L��_O���D�r"�-5�f&%�X���ٴ�Kı?g��kiȖ%�b_��kiȖ%�b{�ߦӑ�����o�8Q���e�ųı?g��kiȖ%�`��{��r%�bX����Kı;���i�131E���������[m���ΤK97�X���3��#�x�5�t��e*� 	��s{�u����#sL��2�h[>;j�n4�@u�����5�'��.���+�tE����ŷY��U�u3����׫plc�}u�A��p�="��@��'�m֓���0��&�=�:�U��Gs�3��l�s�D��!IĄ�F9c�Xٸ��B���b���]����۪��8�8�:�^���b��:c�ۙ���g47��	��e%�0L�_{�[�oq�����kiȖ%�b{�ߦӑ,K��w�ͩȖ%�b~�w��ӑ,K��}�F�i�
Ude�X�bf&bf���ı,N�}�����D�,O�����ӑ,KĽ����ӑ?�*����>�?ʖ��N�	%5�f&%�b{=���ND�,K�{�ֶ��b�%�~����"X�%���~�NDf&bf/z������N��Kf�l�bX-��=�k[ND�,K������bX�'���m9İ?�`D��~�5�f&bf&b��j/öǃ���֍m9ı,K����r%�bX)��~�ND�,K��{6��bX�%�}�[ND�,K�\��2ٙ����Ŝ�n�7���錞�m\&�ٳ��I����֮عn���C5��~����%�����M�"X�%��｛ND�,K���<�bX�%������bX�'���=��f2�F�Z�ND�,K��{6��Ü@�$! !O�4!pS��j#��X�f��0B�1ؠȜ�b_��~5��Kı/�����"X�%���~�NElK���[�d���m[l�X�bf&bf'���]bم�bX��{��r%���@��?�����Kı=���ͧ"X�%�����ۙuq��u��h�ӑ,Kľｭ�"X�%���~�ND�,K��{6��bX� X��{ƶ��LL��^ﾁ�"yT*�2�m�-��K��}�M�"X�%�����ٴ�Kı/���m9ı,K����-��������)�nI[�������۱�m���k�6k��66�=h�^�1+���X�M#QM*J�*u�I)�[130�=���iȖ%�b_���r%�bX������  ��dK�����k�L��L����?cC�X�Ym�ND�,K��x�ӑ,Kľ����"X�%���~�ND�,K��{6����Dr&D�>������dc����u�f&bf&b~����LK��}�M�"X�/�|x�N��aH@$�J>� ��A�J#�O������q����@�]���A]�[�l#$�،�)�҆T�l��B��M����M��Y����H@�XBh����/#BBh�	�HH~.�ژ|<�B���U�\aC�d�c֘�	�~a���l	� �8��#Qu-�5ˈ]�As8P���4H$��>0T~4�AMD@�@Ћ��?�M���B&�(��C�� �����&��*�G�@x��"�:' p�A���;YϾͧ"X�%�~�|kiȖ%�b~�uܲY��L���f���K��;�o�iȖ%�bw=�fӑ,KĿ{���r%�bX������Kı;��9�&�0��0�5���r%�bX��{ٴ�KıU�{���r%�bX������Kı;�o�iȖ%�b9�'���魗t&�����.`@x9��=I�;e闫̛��?�wv�>o�]�N��7��%�bX������r%�bX������Kı;�o�a��E�2%�bg���iȖ%�bt���L�.���Ys5���"X�%�}�{[ND�,K���6��bX�'���m9ı,K���[N@T�,K�w�3
�B��+v�bى���������-���%��｛ND��H�9"^�{�kiȖ%�b_�kiȖ%�b}�'��˨L�unL���r%�b�'���m9ı,K��魧"X�%�~����"X��`�"� ������Kı=�0�i.�k,֬�k6��bX�%����ӑ,K�Po��kiȖ%�bw�ߦӑ,K��w�ͧ"X�%��{_���e�V��`�G����k�4N�]�y�$(ہ�Z�lt�24�2�$�a�5�VX`�4;.f����X�%������"X�%����]�"X�%��｛A�,KĿw��m9ı,O�G]�K�d��[�]k5��"X�%����]�"X�%��｛ND�,K��_kiȖ%�b_w��ӐTı?g�����f2�Z�kWiȖ%�b{;�fӑ,KĿw���r%��X�%�}�m9ı,N�^��r%�bX��5�j�DR�M�m�k�L����,��_�m9ı,K����m9ı,N�^��r%�bX���ٴ�Kĳ���F�c���۬[1311/��kiȖ%�b�k޻ND�,K��{6��bX�%����ӑ,K���*>P�p����(�a�����MUS��\��}qb�Xٟ+�͹@�Db붸֕չ�y���n}6N{v�V�Q�t�8�-�fڻv̻���3��-���vܷX���si\��PX�F�lsÞܧ<WnS�U������Ӫ�ݮ�6��L[��;�\�$ɰL���3���vzꇙe��u��+������ g��6k�X�`�[:.t�����}���O����m�ª�8nc��ps��n˦�M�[@!uy'^v�v�e�Խ��R��{ܿ}�]r��:�MZ���%�bX��_���r%�bX���ٴ�Kı/������bX�%������bX�'s���Yu	�.��˭]�"X�%��｛NDKı/������bX�%�}�m9ı,N�^��r!bX�'��3�&�F��ՙ�fӑ,KĿw���r%�bX�����r%��$��=�����Kı>�fӑ,K��ާ�5����v�u�f&bf&b}���ųı;�{�iȖ%�b~��ٴ�Kű/������bX�'��B%-�\ֳiȖ%�bw���ӑ,K��w�ͧ"X�%�~ﯵ��Kı=���iȖ%�b_ǻ���i�;+�b��oa����t�(�v��kMW�ng�-Ŭ���<H�r����w�%�bX���ٴ�Kı/������bX�'���m9ı,N�^��p��L��^����j�M�m�k"X�%�~ﯵ��(?�(A�C�� ��S��%�bk=��6��bX�'���v��bX�'���m9ı,N�=�L�5ksV�5�s[ND�,K��{6��bX�'}�z�9ı,Og}��r%�bX�w���-������Ӿ�UT��Uq�vͧ"X�@ X�����A={�fĐI�ݽ�n	"z'���m9ı,N��3Ʋ�4][��Z�ND�,K��{6��bX�'���6��bX�'���m9ı,N�^��r%�LL��3��9"��hwF�+e���p�1��3vpܫ�#3��[`��L��\�8���k%���bf&bf/��ޱl��X�'���m9ı,N�^��r%�bX���ٴ�Kı>����f�2�)n�e�m9ı,Og}��r%�bX�����Kı=���iȖ%�b}�_siȶ%�b~��̶�HL�u�5��r%�bX�����Kı=���iȖ:vDH���D$ �U�Q: M�Ȗ%�}��"X�%����ͧ"313'��"�A���E����f%�b{;�fӑ,KĿw���r%�bX���ٴ�K����]�f&bf&b�Ⱦ_Z�D*bm[l�IȖ%�b_���m9ı, =���iȖ%�bw���ӑ,K��w鈴l��L��Z�#��rV:Q�����x����6�u'�>S:���ջs�Pع��Pu�d_RW�����{��'���m9ı,N�^��r%�bX���ٰ�b��ı/Okjى��������eʫ�+�kD�,K��޻NAı=���iȖ%�b_�����L�bX���}Y�
HRB��D�_+��*�\�V]j�9ı,Og}��r%�bX������b	bX���ٴ�Kı>���Kı=�HO�ɬі�j�ֳiȖ%���L��=����"X�%�����ͧ"X�%��u�]�"X�@���K�߳iȖ%13~����a��i�m�ų18�'���m9ı,Q����ӑ,K��w�ͧ"X�%�~;�kiȖbf&b�Wڈ��]d����h:�C��q��2Sŵ�dQ��b�wV�e��6�K����w��6ސ(���f�l��L��]����Kı=���iȖ%�b_����"��2%�bg���iȖ%�bvy�Ċ~����k�-��������}v���"dK�������bX�'�w�ٴ�Kı>���O�3#�L��⿗��:��V�k�.D�,K�������bX�'���6��bX�'�׽v��bX�'��}v��bX�'O�&[���3V�.�f���Kı=�wٴ�Kı>���Kı=�wٴ�K��A�:�����L��L���ߕUH�.U]a��ͧ"X�%��u�]�"X�%���}�ND�,K�w��ӑ,K��}�fӑ,K����(�p 8�B�|�X�@j��A+$�F.,q��X(T^���:���e{���+��+�D�dҧ8��CkSíB��g�KT���N��ɟ3�N�a�s����]m�i�\��:'^�≤�ne�q8�u�;-�)�M�����M;rBzMy�:k ��FczF����sO����;ƛd��ʻ�l6�c�z��&^iݷb��\]q�Ԇ�6;���M�/��!"�(�67g��sҮ+��B�T��b_%������R4���l�Ӥ��y�/tg�ű�˭�C�v�u�n�J��8�Kd��R���Kı;���ͧ"X�%�~;�kiȖ%�b{>��iȖ%�b}�{�X�bf&bf/�A)�0v�k�iȖ%�b_����r���,K����m9ı,N�_��iȖ%�b{;�fӑ,K��ާ�5�ee�).�ֵ��Kı/�����Kı>���Kı=��iȖ%�b_����r%�bX���̶_-u33Z�r%�bX�w^��r%�bX����Kı/�}�m9İ?�fD���kiȖ%�b}����3�-�.I�f����Kı>����Kı/�}�m9ı,K߻�m9ı,O��z�9ı,O�׬�ՙ��F��zݖ��c����.�u����nx}�p��zY��.�!s�:�O���Kı/�}�m9ı,K߽�m9ı,O��z�?�@��ı;���ͧ"X�%�����.]f��3V�.�f���Kı/~����>Q�@ �X��؁�D�Kz׽v��bX�%������bX�%���]bى�����="*�U�w5��"X�%��}�M�"X�%���}�ND��E!�2%￿�[ND�,K�w��[ND�,K��ĥ�LՙtL�]fk56��bX6'���m9ı,K�}��ӑ,Kľ���ӑ,K�﻿M�"X�%��I<g�n����9f�l��L��]���u�f&abX,s�����~�bX�'�����Kı=��iȖ%�b}����ɕ���N]�;5��rU!*d�*M;NƲכ��N��mf�g!�<�b���Ȗ%�b_}�kiȖ%�bw�ߦӑ,K��w�ͧ"X�%��w�ֶ��������= ��#�j:I-�r%�bX��w��ı=�w�iȖ%�b}�����"X�%�}���bر�����<׉��4[%�iȖ%�b}�w�iȖ%�b}�����"X��!��H+��DM�h�7�����Kı?{�iȖ%�bwڷľ�̳FC)��ֳiȖ%�؟g}��ӑ,KĽ���ӑ,K�ｿM�"X��L��{�6��bX�'���̺˫ɫ���]fӑ,KĽ���ӑ,K�ｿM�"X�%��{�ͧ"X�%����ٴ�Kı?w��I3$��JAX+ms۞v�Ɍս@����;y�jN[:��ۦ�b����Y�Gh�5���w�x�,K���6��bX�'���6��bX�'{�_fӑ,KĽ���ӓ131s��h��c#���,��n%�bX�g���r�ș��{�fӑ,Kľ������bX�'}�|k�L��L�ɂ��}��*+-5�ND�,K��Ofӑ,KĽ���ӑ,�"�DȞ�����Kı/����"X�%���_sZ�[rJK�j�W6��bX�X��{��r%�bX��w��Kı/�ﵴ�K���&�~1&C�*dH ~ǌ 4������\�r%�bX�}OfKg���i�S35��"X�%��w~�ND�,K���[ND�,K��z�ӑ,KĽ���ӑ,K�w�����`(�a�Y�{n2���B�a��=Y� c����-�[����Q�<�&N��f�6��bX�%������bX�'s��ͧ"X�%�{�����"X�%��w~�ND�,K�վ%��t���kY��Kı;���m9� !�2%�}���m9ı,O{�iȖ%�b}�w�iȟ˕2%����������,�k�L��L�����m9ı,N����r%��%��뾻ND�,K��z�ӑ,K�]��Ԭp*�U�n[�[13?Ȟ��?�ӑ,K�����v��bX�'s��ͧ"X�%�}����"X�bf.��J¹*+�K)�[13�b{��ӑ,K��u�fm9ı,K��m9ı,N����r%�bX�����XO:~�z i��\%�������oag�l�f�;�f�����Z��G{a�&��x���T�@&�����\���V1H�@������BGI*��B!��t�d'�hd��H~�a	��4��2�B2D���[�Ѱ�-J�!�͵�2M� 2)!{�4��C��fՏ�F��A)�5DhC�cHX�\}^�[m��h ]0�\       �Sm� �� pBF� �,�Y.�K�g*M��Q����l�F�6�:C7]�u�3�o2\��^�N���k�:U��pcZ��h���E��j�%A	���-��e����4Qځܬ�iC(���0r�b4su\�����¹���k���#�u2����ɻ\d�yɴI����&'�ʦy^����w�:��s��zv9Sa�Y�ۂapsF��l��&sؽ�9�.�O^{q��u#�68���a�Z�)c�<)��� ��9�t�Ȓ;�{Ln�z�� y��,.�D��
�p�9��n��ysBv�P�6�v��4��@�m�Wi�'���ix��!�qm�kf8w<��r$ΆtcE�:ۣ:���幆���uK���m���%��@[e[�`�#��5���� �ml�%=]x�EH�4�[f��kGOc9�C�g�'c�z7m�fP`�G�+��j뱐�d�7F A�݆t�O��	MN]�0���-�nX�-'>��-�\+�ة���l��\˞^��Yф����j�8K&��z!t#b�aJE�����D��bó���9����Ю)���wn��;b=�W���N�.�ف�:�w���.�9��ڈ��P90筋q�e�L\B�qd�,��5�Ƙ S��܇��mx�{"$2�1 ݵ=s<�Ƽ�#����3هpy �U����v2v�Y5glA��r����l�[��+���8h�ଡ������b�U�V�@\�Uٝ+7V��`}�P6v	N���p�eb����ٹ7up͓m��Ǉ�]��UA��55�a�Ձ:�KŬ���)S.��a�ڪ�h[N�+n��Ci��7)(%LAŻp��m�Ԣ�X0�����+HAnI�8ZMf�#ˮ�(i�KLT��`�gQʘ���"�P�7HBiI9���+RIL��B*�4R�:1�5�qQ 4��P��՛N�A�W��傡������D�`~ب*����=����{���y�[��: 
�܂g�K��8�ɮ�C�=�ɼCʪܮc*Qrss���������g7;�v�o��u���t�n�4`�Ve�<��b�;v�v�Whp��B��ݛӪ}n�j��g���!w�Er��p<�Z�ny��`M�Սl�NȬ��gn��� Y�h�I:���L`\��m=`Ɲ�*�$A�7Vv��5��B�b^��2"�7Jդ����Nq��8�uq���TM�\�mƧb�+h4%�@�>����8쨬���L��L��߾���Kı/�����Kı;���a��?DȖ%���{��9ı,��ߵ3�ǃ�hv�k�ų13��{[ND�,K�k��ND�,K��}v��bX�'��siȟÕ2bf/�e�1��$q�:I-�-����b{����r%�bX����Kı?g}�ND�,K��{[ND�)���<ף���qF�]���L�bX����Kı?g}�ND�,K��{[ND�,K�k��ND�L��^���O�8;�mR[f�l��,K�w޹��Kı/~ﵴ�Kı;����Kı?g���r%������_�!}b��˒�Z1����p�D�F�x�ؠ���kj�^�sCn�Vc��%��bى������ﮱl��X�'~�}v��bX�%���[��&D�,O����6��bX�'s���T8B���n۬[1313�}��r�|"t�Ӹ�%�{��[ND�,K�k���r%�bX��w�X�bf&bf/O���h���+��ND�,K��}��"X�%�����6��b%�{�}��"X�%�ߵ�]�"X�%�_��_9�WD՚�-�kiȖ%��$��������Kı/���m9ı,N����9İĿ��kiȖ%�bw���Z���e%ֵu��ND�,K���[ND�,K;����Kı/�w��r%�bX����ͧ"X�%�}�e�fk!�m���WcvK˱WE�Y�gl�ng�j2��Ŋ��-��;�6;\�Yj�����ı;���iȖ%�b_�ﵴ�I!H����^Q��}x���5G��M�-��@�}u�f%��~�������ٟ$�����*�T6�v۠<���h�ﮏ���0BB�4h�@���E'=�z�ܒ~��tW<��c�������$�~QUϾ������]�:���z�LI�fL$�$��W�hg��߯��*�|��wu�.��Hrc�BL�-�z7W�c�Kn�t�%b���66�n�������A��H��h�٠t�sX���/����a�OEe�	�94]j{��߾��ߖ�{m�������B3�
H�O@+�]k�9B��{��/�k {�U*I�S�\ݬJK�}8��{�}~�nnOʟG�
&㢢`�3F�
1&�*���G��o�~7$���e̞չe�,$rE���s�����W�z�'���O��ƫ�$WUN���e⎸籗<c]3�7n�l��x�:�F)l�.EH��G��-|ށWuzW�h�٠v^U�FG�F�q��k���L����S'���뺫 ��VL&8�H���@�Қ�h���]���.q,#S�)4�l�;���Ϫ�:���gQ_�)��LIɠw;[�;���5� ?6� ��B��D�_wO~�ޞ��;ݿT%� A��cnō�}8ؘyiG���J�g�xe�-��ka��uP���uҌ۶��Mm͓-��]�:u�v�V��'gf��S�F��N�gwAg���Sx�[DMg�}���mqַ H˳�xV�[K�cm���Bg�b�'����ͩ���s����3ִݛ[����Ӣ�cװh���yI��";b�2��*R[B�Fm�i�t���w����{��ߦ�2�	��j��v=u�ζ�OOcE�$p���Vym�u�x�Mt�&�i�9$�篪�:���ym�����9�}j�A��M~�0{lϡD)��� ��W�6���M��QTu�S3H�]�]���4޵�=��+] zS@��m�LX�M���h�S@�Қ{��;)խF)�ȣR8�}��^���f�{ֹ�{��ɀ�gg�!���I�㙴���JG$�v+�c���R�3̑��8�L$2D��^���� =���(_�;z��5�R���N܎�l��=���X��0Y�S3*P���N�W�~�`�ٜ�%�P&�蛺-
�����ﾫ���@�Қ{��=�g	Մ�i�2H�k�hzS@-�h�k��~��Ŕ_�2'�ץ4�/����_�s@���ܼ�	�G�����oEػv(8��k4"�sb�qk2ޭ�����9"��bc����a#rm� =����s�����7x���<��K#�@=�\��_�-�o� �n�B������Q�)��*�n� �ﾬ^�0���S�aT,��#+"V���Z��C��6��n��������kr��Ě�2D��=��د�~4�����h�נ{΅x��)?5"��@=��������
��=޷s@��z�IM��m����û]�<�ܜ�xtbv
�<�ِy.�v��g$�%�E ɑ�< ���h�נ{���%����<�xS](�fjfh������n��	Q&��X��x�w���I6{�²0M|�E�h�}���f�y�Vh�נr��QTSUTUQ(�uV�:D��u����ܓ��{��*"Hā	�3I$%�g����<;'�))!��5w�����G�%��}^��b�m�@��5�G�'/��_��m=�;lu�:=�8y���nn{b���\0Mc�N��%�ȣRE&�˭z{n�{m�~����r�|�M`�1a$I����w�m� ~�xηY�BQ�U����N�V�Tv��t�߿] o�n��L�}Հ�� #W�\U��
�����}3��� r�� 5�xBIf7߾���?���m��%�������%�B���������˽�?u�XAa�B@�A �R ���!��B�{����{߫��Y!�4�e�d��9�8�ⵔ��
��n�k��1Bcaٞ:8�Ȗ���j�d�v��T���׋�4��E�z��K7-�x'n^��ش�W$�MlG�-���	f���m��FI��-͒Y#Iu���Kq6���N��Ŋ&��#���'Dй۷b�c�N�;n���-�}�Q��:��=r��3���v%ՋX��,ޗ5��u��#����l^'٣�=xm���s;�nܺ�ͬ���7F� ��`���w}�����r��	~��Ӏ9�eEr����DĤ� ���z�4_U�u�s~�ؑ��Q��plbYrM ���h��@�n�[�h��Y�D���Q�"�@��Z[w4޳C�Y������y�G$��mn[+�m��z� ���@��Z�ֳs�]�\�s��7]�ls�����I����j��iynܮ����_���w�|�;��rHI&x{女����=���:۹��οd��d*�[�8��릹�*F8��Z,S&����irP����ߧ }݋ 7��|������/�(!4���@��hkŇВ��^����3EtR%$����@�n�w[4WWf���(T�Ͼ���ꚢ�U4���Z��X���BI([O�����8��4�3��_�J 1�(����s]��%�0iݶ�::��e���NxF��{ݨ>O�#Q61,��'�U�����ڴ��fx��女s��5
)��"�9��M�|��wb��� ��x]��MbC���@�n�w^�s���:�?P���v)��H�p�0dV#0,cE"�\A�%`HP�Q�RE�T�	e�J�P�y��r�*�D�#IE��k�$c8����,H�'Ԍ��	!\1v���\0��H�b�� �CV$�`H�`F	�`�I	��!HR�&&ЈAĉX`H͠��D @)K6�fb�\Pʃ�H�3ZD��A���0�7���P�D�%H%aR"x\!����	
J�
�����U��Cc	#JF�e�8�MYi
[�e�Lِ��F��
RT����hA	����$*�����S�Ԃ�#��P�����2&�+�j�L �q�E*�	t�*�.��]nl�IB�H�`H� T�GIAC�*i!��a�1~D� ӻ�� `����H��#׀��|���mSBD:A�L�泺ܓ���݁ע
�FdY��$�4>���}4��׀y�s�ko F��qUut
��M]��t� ���'�}����4�٠wteL��,�$�q&����=�-r�U��;c:��'7-$���2��c~Y"PB`�snO ��-�������Hl���xb�)�S3B&�����ş�
d�e�u�uj���r��c�x�F�4��M��٠{�ՠu�s@�ڔ�Lr(��G$�C�˝��4���7"@"`�A�@hSynd=7�9�;�4[#�H�[�=����ŀ�� ��x�%����߃�׉��ms۞{^y0R�Ƚ�;���ݱQ�gZ5�n�sK���?p��n���>�����z٠z��4yڴ�W�3"Ȧ7!$����~��L�/�� �]Ӏko}	)����J��AT�Z*����׀{i���Q���4��M�Z�,uB`�s�]�}��� }݋ =��B�!(�g���h���b��I3ȤZV�`���=:���� j�����0�+@�fAL���;��O��~�� �F�N(y׎1��e����"�Fݺ�!�v��7tX����ە�]T5�G6֥3��wjr�-n�dg�@���67\Ku��)�)l�0�#����5�-��٭�.͝����瑷Cu���*v�-������7�#��xKQ���N��\B^�`�k�ø.q��s��y���d+E�xXa�N�abX�mӫ����9b�2b�q`l��cn[�ڭ����q7������W��x�`笆#���sp��������o�:4��x&LJL�߿�����@��s�B� ����ɻWw75E9�M��٠{�ՠu�s@=�f� �E3'����)�̭�˙�f��>���[x��$�f'_u�e�u�;�I��v!a5us��I$��w��~�h����v��dŕ�+�R��.�� {[��J;���������h���eqE����s��Z9�&Pˤ�[�m�Ղ�.��1$�鑩����	�rh���ަ� ��/�BK􁯺�ژ�U�R�qIac�@s��z�Θ�I��I cj��00�`$r�`R�	!�J��(�%�݋ w^ {�Y�{�gǅ��fA'���� �|�����:���9z��l��iHE�����J&|�� 5�����8%=�ߖ��=�V]ܗTI2��I�ڬ�=��h۹�u�@��|щ��&
���#�I=x�F	/Jۧ^��&�H#����ex� 73��r)4yڴm��z�������*�?��H��8��-�s@=�f�{j�@���~ċ�Ɉ|�,�4�XϺ��˼��!SV`%H�Q߳���w�wf��g��`�����@=�Y�^v���`}
"g�u��0�WMJ��&������ֹ�:"9��� v�^ s����X��}򍄎V�ʛR\v=��ɰ���X��'��/c�[)��H�]��v����	������>��� ��f�{z��z���W,�ƞ�B�4�m��������/u��;�U-�2dlBY�M����z�>�m�, ��^ �u��2��˕5w5�z}���x����Q�HIP�H@HD�j?�.[ ��E�L`��i�ܓƦ}��Y�]�v������ ���D�,�h�x������{�������~?�� �oO=�^���f��6�v:v7N�f������{(�s�h�b⒪���� �>nk �/]r���;��X/�����(U"�WWx��sX�z� �׋ 7��G��]��W¡�����:�}�h�Po�����zze"��`��z^�����.�=�����*���|���!9��f�˭O@�{kܓ��ݛ�Q�cH�5���-�ll�D����c�[T�hׁ�u���=�

!�X ە�q�l.ݞ��q�Kg����������ڽ���� ��|F�-���}n��>s����[k���P��DwC"�G)��m�����Y[�����7e�qרI�̘M#<ݧ�i8�N����kXkg NF���h.���TY.��	-\ɦ�%��mvW{����~���믐3�חu3�={�]�{��qkN�+��K�'nܹ���s<qb�E~+�ItiL8���W}�z��^�׮�{�Y�_�k�,q��D'"z��^�׮�{��=uy�Q'���]J����U�\����, ���
&\��ӽՀw�U@kβ��d�IV��I,X�Jo�� }��x��u�k׋ !�n�Ĝı�M ���@�{k�:۹���h߽w��4�ۑ��'"�ov<��λv#�lZ밄��5���۶$�<��N��=�icx��jG�����=�w4�z��]k�;ֿT*i�L�8Iu�{[Ş�!B��r�}��<�w-�]�@���6�p��0�Nf�{�� ��np�&}��8��X�l���meU*蛻���B��>�pu�Ӏ{[Ł號k�ƶ�p��WD\Қ������>����}���7���=�v��m������&5�Y1�1�̈́�F�׶X	z��b㳲��d��Q��BcMO�pZ�n�y�f��s�hs�{�~x����&�nf�~�w���5:�ΟN�o C[k3&1�cȤ���ՠyϪ��<��
P�#�c�}B��x(���r��<��q`o�^��KZ��6��3"�<��h����u���ՠU���,��ƙ�r)' ��� �/��[������p�Z�@;:�L�B"4����(~S	6�{6ݣz�H�Jdm=f[նM���]��+��+�h�r� o���]������-���ۚ\/ɽd�A�%����=Φ�>Jd�Ӏk�ŀ�]�%	)����5�I���46H�k�-�n�BP�d�}xtwV�G�˚MM�G��s@<�@�e�B~�� ���"1ʦ��f�/�&<|�"ĚM���u�s-z����n�����<�!)�?|���{�t(�nw"+�f�Q���y.�v�Q5�dq���ı�RO ��|�Ӻ� �o�/����=�I��P��M)�����]�? ��s@<n��g��N��t��R��VUG�w�}����h�V���@�����\1��Bs4?�g�K��4Y�X��u��|�?��� �>��-ؖF��@�e�@�{k�/[��'��w[�i
0&��e�?&b�F�0"BN�dxa�3H��ă ��C���fq�$�)`B`J2�_�O�6o6RD��|Oچ���]&
Y\����@!#ņ����"'¶�i0����{i�C�u��c1��.뙙��fā�*����~R!f ��B Mms`��F4D�����,�?~H31BX�RD�"@�A��]F\)`[y�P��B����� ����C���[�F��4�f�l�I0$�!�3�t�~�!�y�:hQ��V��MX~�!��%t�<>�Ǝ�@���@�8~6��iV/:#P�]~@���HAbhV���˳;��G�;�[u�k@  5�m       %��`  m`檪U�ꭎ�pm!���\�����,燂ݭ@+ʳ�)	�Y�\<�ڻ1I7V��^�}^μۃ$ppv���8�uf�t�li�k��ʱ6��m� M�[m��QUT�Mq�ኲ�듧�����Y���E���E�y5Ǭ&��s�h����.*6�vb�G9\�o;�ɗ�������t�70���l��)�miᆤdqy융��=r	';�P�x�9�v�%��լ�Y܅�[/������v��zŎA�؝ڴW�¼;�($��x8�/[^�u��-YN�C��yz��b9M�N�!�̎w�M:M�u�ko�베�κ��4�gC;�; �	gk�)rc=���f�R<�N�],h�:tSH�*J��N�n�;=���줻�YM�ڳӐ��.Ϊ�Li�3��x+���V�]��^nZ�k7,m�"�	s��$�n����dlm�;���78�Z;�#�n\v6p�	��	�!�
�)��6WF�P)��)k������V��*+�*2K�ʚd�LO8;8��A$���@&�6N�l$3�7MÝ�1;>z�8�kz74;FS	9Sa����������h�qn.��qn�����vۜ�k�mt�se�m��I���ѷ8 �k��l�5�1d7"�a��[����u��f�Y+��@��EΞ�L:�����xN8x�m�ܚ�m�Rƶ�7��ŋg�4[ke�w<���(B٪��A]T��0Wꀝ4�+G]tn�̷��4��sg�ղĠnu���nr�v�ۨ� dU�-k�����$�gi�q�� �1��.z%X�tf[�MI;Z6�jN��H\'NY�&f�&�z��]�(�!�6�Pi�Bޭ�n�ˆ�,0Y�]1NE�a�d�Ψ����X6�I�5m;����ȼ`�*�pLR9��RfMjk3W1@�?��G����z���"�^��
"|�~Et�E*1 H�B�E`���D��D�pNP����g����I�l��N����\˂�H�2�nݰ�#ڷ�L1@%nm�=YB+V5��;P��Xy�Dq���nZ5�m��t�MVt�'lny̾��1��v&�<���pHv8��x����\gt���L�hТ��7.ke�t������l�/m���-\�!���7N)le��9ě2K�N���+��&���Ь�Y��.�7mnf�Jt����������cOa������ٔ|�v�,vv@���\�����=�`�ǖ�Ɲ��2�� �Ss�=o ~z�~��Gu`��}�Ě���c�-�����4̵�����H�Lx,��E�48�s4߯�@��k�;��h��`j��H��E*����}	B�MwV ��N��,	_(�����=�I��R�����MR��}Z� �"7��/�zy�`:�������5ssjWS�Wd+�y�s&�^�q�n�Qss����4mj���1tVR�QB.�����ŀ~�n��M���5�t�<�&�S�r�.���rO���7�p�&Ј��l�~������,�L��q��&�,��=��|�W��=��h�W�_��Y�"3�@��%`/]`m��6^���RݝՀyW�A��S��G�{��hٙ_���Y��@�z������!�r;�n,�u�v�;^͹	��έu��v�&�[ӥ������c�Ύͅ����?��`t7X��_B�� �v, ��6�pbF8)��e�@�z���X��Y�B�=�I��R�����L�wX�}X�x�S
a"F/�"�P�Dt�B�(
0&}{���jo ��EJsB�(E�wXB�o������<�x�:>J+����������I
	9�+��ܷs@�z����Wդ�#X�Qf	�cq4�����صnݺ�hЛ����#�0�罅E��u�����,�`}���Z��[x��_����67�� ����
�������tBIB�wb����5��g�D)��t���USqEX�uwX�0������݋ sϫ ���E$��h�W�u;ݛ�}{�sr~S�D� lE���h�_�Y�B4��
G�[��h�W�[e4W��=���h���❏<���rgkK&��t=c>7���+m�$��i�Kv�	�sv��[g<��ݳ �z��	/�˻�K�CX#>c0��z�)���ؑW�Հs]ذ��g�����])�*���nI�0=�X�o(P�\�|����y��X��`��FAI���ŀl�� �v��B�.����d� ��"�*JWV���`-��? 绫 �M��*`]
/��k����I�ﮏY$6�׬��n�ϥTCwm��tY�]�.�gk��DM�B�	�X���y�ێ��6M�z�մ�G�Ö��-��f#`^뱶)�m�h{<t�v��p|�6j��K=�m��k]t�tm�G�xkG1�J���G��x�����Ʊ�6Ukvܬa�u�MdG� N2�@�[vݕ�'BX�i�����=���mסΩ��i$ۢqי�<��ێ{^{<���-�==��ؤ궠��m��i8&���6���172��O�@�������P�~�|�ک�Jn���M�h�W�{Ż�^���)���� ����b�#I�z�݋ ׯDD�>�0<����)bo���#��u빠^���n�9)�;�,�L9
	QB.�)&h������in�����bŋ=��A�p���ѻ(������Ӷu�^5�=n����ltܾ�lv.�dU$ڙ�? 绫 �ŀko�x���|h�ؾbؔb�m��z�uټCI � 1D)I�� ((S�kS�s@����������26�H�3R]ـko��tB�s�Հk>���Xٕ���8a�����h��@��)�u�s@���TQ�X�c�����u>ߏ �}�����0���pI�#ɌC�r�o!K��F68���1:�:�A� Kv���(�I�z�YM�]��e4W��<^�8�7�CLS�H`��Ή�{���>�u;f �K� `��f�RL�=�S@�z�4PPqҔJ6�� �X
��,I%�;��� ����ً��-�&I�&���.��`��0z�`�)�y�Ef�l�&��;��hz�h��@�z��hŤ�79�qn�t�T����-��v����h��}��墱�C�nT�&���z�hϪ�9^�@�ܔ�<���Ƨ�9����w>�n|��(�}��@�zd��Ď�P�E��mģ�@����-�M�]���Z�=�)U.fdUd��DD)�fq�>}� {Z�k�(�
b�M$�9u���R���Lb�%	�]X��8��Xz[0P���ʤʰt����;�>����&:�ma���pi�v��m�2퇋���z6v7|�v����﾿���s�n���(J?Hk}� ���0x� lHS	"�9^�@��M�]����=�|�9�AA&�A7��ԟ^����h�W�y�+��63$hHp��:�Հ=�s�l�u��{��`u J��0����/>�@�wW�[Ħ��[��\�����	$�I$JG�0�9��ݠ��d�E�z܂��-:���Im�8������q]n5C�E$D^9�(����mW/n��Ö�d��b7����ӁJ5�=i���;��|uh�
�uM�rd�1�B�r���V&h��j ��@�]�I���ak����#%����]��3,�-�u"*ev������d㨕t� ���:ᶛ<ky�i�����������,�'�"]��m�;�vt���X�捸��KB�^���?�
< �n%Z+~z�Jhkx���:}8�ou�Ae�̈��@��Mηs@�����^���d�pq��EJ��L�v`}ذ��p��U9������0�f6J�I-3���^}V���@��Mηs@�q���L1�!L$�@�wW�}�(_?�|x�ŀ=�s��ڒUu��t��^�q{��x�.y0�b!���ە�P����6�i���i��XWu����������n�y�Z����L9\�1�
���m4��iig��,ŚM,y� 
�Q(�1X�:F��(`E��S�@C��~�Y�S&�>���� ~v��B�= ��u��ZEU��>�ӻ^�}���n�ײ~�UD�nL�\�t%�P�;������~��`�U�m��E"�8G�}���o �����u�}�ιT�IZ�x��Q�g�\-G�N�n���ys��<��:�n�8/�������^3���+~����X��8�u� �� �3��B��#prf�y�Z������otD$�Nc�R����j-�@u��M�z����f�iqN"`i�L�$�Fp�@&�~�����������8`C���M�!�1¤(�	)`� m0�JJ�n�(~h`�"��U����ነ����DwI���BL�d �>�²�����*IZA��!d��X��4_�F��YD��J�4YC4��p��~���5�߀�0�`EC��&�\�3{hE�!���$5��lPn%�)x��E>Q:�(g»@����?D��L �4?'�S�:�q @G�],Ph�T
��w?v�I߳���qW�̒%�2	����<�np��p:�;M�`���*��#BD���Z{��=]���)�{��n �8ؑ&<Y1N3>���Ѭld��^t�^v^�Wɞ��#�J<0��E�����^�}���(^��ﾬ��7��܅��U]�U���u�(�2v��z_u`�w�m��H�/�p�=�e4Z��ď��h����0��ii6�U�ف�)�>���׀zw]`yB�+-Ť��htXw���M�9���ߓ]�Y�{���v�����@�u�@.Z�I2�$ka�sv����[q��h+�����.�-��&��Ŭ��A<P�	"�=]����<]k�/>�@��Wds$�Bj�VMU� ���
>UF�}����^���}5�f%�9��Xդ���ـy�t�-�áB��o� }����VXҏ�0d�h��@;�f���h��h{&0ŕE�m�$�@;�f�������ߖ���M ���31.��X�$�}ߵh[hH�t�zo4�֓f�S磶;z�_�>�s9e�K��9�'^m�n���Bؒ�94�(g����-#��d��ҕ�X�-s�R�y�A�^ˇ9�؛�m��s������&竊۶j�s���[XzsOnx����!ֻnإ��a�׻i6��)3,�ڹk�5:c�d�Ie�g&�b7,K`N{\��b)2�B�k�gZ�g�]H�����_|}�	�1�����Z㷱�k�]q�v �ѬgF�\�%�F�v�hI��1�C�L�6ߟ�����ֽ���������u4�16��'�ֽ�������S@-��U��b0�G����N�?�/���=/���l�%K���nnj���v���u�~�n�Vנy��u�`�2	��nـ|�#����{��|���_s�×�tm�3��d6Vy�&U`����s�P�#�X�jsyz�SU��Z+k��٠u����+2�(���E�r���ٙ��PF�����< ��w�nI��^���^�@��1�,���q�#����5�fDD)��}X�� `�]�E�\�ҩ���K�J}�߾0?�=�k��٠w� n�����&H�4U��
��@;�f�m��=�ǅI�!�N3&6�X��/'4nH딶9ζ�Ҫ+A	�ly)Il��,KOM�hb�#�N? �}��@;�f�m���J#��>��2m��*�d������w�
d}���ϫ �m�|�f~�Y!����R��u��\v��}��)%�G���JbD!�(ȏҔ�ו��� ~��ȪV��ꤻ�0:D�7Հ9������l���/E�A�Q`HL#R=��X�O�u��_�u��B���O�p������K��m��znj�&���n���Hrr�e��Z(�y펍mі�G��女��h���Vנ/+̉�?�x7&���oٙ�BJ�s��`?}�`�n��P�G�э��F6�a1��r��r�� �[)�z��b�FH�x	%�W_�}X��׀kv�BO�RQ�t0*@8,d�F�*�D�T� �ʤ4���Y��rhp^DO����\�@�f���h���]k�=��J,Z}�bcczZ�v,�Ք]��Z+�tu���o(�<-5K���k�c�ÈCtf� ﾟ���@�ֽ �޳@����f,�c#h�C@���h�נ{�h�)�{�әA���� qH`:�`�k�>����*����k���:�Fa�* dCn8�z�f����m��t�� M�Y\��PM"�� �v��/����t��V�7�z��řBՙN�KX�m&�tY$'i��?�G�WWQ����S�0F��t�&�;klax��.esn�Ck�W2�)�yn�jY�ѷ��5�4�x�H��--4�Ɩi�m#���'[v^uX]�՝t����l�m�yX)��;��7A�d^Nc6�Y��x�ɚv�t��J���͜�'DЩ۱��a�ᱞ}�m���2���WC�z2u��l���;�ߞ�ﴝ������5��)<���v�qu/yv��ۦ�Oe����,#H�	� cqD�m6�c���--�$�W�ou�J!G��|`��t���yH���p/]g(Q�IU}x�u�`�79�S&д�EH�
jd��)�{�@��4}v�����ب-j<"i5����-�M�]� r��B����>���M�U���I�l����z���Jh�Z�
IY�ap\�sێ
s��b�E��yN�f5m��9���Kh�CpR+����4�)�{��:�Fa�* dCn8�z��~[
�"��f����;f���|�P�A4���E�\�ҩ��{���l��˭z���_<v�ꪕ���09)��� r�� =���)��� 7fa�
Jz�r]����� {�����M�В���\`�θ����^��N�������{�8|����M��5����o%�7�n�D�� ���h�)�{�y� ��@<��W��5����<� ��ܴO�� {��r��;C���ڪ�E�+�� ݮ��6u��a,�S
&e$%A 5�U  �'d���?/�@�Қ���Јn~CvwW8ηX�7x��`|���T�߾0���+�,�UWWWu��w�|�{���n��l�u�yO����;fŬ;gucV��UΜc���ɳ�k\]h��P�q��g��RM�e4}��.����4y:
)�A9#�U�S@s��5�blr�� 7{� �v��S!�3PR_&���4
��= ��f����M�F �Bȣq�g��3��x�_����J"�(���~�Q�s~�nI��Ļ�Yn�CYNM�e4}v��Z��m�z�<���DԘ�R4�X=�ob�=��u��۔:��m����r�kii^�m�#h�C@�Қ.�������Q��� �_uO�rU\ISV
���6u�ϒ����7���� תcYQ"q�#��@�e4�)�n���u`V��rYUrRƤ�[)�^�M����٠w����f&��2D�__U�rm� ?k�[�`��	J���"~F&8���I@C䊑 �P�X	� ��%I!�B"��d+������&�̺M}8I�����ٴ� 1HM�.J�Ct6̄0x��3_h�u��`@��� �ŀ��>V'��A�yÀ&�~`&¾��@8��(�#j��kEp��I4�(�jHa$s�bFД��t2!"�SNT>���8����##�# �Ipe�D�1�3L�@�P�		��ڻ6�H$��&`��HB3?0i�b���`�D0B��QHB#�(�(B���3��}1,X1�����f�d��9Z%,XE"@�@	$	�/{�{~�~x   �6�      �   H�b�8&�t��1CQ�#�3�r��Hi�t�"�\AWl�V�gH�[���l�b.�O�������to(ly�l\	FՉL��x'S������3��;o! K�7;<�.W�Ω܍�{3f�zN�en=q�j� j��#5*��ڝBu9!�<v5۬m�)\r�xG.�#�ш�]����c]WA�;�r䝸���mJ�mz�N��m���u4ds��a	wl����]�^z='p�^e\_1��b;���>�3�p���ƍ>���R�&��:�^�@.�!:�v36��f�ri]��X�'.�m�N3��)[f27n]�'nrZ�M�j[<�5���uE���mE��:��tp@XCiպU���K:$3j�3��2���g��%�/@��N�����>R:��\}$��.�M���{k8`�JB�{v��a��z�}#�ܘ�/c�y7=]zVm6ݷM)�Z���P�z�牲#)���}�nD�@6ډv��-0n�n�ʈ<���.&ԯ#A��}�v�%��sBv�Z^ϟ9bd�t�����5u��s&�+n3jٌM��]�x��C��&��9��]����/h��n<��Ź�s��v;����G:$��6����`]�'���ƱkI��3m�.�9�P��\�k�np ��6zg��wc�n�lv��ˉΔػ�T��R؍[�+�<qc!����ն�'�`pu�:�����Xp��\�o���l�ځj���΢`ت���������j�eV�GA�����k�^��70�+�e����%�u�5S�/�hu���v��ըX;`�k�C�.��ݐ�ó:�nl�"�p���&�k9�[k6a�:��m{$9m�U��VBUn�Y	�]&��ƙEF �4צ�Zl�H���D�˛�:�#�7B�k�ܼYs�)d�=�kU��]����i�V�{���w绻��ܪpN<�QV.*3�����|��u��'� �����o{���;��?Bt 4�n].⇘�q���f�rƛ;Nۓ�7k�1A{5��]��g��n�+Wgf�<�u6*�M�}�+Rh&BnV#GH*K9��ؗy���q�F��Ʉ}c�5.�ҫ�ݬ��(0�vޏϞ�����6��q0����w7;;����޶Ą��ڬ��rq��<�����/i�t�<,�8���.���ӊu����~��/��y��)\u[9�v�\��6�nI��a�!:^�ym�f]��v�������54E�8���= �����h��h��0h��E�@�����k�g[��IL�|���4�4���;�Ɓ}}V��D˗�X����n�ꪉ�U*D�$��}}V�˭z}�4?�}��h����D)�NE�r�^���������__U�x�v$�)��q��� ��<9��Ɲl�Z�\v捍��Y��D\��ۣ+3O�m���,�=�S@���@�ֽ���Ue��!��@s޾5但|�FI-�Db�I�J�ʮ��}�X ���D���ǉ����c�H�4�ߖ�˭z}�4m��}K� Ǚ[H��]����� ?k���09(�=������>@��(�z}�4m��/���9u�@<�慎�K�z�u˶/v�E�'ݎ�]��퉴��Z{so驲����Nx6�k������ ~�s�l�u�|��Ͼ��}Y7#,�D��m���'|��bI,l���V v����3��=+�O�7dU������ ~�x~��R%	D$��P�D*�yx`ծpz��)NKrUU���`|�S=�� ��� ~}V�˭zYqr�,Ȝ�xԓ@�v���/��_u`���ߣ�����7a	�D}���u�ju�n���*=��s�DƩ����,R(P�;�F��s�-�Z���h�)���p���h�)�@�ֽ����}x�_��u�=�AL� �Bȣq������i���/W}��*�|�/b�-Dh�x�G�@�v�����6u�����JbQE�K�yb��}��9��5;Ti�����?O���P��W��׀y�f��;�J�X�U	DDeN�K0RE��/O:���M8U��a�
�y3��c@j�ΐN8�]k�}�4m��<^������˅	%�[4�w�_�$�ɽ������6u�ϒIDɲ�O�δ�(48�������|����"S._u`���=+Am@��h����@�{k�9u�@=���=�S@=�,�!�Q��"���]k�?�$��ou�~�7XE�i^�t-�lnΤK9��GR�T�j��Q��"Sm B�۵vv79'T�x�m����8��v����F�&c:w8��8�w)nxx#\�nc���&�?���l��xl�[sl�^Lm��k��p���%r=ZEnq��P��� �S��k��mz��j�n8�`^�x̯�q���[ZWiB�[�N 9��<������HU(Zݑ���TIՏ�ǋ[�c��Io.V�`v�\[s�u�&����%�oV�q��iv�vl�7ˏ�-�h�)�x����נy{�LPy� �'&����ٙ����U/� �ﾬ ���}
d��U�!I�b�������נ��h�)�x�ێ�$��$�=��0��x��`tG�"���V�r�g�'�Mě����h�)�x�����hڮ���F�?�d����۶=mr�t�u��8n�#�5��^K�=�m4$�u�ZE�Q�v~��h�{�@�s@=���=Y����b�1�.��?O��!-P�l(�4U7� =�@��M �Ըć�D�$n=u�X�k�?�L�u�zw���l`��4�(�s4?߱.���;�Ɓ��נw[��y{Ѽx�BA�]�nـ|�I/V�W��ŀ�Y�{m���"��Ȍx�,b������<����^K����ع���-��[E����JHh/mzu��}�>�������Dɲ����3%�d��� ��� �����0��� ת������M�܆�{�Y�u�����5�D�J���S��.+�Yb�s�/�)�z���cY�9�Ğ5%�ݳ �>n��x�:���׀r�
����Ls	��{z���s@;�f���M�lxT�2�i(��d��udt]��e��;�<6!��[v3���,1��X�(,liiI4��� �m���4��h��*<CM%3uSV�|��%&�0y���w4=�WF��M	q94oJh���;�w4��h�V�����U�wf%
������ >���rf�'b�#T`��C��ŋk��٠:�_|�ZaI]��7�l��w�~{l�=w�tD.{�On�H�-�&[X� ���yP��nޖ�iX�i�9-��k5j�<�\^��D) /}��<�)�޳@�zS@坋���(�xԓ@����Wk�}�� ~n�!L���:G)�&9���@�[��;ޔ��@����ﯟ��bH�5#�;ޔ��� ����'�����'�R�mbQ�!��f��}V�Wuz߾�f�4��R&$$M`>8�~~�?u�UUN��ݬ�g��.
5��J��p�4V���nڹy�[��6x$K���n�j���pj�qL���|��!���d�mѫ�U�(���p=<���W������8�C�����I-�l�d���2�"�]��qu�u�kp0�u�9��GW��� �V��c�0!l�6��ҌV��m�8��Lv�ř�l�p�7ӊ:�t���{���X�u.k�ҍ��5(Yv֘nv-Ϛ�g�pqCl�ŻyoQ[<.��s�#ǎ���rz���hwW�w�l�?H�׀wOVMMhAt�ʫ��U�^�����_m���Z���Ib�0�O�8���4��hW�h{��ܹ?�⟣���4�]��k�ϵ�)z���Z��Q�%1�&��}V�W�^�����_z�e�1T���z��b=���le��<6^ͳv7N�,�Y�-$趓i�uL���#��[%|�������y��@�����<U!6�qǹ'߾�f�`�E"�Y�!�� E"@BR��� (�$���$���h{���~��H�*����k�� ���@�@�ޯ@�zS@�+�x�B1�q94+��J`�`t�k��;���*���]'�Z��?߯]�����y_U�{Aց���F��$H����c#�`뀳���-U���ݜ�ͫ`8m�Ɛ�$4��4��hW�h�S@����ŗ�	��!��f��}V�}�M��M�1#��*���p%j���u>��m�:Q����8���?f���9�<>�N;]��pJE�Du�FE�T�>5�I�w��Q8��A ������΢p������ݓ��B ��$�Kk$��d0��H�Y5G	�5� � E��V[#�#7]��~�D��H�nc2iS�4�!$#!#<9v'��G_-@�,��A�HE��SE��F���`Z2m�J}��)�&�w�S`�n�@����@����?o\ z �"�)�u��N}��q"f�&�o	#� �
�w�q_��8pHH�3�?}��4��&�\V)1π�]������i��t���P�\�~�$C? Ϡ��	Hh����X*��$`���
�P���@��4�D��|�Ӱ0� U*� 9���Q����(
 |�ٙ�Z}�ƀ7�z��`��c	Z�����%<�q�=w� ?7x�fc���=��Li��i�6�"�h�Қ}�hW�h�S@��%l@�3z\6��3x�0\k�j"{uxx�g�'���m<�=��[w��d�����|���k���9B_��� �򛟞<p�i #�ɠy_U�^�M��� ~n�%2wOVMU*�At���Z��M��M ��4+�������b$$�{Қ}�nI��ݻ���E�0�A���S��ٯs�ܓ�<i�:]:�q
C@/����� ��h�O�\��@��Ie��¡�j�:�+n��j ���uM:D6�u���Yn�1*bhƖG`�5$�~w�����΄����x�`N��$*�-U�\��w��)��0���ε�t�����<_,M�"RM��}�hW�h�@���LhTm���UفТg���u>� {����4=��^,p�i #�ɠy_U�u���f ?7x�ЈP�(]߿����,� i6ˣ��9�npl�IM�<�omى�����[�<Ȉ�<���ۣ��Pmc@�8幵<� ;a���ݬ�hX��[��n7.�ȸ�ی�2�9��#n���<X���Z��ۨ�og<�� �(��i��h��	���	űk�����2�n�r	#���4���\��Bggc6����Nll�6�g�����;�}6O{���%ŉ$����E��-rJӵ�(n��i��cؑ��{�Ghum����r�X�0�#�pnE��w��;ޔ��@�@�zZ	7�?�"A�I�w�����ֹ���>��;c����Ю�5W$ݘ��x�Z��';��/Y�U�.v_��,JcRM��� ��h�Jh�٠x��gc��x�0�Š����M ��4+�
���6�X��l&<<�ݷ�8�ǒ&�^�ae���Y�b����k�|rx��ؒ �$�;ޔ��@�@/u�����I�bQ�!�����oc�!� )����DMf©�= ����M�j2W�#H�rh+���@�zS@/��Ъ��y�ۃr- ��h�Jh�٠y_U�}���/��/�2L$�zύ ��4+���:!%�n�E3�R������H9s�ڝ���9�ȷ�Mm*sr=\�4/��R#Ϥ1LS#�7�< ���h+���@�zS@��\�����,JcRM�z� ��h����lۉ��e͘f,O�
8��Y�r����|>�4! �41��D?*!� ���B�%Qt|���~V�V�J�R�MQ3$��/z� ��4���Y�\�ΘЕBM��I�_m���z{��9{����4,t��M�H}�/c^�/�n1tR���ʺ�ͭ=���t͛6����ƒ8����z{��=��h�٠w�{�n$��'#��f��>�@/���ֽ��U L��I&��>�@/���ֽ ��h���.(�G�nus����u����RP
!'B�E�  ��A2/�1X��^�����Th��uGm��[� z���s�����w���C=P� �����Pv���pO����[�$�=��p@v�����35h�������=��p����C�~��ο��DI�{�l��w�~�n��S�艓���З�I�bPnC@>��x�ק߿~H��Ϧ��ύΨ�^,�&6,XG�@�u�@/�,�=���f����M�#ۃr- �ܳ@��ـu��i��5G�H�(LJR]{�~��: ��̺u�{[ptڪF���[p%��葡L��D6�,r�@�4�����3�t�s�ݮ���;�im�9��R�X^cksˍ�x֭�.zrt�'�6�B
λ]���V��ە"��9�#s���`/�'V���{]�s�n�7#���0ys����.��,3,��q�9�I4�Ѱ��V�C�7Dn�y):�(��nd�u��S�O�z��h�DG��k "���q�b73ݝ��Z�ԐpGY]5������6��6����c�{s�����{��`�w�~�np��x����)�<pJC@/u���Z}�f��t��U��b���)�94:�h����gƀ}o�@�_�vX	�I�"p�s��=��h�f�岚z��Hx�M"Y$�;�U�����h��h��?;���?����W�7��\s;��q���Y�B�i0^��bn=Z�&ݷ6��1(9"���@��M �:ϳ����=�$ɍ��$�<�Sz�SqsN�X��'�!�خ		"	��@����*1	@����G���� �W�N {[��-oX��0�F�$��{�l�;�U�r�^�岚+QR"�c$��$�s�]k�<�ՠܶh{��sS򀛂�-�Z�+�h�-�s�������RH��ϻ��[��N��#���^�^�t p[�-^K��;{rГ��K��"�����?���}���@�}V�˭z��3��0o��%#�n[4��h�נx��@�������� ŒM��[�}~�ss�$����B~{��=��_����LthT&��A����Z���ۖ���Z��dYcɏ, ��@�[^�{r٠w>�@�v�������N8��LF<�;b�Opf�/<�������=�:�C�.[X�#�&�8�n	�� �女����ڴ����R8~1�a�d�@�}V���Z�ڴU�^�ײ~��%�
8(��;��@�[^��k�;�U�U��\s(�7�]���D(I)�_t�<�� ݭs�v21�-K �A#KE�J�! X�)D�2�
J�?آ?���7˹'��Ϡ7�I�"�=W-zs��j�<�ՠu��i��dlM�Y6���'$[�;�L��v��l��k7K�1���LM"�H���h�W�y]�@:�Y�y:4��bPww8��Y����������s�l�~e��TN4R�^���:�Y�w>�@����-آ����*���B�����i���\�W�h.�T�	���`ɒM��f=
!C�}> ��`��� "��Ҡ"��¨�����@EW��_�U�TU�DC��B"�T �B0T �)BB(AP�T �!B,�T EP�$�T"$��P��
�P�B*� �T �AP�� AP��T B(�T"��T ��P�,��T"AP�B"�T �B �P�BAP��P�0�EP�$�T �T  ��B �B�EB� AP�0T"��P�B,T �P�P�AP�B�0T"T"�T"EB
�T"��P���P� 0 AP� �T"��U�,B(�(T �@T �B"U
��T"�AP�(@T 0T  �T  0���0B
DT T!P�UaB!P�0T"�EBAP��AP�)BP�B@	BD	B@T"�T!BDT"�T"$ @T +P��B
�P�0BAB(AP�)  �?�**�� �*����PU����@EW����Ҡ"��
������*������"��"����
�2���	8������9�>����@I &�  h
� R� B�P�T� � UT �� xJ*�BP��
$
%%P@	JRR�����H��PU@R@JTD( �
B� @`     {8     
P�h|[�>�����n�iI�AB�zX������#�s�>ރ����^�A��^�  �y�N^��ϸ h��ǣϼ�^C���g� 0��v}���x��6��������f�� ���@   �A�4�O���{�6����g<�Wy]��6���}��E����˘r�nfT���yP�\���� 8̝�Q]���<��ooW��-o�o�x�>��s�j�v=��{��X�||�  �*�@� ��������x��bi@R�)JQ���B��r�R��tQJX� )��R�� t��14 ���  
R��J(͔�(`M;)J&�)LM�b�Fl�����&�
14��7Y� bh(� x�  @   {�F�)J3e�1��R�}�t�®� ���Y=��<Gz�<MOm����@t������ ��\���2����/)1۟v牥�N����Y�vW�����{9t�� >=J    JP �2�[��g�=q�g[�D�� ��{6�k��69d���`=��9f����� ���{��^� �����M��^l�y�/)]��y,m�py�{j��{��zU�  ��ԓ�*UA���ha��)J��` !��=U*T`   ��U*M�T��d ��M#jR�  �!JP�d1OA?�����k��l�M�ϧ���\���_�PAU�5���
��T�
��
*��PAU�
��z'��A���ҩ�Z���?�ƴ��/2_�ż*(¤l	$�b������H�yb�|�zm������(R'7���B�)W��S~Վn%!d�ޥX� w>S�b2Z�R�&�W���BB����ܼ��y(��i�M�J0��x�	"x��"FF'��n��)&�A$"��#M�rO=�$��X�o�,������H2d)�0N?����(�'�@+��(c�F�(A��$�>A�h�b��"QHXI4|m��K��A p}+`�"�X\�\��0B0#�4�����D�!�,d^sk�İj�T��Hr�:[��2qYu0<]y�Y�Z�#�5b'0��I�"�9�f�Sr����<�H	
f�͙��j�z���D</�
`P&�s�D�!L)sF�cǁ
��#��k9���B5�n��
a�e4��a��:4��|5�Q��%�-�^??Z��hbVJMAYQ���)y\%W;�r�M����x�6�yEL�kbixr9�ޡ�
�2J��X��R���^[���2[����i�^�<�we�SR@����V�T� u;�'�)g�WY��ÿ�2�$c�	 �ܜq��w˞}�؋*T�JRMV�{HA�X��A��+i DH�)@��E�,� �
"B" U[;c�����Bi��J�ܺ����վ��(i!C�*�� h1Ѱ�a�XZ�D(D#�0ie�
S{3˻�up������)��a��`B���.]`J��8��)��L�홄�o�M��<�H ;R�a$�Ɂ0�H�&hN�e��ﰞZjCQjE�F�h,*b�h$�򘒘�@ۤ�\t�!�%��S0���	�� E�!�,`L�s7HRY�'�(LRV�7w^�P�i�.�^Q�d<�8m	�D�C�R����Ҹ��[�&�@&��P�H~?Nd�7�����N
BjP��hW�M5��ըМV��gx"_A1�Dl�%����xkh�H8¹�h��l�!�
��r-�?�
xģ��n�N1�4������BP���@ نR�2k�]!T�B�WJ���B�pw���_�7�k�{t�BB)D�+	!-�QkD��� V1�9�� �#\x��$�L`@�d#L$�,�rjl�9�ܒz�H��.���ha�ڌ)� �l1�"} >1���@�h��Be!%>$#�(@" "FE�"�`���dR, �H,�^B�M$I	���a,��7�����l!Td�`���0���
� � 䐒Hd�HF���> �f�5#d)�����B$ Hbm&��!���Č���"a�(i�B��6a��I%7�R0$ٷk��� �pv���sDf{�D�v��RdI���=cFF�R�sF�@��!BI��%�`��xi�5�|���D�X��$V�!@��$(�T��R����o�� D��¡8 ���O$v�
+	Y	
���9	y8�Kʒ@'P�D�Q0X4p� Xę^p2L�h�%�^�<����SD4�M$H�[X1����j���4��n�o���N*�Œ:Ռ$p((Q�B��R���\n,`�p�B+��E��AF!Ja|�xE��}�0`\��#pIS"BD��qe��7��a�P��S :.��&�I��EIi-��>:%<����V�
�.:�F��6�"C±�j�0��H\5]�B�e1v�d��a|n���)S��Ca",�HJ�bȏ-S��&6�����Hk�CN�w#
�i��l`M��q���d�ݎ�D��"%]ԥ�6�*Ĵ��L��IN�\H1��͌�I,$HH��N-�<>J� �4i��O
o��c�)�-
�kR��g��!���\�o��=@�V>	�  4B���� �hx1(��CcC�+�H4ƺJ)L+��
a��#��:��j��8
�k�;J�ѐ#���m�kl����.��k-&6JI@i��	.��{�	�D��%!���kHXY�	�X!"�;�/����=6��0 B�
C��i�M]D���]�0���y�$K
�a�Fk�3�m�ia\5�n��ָ�I����T��Hni\r42���t%�j~�U����T!8�'[un���Aj�k��Z*�inm�T���l �L��9*�A:hA��1�`,h �D�,�7�w[BF4��\���$�@���q(���L��ջ~u�|�Z!�&�yi�#2�!C�˗%�VR��Mp�# �0�<�d,3����	��f�
��\@�HF�Mq��]�vl���Bk[��q�CaH�Jx�FH�$I`HW��k>jD�9G1�4�~X�Ҙ�*�(!��  n�%�c>߇!##`�T�@�,lh�D$B1HH0bBEl$J��,e	L!��¤H4"�!J��;H50�P�0�'#Dq��jos_��r)�W
�����0h�~��4Eb�H;�d�~kD*��c�#�a@�IJ�d��ѤK! �ɲ>c<�i7Ï�=>M�4��i�9�z9IS����&R����(F�A��sD�\��3Qds4��m� ��-Tc��n��*G3T��n���� SL+�
�k,\��9����ѡi��4�H�Ji�l��k�5�O�A	�$J%����r	�����Ѡ��1��5�,ME�dcH���	����1���h��cL�:a�q��!B8h�)�y��U0cBq�r)D�0%1q�{�g��s�sP�Q1c���X@�:aR$`�v���|��&�h���bHR�,hbB%k��ԛ1�a\52��欼.����5��*A�ɛ�|י�ٌa�$r��m$H�F��Ywy�9�Ii�|���D-k�s�Q�M� &��]�%<��r��E)IT"�'s�VF�K�h!@�D[��w��|(IXD�$H�r�|�Y.Zk�ژD�1��zԌ�)�#��F�C�!	NBw��.�yĕ�o�fۭ��y��j@�.���.r21�B�7��щ�6h��!9�ٓ��tJn��>���	p�.0�H���ˁLfa.��
�
ć�!�Blaa�|n$��ևI��i��<]0�[�hM��o�Sg���[v�&ī���}�g���}9��8Hnq�^1�t��u�n��MY��!9���;��G�r�=���'���=�7�w���.�oT�8~�z��.����4��U�#��%�� C]	�H{�����!H�<��¸C�8D�ƥ �U�Œ5W�r��y`�UY����#� ��i�tLR_~:��oZ�6���HT�컼��s1��r�T�i���ԇ4B䆝��B74^�P�!�Mʨ-'iZ������&�C�f}.B�LB0����ɉ���o	XX\6&�\��dk\���~�&��H�5R���<�4)��T"�S^j���<��o���B�0�J�
{�KD}�`�,	$$���(��Ho9���`x"Č�B!E(F&��My,d��)Ĭa���,!���D�	O��~ۃ�"Kϒ|8h�$ X6����= ���0��\�!��8q4c��K��h���C$=%36�X�CabX@��kpٰ�L	v�,����la�H����{��_�5��v;Œ��FD�y��U�/
*gm���5ԬNiZq!A՜���'��XS0�0��[|L5���Ԛ����G5H�� @��%2�`f��y��iÁ��F�᳁�ơ�rf�Cw{�}	B���.�����F":v��BE���E���B� q+��,� ��-�ō1�$)!ƚ����Ͼ9�y�zXHЮ0,��V@�(��!ᇱ���cc	 R������n
��e��5�\��~�0����@�|�4˳�����}�>�  ��    u�   h�    ?P|          p   ��     ]W-�  8        [@�-� 6� � � ��        m�p �JM���$8޶۶�ga��l-�	��V��=�m�r�#U��v��讆q�k��?w� ��|�1���)\[e �VI��W����ڶ1%��g&�R��a�U�:�o�||�-$Z�]�ڥn2J�T��-�mGZ��l[\-�����t��8�z�Z���^�� _Z�v��ے�}k���9�z�-R{ciU�p ��-���j�$�Z���N�
�֔)l��Kv�3n욜�����.��@�eG��ã\EL7kr��5<++�ʤ�V���n]u�Z$
�wl�����V�t�ep׵�.H{m�CGk�-��*7GeI��Jt��5�Y�m����Xv���M��y���hLI �Ui�[q�=�c��9��@$$&֦��m�A'm��I2;m�a��p�a�^�����WnzV�m�H�8      �� s��� 6��2�6صz���u�^ l�k$���֓��Z:��k�݇� 5�� ր m�p�	  A�F�$���3���]WU����v��YZ�?_ϭ�� *���e�sM),�UE�m��m� ����p��඀�OER�[R��aUU�c3m�qq�Uy��ڨ٨�ӶqD�[N=���   p       [A�Ku��p��K��@l63��� પw@A\�t�-�m�ͧ�!m^����5�j��P��G(MU�+��b�A>ފƻt�Z���.���i�hS14��� �"�[��6 {Y�V;v��c�S�,����٪����Ul�x���J$�nV�V�%��2r���mR�j��b�ѶP���54�qr:'Un0��⭪�����+�EyV�[\�T�Z��m��. y���RLi �Zݝ����SmG��N�>~�Wնb\;&ī�uR��-�P��#s��G5T �Sf�I��᭠'@ �� �%koIz�{wUV�& �[��y��89V�^P'vJ��P�bn�ݷS��kJ��P|�zی����q�2.����b��ڂN�uv۔��;5̍�!�'Y54����ң=��K��ޢB�1 �ml	l��2��U[��-[TuR9P63Ɗ����q l��0i�rtհm�I�� 9�KZ���67��*�vaê����n� 	6� l��� q���Ĝ���$���kC�Ó�Z�kT�`�
3�e<	�Ps�]J��JV�xc�r@7k�����}�;��),�Q�V���]\�����n�'e�0����5��;pj�7R��W%T���f��Wf�[��mV^7U�ձv8����u�d&�����L����}����d&��6uɴ�T��8	 �m�M���ځ�Er�h�	 l�5��k&u�e�q�m��Y@��$ְl��K%�I�@[M���:�y�*m�N� ����N�[p�m��m���ݖ��ۛY5��6������ų-�`۶��U�����ڙv2o�յ��@@UBti�Zv�4Sl��I&��r��6Zm��'�l[�i	m�����U	�eZ�N�pS�\����k�ɰ�^�	&�\�ⶐ�Q��!gN�K3M�([!�8-k�j8�j�)=���ҨmvM��3 "���s��z4 0e�Է�*��[�݀j����[J��UW[uʼ�JյKkm�������&PJ��m@n�C�n�W����Ğ��a�N{/=X C�.˃J�4����[��	ezM� '��)Ie@h�X�z^j����-�	 ��6ۖhM�1m��P�0I�©V�&�5A*�j���}��H�i��z�$ m6�H�I�q@.�n�Vn��8 �	���#��	���Uj�yf�a�փtIzvն(I��V��kUT�J��H�	 ���-�I���	-�iq"N�����%��j�caS2i(�U�5A=Xv%�P-:6j��-�V��ܶ� ��6��iYm t�� �I�m�m�lB� �� -���u�I� kXl�.��&[)��' Ik+�m#+��Y��IA�o0�   [%kZmpH���l�۶3�Im��  ��--7bڵ;]�m$�"q4�^���rI����u	p�R�ʖZ�Y͍=�R[-ғ�t�����J��0 ��Ӗ���l$�M��^� ulHF��=����4T�/#A�m�)Y+n�V���v�p�m�g�.�ur�hņm�\�r��[weUNRVV�a���WM�N�d�n��a���oG\n�/)-�I� dֲAt���\�z1�lm&m�	�m���6���fٹjDۮ���m����m�m6�o����\�h�P�� �e2V1��P�5PS�ݶ �$  #�m���88�6��EbZ[vձ�n�hFBU�X�V��tR���Xi !���H$�M�W6Ͱ 2[��m&-��i�l$Y`  ��6N�LͶ���`�Wl(�I�.�$�V	8��rM��/Z�-� ��۽��7mͰ��m��t�I�J�m�����)�#l��m�L�m��D�R m۶m�k�I�\%��8U[ml�6��+�)l�khXͶ���m��+#2�ˎ��T���8	�t�������ɜnٶ�@6ض�T����)8�UVQ�>��p�#icn�Sm�ꮧ��+[@]� ۵V�z�&U�6��D��U Uj�-��GN'i^�Z�]7*Ւ#�SE
\�TR��fQ�*�O�7��~��m 6ʹ�l�����I���7[J�U�q�rpΖսI۶�A��kdpZh����g8 ����	e$�m�m��Y�u�[@$m�ֶհ:cm�,�����Bۃl٤ZM���m�m���m��&I%ٷ` m]Z���[M�e��i
)�*�T�PmFJ����� � �na5Q)wK��ʥ�.³kaC��n��P�8�L�j` ت*� $���Ƈ[m�����ӡ�m�&Kk8�I�( ��gm�6�!����kh  �.�m�h�0��ڳ
 ,0�h ݶH��'l��6� ��kkn���꾪i��TT�R�F�(�ep[N[�N� 	�=U�t�m74�� ��%]��R��5U@U �4�ZI-���6� 9<X;H �]F�j�� �m� 6��Ulr@m�d�I���m�l=J8 �����m�R�*��,t�<��P�D��V1UR��MJ�ԫ*J�T�-PO7�M�0�l�n�m� 8��� m[֒� �` iX����  iʵ*ʫ�K9U�[h��m�oW�Y��0  m�ť��m���� �&�֭���6�lm  $�  �e�mk ph�-��5�$m�8`  6�! Im	�^�d]���e���v�:N �P�;R��v��8 �l -�� �Z��ޤr�	�[@�ͭ�͛bA�͛`   �`m�$ �� ڶm�u��*Ҫ��T	�5UM�\��ZU������h 궪����W�@t�J�l�	 u�ѵY@�Z�jU�����j�`HH��M� 6݀�6��"H;-�-�[%$��붪B�]0��۳l h��J�רඃ�,SZ��l� �`֛bA���v�KdI�Ŵ�[v�& +��`U��]U$
ÕVm�Y��  H�y��k��*NW^�$l��h��T�(R�UUT�

^������$嚠*�h��m��L����[.�̪�UUJ����  ]Kp6̴$ $Hk�7m�6�m�h�8p �����ݐ�   $   ֵ�8�h ��m�kymŴۗlV�5Q���Z(�v9�j��
�GM=<U����չ�M��8c�	e�cm&IĀ p6�m � ���A�[j@���͖�8 m6cm� ��|  �[��r�M�� �� �-��  $�  �	H [@���EI�m�m��`�� �]�Ŵ �!t���k� ��d]���]6��a    -���հ�`   �����!�ll�m��� -� p@$�7J�*���P+�X*Bj���q�+0�m*��86ۀpH  ��(ְ�l
P�lձ��� �u�-��:�p6�l�Q�Im��6L�P�R��i�V����Cd9�^�����ٶ���^VU�)��ڶ��UP ��'l�U�n  ݛ`  H�6m�h -���� ��`ְu���m���[� � @6�0[uvŴ��I�6�t ��w���w����{����<���?�� L;����O�<B�H��bm�WJ�A��x��<SГ�J��|}��%�81@� D=Ј�Q�EY��� �ҧ��3���S�	x�r��D=�؞�S�/A�B��b!V���1@tJ�����/�H(E�"���J� �O��	�S� �b��>I�c��(x'H A�B��]����� ���Q��+�����M�➆�+�F?)��@8{�!調 &�(a��Qx�l~__GA���m�~{�  ��ڶ�D�Phа�A�UB&EA��B,RV �	��P�*|�=��LC�T�D	�E_�P�"��8& *h$ h���(:���C *	�|�Q�}u��0�0H���@P|�&�L^8���8zD0�@"���T1|��(���q��)��4��ӊ��"ߔ7h:'�~
�`�(@�"P�D(���DB8��]����>V 1CT�"D��H��2�"�$���<D�
	D"k@�a�(�>�� �)��B��Y aB�D!t ஓ�HC��Q}6����^@�XA�|Q�I���!�� ��~~D�@���"H#1�)'�����0� O�}`�<U� $B �ja�~F*�i����� 1B˱�U= � ��Lvx���*�Q���)
Qe�H�N(U*1���UTYT:T�-w.�$�I-�����` d M���l�E�6� Y��*҅�޹���+U�5�[j:��(	�xEc�v�5,�Nv�p���sl���Z�5J���4��+O^�nU�c`��� 6x-� �@�m������2�t]n���.W��P�@C��	�)d8k�JB���6�֞����*��	�E��<�s�P`��cqԥ�&8���v�mv�{/-�������0���Aug=t��K����M���eu�!�t��/���S����W2c��[+�:+1m*Q�Q�ή8����,���&�O�֮0nU,u�N�]*�dd���֭awe�&u����F�nI�U�Hv�tGl\nBvv�j�T��v|�a�YĆ���h�$�N�-0�ۇ�� �H��Θ����̚�R���ng
�<hx��[�gH4.7m(Oi0�F�`.�S���¥T�^!m�U�QڵϢ�V�V�1ٳ�єC6���:wMt���ɷN�E�
�������Y�]lm�*[���y�v�  �h���{���j��v�.�@v�q�e��Y^�٘+r�2�
��e�S�k9�:aȻ5�w�8�ð �'@�k��5a�f5�n��u<��;)����ݍ�;�D��5Ѫޡ�'�3�A�Ԯ���x��m�۵�ź,Wn%;&���n�`W�����Qt�++�V�Ѷ�G��*�ٻnI�WQt���c<yzK���7m�UԫÞ��M9l�[:�8�4�bR2����kT�v�9avV�p)5=�]����GR�;AX�kM�NР4�p4��xٺ{&WU����N�zuR�dxE�s�Z6�2-u�EablFP�Vؘ�OS��fN��n{t\�̯N�p'@6�Sm��rל��zMu:�da˃M۪���lJ Ö�u+�]�L]s$�����Ӕ��ʶ��\����L�� ������vpl���۵E�,\ܖΎw4�\��[Jݢ8�q�\ڭ������*O�~Q��� �#`���)��`���C��`�;@_��J�x ? m|�AGB0��sW32��fd��ۗ%�����v�CD�kt�6t�.t��'iۚӉf�w7vٚz8��]gl<�Zq�]�ۉ;pٶڻv:�aD(b��#om۵��$X{[�oGm�+v�6l�"��ݶ۵��$8��A�nt�U��'G�Q�f����hRWSۭ�nݺ�#��:��t�՟j@I:O;i�^��9�k5�7u��a���MG��w�����ww��w��w��p���)����vG���8��6�ۃ&^���� ����G3-��J�7��6u�������q-|�rҷI�ـr^�Y꯾� ��x6y��� ݩN��vU��N�Ӧ�nǀݏ ��%�E���`��+�wCE]��{����r^�X;���֭FZ-QV��x�`�� N�x���T�v��`����b{Q�8�oS�K�n�4qm���d�f�\,I�j�^]<��Ͷp��y`�ǀݏ �� ��W�&�*U%32��{z��^��j����!�I���nI�=�� 佨�Q-W.�cT;T��x���	�p�9/j, ����m�	�i��ʵj��'u� 佨�wc��ǀEKU�էJ�f�{Q`�ǀݏ ����|�VZ��Nd`Z���A��1�$yc�F�e�ج�M;�����v������4� {g� ov<w\0Kڋ ;F���Wj�m��c�'u� 佨�wc�}�$v�jיh,�6YrN�ɧ �/�ݪ�RЬB;��\��D�9�/ 7v<�E'Ɏ���1���`��v^ ov<w\0jV�N�Eհ����"����ǀw���3�W;��G5m|�(�%C�Z���[uV#�Sh��8rQGS��ô�Q���Gi;?Ͷ���~�lN��{Q`we�Tۥn��r�V�ܜ?va�I*M���k���x���@��D�wui�lM�%ʋ ��/URD�� ����;��%We[O���7�uwe��Ǆ���}7'�@���%D�D�T�B��.I%i(���U�o��┡���[w���� ����|k��V��w$�V�����ga溴��[;]մ�"-��sd\CX3s�	2�U�[E���6~� ����~T�����;���8KWv�#�;u����:���wc�9�2��V�N�Eհ���o ����ݏ����N�oV�����"�%��Z�+w��ꤤ�xg���r\����xU6�B۲�N�Wv�͓ ��f�י����8�%UąL�����r�K�K�6ۖ��r7XZ�nyƸf�)�/b4���+c�.�qq�V눥j�ާWQI���l�lnxv99�I��c�9�t:���<�n&��b���������6-�>�8�H�Sb���M6-a�8ţs�Ք�5�:e�[���AR�dd��{'"�ӝtA�* �%��;9��2�XL�n��m��Y��quc�DΊ�pf�x��?�������;r�`�H8�;i�.�N2NzW^�:�tN�ӥ��`{�Eq�tr��+��M�ۭ}{^XV� ���l�XvS��J�i��'n��:�e�ﾤ�I�v{�X%ʋ 7EF�WE�����cn�wc�9�Z�3��;�w��ŻN_Q)�4RE�����v{ܬ��W�ջ/ 7v<v�I�c���Lk�u�r\��۽V��Vou��	(^��?N�+r,�Xx��0�|�\j��<ې��su�e�x�S�6�.<�yW����<�wc�9�e{� ���y�{"�.��-������9�mjC�M���1HE�;b��a�K�I%�
a(W�z�Ձ�:�v��xU6�KM��N�Wv�͓+ �Q`wc�ݏ �MUj�i]��DK�����?�5k�s6p��<�&Vݔ�(Һ��'Bi�X���wc�9�e`�*,{�m�?;`�X�u�ň/S�ݸkf�Wcc\F�/#�J�CͰ�\�U�eW�ѹ��wc�9�e`�*, ��x+{�����6Y$���qsj�6~��y`����ǀn�$��wWwI��4�����=��bJ$"(iC^IBU�Q�'c���7{�X�q(BH��]��X���wc�9�e`�*,.�l6cT;T���wc�9�e`�*, ��x?��û�Ӄ�٭������&v㬐u8��kp��m�e�l0p�<Y�a��N��0K� wv< �����V�i]���?�ـr\���$'� I<�lp�;��%WV[O��M:k ;� n�x68`�+ :���Eh���h��I|�T�fl��f��X��$�%HYI$���)��M��N_Q,$�M�So ���_w����5I��ݏ�?����|Ɏ��~���[��l�8��&��.�M��\��J&�-�"����n�6p��^XV� ���lp�1�e�	�-\
��Q�Ͻ�璤�I�vy��9.TXU�[���j�j��� n�x68`�*, ��xU6���[I|'v�͎%ʋ ;� n�xZj�E�v��4�`�*, ��x����\X/R�q���e�ڗR*1�n;��iz��4���+[q��$q�s��u�(�\V���p�;fD�]d�u���� �d���6��6��!Ɇ��n�1�3�X�=��i�s�n��^��Fz7�7a3=s7�Z�*�um%SS��M�M)�b����yT��cW[���a��j�*�۲e��/!ڱF�E�Ŷ�l:�]s�k�5��d�*�'b��f�YfL�!�s����u�\)�mH�� �-9�J����A]v+���b�v"��������ݏ ����E�mm����v�]	m���͎%ʋ �ݗ�r�Z�t�­�"���9�� �Qa��KT��K�X�ғ�t���]6|4ـr\����x��X68`mK�t�.���wt�ջ/ �H� ���r\�������ϑ�g�=V
�ʇS�s�]�Hf�+[պ'\�h�er'gDt����tv�hnjl��voWt���D(�����U�h�m0�i/����9�_MՈ���Cy=�l��I��^�{���q]��M�m�%ʋ �ݗ�n�ŀsc�ݔ�(Һ��'Bi�XV�v�,�0K�����N�Wm�Бcn��ذWg�� ���un��=UY�P���]���mb���N���W�=�����<ֶkitݮ�zN(J��ͤ�m��;<�`�*,�v^�{ �m<ʖ��v�HQ� �/>j��#T��K�X68g��)^�|4�J���T�}�M��;��Y������@>� &���jTM0W����a����<��χ��@a#��o����s��z�QC^����>���20I�$P�d�J�J,n&�:�0db��	&�U D����� �`hK�����}A:��!�A�a$��Y�����Q>3���'�dR$dd#M�F���Oi�'<6���~_���+��w��"H�G`�h"x���tn,�M��|=`��}��Ł�#�jaD����@4����'���`;����E0�q��#��:QػDSG���Xz���P�(�O��QhBPuX��A'>P�D����G�`!�x |Z� ����~�^��=�6��"ꭅ�av5M�J����`��r\��=U�ۓ׀yW��ɴ���k ����E�un���� Կj�0��ے�e�p]�Ε��Q�n�:�'p�9p��k�]�n9.ݮ{���ڻUi���w����:�e����R���٧ �j���݊��N��:�e��.y`�~0K�6�$ًY�EmۑZ,�_ ̹�oc��r��:���9[�Z�WJ�*��)����%ʋ �3rh������Q0#U*�t���=DS���}�k�\ݺ[>v���]6|4ـr\����(]]��7��vl�@^��h� ���g��hr�gɶ{jw[�9�گ/�d5�]n�Fx��W���m�^�����z^ݽ� �c�͹Q`^�F]6
ʶ]*�xv�,�0mʋ �ݗ�H�KG���[I|����͹Q`[����X��TĬISMS�m�6�E�un��;����ɇ�K��Q7��V\r�.(�R���m�*�پ~T�0�{�\���t�ܓ�$�b���/u�fY������C8g��ۮ����:�8��/Y��3�3���˵Rc�RO\�'I�n{�o��P|sm�����H�	�Y/��Ӷu�N�`����H�όX��Y�<-$n8uv�p�eK[�����'c���"�]K��'ggDj�����m!�6�����hJ^.��/a�u��B���m71����T�s��Zj@ ��$M�)"�Ir�J��������Ņ��r���F`N̯SՎ.�mm�6��F��%����]r	\������,��6�E�uwe��֭\�UaVƐ���9��snTXWv^ݽ�?RF˥�|���φ�0��y`]�x*�]�_�,g�����)�l�p*��G�l��m��潤�a��4�}T�욵�}հ� ;�Eh�r���q�R�T�ws� �W�ջ/ 9�U����o���G)��,�W^��T㞗����i�����V�峗"��&�	w�~͚p�y���{��T�ʒ�aݽ�����Pn�݊�jQ$8ݼ��9BH�B� ڇ��zy5~�ٹ����sʩR�UWf{�&��e�)�r⏀c���ݾ����W}�O�~^|����Q[v�V��$���R����� �ܨ���x+u�W,�V���6�͎6�E�y�����v�(J7~E���6&���vOa�D	/7r;Jn�^]հ�L�u٠T�l�Wr�QڻV�(�C�?e���:�e��ذlp����i:V�հ����:�e��ذlp�5w_<ُ���b�H��ݼ۹'=�_M���2�D�G*�@��L�p{�����ܓ���7$���fIq��q�5?ټӀc���|T��5�݋]F\��[�J$� ���/�yyn�|�����fL8��>�m<��	v������s6̀ݘ<��b�D�zx�lOUs�v�����غ�cJ�����5n����׀v^ŀs�0�_0��[|�b�2܊��q�����W������5�~��6�6~]�[��uj���	q�ٳN�d/}��l��w��,v�\��;Nթ
#��j���V� �^k���ٹ8�*�D�
�� �~DU��$��Q���,���7I�r����R���q�T��n��~͚p}ŗ�<�W�F���.�]�7$vFH�!z��g��-�=OZ۫�^Jj�/fPyK���}���-H�p�Z���}��w&qe�I/�w/5�krٮG�Ch�r_ ��0�y%T���^��{��1�2����6n�F�2�݊�jQ$8v�k��}��ު�����|���}܉��ڲ�r�.(�UJ�rf��7o�}ܘp<���IR��<����o��2܊��q��_s/�yz�w}���g��π~�� ��ԕn��x����~~~e��ct�� Ӹ�Y{:�kg]�xTD�<a��5���n��Y�Af�\\�`�:�{��ƥK��1�[v촧m���5��uĩ^s�u��6���d2k��Dn�v�b�5J�o%����t:5�]�X�6�sv���՛j�sh���<L�g-��S�u�lUɵ�8�3ۨ-��%&&�U������xX��f絮֛��]:6�X��@ �&�.���s�Z�V����;W�孋�X..ݞ��i.D[G͡qa��Q\�n�hui�˱\�}��?��/>����U���^���7mz�W-��RG!�?e���/$����>�}��w&�I���4N7��\���e�,V�xy.�?��^\���Z�.+Ar>�K�{7޾����?e���ԟrf��n[56�+t���ۼ�0V����˞X������WI�Ֆ�_=�H���pH������sM��#i�K���/Z����]b���ݕi���o���wob�$�[#~��K���I-�t�cJ��b�4��L�m�mo<��
��j���(h.�����p��U�"> =5����n�o��}���w�.��UWv�,�͊ nE`6\r<��o��o7����$�g\��sm��9��$�km��]���ʶݼIz�Dϻ���m�s��Ͷ�����m�	)w��8�o2-����Nթ
#������;�m�/RK7���[l{����w9��� �??0`��|�Yz�M<��R��+W�t�+�!�4g5��D+�M����q�\�*���T�m�W|�l{�5m���sT�����Z�Y�� ;$R+Ar?�m���s���K�%$o��x����~^w���;��U�z��\��I*N��x�K���I.�Իď���RD(���
"`+�8*?%ߝ���^r�m��d�m�Ɇ:���ڷ�I�m�%�T}�=��z�IMs˜I$�cx���w���������q��sb�؛�� ����m��&{����~��1��3˦m���1�ۓ��d�X�,,�)^���k��U�jܬ m*��n�����}���"�mw�$��oIsfC�I.��韡d�o����z��I?JJt:�*�m�I.wr�}_y���xOIl���6���si]�}ض����;V�(�C�l��q�?�w�}��^JH<�\�m�����6���q�����H��I��Ц}����=玲��{o��ޭ��y�;$9��<D����Gx$-�ļ˦�Yln��M��M��r�m����R�K��m�����o=��cm���5 �nmT�3URK��v�Է	�����S�#��ic6Ų�vãu߾�n���-�Y�� ��Ͽw����8�o����]�m���8�ooƺ���j�jQ$>���ט9�*�%IUU7������}�Um���|f}
"&e�7K�4���IհlOIwfx�m���8��IR]RN��|�gots����܌�Y"�6\��m��*��J��I���m���<}�m��8�~�^�IU\���>���m�/֛�-X�\���w9��6ߩR^�IT�x�Ͷ�w��cm���V�n��ydxP�p��>8���4@5��A�>�@��i�Z���XD�*BJ�%��S�p���&�$�@"�!x��	!"���@�@ 2PѲ��Bx>�a!��" _ЀD<X!a#VNz���D�xM���"#(F+�qi�W�EFB$HA�<Ĉ�@8�0][W�b��^�S���`H���s�`�H��L�@�@���'�Q�Hq �!!l��8	P|�B)G��˃Vl�"�q��<P�*2:DѮy��:T7��D=0��!��a@"F5�,����Č �y�浭kZ�D���  � ޠ�l�E p��r�]�rK]�vv@��˴��u����lvIz�]�v����t"��N��!��=�*�;t�%��3[vW��ue�# lPu�Iǡ�pe�r����Ҧz�qy�<sÃ��
�:VU�m��c�	y�vnVQVYZ޵�_�u�g���a�wM÷Y��I-\���@y����q>x�OOGel��-:�,;s���@� ���	lAq�lp.���:P�=k����d���\:�o^��;����h{�]���e�l	\�φ�5=���td�I̖v�/\�[I�M�n�/���6�M��u�Y.ݺR6�G��Q�j�,�mΔ���؊7���r"�Ŧ91�;Vx�k��d�r�ϋ�N���ovc�M�I����,�kX6��v���j���QH\��e�{)4�̖P"�M���nLPB�٧K9�.�����p�mM�--Ǘ<���-],gm��qe�i0*]��ţ�5�,U�6k�n&�ڛv�v@Cv�*a��MU�h�$�k����5�����8��b�!�[�a�n��(ܫ��Ts�K���&��܎٠�4B�I�Rs3xrPVŰ|�}�ܚ&wC�Z��neۍT�x��>z��M[omVc�J�v״P3��k5��cUd�=��r��e
�B��e����z�;hڢ{
ˍ�I3]֕n
Z���G�& ��h�톕���A����Փ�D��b�"�ۍ�5�9�5�c�uQ;-�(�UtUk�lG��Y]n^�v-6���$6����h�i �4�c����k�t���t�uO`z������V��� �bj$Ժ�h�qZOl���&��r�#�ղ�ݚ6�R�}����i���s2��pv���}6���rK̭Ί��6A�v+����	Dv��)������0u��;:n���J�̻07`�=�N.ݭ�q7m*������g���d/VGeI�Y��kZ�4\>z��v!�lC�<�1 ^����|����P��> �����(�Ã������x*\	G&wi�j\7Ba�7W�2'$R�-:7=ktPN�9�8cC�x�М�@��GPI�t� r��;���O���v���9zi����D�����qSnk�=]m;d��uή�l\����eNpZڴx37`���Б�ا��vD��'n�*_2���x�Z�v�8�l3�rD�4j�*U�:��2��-OY�n��;��7���u�Q� ��q�7p��I��g��jY��2�[��*���SG��q����B�6�����U�E�jԅ�f�����q�����f6���5�D%�,~��1��S���N��j$[R)����a����*��}s����現m�׋9g5$�ݷ��`�V[��m�ĒJO7�$��!�/R�UUI1�{���o7y���Z����,wn�����I'�~��o��6�o۷�c�(J\��M[m���q/\n�q�D�������Y��z�$��s�z�B���K�2Ē��!��K6t���]�Mf��"�u�\Zs��%��̃*��߽�w����@�.-��m�u�f6���j�m����D(�z[yz��q��,��"�Y"�6\��v�}�����D* ��e"��(�`�lO��W�BW8����cm�����~ݾ3>I%3o�.YzZmZprՊ�8�o�o4��������(Jfw��3l}��V�ov,����Nթ
%�_|�ڤ�&���6����>����˜m�U%䔝��W�6�Y~�8�Wn�j%m�,�m���a�ͷ�'=��X�o��b�m��]r[m�po!헓?Þ<�5l�Nd�����ZS�8��L�BF�+�0/_����}��ul9�s�UQ�6��玲��n�,�����'�J#�~������ͷ��둨��ۅ��%[m���W�%���}jm�߻��1���d��*�7��][�ݵn5(r/�����홻m����9�뇎����7�U��x�K���\�Iv7JX�JƝ&	Z����*�Iy);����6�{�I��w����<�U7��pm�]��"�Y"�6MTј�c�sM��!f�y{ͷ�����m�ݾ3l�C�>R��9h%��ku�:�V���K�Yz<�k�ݕ�v����º�&�M�N�R�SSSX�o��b�m��1ZĒ\��z������޷�$�u��MJ%9R��*f�cm��[�DD̷����m���M[m���Y�D%3/d����J�V�I�kIvL��$��%�K�BJf}��,�����r���+}CS@�H����ߒ^�������6���9�m�>�w.�� @"D:��JAE� ��O��7�~��oֶ֯H(��ۅ��.q���������w�yr�m����9m��%�I%�M�XF+M��n�Ӳ���"v[�����F\5*�ӷ]�n:/n�����wt[���M+�bwO�7]�IK��ZĒ\��f6���5�P�d�o��b�m��i?���a�������0��$�IRRF<�\�m�����ͷ���-�RJ��]h�?��+m��I!l��I%��Ř�J�����v�o����z�jI���NZ�\��z����f�_|�}���$�7r�仳� �����]�HQ.��gs��<�%^Iww������nI�}�f䈏��GK{�����v??��C��:�j���x�)mP��	4� ?�O��?I]���c!)ׄ'rs�X�s��n�9vr�ڻd\cy�����-=<dQqu��������GI����y5�1⶞�{@�s�v���̲�����y�F�k��r�\ں�f���ˮ��n.��R�"ꃡ�V� �]���ZL�Н��S@���⑧[V$�Dȅw�*K�Ie*�J���Ƌv;�n��i�Q�O\�l�.��Zm�G$tyZl�-B(��k���?}�.�u`�;a�;��0{#�9����������7}�!E��"�ـ��ٕ�N�E�su�=UM��Z�[.(��ۅ��' ���\v2,=��R]���Oy�i��Q4�ݎZ�9RI�o|�dӀ���ԓ���.ܽOl�e�8D���Ày$��~�z~������`��b��$��:K�J�;$j��hz^�NML���Kڣa�F��[����o�������R��8��<��+ �!�i,�a�ɧ ŗ��F�Zpr��ֵ��9�l���Hp��]�o!��w2i��d�J�/Uٻk�ꌎ�թ
%�\��y��ه����<�{+ �.O��v��T5c|I?ٜӀ���}���K�W��ǟ ��/���H���w�8��V�ܮ��<�n�`�� ��غ�DQ��]]���;v��`�!�p���a�n�}�N�羛���->�=��Id��su��UW���xc�z㻲�-J��fY�|�%IR�%Wgwg� {���w��ͤ����]z��bWI�	�ln���`�=͂�DV DB	���Wg�@О�Y�6nI��jv�I����DR�$V4�IҤ�&�3g ���\?d1�<�z�%U}��� �������b�rp�3��jT���Vπ�ɧ 3���=T��G5�������{*�`����7W/.��J&m��4aq��NDK�(��jԂD�� ����3��p;ܞJ�/�owx��/v�!v�V&�8w�m*I��͜{�����'=I$��Wfe�@R�ԑ4C�����3���f�W������u��'M'hWm����w��;هR�T��%�T6�t'7����<���^�\̆V��պ�	�Q���v<�L\ʫz������Z��bm.�]M&;h�dts�	r��F��OP.ʛ���{�\|�%t�`�4�7�=�?� M��I2�vTxt��C���n�T��� ��'5RM��w���[8{ه=T���I]����wᡖ�#�\�8}��X;*<=_U%$~0�y��R�)jڵ!A..�I7�ճ�fd� &�x$�X!r|��i]X:���x�`�流��������d��
)W�؞~������nEw�M�,u��S6�1ka��؎h�{Q�n��Z�L7���6�B���Y�
muW'e:�NnR����UN:��Xc�5��
(��v*[����z�-����n9muf��
M��;m�8�0Y!,�Tv\�]�lPv�]�Vw�����(�r�Γ�	�X6r�K۩l���Du����slɗk�8L�Om�E\k4�=fY�|�lz�e')�r�)��4\ֳ-�{N��������tu��䴖���H��"�ꤒ��������� �� �+ 'd�靖$�����ם��t�v�v��9$��}I��6M8�����*lצ:��;���(�� {}���p��W���w��XZ��^6�8����N�I�s�p{�8����yR�J����8if�8�M��;�!��ܜiR���� �g��8��7�+clw�3�W����jnK�����ݮ8S�zK���skhn!��J�#Zp��r��}�����7��������<����i�mZ��� 3�a8�T�!#�_�8.ة���I��8��r�X/�y��9��rI�����gs���%I��^�B�vݫ�r�8w&� �ٓ���%�R���}��o�N��⼀�e�"h�C��2���V��U���!���X�5�d��9lww' �;�\j�%I����&�� 'dx���U�wnqs�ݹ�z�8j��#U��絸F�N�l7��[�������o�'ĊpE�Cw�lnn��w�f �ٓԪ��UU/�����wmy;W�ݧ%�F��w�f ����2�l����~�ꪫ�x���2P��;�!�g�8�����^�dd�F@"���JQ�3�M�$��FB @��C�������$��|��!B{��H���!��~פ�D`��E�BP��h>�a��R�CE�/�i���k��xxF}�E�S��a1����H�������͛I�S���l�B�詁�|>���
j�j m`1CjE}6��&�tQ�@�S�f�o�Рi4#���������"A��|�m�^.���`"p����2..���@|� .�im$��;���7f�2���&�i�:e�'R�����pst���0�� ��#%j�U�g��� M�x���3� =���96e`���{���O沌��+�;T�Y{�+Ws&��Q���r�W>�/���k������;I7.��<p?fN�w8�I/RT�X�x�2���Q;-IA$8;#�9$��	� ����UT������NЮ�����l���I/%UUw��� =����uռr��MƥGqp5*T�{����4�I������� � �P6(�ן\�`�ԥuq%t�c�)�lx�p�J�=�l�ۓN g��pRU�����nL~�DO�m�Xb��6͢*��8:�;+<,�m*��7�����u�>#^�n�T��΀~���Mp�	����$�a�ɧ ݬp{L��2�ɀrk� N�<{�;�羯�侀2��F�v��R����8va�RI$ٽ͜��Ӏg�y�-�m��"M˄�yR^I*���� =���95� 'd�ܫ�)ӥe�n���~�N��T�}�x�����;��nI�D�r<\�@C���ߏ����1����\��1WJ��iN���W
��ð�K*�cl�&"�U�s/4Q�k�I�h�8G]�GT+��qi:ɵj0��{c=e:�.�m&`���.��<��k�-��N�۟A��s��F皅2=\&�(��6x،�<�sn�F|�j�r��)�4JW�r%-��Dp�^�$&�k�Y��q1�Ɋ�5p�e�x�����߾Mu8"9o�.BY�3$ٓ5�˗F�
$�k`�x�S�S�'��Z�uŲ�(v�Ѻ�����<��M��hWm������ 'd�� ����������v�_��0vA�H�� ��<�\3�T�ܵ�ڽmږ�"n�8w&� ������Ԫ����x��u�%MՊ��ـ�ɮ; �IS��4�����M2�W�&ɮ���{g��&�� &�x�������{=/�_#�u^:�i���E��nR�:8���-ش�ś����������V� {g��ou� &�����;��`ڹ�n��u`�vǀou�6z����� lt砉�J�}����� ��<��WΝ+.�t�f M��Mp���|��6?Ul��M��hV�x�_^���=���9�фJnǀyB/��ݢ���`����p�	��&Vݱ�diӪi�)��jɔ�yQ��F���]�%�8ȸM)͹Һ�%t�c`4�� �� ���fg����p�nY�J%��m�`ݏ �+ 'v ���ɳv�X=��Zj�b�$��w��y��[���qB�0D/��V
5�A����_��I����j���WM��X;�x�`ݏ��R��V�����vݫ�r�8{ه �J��l�����	݃�9J��Z�����M�HvS�6C:��<�s�N'��S6Б���]���SSm�Ҳ��]l�	��&V g��=UU�T��ݞ84i��@q��hV�x$�Y���� �� �?7c�"�W�;��v��� N���z��ꤏI�w��V�k�x7jG	 ��'iRT�3�p�wﻭ�9��lܟ4a�~_����l,�c��!��R��0n�XB�����X���X�\X��l~a1��.��m�\�C�=^��Э��Gie��4O5��l��k`�}��O������ˤU�� �� ��<w\?}_q��8e�Q��mZ��� 3�p�Ԓ�$�ٹ�� =���>��<��Uv{��d���XD��	�76x�ݏ �ٕ���w�*6�t��.Z�.N��߷}8}���~���J�w���4�� 8�N[�' ���`��}�V۽V(��|�C�A�5 �0CI������~gx+���&��>U���n3�:��N��MX�j5�wdZ��3v\��8p�a��d�h�n1y9ptl���m�.1ϴ���m�۰t�8���)�q�i�l-���v��n�����b�V�K7 ���a^������6�l49|ՠ�7m��9ɳm���@����v*�A!��ㄮ�C4�c;����k��pL��]�nĕN���қ7l��q������ᵷ;-˸����җf��X�uۄ��pԵmd�v)�t�����?nI�v��v����{���ǀqM��j�J}pJ��覕���c����=���:��� g��sj�;���:��CvR�jۼ ��<�l� ��x��J֭*Eҫ"ݷ��I?׹����8_���=T�*^T�]�7ӀfߏA�թ
-�| ��<Wv^ N�x�x��F��߫�������݂����2s��^��	����aP����{�<�o�;]�˄���_ 3�rp�w/ԕUyUW����f_��b�+��Ih�r���~�戴$B
D�
�sۯ���v �ݗ���#U���N���
�uzz�vA������� =�g ǂ��[��ܵur��<��t� �<�wc�8���5T�*Ȓ�m�D(��p����yRO{�>����	���Ij��t}l,������GV����ͮ݁���m�-9n?��o������J�v���y�Se����ǀIZբ�H�Uo�[��)��wc��ǀ�z�6_�0�����w���ݏ�T�X� @Bt�!@a# ���WV�f}�nI��~́���S$M�j�$ܒp6�/*���< �=��Se��ǀw�*6�t��-��Zv� N�x���~�� {g� ov<@"�iU�T$�bOI�a'6�/OF��,Κ��)時�{����7o��lun���
��:�=x;���c�	ݏ ���ZwJ�݅[�| ����*��s}8��N����U)O�$���7E4�x���~�N�^J����� {7Ӏw�u��Wt�%��]�8�$��6p�so��ߵ�4qGJ�F*! X&�E�GBδ�F���X�i�&P���jr��<�_ �^�I+�o������ǀoe%b
H�tƮ�ZN�u�@��uR��Z���˺�3L͵��T�C�vի`t��WM��� ���]�x;2j�U��so�n+�I�c��rI�:�w/���yRUv��p�o�����RT�g{z�T�������/����|�|=UI6n������?4t�BK.(Ӗ�r��=T�����f������*}�ݾ�@�W��-;���ۼ ݑ�����%�Se�I�Ϲ�8I4D+$'ڟ1�>'��8\N��b���,��6���&����R"k�G���6����B�υ���X�OB� �f �������5�@�ڐoO��!����H���	0/�ސ4'�c�
���������ixI�xz�p0�r"Hc�<� V%�6|%�0�FH�niS�Cy0�!G
�&$BR�O()(�"""��rff��()��  d ��� :��֥ ��4�i��$;k��%y�]1��Y9�����X�4��`�7g����� �秺��zJ�Q���c&,8a.x����\�d�$Mgs��٢&�泝��c/]����U�'L���l����\����N�6��cU4 l�󩡤ݮ쇢F��&��M�\n^l͹��ꃖ��LmڑEmu%��Γ���+���,��j�j��n�\��q�nz�)���ϮsJ�����۱���yW�xwa�/&�m!G`�^|Ft
V�/Z�ݪ�Xwc�s p1���YuMc">�,v��ko1q�������7S«8&�X;[qӣ��*�I���;g��v�j8��c�ѝ%��.�G>|G1���Ħ��*2B�mav&;]��;ӒY��!�;��Ln�{+8v���P.��d���;,֍��.�x��B.£�05El���x;cjt��z��ogpK�-m�6�أky�)4����ND�Х���x$٧�8�T��R�s�MB�]٣Y����y��.��p˸�.ͺ�Y��H+'H�VOU6�v�<6�&)�SfJ�9ۆu:8M;Oi��g3'2NW*,q�lgs�q��{[�+n�k�����k#m��hU5��,��9�I9r�$έ,���Q��lU<,�T�s�$q!Z=9�]�ӴN�����L��G�P"w<�ؘ'���Ӧ��Վ[w$3�������)C�� J��U�	�Hm��Νo$��!:��6�{#�N�j�N�����8)Qq���jG����fڮn,m���QU�5����-�i��Y���uH+K�]�t<z;�ٕ�تU��4g�9ל�A,���ɵ������CFUK�ˎò�+:%Y�W\YZ�۩i5��s���l��a�r�5pm��r���>4�3���Hg�웡�[T�A�n
 
^�a[�"�R���Zԙ�Vf�� &��+�OT�N�:�X$@>h*�Ep>�C<��J���~ Gux`��{�\�Z̹gF�n^4Bo\;SrQF�F嵛6�%��h\>\i�WS�!�ta�&�=�m{�	$��r{ad�;PvusŨ�P�G����Jv�M�۷n��6Nãm����v��u����.2a��Q;4�=
.�݈�}U�m]�"9ĆyM�tlШ�j�c7=�����ɛ����u�s��[JR�E
f��R�*��I�b��ٓR�����;\pݨ�-�۱�ۋN�9��9�=�2쬝�︺��?�-;hZ���so�|�|���W���`no� ͷ�����!&�Jշx�x�x����:�w/�T�^T���^�մ/�����w�j��׀ݏ 7��6^ݸF �Yj��>��x����< �<�)��=UIw�� ��{�i�i]X:����5we����M� 7�<�� j'i��t��n��jҝ��w9��X�k�1��EN��"r7B���ayO�N�����n��^�� ���{#�\@M�x�4�cv[��;C�f�rIϽ�[�ȼ��7�j~Uv������~yܾy�^���Ei�+��m��y��c��}T��O^ w�� ⭥*�+�4�`5m�R�����׹��>��>��M���e��v�vR�]��Se�B������}�U�g�����:)���:\GB�bdnVfҬ۵�t�%ɕ������sss'n�Ǜ�e������| �w'S)?�͜KԅT�/�+)2�)m�}|��I��I���ǠN�Sj2f�v��bX�%��w[NC�
�șľ����r%�bX�����ND�,K�u�nӑAlK���3j[��vXD��')|Re&Re'��w[ND�,K���cvQ0D��@S1�(���B:8j&�}�s�iȖ%�b^��u��S)2�)w���J�+��Ij�9K���+���~���"X�%������Kı/��u��K��L�������I��I��h�}	,��N]�5��ӑ,K��>�siȖ%�b߻��iȖ%�b_~���r%�bX�����r%�bX���۳Θ]e��\�v�j��]h�0�-9�n2ک��-���F�=�mmٞT6��w�{��7��{��[ND�,K����ӑ,KĽ�{��"X�%��}��ӑ,K����Vh��!l#�')|Re&R�/���m9ı,K����r%�bX�g�w6��bX�%�{�m9ıK;�ۊ[�i�rNR���L�Ľ�{��"X�%��{�siȖ%�b^���ӑ,Kľ{�u��Kı==���va\�f\ֶ��bY�BD�_w�m9ı,K�����r%�bX��~�bX��Qk��
� �|8��@bҠR H����~�<E�=�����iȖ)��K�ȳ`�n�R\��K�(�,K����r%�bX��~�bX�%�{�m9ı,O3߻�ND�L��^UJ�s�v��k�d���r����m,�;=p�n���q�v����mW �s�b�o�ﾩn"��an䜥���L��O���ND�,K���6��bX�'���ͧ"X�%�{��[ND�,Kﻹ�R���.Z�.NR���L��[{�|NC�Aș��>���r%�bX���ߵ��Kı/���m9ı,���3T�Wi�eܹ|��I��I��{�siȖ%�b^���ӑ,ı/���m9ı,N�{��r%�bR�ށ�Y�-]�`���K�)2��{��[ND�,K����ӑ,K��w�ͧ"X�('���ͧ"X���Mj�4wc��˓��)2��b_=���r%�bX������Kı<�~�m9ı,K����r%�bX�_���"�_��cq�0<9k��m��n9.q����l�72�v�z�lԹ�cn�u���n���5�#q������׵�Q��� Xh��M-���9�ȧI�:�8�lbκ�<ڳɭa\	���f�k�Q�i�,`���5���Xr]��=vܡun��ՙy9�언�ZŸ�HJs�M;����9����nbK�˒�Hԟ��jU�RG����3�l�z�)v����m��vpu��,sj6�	uv�ugn8�Z�{ı,O;��iȖ%�by����r%�bX���u��"dK�>��r��&Re&Rő�[c^-��O&k[ND�,K����Ӑ�1șĿ�~���"X�%�}�����Kı;���ND�
�"dK����@F�ں����_�I��I�����bX�%�߻��"X�b؝�{��D'���mI�>���&�L	s4��H�b_=���r%�bX��{ͧ"X�%�|���iȖ%�b^���)|Re&Re,�8^�QK��Ijܹ��"X�%�����r%�bX!|���iȖ%�b^���ӑ,Kľ{��R���L��[���`6]�+�.A+��:��kS��4t[jqբv�9�X:��[7�lK�E�4�j��_�I��I��l�r%�bX���u��Kı/���l? �|��,K����ӑ,K�z����j��9')|Re&Re����r*�~x�� �m�Ȗ%���bX�'s��m9ı,K�~��!�2%�O�ߌ��]�!l#�')|Re&Re'��NR�Kı;��siȖ%�b_{��iȖ%�b^���ӑ,K���^�2�E��$L�rr��&Rg�IYK����r%�bX��߿kiȖ%�b^���iȖ%�b_��u��Kı==���v5e�%�m�/��)2�)2���ͧ"X�%�^���iȖ%�b_��u��Kı;�����Kı;�ݻg��Y��������\4����YzF�M����:p�D�\���Ϩ<��q<�bX�%������Kı/�w��r%�bX�����'"X�%�}���_�I��I�SͨD7,��7zֶ��bX�%���[NC��r&D�?g��ͧ"X�%�~������bX�%�~����"X�~�韴I��������)2�)2�����/��,K���[ND���K	UcS�(�LX�Dm"�G�/�<>��K���[ND�,K��9K�)2�)e�{N(���ܚͧ"X� %���bX�%�~�bX�%���[ND�,�"�=��R���L��^����-]�rY��m9ı,O��w6��bX�*���m9ı,O��w6��bX�R}���_�I��K��hY�M�(r�U-��N\���Q��e��"T/]`�k���ݻOny��T"�M�g�w�{��,K���bX�'�߻�ND�,K���[A9ı,O��w6��JL��]��n��i��.\���Jı,O��w6���@#�2%�~������bX�'s�fӑ,K��>�siȟ�`*dL�b|}����ɔֲ�mֳiȖ%�b_�~���"X�%��w��ӑ,K��>�siȖ%�b}�����Kı>ý0�.��:�,ֶ̺��bX�'�߻�ND�,K���ͧ"X�%��w��ӑ,K��HG*a��%_�D���5��Kı=���]�,"Ww%��&Re&R����/�X�%��=���ͧ�,KĿ~��[ND�,K���ͧ"X�%��ݿy6����v|�jx[��Nt�q/fk�*q=��$n�+�r0/SGUƺ]�S�.k6��bX�'�߻�ND�,K���[ND�,K���ͨr%�bYK/7o��)2�)2��0ǱD⎜,��k[ND�,K���[ND�,K���ͧ"X�%��}��ӑ,KĿw��iȟ�.DȖ'�>�����50˖�s5��"X�%����ٴ�Kı/�w��r%��"w?w�m9ı,K��ߵ��Kı)��:[�G[�r�K�)1S)<���\�bX�'�߻�ND�,K���[ND�,�̉�~���r%�bX����n剴�i�.NR���L��>����r%�bX~#�~��[O"X�%����ٴ�Kı/�w��r%�bX��@ �$��J����1R�Z�#�TRMJ��/_��aw#N�m�q:*�k)ٴש��L�&{qڌ��n�,���)�oVyN�Ѹӫ����kǷ�G����Q�����[L�=kNg��9͒�8�=7��c<v�h�H��R��g��:�'j�8{���:4ݱ]�� ��ng9�.%Q랻K:㷧 =��ʑ]p�$�� �]�X��.��[rHlx�m9��{�C���ф�yL��L֬.I�����'b[q����˩���ԽL�0�[1���%�[-�-�m�}��&Re&R~���/�X�%�{�{��"X�%�~�����Kı;�}��r%�bX�aޘv�V�jf]k[ND�,K���[NC��r&D�/{�����bX�'��fӑ,Kľ���ӑ,K��Y���&䓔�)2�)2����iȖ%�bw>����Kı/��u��Kı/}�u��Kı=��kdL�]��KV���_�I��Ko>�m9ı,K�{�m9ı,K�{�m9ı,K���bX�'�cآqGN���_�I��I�w��r%�bX�����r%�bX���m9ı,N��w6��bX�'�4o÷;~�/D�R�[�U�Cn��/#єV���Sp�{u�a8�Ύ͞D5���ӑ,KĽ���ӑ,KĿ}��iȖ%�bw>����<��,K)<��9K�)2�)5�Vx���.ɫu�m9ı,K���èb�N��e>C�4���<C~>��KY���ND�,K���[ND�,K���[ND�eL�b}�~��nk!iu�R�f�Z�r%�bX����fӑ,Kľ���ӑ,KĽ���ӑ,KĿ}��iȖ%�b|{�Ӻ�S&SZ�e�5�ND�,K���[ND�,K���[ND�,K��{��"X��fD�����ND�,K�~�a��j�#Lv�R���L��Osvr�D�,K�Ǻ��ٴ�%�bX���߮ӑ,K��;��ӑ,K�y$�x捍�~�!�%��Wpl�mW!���\��ŹZd�ͬCΪ݇�q��ɒh-ֵ�'�,K��w���r%�bX�g{��r%�bX��{��~y"X�%��ߵ��Kı?}�w�����K�nI�_�I��K/wo���"X���߳iȖ%�b^���[ND�,K����ӑ,K��	���F��U���ֳiȖ%�by��siȖ%�b_���iȖ4_S�=@���U6��&X�P���1����"Ā$d�Q�D���;��ސ��5B%Ŕ44m)#�X"A�V,"F	P�XG7�E�&u��NP��o��B�iN� �,Q��:<0"IJC0=>��#It~F%(�`��KIT�HPRX����d�>!����W��<B�����jk),������H� sy�e�X��"�%d"@�V4R6V1`H�e`�ְ%�������a�(]��.h�M�N9�xE&9� �`"z��E"P��AL~@�TA<Z��?���><"��Q_��	��'��AУ�l M��%޻涜�bX�'���6��bX�'�1�5��jݶ�_)|Re&xJ�����[ND�,K���kiȖ%�b}��siȖ%�b{��siȖ%�e&�w+c��G[ܓ��)2�)1/�w��r%�bX~Q#�~��6�D�,K����m9ı,K�{�m9�2�)=Z!��6�.�\c�M�NE�Sv궣ꦍ�bykl�����q�dťֵ
Y��kiȖ%�b}��siȖ%�b{��siȖ%�b_���iȦRe&Ry����)2�)2�.�n��2e5��ffj�9ı,Os��m9��r&D�/~���"X�%�{�ߵ��Kı>�۴�Kı>��cN6��4�nK�/�L��L��w��r%�bX���m9ı,K����r%�bX��{��r%�bX�饛Wr�n�nI9K�)2�)<��m9ı,N�{��r%�bX��{��r%�`@�HE@�P���Uł'��O4��y�߾9K�)2�)wcY�����Ium浴�Kı;��siȖ%�b{��siȖ%�bw��fӑ,KĿ}��iȖ%�b~Oߤ��r��-�K���ؚa�^-��S�;�htN��R�k-��@��R#�"��8Zv䜥���L���?~��ND�,K���6��bX�%���[ND�,K���6��bX�R��3�Z.��cwrr��&RbX��wٴ�Vı,K���bX�'s��m9ı,K�{�m9�VRe&��kĻp��.��I�X�%�~�ӑ,K��w�ͧ"X�X�%���bX�'{��m9��I���vX�X�NH&�r��/�,K?$��_�~ͧ"X�%�~������bX�'{��m9İ?U��wޜ��I��I��ƜW�F5e�$.\�fӑ,Kľ���ӑ,K��~���i�Kı/{�����bX�'s��m9ı,J��#��(#>hP�	"�I�iC]���~ݏ��7!�m����&�v�(t8�j���!�JS���;v�`��Ͱd�Ϩ�%Cml�mF6���n��%3�
:��ƽ\gn�r�u�5nM�v��p���UG,jq��/kn2j���\�ކ���!Q%���i�� [1Evw.nB;qv��	c�-W�]"mn���E����ɺ�\�P���K5�W6�1�7w���~�� �/���%���Z��,�D����;�j�q4�"��3m�6E�3�ߞ����'8D�q���;r_)iI��I������r%�bX���m9ı,N�{��~Ry"X�'�����r%�b2����Uܻ�-D�$9K�)2��~���ӑ,K��w�ͧ"X�%��w�ͧ"X�%���}�ND�
�UI$��e&R�F�҈���IumܛND�,K�~��6��bX�'���6��c�Aa�2'�߷�m9ı,��}��_�I��K��1�Q8��3.��ND�,@��;��ӑ,K��{�ͧ"X�%�~���ӑ,K��w�ͧ"X�%��tߣ���L2�\�fӑ,K��{�ͧ"X�%�����[ND�,K���6��bX�'���6��bX�'{�.�ٙ�)e��v:vqiڎ���6)ӝ�m͸�=����y��t<E�N�M��7�ı/�w��r%�bX������Kı=�������"dK�������I��I��g�,w,M�r
�.^���Kı;��si�oЈ�����`.�J��\4� )�+����<�siȖ%�bw��iȖ%�b_��u��Kı>��lΒ1�-�����/�L��L������bX�'{��m9�Ŀ}��iȖ%�bw;��ӑ,K��;�țN6��4�nK�/�L��$%e/{�?M�"X�%�{�ߵ��Kı;��siȖ%�؞�{��r%�bX��m]˱���H�C��)2�)2�ϻ�m9ı,?k��ٴ�%�bX�g�߳iȖ%�bw��fӑ,K�w����n�~靥�h��D�ˎ.��(���u��V1�ܺ�:���x\]�2u^�C�mk�5��"X�%���{�ND�,K���ͧ"X�%���}�ND�,FR}���_�I��K��1�Q8��&�Zͧ"X�%��}��ӑ,K��{�ͧ"X�%�}���ӑ,K��w�ͧ ؖ%���/���Y0˖�s5�ND�,K���6��bX�%���[ND�߄#�@��b ���������Kı;��|��I��I����Z(�8�	,	���r%�`ؗ߻�m9ı,N�{��r%�bX����m9İ?
�e/{�x�/�L��L��=�c��mK֡���k[ND�,K���6��bX��c����m<�bX�'�߷�m9ı,K���bX�'�@;������r�m��:-�l��KF�Wjk�.8u�)<)d1����knl��F9�Ջ�3Y�{ı,N����6��bX�'{��m9ı,K���bX�'s��m9ı,N�zwD�մ�MR˗Zͧ"X�%���}�ND�,K��{��"X�%���{�ND�,K���ͧ"*dK��G�����.Y��kZ��r%�bX������"X�%���{�ND�,K���ͧ"X�)��w�r��&Re&R�Ƴb��\��9.k[ND�,K���6��bX�'��{�ND�,K���6��bX_�Ĥ��q/�]���H
ke�p�!�S�*x��Nzr��&Re&R�G�{N(���eֳiȖ%�b{�{ͧ"X�%���}�ND�,K��{��"X�%���{�ND�,K�����32�1���8�3�vY��uny��ê�g=��4� �	�u3�7�\p�n�r}K�I��I��~���iȖ%�b_~�u��Kı;��sa�H�"X�'����ND�,S)5嚼)v8�	,\9K�)1,O��{v��bX�'s��m9ı,O{��iȖ%�bw��fӑ ���$O�?~����B\���A?_߿fĐIϾ�I�$��'��xm9ı,O��{v��bX�'�N���֬�L���3Y��Kı=�{ͧ"X�%��{�ND�,K��ݧ"X�%�~���iȖ%�b}��N�Me��MR�5��r%�bX�w���Kı>�]��r%�bX���bX�'��y��Kı8�wU&�����vK�[dAl��VWb�ⷭ�n���vӝ���&"�lv�͌>��$Qɷnu�c����筮���7Z6�v�.�X5h.��&]���n����a�S�[�۞m���v3)�Y�f7[)�ϱ���6Ƭ�����<(��`(;fչ!Y��[*B�2��)m��Y8 (��۞�)�&�l哧�2�gl�R;\��Uq�3�q�{����{��_��`���y��(�0�ں�#��������틣dkj�+ϕ���nm.[0�MkG��Kı;�۴�Kı/�}�m9ı,K�{�m9ı,O;���r%�bX���}�kS2K�j�fj�9ı,K��w[ND�,K���[ND�,K���6��bX�'�k��ND���"dK�'����'t�iےr��&Re&Ry�zr��%�by���ӑ, C"dN�_�]�"X�%�{���ӑ,K��/���Y0˖�s5��"X�~A��=����ӑ,K��u���r%�bX���bX�%���bX��֮��Gl��"�mȹK�)2���ݧ"X�%�~���iȖ%�b_{��iȖ%�by���ӑ,K7�����}�'��P�6瞬f]M6&��j�GS��:�.�j�*�z��w�f>3tCY�C����r%�bX���bX�%���bX�'��xm9��I��&��/�L��L��4��e2e5�Y���ӑ,Kľ���Ӑ��4���Ñ2%����ND�,K�u�ݧ"X�%�~���iȖRe&R��W�Զ5p�2��9K�ı<�{�iȖ%�b}��۴�K�ș�����"X�%�~������bX�'s��a���̳$ִm9ılO��{v��bX�%�ﻭ�"X�%�}�{��"X�%��{�N�I��I�[[��B���]��_D�,K����ӑ,K��@3�߿ki�Kı=����"X�%����nӑ,K��߿_�)��̤�d�B]�l��a�k%�Q���p�Qtj�*q���k%u����)O���oq���������r%�bX�w���Kı=�]��r%�bX�g�w6��bX�+�D�
�4喭�cwrr��&Re&'��xm9,K���w�iȖ%�b}�}��r%�bX�߻�m9ıI�]Ťn�e�ⰶ�\��I��E����nӑ,K��>����K?z~b�!���AO��]�(�(�� <A�x�5!!�Ut,A���@��O"^�kiȖ%�b{�p�r%�bX�߉ܽ5��R��%�|��I���HJ�[7}|ND�,K��ߵ��Kı<�{�iȖ%�b{��۴�Kı=>���V[R	ۻ��_�I��I�7fӑ,K�<�{�iȖ%�b{��۴�Kı>Ͼ�m9ı,O�;���5Y�ynlnX�q��g��7l�o%�i��w`�HB.��`z����c���Rֶ��bX�'��xm9ı,O~�{v��bX�'���͢��bX�%�n�R���L��[z�ڸ�ݻe�H�Ѵ�Kı=�]��r�#�2%���fӑ,KĿw��m9ı,O;���r'�*dK��Y���jfIu����r%�bX����m9ı,K���`"X�'��xm9ı,O~�{v��bX�'�Ogoth�Ԭ��2�Y��Kı/�w��r%�bX�����Kı=�]��r%�`E8k�8"U�
xmN*�M~���m9ı,O�h�a�ճY)�-��k[ND�,K���6��bX�'�k��ND�,K���ͧ"X�%�}���ӑ,K���Kl��&ߦիc/c6��٩g4��`�ӞD�^���h�E�ݧ��n���nv�]���ı,O~�{v��bX�%��w[ND�,K��{��'"X�%��{���I��I��p6�a�K�V��r�9ı,K߾�bX�%���[ND�,K��xm9ı,O~�{v����bX�v}���SE2e5�Y���ӑ,Kľ���iȖ%�bw���"X��Dȟw_�]�"X�%�~��9K�)2�)m��`��� �ֶ̺��bX�'{���r%�bX�����9ı,K����r%�`~T`��3�����"X�%��?����f\�ֳFӑ,K���w�iȖ%�b^���ӑ,Kľ���iȖ%�bw���"X�%���|`F#	&Җ,4J��h�D�p�@�42����jjPC� E��!���~(+��$!$���D�+ � ��U>�1-��CN�	>e��E���Wn���>T"���S�6�R�?)A�# �U<�p�i	�k9���B���	�穵By����2PH���L���� B V1b��A�&�HA�!F0$IaA��Bi���I�!G
�N(��V�����.*\XF@��v�<��H��!'�bD&��}4ht�z��8&aH8x�`�H0ci���o� rE�%   �6�	��� &�j(@��l��s�Z˲($g=��[�1vY����r��X�eQ����-���9��:�=n.K��2�]N�m@�Λ�}uC��6�;��ѷ\OS�]�$|�J���Ai'�ϧ� ���j��֌�h��5��Y�I�!���.��J�T�m�sƛ�`W��d,[��F�y��8�m�et��2�N�\��!q�狂�\��Ξ�K��;^��vylk�a];�sٸ}IϞ�;�e<���;c]92�e�&�N��� �K���˪焈}U�۝C{uv���=
�)@��՘^�"�j�eڗ6�脧DC��r��v���tr�ʡ'j�V_!�9uh�PWL�vG.��"x�t�f����ݒ��a�cmgv�ڐ^�m\�"�om��v�0�4Î��{rl���U�x��ζ	#m�(��3�W"mӧ@��ܡ�u%$-�6��N�5����ѱ]��*ݬ�g���/k�v�@X�Ƕ�[���Һ65��ËAs�q�ᴽ���˹��b�q���P��B�:�n�N`�W�����h����S��l�ρ����ZVn���a��]=sWD��K��s�����jRP3������A�1[v��94�ɦ<]�s�T�ۍu���;��6�s�\Z)�2nP[���X�C�l�����5�R�r6�p���]tTf����^�w]0�pۀlVΚy�vV���n�[MD�����61: ��55@nS�n����:��%Km�d�5�5KI4�
Цf��eS.z�*uᐝ��5���ѯaࠓU`9����*�:%��55m�	�Yk*����H��r�5J����s��V-ؤ۵��9J(�p5WP�+�8j��\vv��A�un�m�a ��a�p02�#ȝ��u-V��,��g���W�&�l�l��j�V�v���r�n�@��VZ�-��ǽ��w����C��<@	�'�F�z��|3�@8 �P� E��`��!�
-T Ћ��x!�`�<D��ZK�U]�S��~�˒K�4[n�\����볥�y\�m�6�v�ݭ�6�"ʻ�3�^ݶ�3:ۧ�'�q���)�[uq�,+��Ō��7:*�.��cV�Y��lH�m�l�B=�,��|&�5m�Z`�i���&vdmݭ�֠xЄ�S�%v�Әph�q�6�Dd�9��v�Ϭ��X�<`'��-���q	�jۮ�&Y}�tON%��7/�HhK�4���ww��n�V���e��rrn[�y[��9ݫ�%�Z�W���ժm���|<��b�\�
B��R�=����L��O>�u��Kı/�w��r%�bX��{�a��L�bX�w_�]�"X���Yh�_���:!iےr��&RbX�߻�m9ı,N����Kı=�]��r%�bX���u��E�I��dM`�cd��v��ܜ��I�X�'{���r%�bX�����9ı,K����r%�bX�߻�m9�2�)5���r��e�*�I)|Re~`dO��߮ӑ,KĿ�~���"X�%�}���ӑ,K,N�����L��O�w��إ�+NK���,KĽ�{��"X�%�����[O"X�%�����6��bX�'�k�ݧ"X�%��3��Y��,��ji��I��;���W������S/G�h^&6[#7j��{�\���ae� �wrr��)2�)>���m9ı,N����Kı=�_v�?O"dKĿ�~���"X�#)z׷тr�j�eےr��&Re'{���r >�J��~8� ��"y����nӑ,Kľ���ӑ,Kľ}��iȥ�bX��Fm�r�v�Q"K���)2�)2�r}۴�Kı/{��iȖ%�b_>�u��Kı;���ӑ,KĽ�f�hR`��#�/�L��L��{�m9ı,K�~�bX�'{���r%�b�'���ݧ"X�%��#{NA�Nܓ��)2�)2���w[ND�,K�G��߼6�D�,K�k��ӑ,KĽ�{��"X�%�������7��ݿ�T�9K<��R�n�c�=c�b�2�ˊ��Sq�v�;o��O����,jݶ6䜥���L��^����/�X�%�����iȖ%�b^������&D�,K����ӑ,Kħ�5xr��V9V�nE�_�I��K;3�iȖ%�b^���ӑ,Kľw��iȖ%�bw���"�%�b_����i���%��K�)2�)=�{��"X�%�|���ӑ,|`��qJ��
�6�.D�'{��6��bX�'�k�ݧ"X�%��nr��ae� �wrr��&Rg������m9ı,O߿~��Kı>�_v�9İĽ�{��"R�)2�����9v5p�2�I9K╉bX��{�iȖ%�b}���r%�bX���u��Kı/����r5�鄱�Ӷ�Ӱ�5�.՗j(ǠH���-��S!l�C�U�O_���=��޺\�t��� �s� $��&���� ��������˰�J������UJ�&�}ݾ����=ݙ��RM�!��[�]+M�-�� �L\<����k�����i���6K�j�ڷx�e`vK�	$x��}\�D�}4�����nI�:_���wv'��I7X]��I�I2�aI#n4���A��.�ہ�Ⱦ2� �n������f]Q�£#nV�9�[-]!�e]+Wn�I�L�-�I/�k���[����mH&]ܜ{��*I�ww��k���32siyU*�:׷тr�j�b�����qp?fNIRl�ݜ^f� ǔl����h�uCv� ��^��}�_j��*�{����3}HۻuV���"�^�I2��>��?�� ��D���8{�}�w�����q�a�� ��"�9ځ�s�x緷$v�N��C�y��g�x۳[�� {:$ȅ�ٻh+A�i�����Ķ�]�Xҹ�OG��g�ֵ�&���ţXi3�>��0s�L:%4c�8+'Z���z�ms��5rWo=�BW5l�c����i�Za�L6�^ї`�K�Л.�3�C:ݑ���}�����c�ɵ�b;le���l{M��g^��g�����#��Ih��u�R	��vI��f�h\�yfz����iݗ��W�C�S���O�﯀ffqp�/��%�{�|6�ZU��;Z����x�e`vK�"�^ vly�H�R��2�����i&� �}��"�^��H�O<��������t�*�Z�w�H��G�338�T�����r]�q�[�"�wm��G�~�{��p}<�I��mU$��Ú�e�l�����vܮ'���T8���/.���"�u�͑q��5v�H�7vڸF�v�O�������N ffM�%����� �������-DMk4nI<�ߵ� /���$R����
����*������uXI��Dle����P���E$����|=^T���{���zpΎ�N7I�|���n���x�e`6G�E$�v�T*�Hv*�i���$�+ ��K��|����[��	"�/��e�a{1�Ol���ͧN��6sbz-��Y,W�x�ŅL^z�`6G�E�^ջ/ �&V J�R��n�h��x[%群�Rz�O{+ 9�<jk�Q:�Z��9njl=ޛ��Ֆ��P�E(�� _�!0�  ��P�t.�	5*-K�gٕ`�uX~;��n�p�2Ir�Osw��ٻ0l� �ݗ�v�w~��tZ.�Pݺ�l� &����x�e`��_����,�̈L;b����<�;X�V1��Jj�y��$�~�#}��Q��5P���{�xV�I2��#�5|i��t��]+v�ջ/%z���ؠ�ݜ �{s�*l��i�y%��ZE%n������#�	$xW{��>k,ݱʵ�\IR�J��N {����{����T�IT��#@�<7��������jL�n�h��x$� �ݗ�M�+ >�d����,��
�h��;�3��&M��q�A��c�M���'�,�y���F+��,㈗jݑ���N����������̟ʕ%�svp�����n��Rv� �&V sdx6G�un��&�ԅ[��$��T7n��#�5I/ �ݗ�l�+ 9���6�]���;o�_���5I��6I�����ҍ�l_5+n���x�2��#�5I/ ���N���̇3�sB�v4[s��2W�ơ9x�nơd2�]5o6W�<��J�m�mu���e��۰��_b��Y�H�c�;zٍ�p�nң�mc�6跞qr��rƶ�ƞ�m���`I��5nSM�B���b��&��#���u�+K���C6�i����W��j����q��.k&gO'���pu��us��Y+[v��n.�t�����珴�����l�kn���s�zK�O�j+���kp�E(;-��#�����K�����m�?w8��;��u�e����`n{Ӏu�Ok��	�t�M� vlx�%��̜����U6ժ�ڎ�$��9/�c���fNJ����� ���������ի)%v� 7�<d�X�͗�5I/ �V��di�n����.��J���_����^ odx{�]/��+��M5m&��q�	&|r@7O�K�]l]p�Uʡ7=��mu���݉N�n�`�˗�j�^ odx�2������"�-�I;w�=�}�o\Ch�B"<��)�Ph T�D�LX��_}C�\UU��%�����w��}�����IRF��J^n�b���[w�}�l������� ǻ��2�Zx^Ivݶ���'kʩU^����r�~�י�`��1�OW�3,u��T��˗�j�^ odx�2��U]�,o����v���7	2tS�:뇦)������v]V�py�(OWb����w����5T�T;Wn���߯ 7�<d�X;r��SS�'M]�V4RJ�� odx�2�v���5I/=U�URF���	
�Ulj�v��{���9ۗ/6��*�D�O�4���������#0�k�|X0��5�NR,!9JFD��%���� ����bb�����1�� ��#*^��`1�c�� BD��8��>���^D�by�+��iY�n��D�����6\ӂ�*	!āF���wx�������4��B;�᠉���I��V1�#"!���> �z� �\1X
�Z���p�>E"D�N��U(�����ӵQqd���<�GV6]���T7n�v���5I/ 7�<}�}Jn�ˀ5f�$��ar�r���̼ ����e`�˗�~�'���o���.�y�y����&icn��`�Ѣ�e�ڷ\�x��ǡ����o���g �fqp�_o/UR���_������_��n�We��I�;��\�l�����{޼ ���*�[PTիB]4�u�s��/ �$�?Wԑ��<{������;L�([D�w/�������ݜ������UP����������5��y�'�����;�ݑ��w/�fd�J�%�[�~�t^��x���JةU�;Wv��_��7B�ڞk^�X�)��y��ͳD.�o �m�E�!ZJ��R,�o�OOe`]ۏ �6^ sdx�QՖ�h�$����o'?�*Wf�o����8s���UR���Y�	,e�\�9q�zz��G����䧧��ғ׀u|i��Ҷ/���ۼ�%$��'���R�^�l�~����wiZUvX�m�6e`�W=��zz����I�R%=_Q��A�+�t,��Gw{�?;��Qүl���[�eE���9��!\O/k�S�V�ܦ�b�\r�z�D[u �<������W)��W-�ö։^�����N�cH����&�jU�m۱�b�p��TO�2����2y7Ӥpݵ̽
�cb�<�ʴ���e�i��հ��]v�f�6���:��lO���Ҕ���^��\ͯ�n�S�zNs,�qL�����$��?|6�����Q�V��:ڈ�F{:[n�sȕ������n-.�=��1SV�	ՃI7P����Se�wc�}���Xݡ����e�n�Se�wc�6l��9Kd�jjN�t��%cE$����ǀlٕ��.Ҟ��zz���������"���}_)��V�S޼T�x�ޫ�}JI�%�%RETҰ1=��Se�wc�7�e`J.�^����n�+�r>&��]����=�6��Vw/Y�U����7{���	������2�U��A�S޼/��D���������ΥIr�AI%k�T���ќ�� ��n� ���|��KK��wm*�,I���X)l��ʩ%M�o5���8溟VGn�Ⰼr.Ҥ��}S}����> wv<{&V s�#n�؆�2���xe�X����X)l�������ڶ�k��f��1�In�̜��je�v��:�E�Pe���:��?7"�:2nf���}V��Ձ��t�(�Kj���ہ�I
�Ulj�wv��g5R�I��y�|�� ?w�9�U$�Wg^�?Ee�-�...��޾������a�$�W�b���*��(X�!DFa�}u`w}֬N[�	,e�\T9/��T�̛�����;$��9Kd���Cj7Jؾj�v���ǀ~��r�Q=�wnE��N���qӛ��g���\��t%U�9�$8Ȓ�F f�۴�N,����X�m��2�#dx��X���*�-�*jա:�cM��<�T�$ٹy�����3�L9�I&�}�#�N�Co��av��s� ;�;0#dx����ut��*l@����K�w���}�� ��̜�ԅ�>@	�
��&�P7DZ)TĠ@��}��7$��h�wm��i�wrp��8����>v� wv<t��P�j�]Z�@��6�^GUv:MM��9��l-2�<�[�o����X��vZ�[����Oy�^ŀݏ �\0I[:E�[���x��`fǀI���	Q�V��WL�� vlx���䪩z�_�8�{��1~��^I$�ҫ�ěo �\0-R<Kذ=T�}���?vО��n�r�"Hp�^d�������3���3;0���4r�"���;��k0��R��5�.8��������ٛ���÷�.M� k�5���c�O6pe�ѱ�Qۦ�L6!�%-����lp�fMX�p�<h����m�4���n�5nwg���wk�!;vQ�yւ<F�\�Gv���9�rⶎ��Y��M��˵R�ct[ѧ�[;'IR�GP7��Ȩ�+r;KJ����`�u�]�v��K7&t�����Z���.��u��{�������ͻ=����{��,tW�4�Ƕ+3�e�L۫��v�Z%�nIN"�O�{��| ����3;0�*J���=��1w�n+M�ڐ`����ܜڪU_�]����_�8e� ���dN���i�wq�k�ŪG�I{ vlx[)GV[�J�[M��%�X�;�����sN a�6�L����x�p�͏ ����Q�������9E�"v�U��dc���t@9-%��t�L��;����lzm6`fǀM��T��A���z����v�UvX�m�u�6��*!E�I;%����� �oU�BP�g�'�F�۵n&�$� ����;0��F�y����'v�D�L��t��m�~�^�<�}<�	�p�ڪ�����W��v�R-��ٱ���qj����`�������v?��	ݗ�i���Ky5ɭ�^]մ�"�[6E�3���x~�o���iwv�@�<��;{� 7e�5v�J�;�+E���l�9�Z��� �����꤂Q�eG.˔����7����s'j�WCZ��A�R*����s��/ ����+i��m����`w���3ӳ�a�	(���%>�o� ��=/�I.���N��0�?W�]�/��=�<��#�7�]O�y{E��ts\:��v=�ɦٺs��sh�n�p����\v.�]c����;{r�	�ذ�#�'u� ��"2Ӆ�$�#�/�g��>z���6���=���9�ۗ����"VƋ���E�Z�@%m`g��	�p�9�ۗ�E�/ �ڍP+�)1�E��x��*I�w�pݼ������z�N� B
E�C��C���kzܓ��=�cwuj�[M�V�K�"ݗ��;0��1�5n������a�=���&:oc�X�l䱜��<	����l���v[�J��n��l� ��0�U�J��{���<��^�;��ӻn��#�'c�ջR��e�JK���We�6�;0ϽY|5*I&��m��n���ʂ��]Zt���0�ڗ�E�/ 9�<v8`��:%�v&���e�w�E�/ 9�<v8`[�/ ���ߺhŔJɵ8�!�X�CL`&��h�Dd�!Eլ���&�K�Q5�� ��Lxx��H	C B%���u��<A|��61�Ey>��@�q@�ͨ�H��"20"ʠa� ���ϊ�oB�"�H0#�H��0�#��͡���)yƞ��Ϙl��P�_4|*V..8�$X�JJLCVlX�T�;��l�V$`��T�X��+$�f���|�W���B��9��&�b�)"�B����F&��QF ���f�`�y[�J�!0pwd*���A`t��t��w��v���z�@  d ��� I��m�@ͫ��$��O<l.�k�ꥎ�RX��L�&��o���`d�����8�ul�c����+�n^�v(�l9
Iz6�B�)�sNms:KRe�n��I��M+�\��5_�}�Ѫ�mU@����ݜD4�^�
�Tbtl���u�-�ĵUJ���e����*��v�tX���+l�m��39����n&��N�s�A���W=���=�HeeR烛����S���9�o�&��ˠ^�n���unZ@�xƹ�N��fuN�x�3�bu��j��%�Z�Z2m��ŞtsD�K�.2��ɒk$��'6�w��uĭ�َ�2 ���\��]�:y�,��nغ5�ݖvۚ61�U�kq��{�wq�rr�n�'�����7uQ��}��F�v����<��6^�l���w][l&�B�P˖���]l%b�9*��5ppkvspAE���^5�ƭ�CP*�ᮋ�靻��BV��J�� �p�c�65����c�l��� �U��ɩ�(�cr���jmv�{u�6���MV8�Z	˃V��.��=������`���t� {$���)�� ��V�WL���x����A��-�su8����P�P �N�`o&4Sf�`�t���7o��]�ү�/�܃��a�.�W^ӊL�������Ԁ	­V�r�X�����j�7���c�0U���;Q�Z�	�qdf����J8@@V�JD�d�[�öoR6)�Z���}��s�۬T�s��$�Ur�V���j�a��in�ຸ�$yt=�fsj�Ct���[��]��%�U�̼9X ^���Fm�\�O���� �gtJ��5��)Ċ�UWR�YI$2�u��;��4���=�V�)R���r㰣��꧕�Ў��E��*��G-s��hr&c�`j�m��4F�pn��A���f��u�e���c���Tk���h�eRPhٙ�5�PxE}F�Bm�`|��b. mQ�t�׃�z��i@�*�y�W��{��?��݋�J����Ϥ�nށq��������6&�\&-��pp��+��L�۞�m̀���s�t-��:�eop����냐���AP��-�t�;�8�Ļdtr��졚�[W6��/0S��T���3��k�fYǪ-M�ѱ$�j��榸w<1�6*V���]e�S�9"��4Mm�2�=<�
�rt�c�u����/Ll����{�����3�-.'q7d�ѢEw��M��â��q�O+�J�i`
�������}��
��T:@]�����N��v��n��:��gµE&5H��o ��V�K�"ݗ��+���}_W�f<F�Y%ڷv\
��8��Ӏc�r�yR���7g ��ӀF.�Kv[��7�E�/ 9�<v8`~I*o��g ֵ�V��أ�.� sdx�p���x[��u%�|�����F��l���R�x6�e��9�n�he���<r��U6yw&��	��ݨ��e�6G�n��`Իv���D����d���J�Pxa%�+�40�S��,��޾ o�g ��0�I�{�ۅݪm��v��O^ sdx�p�n��V�{�)b�R�LA3Sa�BK�W}�zpg�� ~�VN����f����UB�E&5H��o ���ڏ �v^ rH�	 �|��]X;�Э�n4�5'�l��$�:N�z3����E�a��W%\��vˁW� ?w�' �����ٗ�/U~��zx�-g�Ic.ˉv���ܾy*T��wo�ovi��Փ�T�5�hձD�6(�K�/�c������$��Km$���*DD�<J��7/vy��:�f� ��}/$�\-]��ܗ��R�����^x[��]��ۡ�tի��*t6� ���.�x�p�9�!�PI[E_��M�T�z�z�3�����q�uX��y��'�w�{�]���˻T��:*��|�O^d�v8`ݨ���ڎ��.��h��w�E�/ ��7j<-�xT65T��Rc_"����� &�dᴩ&��m�}ݾ��gr�F�2����C��UM�b��5�m��}ǹ=\R���qM��>���7$��fdh���.$;�' ����*�[�<���� seG�s鲋�J�Yg���nP��y:��m�1�OG����tf��dΜj6�E����b�Ի����q�	���Q�n��%(-.6۶Z��w ��0�%T�a�5l��6���q�ʩU6fZ�KD��q�D��wV������IS{����g���Q��T��:*��x[��	��`�� 'eG�n�u�:��.���_ ��q�U*K��4�{��5���B��P!��@����Jd�0=<�3���V;lFB�-�޶,g� 49�-v���������=��٬�l�����m�rh�vB�a�{�+�^yֳ�\���n{R1cp���Ձť2����v��)��877e�\��;
��5=�tV̕�haxrp{]8�=�p������4	 S�Ӛܙ��7M�f����a,9�m�:ag?�޿��{�s���?��Ga�����o�-�+�U�7;T:T�����;u����=4�7�ͣ�m��=��� Nʏ ջ/ �{��އTܦJ��uE�w�u_�DG�*J�׻����>�dÞ��~GV�@݈�-�
��"�׀M�� �;*<U%Jt��E'j��w�M�� ��;*<}�Խrz�	K��ݲ�Wj�v8`���e�ob�"�tF]��B��t�`9n)�)jh�m���"TU��u�頴��hv�ȡh�Zn0�� �زp�e�ob�'c�݀�(�ݪmä)�UV=ޛ��I4�/B�t��;�����7J�ڎ�]ݗt4P]��&�ŀN�=T���y�Rz���]�]*�5�m`�� 'eG�E�/ �{�GvU]���հ�� 3�,�UR�������|v8`� $QwIV&�]��[��o%�.��j�.Nt�^'��U6�!�eSc��=�h�E�n�Wt��m�X�xj���ճ�k]kuZ�+���j]�x�ذ	�����"ݗ�m(-.6۶]���]��N� ����uѡ=(��f�*�i���M�Nh�}�ۯ�����|��3���j"HpvTx[��	��`{�^�g�exn�X��:*��x[��	��`�� 9%G��R�`�t���w��0D5Rki%u�ϓS,��/j�a�Z5[�t�t��WCEۼv�,v8p?bɩ/�k����z^Ɲ�M\#LRH�~ɇ5USa�ճ�k���ob�8��ʫ��Һ�6�0vTx[��	��`�� 9GjF��v\�;�8T�R{y�|r�_ �>��rp�L�.),$�1�P�o�z�kZ�R�R��'R�L�M�6�,v8`��x[��W�_?�٭-h�bq)��ˌ%���f������NH�*2Ɉ;8���Ś�l��]�������mǀE�/ �{�t"T.�e�N�:f�mǀE�/ �{;3�|����7v�m���m�Rz��ذ	��j����j:t��WCEۼv�,v8`$��=_/\��t�k���]][GͶ�	�����"�߳rO}�~��|uN�|C�� ��K����ݻ���_���f��쀈&vb]��\����CO�i�v���~;o�3�[nݹ����ɭ�`����j�fۛ��phs�m��9ܼ��'����9��z}]���G=5p����Ur{&{n|eQ�k`�`�6�:��93k�pV�q��+va�뢑C]fk���9�Q�̣6���@��̙nq�q�ݺ��`�ѢCm]�����tc�ۡ�N�X����u���P�5�	煹),��MR7Y��9F���h�ڟU��[ajh�vh����]��e�WJ��|�l������e���`�� 9GjF��v[��7�E�/ �{;0�TxUvTwN�[h��S�n��ذ	�����"ݗ�E���n�uvUڻ���{������>�/���>�n��hf�-�M��D�����|-�x{r,v8`K������N�m�z�͠n�ܞ]g%q�.YG��+3�e�M]@�����Iv��)��W�{� ̝�`fΔ<�S`n��R��2�Vfk7$����
� H�E�! l�,` z�q�⠇�BR��k��w)�9���Т"=�yn�շj��6+$��ovi�??ي��e�{#�8��Ϭ�j�][�M�Wd��"ݗ������v�׼�Н"�T�n� �v^ w�<v8`]�� ��5�ut:���Ρ\GXϲs�=U%��%�z^�L��.ӸO]sF�N������??/�ӱ� ��x[��Z)j��WeZ���	��uvJ�-�x���ۡ�tի��*t6���U��zl�#$у(������B����9��˲3Bx�D]lHl��>��S罹�d��>�������N`!��y9�`�D�j	|~�1٧�<�>�p���O�`��T�6�&��x�ہ#����ʹL�!���)��oau�'��%����^hM�&h]�9���݀bB0Bj�&����I℡��2Ʈ	�x,,�B.�b����n�M,�5n�B�E����ڦ$RI�B
:�P��i6OPW�P�  �S���V	�+�F�*b������*� C`l�)��Q*�؈IE�=�`ouq`{c�#��Z����n���'� 7}�N���I�۫g �-�+M�e�1ۼ ���	�����"ݗ�sG�a��c�l�y콻,=fv�d��7˺���E�vl��4&�ά����cm��� 9%G�E�/���U��� �g��ݫ�ul>m6`$���e��G�N���ʻ"�~��I;V�uE��x��~� ���	���Q�n���:ul'j��w���;�\X�WU���
?""5@��Tҧ�A�QR�.;��GHؙ�.�j| $�<�;��E�Pm7l�-U�M�v8`�I�ql�y�| ����<��u�v�v~�C˵���h��qƜ���s��sha�s�`{�%qغt�#�q�j��`�J���c���}��?��Dl�m\���;�N ~�ܜԼ��7=��;��8�:�s�6b�O�i����x7�x;0�j< �{��~�_K��e�Wq��eܜ����wy� ;��p����j���� ƍ����t���ͦ� �ڏ ;ݏ 7��`g���%G�DT6�!$�n�w���o����p%l�i;�#`+q$S˫ϲlEҗl�j9�ܝ����kkmXaDX��K�]a.��n�v�����X+9������4��#����TK�8��%�2�p���h����t@v�r{t;N�l���j�����3�t]�W+q�ueꍴ�Un{<�A>ܰ@��k��x-�]��<r��襒��n��0[:��2+;��ύ:�g�h�nN���w����f6e�l�Q�ԋ܄3n&�v�屜��6Q���� �M[��������� �ڏ �t���ӫc�;T��x����;�4�w� ~�ܜ��M��yoI%˃��Z���;�~0�j<=�|��<�;�8e���Q۵n&��I�ͨ����{#��Iw}�M���ݪ����n���c�� 9� vmG�otBE�(N�wJ�W�6>��H��Y���]�e'��ͥx!��n�h�Ei���1]�> ��� }�2p�j< �v<�/m\E����I"�fk[�Ny��ߋ��{��|(��	Z�Q����U�n��`��<��*�Ʈ���|����j< �v< ������R�I�V�uE��x��x͑�;#���xv���Q\%9m7w' >�d���w�| �+� ;ݏ �}��}K�(륲~��N+%v�/k���]lh��u'N{[�jFضX��$G<.$�L��ܙ�����y�wj< �v< ���	.���]5j�ӥN�����x��x�̜ ��d璦���D�K��INН�U`��XouY�bS8J1DE�~�Sb`������A�+�'>�g 7�[8zZ:�+N��h���I�� s�< ��G��ǀw��/�i���b�w' >��8�U����'�< ���	6���W��B����;N�4p���n2��.��M�q7=�*Ir��ڸ�8��Y8^� ����G�uJ�`�I+EӪ.��5n��l� 9$x�ړ�ٹi�{j(�%9n��| ����I s�Q��e�TZ�v�L�X��3���3ں�{�6Dp�>�D�H-��`�'���Aɼ��ܓ�a>�O�Gnո��9' >�Փ�z��ٻ����N }���yRUY���X�~`��sn�te������S��˦�m��С=X$��-9%�WrQhN��1�m���x�#��qݕ�
�^ut��WCCi���ǀ�< �v��7��|Խvf#b�A�i��lWr������7H��U_%%�, ��<-�I�]]հ�7m�7H��ذ�������ݜ�Ջc!�e��ݍ���`�wg� ;�y�7H�'�P)��I��s�k2̴˩�b�\��Uz��=E�e-���������'��9��pu��a��!Ѷ�%Vݱ^8�9w���C���ݞwMnB�ٴ�%hk���;\���#�]��-�!�9�F�׻.��k�uʶ8�⬱/l�&�DKT�- au5����z�d��\���ŐmF��@WM/R��'��ɪ�)�2���YRv���D��#�z3Z���h�� G��uP� ��������vy�;��oTi�IB�ؙ��
v�ϳ���U����es�gDtc�3�\��N�¶����$� 9�G�� ���^Q/�v�WeZ���< ���{ s�)"*�-*�Q۵n&��I�ن���q��ISg��� ~���3"'�]�.J"lo ݽ� 9ݏ 9$x��< �Q��Wi][w��ǀ~���π?w����_ �K5h�v�����4y�����n�`�Q����^���\���u����Zsr��A���m�������j<��/ 7�բ�|�ݫ�p*G!���'-T�B�K���ȴ��� �A&dA�!%	)����7���v�V{��ԫ�i�J�tꋻ���� ��x�����W�6�ir�l'j�v� 7��� �ڏ �ݗ�ESmm۶:�*իo ��ɵ M��{���h4*�1X��=J���Ӆ�(�!���#14n��5c��-���[\h�j�RC�ۋ� &�x���	��nԧDi�e��N�WM�-�x��x�p�v�x�*6���Wjw�y��ܓ�>��r)�mC=0�/Ⱥ��S�J��͋�N����>_�K/*�j��4�-��N� �jG�E���z�}�l��y�HGj�\���v�n���ǀN���R���mX�л,v���ܵn�n�H��;]+r�a1���9c������E�!t�V7�?/{���c�'c���K�5TZ)t�;iRv�J���c��|����uo�^ M���m��M�WeZ�m��� �R��|��<�l��"��-TLV�[���l�Ԫ�W�_g�z���N w�rp&.5XP��H�A��#T�BIc�����R:��Өt�J�� ���{���� ��Ix�JN?�6<\�e�s;1S�C����S4m�W���ȵ%��c���"��74� w�;0.ԗ���v���~xVi,�VЮ 2I8~ɇ<����k޼ ��x��yﾤ�����c�.��U6ـw�+� &�x����� ub���l�j%wv��m5�<�l��'c��w�W���R��r�mܜ ����j��~��'�ΓRI�{��?��
��E_���
���*�PAU�"�
��U�( ���E����@T ��T"�BDX@	P��T"@T �B(EP�B"�T �EB$B!P�P�P��T $B�T �P��B�B
�)P��T"�T$AP� PI$B*��Q
 @T *�E`0�B dBA�AaP�DX@T"E`0PEB �DX�(Q"�B0DX��b�B �b��QB"E`�DX�Q Ȩ"'�
*��U�����AV�*�_�( ���AW��*��PAU�"�
��U|U�b��L����p��5� � ���fO� ���   � ��   ��    �     5l  @��UTU(P��  T�P%��B�*�AR
�(�P�*�R@�Q   �	�     �    �	H� ӟJ�|�f��彵�x�+� t�����^,�n�C]nm)o���_M���Kż�  �׌9ynOK�xz��>��m�=3�,�]��r��w�({�COy}m��Z��N�����^��h8 ��  (P
 �X@��Jq����W��Wzo&�������փٞ�V�'lё�0 ������X 1خ�_J�{�N���'���M糼ssz�X�מ zW�-�y^m<��׷����^ ��(   �@�� 
}�9>���wW�{ŕ�g��/�
'��m�S�����t���wJ�� �=R������k�  /v�i�g��V���=K�6�ҹ5ֽ��^[�)w �{L���\�w���N���m)p  ��@   �6 �*d���x������hi4` ������� bh � �;=:z� ��J '�  @�:=��� Ģ�s��@�@3�Ҟ�x =;�i�c)�'Mtq:t7��� �<    �P�=����=4��f�)�=�t=�g��[� {ޕ��m[ru���.���OR���{ʖ/��J�c� �������� �����y�yiɥ�<��ۀ��Jd��x���y5{��6�W�  =AM�R�  E?�53J�H��<z�RLL D�*���*Pa2 OД�)*D� �"�b� ��D�����s�c������g���x}�~�"���o�A\�������*�����EV(�����H�D�,BR$���@���HMbi	�LI�$���839̸ƥ��f����+���0���k�����n��BB��+)��1�HU7����S'�.�����ֱ���GR�ӡ�x(F����6�i����a5��8��Ƀq�}��醰#T�i���)�z�F��HP�~	k�1��.�%�,Mr�B��eb5q��
� �F4�!D):����� �*Lb��A�L��3$��n����rvg/�H��E!��:�5(K�����5i�����>;�Cq�t�!%.Lt�1��vj$���ep�� �!��B��9��sX�HɘgHC�F$��Si�� �HcY��1�L��q�k_w��Bh���B%H1��!
��a���}���,�#�7��$g�.)��u��q��S�ƾ�Z�	�Syf1�f`��m�ƹ���@@ƹ����D��7I)�4��Z����	��Z$Z��%1�!\��L�)�r�s�$
���93��^r�HA		ӧ�_�2�X�|�Sp��E	�O�g�s�Rt8ay}������2�D�g:�����&|�1S)RT*�[[�Lː��1���Hc�%�B1��>4��2j7:���S;�a���wY�Ӣd��, �9y�@6~v��:�
�i�Lђ�i�"1�����&��n&B�wm&���یˉ�v\_�u��8'�l0kn(@�!!# @�$d�X2�軤#�j�p�%��.2T���.�����L�%�0	��	��ٌ��7�Z4�Gn�"3��3�[���:���gD�]��lL�hF��:�.~�VCl�hF���,������-��eʜM!	��y����*a�k������>>da !o��jm01�����[2>�ʌ��2^�E!�l����S�d����w_:�B�� ���)�����Fh��a�����b>���P�1^�lJ�N�d��|Rr��rj~�D"j<��dK�tBC
@p�J�H��E`�bDr�-juҟ8��RMi����
H� "**G�>*2
E��#�	}M80d�$����fcB����0 RH?a�#`VF0�T��WAK��,h�0��>��$!�vc���.!L���VM��pl�������00H�n ���rc�3.AIoq!�
�H�
0�(Ĥ(Lh	I@nY�CQJ�L��HB ���ۮe�BE��)�&��"R��Q�t1k�N?k��K�8���_����w�|c�7�9E�"[�Y D$H$�p����!f0P��)�C��k��˜�de0�����2�]a�"ňa>�(I!d�9�� j<�޵�p�A�
�$�PH�!#�VB)A���1��$����l.�Lk2��@�t9�k�n�|٣<�ܤ��.���+ "|рA�hı�o>1�!�2�_�dƳ���(��5q��XU�\	�ɓ}	!)�I&��,,�mHA�P"���Ꙅ���}�g��d��,b��j���E�!�SIl��d 0 ��cf�����yfO��U��# �!,Y��8�IQ�e�jopރ	���0L,/Q�5]�xK��`RV%w!��lH�!�L�C���``��BLg����!��%#��j�`��<bo}�H:y�(W�L�K~@p�00�!�%$q�~zkD*D$�>9�%	��J�%'W�AY��_l���e C,�"B����>.3y�ϟ�RY�v��s	��]��uCN�������7Yfk��G
"�8�3��d6Rt�!�w��'��P��@1"0�nF�M��d��Z!�� C3����
�!��!RT�����#��(
x��!p���pS44��}��Ye��9�@ F@�p�2Lhl�&#HS��^��7�x�&v�h�(J��oC��y���Xh��\�d���Z��`�	I�g�"D�El���0n���B�"���)D�d9���3��+
$jJ2�131���-I�1d/���F@�J!�A�Q�z����Ơp� 0�!bZ�A`t�)��!���J0��aӴ�$�!����!�2�B}�S� !"DYj9�$>�A�B��\�"шD�$}�$IK�Bs$���1'�i��H!I3#FB4��\C|��a��cxL�a����Z����ns�	XCL����8�9���S73:6���(�c�$\�K�
��0�)�S��&���k��,(B�-�!�@#��}	�0i�3�>X)D�Sl"��@p@�Yc�o"dȘ���2��XЃAeB6�V�
�}�)�@X0,��6$ �	1�db������!�+������@����*� �ƌ�Ʌ����#!n��k������i!��S�$L��ƒ��ȕ̌�3]��8��S��:d�a�d)� ���b��`��dż��ص��0���������`o�{���?5����
9%
һ�p�,c�5��K�cSY���ƠF	 ��t0
���B�,
a�˷�)����4CXe�Y����sϦs�\l���¸L�cH�C���6�^h�� %���OҔʓ����G�K�}�����㯴��mBd�5s�l8}
����p}���x�$V�0}R%H$&���5ɃH;��'cn�-����T���g}%�8FĒLI 1RcF��.��t HŎb�'
BIA�şi��$7���q���R�D�k����H�������BB9:�3f�G��;�C���ɭ�ε�RB�����/>��H��Bm!~�p�n����aX� R�8a�H|h(��B�$������
H&�qN����I&�d8��)H|Z�7̆Ζ�~�!��e���P��&�5�\��%q�A7@n)��@i��Q, ���4�%p�4WrH%)��RS�ѻ��&9�K.K��I�}n31��܁��K��.&
��.�#���Iqe�LYHGN�n�#e�&~�%��q	'�3H����^Stj7Aap���lC�pV3#!e1�J�9>�`�p�(a�����Q���A,������d�Q Q��x�w�H�V9�8ȲHO����	�glC7�c(�`SXYL)�-@�b
ԉX4�KX@� H�H�#�18W�B�W�f(��L�@�A���GZ��hl��N�"q������#L�
�ĸ�ޞ��# �1M���H���"��ƤgaO�50R�fD�d>���,��:q�X�0F��>��1Y�k�w�'/O���F��pg��!��,��ˇA�!��9�[����"���N0�Q`�0�.�"C deXV0d� �Ôb409HU�u�Ja�-i0����t���.'O�cZ��$ab�!q)����C�Цr�8d�����;3��ÓzHP�9����}�q5�d��}̄���.xϱw�&LCF��BaY���K̆�+�y��<�ėi����2��q�Ʉ�IR�!���aqe������3�LgAi��."�W��ڭnKj�(�N�'�h�6�3T޶i�7��]g:�1�|]�W��`���8�Ϫ�O��9��AM���vB�57�i�{V�����p����)��d4�F4�"A0� *E*�oq����ɟ�M`�@����$�d���~"T�v@ �q�s��L�}�9W�mc 6#H���#����rR|t�@�Ѝ
�D�B������g�W��*]���%���T%5��C�9�8�"$c"�?s�st�)�4 �02��8v,v1���ŷ�s��4�1���I�\]��h��+��٣%�1l��_N���:{����g��8  �c�l                         � �                            6�     	    �` 8l       �� �   m�      �` mp �	��  N ,ڲ�;d�f�5��ЭvRSB56�Wf멻lְm���r��2ֵ�� �Lf�=@p�` m��nV�m���[��.�H�'���ρ���cɶn�k՜<�%�&�ې	��$F�VS�7#l�B@�bk�6�eZ�*ڕ�]���P`�I����N���dڧvnƤ���T.�����r�$[m�5��t�c�i9.$�z���f���mU��U8ݮ�`��!�6�qoT�a�]���̼J�Z���ˊJ��`*�mתVU[�vuO��;L�ně���1�=*�zt:�s�����۲&��Ke���Si�c���n�i[�`@Y�l��ݣ��Z+u���wd+\��)d�Öc!͖�@e��Ub�[j��w'ER�Ā ձą�m���`���j@H�e�d�� �9�n�k5j�^V80�y����Q3hq�-���~kZO�K�%�@Bh *���hӭ�[v٢�$�   l���A�@ u.��*[�  o  �[�L�rD�l�.�@ l6ݒh�I6 �6���m���� $���Zl��'Kh6��m6`�A��ۀ ��� �` �un�ܓ��O;*���UUT��n�>�'O���b��� ��amp��m��$ ���Z��ݶm�[Km� H	ke��$�E�  �� @�8��í�ے��(�\�:
��<pU����R�ɴ�  �-��6�K�PZ��f
t]K��!*�;�y�
�UnժUv�]�Ɠ6��[i���`Wq�%^c]�dǮ�gv8�N9�@�i᫪�e�s����a����c.�إ!Ě)jU��Fu��r�X�rkE/=��#d����vh�u�m��N˒�m �Zl�܃�gc�@kN�3�]q��Y].���ܖ67J�MZ�uLZ�Bޥ�cl�t�UW��Kk�*��]����jX�Ȧ��$�`8���fq�6��1Ơ�q�+���B���]�Gky:�4�n6\�le!L��.�l��j�n�R^��,����t˱�&qVK��e�yRZ;t'D��eh�U]��+*����: ���-rPUR��3�e�vZ�[Nieݷ�W�r�үU))T�T��2ł��s�W��͍=rݠ97S����9�	X)��!ř���iV���sJ��n6�5 �̽�]�
ջ%�T˴��R�z�[Jd�jYvyWjs���Y��U϶��U+�Ӏے�ʵm���b���Ѻ�zo�\c!�W�j��T�	ؕx���m�-�uד�8$���+'G � �M�z9V��Br���A�-���W �����u�n�����Tt��th��UR���Y9���l��-p��Æ�-��,sT�q��|%�6�n�]�6Ͷ�i�Ӧ-�]�n�plt� (K�ĥUJ�:�n�C��  �䁶ΐ   ,2M�d���v� $�]�9�{d�-�jͪI��k� �cm�D5�jV�v��D� ������*@6��m�j@G l���U�m�W�;^���v�M(�tS��0�AGOtm��ʽ�m˭)��c�l�]H��:t��B�#j���*��.u<ʜ]j�-�9Z���
���C*oLEq��aD	V�V���^�)�m��8$��p��i%��-���� +�V`�5U<�4� �T*#j�����v� 	8	%�  ���m�!�i"B��n��h��m�	-�-ַ[v��h  6��'Bw9hl�1u�d�f�
�YVٶ�ٴ� I$�4WX�YK �.癥Z�]q����\���   Z�f�m8 r4��)��J �T+�nT��wf�ڢ�[�h 6�>����9  �6�`[A��m�l�tцջ .���D�G��3*Ym��T�����L�BXf�B@ݳ- �[�x���n8I+�vNT����վ��k:`kX%�����[vU4�v�r�e@��V��Ao;�vWYb��X^�p�$���������-�Ff���84r��C/= C���`p�M�ӗZ��lY�'�X �����z6x.��5RWl�6*���n.��h�h㤐:L�8�5R����0�+ܽUJȓu�`  H�d�(
�]sse�GYHHju�V�ᵵJ���RS]���8�j���@���+�V����� i�	#c�ٶ��vqI-� v������T�X+���v�gkŷ�q��. n���b��v�����# I�� ��6��6��r�6ݼ�`p[PiR�p֎��;���UV�5UC��n�8D�� [d�������Uj���kխ�k��Ӷ̭R�*�R�mh� ������ܴ]�n�A�ݤ�۷���ͮ)[-M�$�e�Tv��pi�I)l��l��I3�a�����ӓ*�O%ĵ�V݌�N�N� -�h��6^H5T R�:ۡ�R�p�dଝCl]h��`���UUU\��W&rl����R��$HMJKCm��i� $[@�����n\� m�l�[Amm��,06�6 �6�t!�[P ު�eZ�Wn��.��o�}��@ m�E��j�$W[sE6�@ ����m����vCaU����"e���B���I6� �غ@�@H�ti���ţ� �٫` �I+6�ӆ�ۉ$m��� H8�[i(,0 H �ma]6 [�� ��YUUYXt�+T���[@�� 5��kKh��ֵ��l h�mm8kX�$H  -6 -�Z��d��t�ʹUp���m�d��.�LC�]n6� [��h��*�G�꺥Z�����^Y�s 2�U���ݪ40��0U��	�V�D���E�?>x�|��`fm�� �d�J�M�l�QRZ���j�`�v��h$ ֭�K	$HAͶ�S`�  [F��l�����0�	 M���ln� m��  �  �lk������3�L���`xK��o+D\Ȓ������ƽM��}����K>�ﭮ�;]��ڭ�����pu��<�W@u.��Օ�QrCG^:KPf�`��T� G$	v�IRu�m�� �b�]�m���4ѳ���t��um��.�m�խ̀ 6Ͱ���� ��C�.l����e���%��Ē\sb@Y��m�Z��˻��U����}��m
�`�!!���T�Unl�^֜L�iʻd��n��1��U,��*nJm�avW`m&/Z�m��j��8�ll��m�-�;E r3�l�m��ݛgZ����&[m7mj� ��� �n�l�`  (-����RZ����@޲[@�` �m  �x��p �l �3��� ��<��$g�
%A����n@y��\ �`k� \ݤeZ�j�(�ۙV�) ��+�H5UU*Ԭ�ձ*��r�WU]t[v� ܱ�p��}���P �HCv����%ɮP඀�В��c5�����
�U��j��eS� �M�UP1��g���g 8 � mm��T۰�n�H���t���׫� ګ` l�p�� �� �   ���q  k[: �;l   $ m�6Z� 	4[j@ l�h�kd��6�96�l�l4R����P�� �  6Z  ��l�P�,�l�m��kh �h��$-���h� �n� ����a����8����     lX` 4u&��[k@   �k3 :@[����H[@m�#��6�Q��  �a#��p �l�|m������ެp � ۰��p��۬�ݥ�O�}�yj��%:Xr�\R���e�ګi��'d��0G�t.
TH'���b�MA��~?��ёL��z�6�5݆ٶ p6����]XjU^Yb� �UtTWf�G��0u�(U)2�T�dvj�ˑ�j����%�Kk�إI�KX[T�m�m�m��` ��5�n�[Z� ����p�m�5� [@�m�  6� ]UJ�#.�	\-<�� �m��!mm� X`�]�  m� �   m�}��n`V���H�wgf�� 6�ګZ���n����{fV�	�iV�x)R0� �U*�*U����R�����������V�
��:�]��e  Cm��`��i  �f�i:���(��i�y�v&2&�#��Z(}���r;S� ��E�)���Q		��A��4�L��w�. �GO�&AM	@°� �U"#�N	WH��!���"L�Di�	��Q(�uM���G��v��L*uGg���������2*:`�+��Cl,p��X�F�2�|!�	(�D�b�B @��N�
�t�U8��%�)�+��_�/Q]���hE�������:���*����b@r�2/J��P�d6<W��@(t�AD"�!�@�`�Az ? �pBP��T�S�:C�l�X���F��@�$�U�X�vT��Y�� ��p\�bA�+� ��������0ŌZ�\�؀D�Q(�����@�E �[�kT��*/#�SjD��v?�8�H@� C��9��\A؃��U�� �@J (�8 �@��V���GV""�T(8��v��E����;Q�E��>M*�l*����ѕ~N��x�X�H0� X�b���c	!����� � A��(1��X� ��(u��$�- ؃��~���AD	!$	$0ID�BDRAa!@�]<^EC���|��9Pl$PlPiB@$c�B�����&�@�u�[��H� m�����hW���8N���=
�WJ;��2��8�8��A8��O�g���*�Q��zԔP[h�+QD#�j"[�{����t��{�_����5�  � �Mm�    ���u�m���l�l�ɦJ��h:���c�aݲ��
i�3]�&��t�Pg��n��{b�L�s�װ�x����9�Y�v�z76ն� �Ӻ�����g�:��BҠA`x�8q�x7�!�Q9vu�y5mٝ�!��(53%d,���mKS�ݫ]$�^Hθٺ��\V�9n����U}�^�ȡ\t�'��k�vΞ�آ��o�Mv�3�ZϮ��:�J��8�%�l���L�`�On�;r��ru̓�9қ����-�fK���]����	���Ƥ�j8��E��agB׏�h�W=��k�7<��݇�-s��B���g��a͒�\UYuN�U��l�Kz�dr=7mvyѷ�ƻv�*[d1��qɹIU8M����1�V����6���P5�wC��t�q 6�c@*�M;77浺���I�nG9z'��1p5����n�Ͷ��]Z牣��x:6k'����.v�ws���:lˌ�N:���si��$s��4M����-�c��;]�#���D*�y�o>2n3\v2�Z����ok�X$݋�cJi���h��A�ym�\8M����fn�X����;�������K��庠��u�r�)�դ
5b�;S���Ͳ�z�Xŕ8�q"���H����FI�Ln�#�d��<�oMs����S�Wnt��d�yf4s�(����Ud�'@z����&��n8e��k/q	����N�4�����ձ��i��ܽ+�j��W!�Ksfˍ�A[��vU�"1]X�4�U���ZW&�N�e�i�@4���HE�+�n6m��p�%�H�T��Ыt�mŴ�MK%h܂�ޕٶ�v�G�Hb��T���MΩ-Y��A h�s�)�������X������8v�OUcRʆ�[(6��q=�l\jj^t�F.ܸW6��W+ɠ��ڬ�7�Ք���~�����!��@2~J���?)�@~Ej`]*@4p���'��hO�lL���������#�9�N�u��`8LV���p���,���0�Fq�,�z�������i0��ݐ&{Vb�6��YvӇ���nc����6۳���ʌm�9�.�	�ݣ���m���ܹ�OQ�$�K;�=�v:�M[],
��K�3��u�ѓ�g3\�2��g��n�\d;����RlU]�[N�!��)�]@���!Lf��3�2��W@ڎ���c�m��A���9��۷��w*�����n��I��u���ŕ���� ��q��U|���]X�i��h���N4e7+����Ԁ��P���n�������	��"�1fk�;�۫嵺������M��M�18
��@f6���� 3)�A霦���3c��8�Bpqʰ:�[���Sr�����Z�wEã�&..jg'�v�ob��̔�(.�ے��'�8��n�g�u��k@�e���4��=O����~�>��������p�Q7Ws3("�b���2*��}���bQ���>�It��Ԩ{[�@|�� ��c)�Ҋ�H1G��ͺ�:�[��%վ�1g���FSԓ�I#Sw����Z�����Z�k4��%M(�t�3�5XWZn��� 2r�G����]��`Z\�ݶ���l.�K˟;��qM=�v��ЄeSd�8�*�#`ӤDA58� �����wn����;ך��#M7[%7RQUWWhcj9�2�� �ݗ��RGUg�|i� �H�X����'�c���|�F9�#X�R ZUH����)KM"�U���;�`w7n��;����	)�����Z� f7hcj9��8b�R��I8�M���ݖ�ݺ�:�[���^j�=U�]��
�)M�&���8��N��m�#�[k����e׳���[������(e6S�J* �}7��'!�@fV�@d�t���H�"����30�2�?�dW&L�ܻ�נ-�v,��u`wY��FpCD��:q��n�8�#�}U�������Ɗ��M�nG`uwu��۫�}~;�jO�|�h�����9�+������F�n�������q��� 2r��[�N7H���߽��On'mO���[�F�C�����n�Xx�ݖ���h�:���_;�ϓ>F1���.�� r� =:� 2q��Hk}u`b�6�I�A��j*��,�vN7H�j9��8d�����9��JG`uwu��۫�����n� ��X�zD��RQ�a�UrGխ�Bˎt���t���� ���8�Qʍ�*���n����y�I��{�}�wF��<-G�`)PhREe�q�ə����9ɚS��.�R�T=16H�mý���ԜnL�M��oۋư�@%�]���M9�f�0�t�4�u��� �[:1ۗ�#�lo55���=��=9ƣ����;z�k��s�v7����vp�hB�l>�t��r��-М��{�p�\�&�bq\��\���{wn^�=n{p�R۲ib�q�E�jݮ�\�lf�.�׹6@��{����)o��7"�E��u���!=K��p���oY��kY�|�^��;ΛH�JH�8��}�`uwu�s6g9��,��`w�lh�PM�I��'�n����������M�cn�ct5vs6����n�囮����:�ǲ.� �LĪL��b����P��4�2K���X�̭�� ��M�H���H�n��� 2q������}���c�뭀{x��ܦ���%��{r���Ϸ0��Y�Ea��&�\\5�^Q
��{���B'뾈�Hd��@�����T
A��s6���s��P��2Pbq��
�fI(d��׋.(�7"�/ٓR�2I�"���tqG*28X�MvV7Hq�@f;bue�3R\Q������,y�;V{���vi`uwMvf�[��JnTr;7H������ r� 2q�@{c��<n�ɓ�#h]wfrɸxdug�^{`�/�0{.�x�-��(�"-�S��Ut��v�NCt�������'�"�b:�NWku�]�v�{���vi`uQݭ��qƛ�0�b���2(��3�JR@����B��V�Q�p�Q;�v K{sŁ�����n��JJE#�m4���Z���K����� Ӵb)���H6����vi`|��]����`fd��՘H�إD���+[Սmqp���N���n�ǳ��ɵi����U5R�v�(�FG����vWw]���K�٥��3�F&ҐP��vWw]��#q������`umf��F���i��(	�Q����c� 2\k�N7Hn�IT��!Ԍn����UWT�=��W�����{�I�1�*�(��~ξŁ��"�' �R�Ӆ��+5�[�^'����/Bi�s2[mѼWlwj��{
�ol����=v�S��n�<@��T�7�F��8G`uwu�=/] 3���:@f��P\L�RI��JG`|�5ߪ�l���`y{ƻ����;�(�T�J R5#�3�����8� =-�@=d�3�A�����`b��vWw]����`w�4�3��lQ�I��#��ƀ����]�^w���ƺ@_�o��{w���?W��H��c�%1�K���\��LK����-���7!vv���!��]nregW6�l�$�;]6�1YWm��6MvD�.zNc�p��Bݹ�[���I�.�EM��壝X'
�p�8��۰p�mn��l�ҽ�+\Wa�]�t<��\-:YawnD��ۓ-=/R�nٳ�-���|�1@��1���@k0]DuZ<�N��,�0 ���� �ٵP�����s%���������h�s��]�Fӷ�;�}�f�Iz��9��m�l �ܨ�v������,YY�����3�F��ƇR1�"��@f�P����H��(Kn�]슈��J��U��+5���z9�;��v(^�*݋Œ(�w���p����V�s]��٥��0�`fn��m��M'$,�����\x.Rwm�u��B���'�d9}�=]��#�n��[bs������dމ���".���F��?6ߟ��������:#���Hd��@6��F�!�bT�1% ]ٓX���$�b s[��s�ԓ��w�o�4�3�ծ9 ��R�2K3&�K�H7l@�;@n�T�D�!`|�5�n�,3�fM,�lK\hu#�$�>m�@�;@n��z��G�F�sat��-�]���m�7�nY���]���]*�<hǎ�-O@Γe�< �:��l@z^�@y����[
n%Q5#p���ɥ��^�:ۻJ�.�ɭI2w37\�<�����g!�fU��ؠ>��Tb�a��2^}�����B!�u��'��dB;�`�LS�4�"d\��B��V�q5ϵ�q�E��`P`BP�X��Lx�`��c�,p�"�pP��f��U�A!�? �		$ $��u�: ��٠�=_'ЛM�񁐉@�@�/ 'Khp�B)�;��c�3$d��S�t,����" `����*�YIl�8��"B���љ- H(�
D�f9��<�d>�'���0:���2�|�
nN��X�L�P4��]��F2�!~>Ag�����6���hQ�"���:�]1�5�tp��Ú�({ |
�A"���x�U:
l�4@ި18#��m�B*d(���-:�v��"`@.���7�=,���� �+RT�DJ!+���������B m�}�m����s��@n��yh����YC�R��u��"d��z<{�g'�R;�Gw{�����x�?7��n��p�,r��cg����v�6ۢ�v+�9�0c�c]&I��'�w�&$x&~�3'swz��L�z76>ۻK�_?$̓���M��'��>P��*"$%P�6k�&\�J ��G�'swN�36���&hs3^b_�hu#���a՟�~��wOK36��>��`b�du�#@�7TwfMwyJ�>�ɠ�d�3'H~�8VԦR��FP2a�S-����b�=�'�>�c6��x�f����@|��&�͏���Ҡ� ��WQ����dqp㕷V�m^i�+������|P>q���]�>Y�m��m99'ӒW�~^�;�ݺ��6X��Vӵ�*oQDBR��H��ۄ���z� =/] 7t�.�� ��Q�V��,�۫廮��ͺ�3�ԶDJm)M19,�j�� ֡ n��.ԉ����x�@|��$�w7��fl����f2g0�'o�Ɉ�2�4��N��ԛm�$<G �[s�h�(t��v��L,U7"hG�[�v� O^��3g'Nܛ�cgmI��F�Ev��%⃚��Oۻ��466��j��$�EG%A���E�Jtm��m5�t�lM�铢�p��7d�q,��t��F(������7;OY8��u(�%�Cɲ��!�k���D��8a1Tv�nv�9�n3�fb\f�ۃ$3�d<�@ʦ����*8x�E��۱��X�«�c����b���W���{�;��UvJ�)�ڙ��gr�����P������͒T��t�r�36X��V�w]���u`b�[�܄�Ԙ���3/)P>fE�~DwoR���`n�AԔ�CNIV���y�ϔ �v����ބ ͇31\\� �*\���2��33tn�O���� �we���T��`��N5���n��/N���rF���u��p��.�{bC]��ρ�FU���*9+����7sn��3#�2eɒ^��ޥ@nA��2�)Q�$ď4e�*����BL�NG� Ⱦ&滏n�I�w>��O��Ms&MɔA۪W xq<�����z2��D��@woR�/�-�����P�7���u`��7sn������r'�mIW1�@7�B2��z� ?G���~���}���_1�]���۶"���&�ny|>��=�X{c�v�=��>�t	�仪����B2��z� �����cNI�4�`uwu���V���w6��0�$��J	!)R��e�* ��&�!	��̒x4
`�Lb`X���"�_�fJ����=�Ewn���HB������@���j�v�o]Ձ���T�
t�NTpNKw6���O�ݟ��ͥ@w�@jI�yF�ʍd-��n��ok��.�.^�޳��-�z��//	`Ƕ�l&�ۮV�n��l��@7�B ��h��@nm�PT��$�7A���ͺ��ăw},͞,�ݗ�RF���8�H��@ڗW�ր��b:#�d��s�.�Q&�q�SR7$��r��ߋ�O��gRM��ѩN0��
��K��V�)�� �y&�L�$�������)D�("��j��ݠ:#��ޏ 6���zX��K��Q�)����lI�0�s��<����ۮ���)��u��:�hL�y�N�Dƿ��uo��%@������~�����`gnp�o�n�����`Z��'��*beP����rL�͞(��h��z�I��椀:m'*8'%���ŀ}��G732��ޥ@��@g����	Դ����2PjI�ۻ4�6� ]�M3&\̣s~��و�㠂fQ�^&h���.h�ޟ��J���{�I6R |U
$E�H׻������|����͒&^l��H�=�h*7�ĉ�94;2����[lx�̇3��b�bb���l�Yx�4��y���q�)0FM�n-ϒC%���`���볹l-�g`]���$w�-��:_�L#�]*t�4W�ʬ��ҵ븍���@{A����@ъ�LroFU������CnuFI��n6,�8�cpv������݂��-q�H�8�xz�� 1����9�!2b�9�.n)[õ�4��09����p���{p�ůn�f�z>|��0�@�q���~��mՀ}������;��P�n�xyx���334e�*�I���D�t��Ԩ36_�I�z��m7�m9� �wZ�w]�6� i�31T���������^���`��`os)Ps'n����
`Z��'y�2M� �v�ﳻ� ��c� ����ͣr-�,��x8���)�	�;��:�Tq�����>���!v��>�GWīl�k�&���r��ݠ3u��H����^�7�:�ۈNU�}����HG TpJ�S�Q�	�4+T����g[��I'y�gRM�v��UUč͉�M?TjGCt9,o� �v����&^�(@�ր�[Od81�bԎU���T���X��T�fM�d��3~T;c�w�����*��� ��>����� �͖������I0(����ټتP���wa��ۘz�6�a9�l/`�{�����#�)��r� ��`nf�Xfl�W>A����L�*kȂHJA<���w���&�szh��T����G��FW��J9QI*�77�ԓ�w�5\ E���� +���b&(Q`�X��3k$��&�d���T�d�<́
"f캲��D��� g>��jt����5f��D��N�����}����o� z�����jbH't�v�����ȓ6�yv��/uǍ�v^�ܲ�m�U����S���)콴5�o� �v�xڎ���s�@=�QN�
	�"bbU _�&��4A��J�/;��˼�Z�ܷl�S1��1D�L��{���fMɓs(��� ���`f�Һ�m�9�NG*�S;��f��ͥ@���;2��|�a�1a�W��� |�����wۿU�t��TשD��#��˼�@r\����;;�P�̚3�ڶ�sڥ�e�wZ�[Dl��{)�iu��pq��{5%s�����A�N�g�2�&e|w�4{2� }���̙7�;w�P����dP��TL�4{2�srI2M��@v�R���ֲd��$j����R�Q��JJ��},��Tk32I�̼٠6�iP���8<b�x�DB	x���I$�ɒIGn�� noM�̥A�ɗ$ɚ"�zh���A� "&&%P��hfeɒK������@e�R�)K2W�CJS��G(E����km!,#0���g��(������~��ֻ�_�0:$ �1e����D��a�]�4�TS�:C
]�RQ@#��O��>�$����E��`EbR	�����S-7L�� d$n\��qv���T$� CF�?J �(G����DӇ0xA�$I�(J�S�t�Т%��;è0R���+�0#6@Xȑ�*���X}�����Z�l���4}\�R^�5�jE�H�m0�\+Mh�	a#X\�2�u����q��`&�Bl��,1��c��CR>�����:1}{������kp  h���     4Pغ��"N
X*���(V!�p�����u�ږաL�#�\U.gq���r��iɴd�5/a�[vt8�3� �1�kW ���9�ݎ���k�r��Ӎ�|���fᕷZ����r�-R;9�����m�;P�djUiGk���1��z��QƂ�3��Ͷ���ʥ���/mt��At�A{=�p� �S[�(�q۷9�^��y��K�>��5�ݳ���p�b�4^1�6�O�E��s/i�5����v�v)�W�:�Ah�6k�V�:��m�Ě��t��hǳ�%Ֆt�g�n;I	e����Z4v�9�=@/���ay�����[F�*�]��7h��Ùc;O;ts�X9�m���
��MW[�7�mHGY亳�l�M�x���`��%���/;N�!.(*9�*�\��]�����_�l���Zf^�"���e�.��U�\�]l��B���|r��.�����H������`E�Ίn#ѻvG6��ؤƩ�D}z1��-�A�9�F'9�
k��(��³��[�O|h����r�Ҋ��G���jS�{������[�{)��S%�8�^sr![�2l�7�H+GQuE���a��Ƶ�YbZm��UŇ�PVm����#��*m]���s�H�nz�:���p�&���NiU�<���pӀ*���7n��[2f���vܽ�'v�ӌ�]�R�aL;26E�x���P=/���j��0V����(�Q[.��S��T�Ҵ���gq�F�ij��I<\����Vl�W�<����3��;a=lky��m[d�c�^�/YI��G:9%�ʴM�e�&��k�1��`n$�e��M���9���h�V�d�.��X�΃m������9�����H���t�O/(ܠ1��!��ûp��x�d��m�6��2\�z�c���U��kbY��9�q��
:Á4�#�U0�'�R*��EL��Bth`
$U��@ � \jA3���L�\��9�L�Ob쑬H.E�z�z�3��W���UԪ�;FF�d�>�N���n��.��[>���O�lm�	�������&sۺW��{a�s��C�v6�q�uΟ;8�� �� .��2I�v�i��z���*�[<�]t�!#�/�����g�an,��cūsٌ�m�l[���em��9��̨��1c9M#��=I�X���0b��&�)��[̸ݙ���$`8��8��[�sA�3�
�������z��+���76	������y���ٍ60~䟮��>�d�e�-L���6h���Q��I Si��`wv_��s���{�P����
�ɓ�ix;�}S;�J���`u{|�Y���9\Ksg� �����Ԃ�+j�IIH�;W��flPy:Pי4̙?�sb������*�)R8��M,W*������u{|���vnm�Rn:��c\c��z�r��d.x��h�v��`������Ctc˷7����? ��k��師~m��7f�3ד@y��;�d���<P��6��ED�S�%v�͗|䣜����QZ� XE��"$D1ehP�����8�d�T0�fr��cRO���j�ב\˙�h�{yDE;@��bfh|��FcѬ�����b�.�f���SrrD)$V�UR�OyP���^M332�d�򻞀��u���6��VWs]��,�z|q����^�ͦl�D����O\'MYw��7q�c�=lO�cq׃3��3G=�}��A*v�HJA
8� �����^c��f?2f\��>oE����E$��nK��~�8�����ś�`��UU$fz�nF��DqDG/@]��@y�yyZ��!2v�Z��|M�e������x���:T�1��qPs$�.e9���4ތǠŭ��嚛`��%�	G�w��ջ(ms�Nk���
%�s2Jm��Ms�5�˞n3�s�{o���ob��̦�:A*T�w)7o�)��Cc�O��?zPtܠ2s]t}�}h���w�j��	�RE`}�u_�UI��v���˻��U�Hͯz��p�N6�7r���Ԁ3�w�}��N�Rv���0�	S�F�������U~�+�q��4�wE�Fc�y.L�jfa���	L0!!B �2�d�2I����(�w0.RB�̴�L�?�"��\�̖g}ǀ����vX� �gu
�nA�#U�۴u�D��r����v�Vn�{�(������?>wύ7(J���������k��v{��r�A՞�7^�0nF�F7��@y�yܒf���-�({'K�9\��Y��5�' r����3{����D}2n�Ze���q-��ڪ����a�W8���v,���ՙ��^�*����-$�]{|IQ��9"�)�$�S�N�I~�s�r����1[g��Fum�x�{���~(})H�x������{����z�Ulqƭ���o�V"svjMY�Yi��m{-�ԍ�U����5����pu�,��)9JSU:�"f��S��I&bw;�r�\c��q�mu�ӛ7l��;��ZU˛�v��,z�����u�l���uw`�m�e��C������ӭ�Z���5:H�&�q<�eʝ�ٶ��x:�\�+�X[d.]m���O�<nݝ�%QtS�g���C�Q��S�n���2�̖�x�v�Z��r��Sҏ����������J��s��%����>uq󋕴ה��� ��}������R�I|�u��ՙZ����I%�|%O�8ؐ�����I�u/�m.����$�'�'i$��5��ꪦ��D�W��B��9R�I-��}�Is\��UM�~�?�I#��i$����D��C�����/s�����I%�=���$nmԴ������O�I-�<����Q���M;��ǳ#���$�s(��)󻻾v���[�b��Y�f�J�)"O�R��'�6�Uw:�m�႟���s�*s�Hm`ʭ�G%) r����H�۩i$�w6}�I-ɱz�m%�=���%��v��(�1Iq�c&um���w;��`A��\�s�\�/���i$��k��$�6����w�z��������I�[-i���$~��KI%�s_�/U6׷�I$�����%�Oi])M�G'Tㄴ��M�����I/o��If�ϾI~�W�T{��Ĵ���$����Bn?�I#3n����O}�N�$�zz+I%�7W�$���]~�h�8��]�i:v��K؎ūn�����Zl�{����Hk���|�Y;�Y��+Ē��$���O�I%�6+I%�7W�\�z�G�x��K6��H��U)�*H7'�;��\�rfd�rfM3.����|��v��I-���ޮs�T�[�y�IR!S���ZI/z{��HܚKH��:�(��-F�H@B$��"1Q$@��N�|���
�}���ϾI%�=����i��I$m`�%�9��m���/��L��m���w�]�.r^�ߗ3&L�;[�|��<<ECC��6�N9	i$�ۻ>�$���r�Oz?�Ik����3&��I~��m]k= �qs���K�V���7(����|>����Y�u�̸ďUk�����_���~�;I%�3_�$�,�?ܮs��K����$����7J1AI8ڨ���Ic��������}1�m��{������8��S�9�?w��z$�U~~ }>߹��Iw�����ގ�I,�z}�Ik�i�HtR�	 �%��g�>�$�1�g��~����m�*�&(p��UW��}��v�K��{��
�4�I���]{�ZI%��ϾI,y5�I$����K�UUc��
�� Ĕ"�9��ݭ��COg�w[��!��;��t�\l�`�m�?y�IISD��n9RI,����KM��]������?z;I$�|�^Q�$IҔ4���KM�����O�I%�vb��������I�74̾l��
P4ƩT�A�I%�����$��c��U~�$�=�������;I%���)I7 ' ��|����Gi$�wޟ|�X�h�$��fϾI,�6�����M��H�$��7g�$�����$�Y����$��c��V����^��$�IQ��C���A�Pe�k]���g���]ۭ�q���h@7k;7L��nϢUnf�)v�B]��n�έ�M���!6x�H#������|�;hv�R��`�$��s�F��v�)q��Nst70�lvKo�> n{|{ny
��`f��p��t�۞;�V��k��v���6��n��@^6���v���ocN!�f�K��|��X�^��m�u�ܢu
yW7{Ē����q�\[�vວ���3��ߊk�]{9ͻ&K����"c~�-�|�\�U~� ���~ ����Iu��ꯛI.�}>�$�����!�HRT$����w6}���F?yKI$�����ǓZ��Sm/g�}r�T���$�O�I#����_nl����z�y�I$�7��KAm�	�ۍ������}��|�Z�y�I$����_���������? ���]��d''�$�<�դ��9T�wӽI#����_f���ݩ��)���9Q�����Vv]�W\�s�m�/X�Bp�=��m秴�Y�.6�2�I$j�I.�l��:�T��K�ݞ�W+����^��9"c��)%��G^ꗕU����9UE4k��"P�9VbC 5q2�0'A T_
?s�߷����o/s��I%�͟}�r��6���St��ʊH�$�����Ic͎��\�s�UUs�E�����$�����[��fԑ�ؔ�D�}�I,y��I%�͟|����-%�W9T�����I/? �n�HtR#�E$v�Iw3g�$��U�r�����$%�����Klv�Kp4p%1D��^0:�۝���G�wk�X�u���Y��s��t}���w��>ݱ�#uZ��� ?�߱�I%�nϾI%�6?ܯ�UUU�K}���K����"�(i(��q��$��7g�$�ǚ���]����Iu���_�����}��)�	Z��_��_���m��s����
�DH1���f!�.)a�+��z�)��#Boo�HB$H���I	��9�`x!�f@�d`D���
S%5§�!�,�V	�>M�����2ZP�X@`1!5���:S�!������RA,�)��v�M?a��> �4�\/�4,�vM�s(H�cm�w�dXH��?fa����T�@9�(�ؘ�����!�q �P�D�C����/@r��0�b�Az�!�]���/_'9��O>�KI$������4G��iڌ�RGi/r������|�F?yKI$�����%�6�i$��*�q�$Lrl�O�I#�uKI%����ӽI-{�e��]����%��U^~���TI$��c6��7;SQ��9N2n�=<�s[c���'6�;p퍿}����/�l�tQ �����w������뼞f�L����#�b�$��ߚL�RF�iH(Ғ}�Ibͺv�Iw3g�$��ݎ�I/�v}���r�k��*6�ԇE"9P�S��K7}>�$��2b��2\�I�f�{������E;��wM�D��M9RBI>�%��UU7�ޘն߱�{ݶ��1�oM�P��:�s�K�L���KS�m(�)4���NI��������W9�k�}O�K7}>� �ݖ�Uo�^�R(Q��NTK��Jh�40�C�\�i���s��ܳ]��*�~򪫕r�6�Lrt�Q��7��u`�� {[����>�K�mI/�:iڌ�RG*�;���>��`|�u��۫�*����J��8܃���������n��DDDL�|� f論�ٴ�(�$2��X~�?s��;�n�* ��M }y�@fd����m6% �I��ͺ�=��8�wg�f��=�E�0&M��C�d� ~���ŀ��%�v�ǻ�{{����-��UN��yvU�&��S�^���k�2IF���q��+��6�f�'��ۂ�6�Kturd�V �9�,t,���q�!aԝ,��tp�n71u1�f�}6�����F1�,��Mӳ����>35�:�,��n.H�!�&��s�t���NL왍�n}���O6۞�-��v�r��UG[_��8�pshv��ή:Lw8� Y<'�;�DړWg�9�2b`�2L��*�kX�h���s��[�����\��̕��UW)H��j���G*J����`9����� �Z�8mU�\�RNR��KWs]���I�|�f���>��~�*�76ԈԤ�R��nG@[�lP��T~&M��� �� �ޖ�`�ct��r�ܑ�w6��=�� �k��D�7Ԁ�*'���T��ڧQ�*�>��`{��]���sޖ�ͺ�5wS�4�%0�Sr�n�[˷U�G<s�n�={�[c��^���v�m��3nA�@M�I`w6XwvXwv��\�����7�=M�m() �2��s�$���u��~
>��@r�U�&eə���P�zh޼�3%�[I��bR	I`}�۫ �f�=\�����;��,]AZڭ�:)ʒ9V�s�M������>Ǆ�/���X����
�NBB9,�͖���� �v�mۙ"l����Ň���:+.܅�N�1A�&˷�m�"f�����;�s}��8�0�p��~m���cjn��H�� ceL�U�TpIsV =��@�� fk�wf�z:Z�����ۧQ�*�;��u$�}��S(��6���@-BXZ�`�.mQ�~IBI�j���N��v� ^'W�11$LrP�$��;��`gvi`}�۫W�o���~�ꍥ$t���`n;b�#���G�7�Z ��h�����㇣8�<F�>�΂��p���ힸ��<[���^�ݯ4��m�0��"�Z���ٔ��y4�^O3%�3/@nt�@s��\��'&%L�J�e����}2�� ������mU�@�M�*HI%�w�������Us�T�s޺���X� ��PIJND�&h92f�L��s�‼�@�ɠ��j��DȎ�3�gRI�91m���C�DJ]�J�fR�5�2g�͟�/7��������1k"����H���gp���`Gk[om�z�����z��I�8۾�����+�Se*r7N�F���3��`�d��9��p��Ҡ��6f%�e����33@��֤��(�s��� {/&��.f�7���yfGxW5v����cj=v�=�� �b[6�m�(I߫�7߻V��4��&��d�7;�(|t���I� ����qw7��7==5$���I*�J�z�h��D0�Š%
�E ��?�md���8%�BZ���f�<R�U�g�٦�c<�j����%)ڑs��9�qls��Y&���Q�!��<�v<�����̷T�OQ�n.�^�7[��=5V匇1� �֧<n�����*��]�����^u��\�=���z��{e� �j�s���ѫny���w1m��e��|��lP>�oh�ԧ�e/��|�!�[��v)L-ʀ�4�\��w��w���7������9�����:��ɻmr����v�V�����NLT`�+�0�n'�6��!���ր�v��Z��]�75�*���M(��R9,��/��_��3}���?{ߥ�}��~H;�i	��N�(DN���w]�f�@y�b�P�aO�TQ���jJ��[��`�zXfN�32\��3{ʀ;���^&&9)&E$���,�f�{�u`����ܕ^g�*��A�)���o]S����nCӎ{u����>d�;���c�ٸq�ww����Q�
H$�Q$��O���sn�.�3$�&^�/;����S���C�M�1�L�9��}�;�XD�0�Ȥ��I�̙��3=4wy4ד�k&�F�Tc=HtR#�$r�7},�ݠ=�؀�֡ �UsV1U5We���"g7����@fkP�;�����J��M(��RI,�f���� �����@fm�븹��}�[�շG�ۄ9Q��u�nj�y���&���q�
�
�hm:�tJ�����sT �v�=����eD�?�ꘊ2�:�IV��,���_�wޞ,�����Kv��D&D����ԓ}�{5�I d��$@�
������	���F����K5�kb��	19��8��.�� �v��g9���\�S�cM�ۂ�$,��u`���>��,�f�c�ŪTdJ��)��b��Z���%����#{[���n�1�lHj��\��G*H�Xfl��5K�٥��sn��ݷ�I�Mʒ'%�y�_�"d�����B ��hz�P�#ID9p���vi`w��V~�nMn�M _i�@aqD>J^qR\Ո:>�w_zo��[.�}	��rRX�%"PK�~|�ReL�TfO��B{�x��
�̪ ����rL����<�O{�u`}���:)F1TB�NSjC����8^ۮ;9��}�۪��6뷢G��F�D�""rXkŮ��vi`w��^�r�_ 7w���?W���$�E1@}�8W33rI&�37�P���cŮ�r���y?Sn&�I!`]�Ҡ�ɣ�&I����gJ���H`"9RG*��*���K��=H7lA�""'u���w+����7*H����k�>ݚX�mՄ��;�I8�&�$ �Ӓ7:�GXs�Y[]}�kA	�S� }��i��h�S�`4�b�#�|$ҟt��]Q�����X����4S?&x��%�����tA#�)0�z�Bp'�N�98�X��΄���M!�t�5!�)�CQ�m�B���|dHM��Cg�� ls�0@�0�	��}d$7�!)�E(`2Y�07��ā"�ka�Hw���h6��B���D�lƮs��w�??W���  �mm�l     $ �׶�	pkkU�� 
�+�t�m�b3��5��L������Fn��)k��θ.õ��6�;��\6s{Cּ��Q��
+=+��t��lڹ\ڦU���E�Y�A*5��@��8Z�A�l�Bـc��0Ў�Pe�]«ԫ4E��r���kI*V�n-Zzu����N�yԤ���� �L���T<��XR��G��;�6��{V���E�������z�va\�mۛ�a��t9�I���Z�>x�M]R��+[�we��U^�9�\Yۮ�xV�۰�]usrv�C/v)�:ېe�!S]8��h��F��m�R�x7R&����2q�Z2!��O+W)�s)bت��d���]��M�t[��݄y�r�'=�uʊ9JǊ6�5uV]��ڐ�	�<��i�J��<l�T(��M�i6���]���#ud�ۥ�v�6�Z��j�UԱ���;�;p��<��M�].�v=���Q�mqj�*�Z69�m����ŎVj��Vy�\�2��%U�fƃ�݈�,����e����K�ϰ�wbk���9�^���j\�%�b����6�zn����e����ke��Ѳ���&��(�$���l-�̸uR�s������I�3=���#�gv�|�n�6��nL�,X�$s�w�y@�̆���TXm�n�h�h��ͦ���q�K AȪ�ظ�M *����nѢ���d�x�8 y��Ƃ���*ɗ�U��&�t[6�.��gb�;yQ����;a�; =6˘n�!n������l�Ud��-
ey�iĳܽ�K�UU�/0t�[v�U��n�Q��nYMש�c�l��Y��5�C��EҶ ꆴ)E�M����[$#�;Am�κ\ډ�4�ی�Oh�7)E�&����]���2>��$�m�@dV`�N�K���V��U.�v��6Y�p]	��`A���w��w�Ǝ��hC p]"9L"I�4D���|��= ��0d ~@`��©���aF{��Η���kl����LaU�k9��s���h�+7WL�æ%�
b�'m;[��|�\�3'W.xٸ^l��f��:�hKSH�G�<ӱ�O#��	,�"'=��ƻq���W;c'iZWlOGm�̘R�l[��]]n{#li ��E��qѪ��ʶu��n��d4�^�9�Ŏ��ո2���%��dJ�C�mU�k���`��=����;U��{���q�9��/L�i,y��{vs����C�7�������{��>e�r��fa�^c ��Ҁ��)P���]�����?y6���B��)�'��� �v��uH7l_�&Lډ�ₒ��)Өԕ`��`}�5��٥��sn�uR͊*r&9�����[�w_f�w]�5�(��5#v۳K���Xfl�>ך݀ou���)�5*Q��ay��M.��Ӕ��w��Mw�׵����7tnD���.ЛwLM��pU$�@��� �͖��[��|����`m,Tc=Hd�\�q�RI�s���D��*d��C�~�@gu����P�}��&Cw]5p	�4�$��`w}<��������]��Հn論�������HR�Bq+ffO��Ҁ�fҠ�ɠ���ͭw��Zm&�(Q:%4D�`}��V}D���>��@{]��Ю∎��..�����.��wJk��'m�/[ t���O%����l�礮�������^N;�fN���^��ޥ@Q���c�	�'%��lԯ�+�UT�{vt�.�iP���$�;��:��)Bl��MĬ��Ł���X��S�T�$`�� _��Ͼ�ٳ�X�JM��&�m�*�B�S$�.fJ37��wzh�s��۳K���Xͨ�
T�ʰ��@{6������ 6sA՗d1�^#Ox�gfҏd��g[����{'���vd.�;�İݰ��[�����o� <ݱ��Gz@m��5��EPU�$�*D'�>ݚX�mՀff���Ԭ�ƛM��&��"p��v�7u�?D�k��@gu��=�N�T	E��G%��UT���X͞WRM���Ԟ'P�z���c�K�&�I�$�^$�ͯ�h�]�y�c�	�'%��rjV۳K �se�ff��Uʪ׺�J�RM"�I���wCKt݅7[��������h��{����r�b�&���K�;�O��� �͖�ɩX�JM�i6�6�&.�����DD}��6����e�٥��t�e=�`*%F�,36�ͷ2��v�f��ۧ5p�ܧ"rXw&�`}�4�;ܚX~�[��`f{��I
T�N%`y�b3m�w]�=������ԝ�{�ӽ;�?�čl�1��sFlJ�<v��Aq�w>5f�gC��(�b���O�\��ݕks�<��nKqש�{-g�{q�����7<@U��ar��Y�Ö݋m��9*���'\v�e�qƺ;u��	�s�I,�:�$γ�;��������v��y�����S�
��w*�ă�˸��Rx�K�ݬn��<^󮀶6��2��Jʪ�s�__�$R �7NSbu)�Nz�f�I�N����F�v�"k��V�TZ̊6�b�SDNw&���,��4�>ݚXq6�Q*���7 ����L�3���:Pݝ(�s�j���A��TjF1Ȓq��`w6���٥��%�z@��`w�)1!А�
� �0�>��,36Xw*i`f�)7��ۃi�S��ɢ ��hfű�v�=h�,(���.ܜ�y�OX�8�w��<�-���v뱖�ԍ��P0j�"IQ*7!`w6Xfű��g}�zC5��s|U�L "&H����>��7���d$̦L�� 36؀=��tG�2n�J*��*DQ8X͞,��K ������SK �5��i�I��Mp��k\ �ր�l[Ͷ ؝�MGE:|���>�l�?w6���w6x�>�M,����$ICD)FF����l̾�xv�t��=wcY��:냊y�7<q�ۄ�H�c�'NO��mO�ɥ��ri���@w7�����LR��6�ۃ(�s�s&I;���(כ4޵8V�.I��҈�yr"�DH�&d�/6x��y4s0�!�2�y	;R5�#W�A���P਼̓(��=s��bsLÀ�1%$�;��f���(�s��ri`}]2h�tr$�>�ű��ѭ�<k���@n�rn�ru<99gx�Z��]��b��M�o^8ی>��n�=j���nm0�֋��k�����m����}��� �-m6��LTԨ��V�ɥ��W9T�=��@z�N���k2�5͎@RR7J�>F�`�ߥ��r��s6����4�+��H���"I�ܒ�Y?�i@^fҠ>���!�0����T�.�b0���QnM��{�ԙ��#h��s��y�q���>��/1A�����|�ϛ�ӗ\��\� \z�=\�n:�����>b{���b2�*���m���b ��hfų�=!���lǩ�#E*%F�,�����M,��
�\�\���rh��Q��(�I�`g������?U%��ŀw=�`w�$��$�eJ���qX~�̙�@]�k��̚fI�?�N����i��iSR�qX��V�����;��^(�zދǠɓy0�$2�" T`���)Q##!&�$#�z��fb������qt�:`e�z�Z�Vv�<,lv���^s�bְ/e0)pm��wk��v{%��W]s�Ή0�I�vŴ5;Z�+\�ۛcr��^��1λZ��n����Â:�k[v�dS�n[��������a��jznV��.��!"��j��QۗXX�K�a9�n��r��=5���m��i���1q�Ō\�ĉ����8�����LYm��P:
o3Sf-�&nq����g��������{\6�ݭ�ezq��!�8ےR�H�:t��� 7=�����U�޼���A����<Vy�H���"SWUWv��E7(��(��(滿q#wc�8&Ҕ�$h)��{�`fV�@5��ܠ3(�*�aT�6�G"�;ך�{�,�OuXz�K�7��0U�W���J�QI�<�hdSr�yM�2�����OY�D�Et�����K#�m�Ço'���4�7g�8�F�����l=�,�V��Gu Sr�̭r���[Vq2�FF��7�5_k����Y�b�P �1T�ąH�>XD]��ś�z�I=��:�o�n��\H4�4��D(*jTCr+2�J {����g6��@v�(@nEk��U�N�>%"���`}�n�{�A�.d�2���8[�/2���.�33@}�3"��L̚�w��q��������wӚ�JU*$��Cr�R��U�uyxK�@o=��w�S)��N���8ƅ�J��ӃlR�D�D� ������� �wg�9U��=�`n3�t� MA����*�����WDgt��wE�fR��a���#E*%E$V���bw���`�@��	,2���2�	(±#��H�(`�S2���Ѳ�\�b��,ƖL$�	T�Q�`$R(a�ی��D�,V	�f��,@� Kb��$IP����� <3����hV���&�P�B��X� A`�V1����R��M��Nd�H�L�F�/�, ����M`G*G$!!4
�*�0���f0V�b�a��b� �F)`G��Pv�C��Vc	�Q��с�!G@;؇�	��@�H���$B�*��� HB2V$ I$XZ�����Q�&C$�L�fP�c��%	�A� �aa
g)���J�*/� 1V�u�(j(�|� �|��D~_��ъD�X�DE�'�'�lI��"<DЄ�7��F����q�'p���@�'�NK~{�{�7~P���t�3�t�Yw�Q�I��J��L̺�;����@w��v�Cy%Ed|I����˸X���u����v���r���v�;jp�8b��D8�X.� �we�޳5���Ձ����TR�N�N; �w&���;�pf�w�J������4Y�E"jS"m�,�����wn��w]�w�����{N	�J$hh��Aӻ��@d�u ���>���;�0�&#�"$b ��b�"��&�N}˩'>���PcpqIV˻��;��`w��U����X��&�/)Q�PcR����z�=��q���^�t,ogq֛-����C��}|ݢ"�����Dn>�n��,��j�;�۫���`w
{��I�B��	ݠ3"���7{� 2w��cv�Gҏy��^�I�ʕ��3=���ȣ��;�{�@]��z ���2aݥMJ�qʰ����v��K����9�L�{�*-fԸ��^T@:���1@������[�����n��j�H0�_+����LP+�iT�4h�%)��kɘ�UV�j�c�L��r�I[\T�-g����%�8s�[��H�z�R!{uk�l������k�����(�k%��0ۃD����-��`�6�.6Ƌ�z;�{&�N;t1m�7*�m<ʜp�6S7]˺��}���ͅ��<��^}���Ӣ)Q8�<V��QUʺ۵��n��qns��(���x7a�Σ�{ ��q���ƥ��r\�8�ɋ��b�O�� n�\�ór�[�պ��Y�\���w+��8'�Ug�k]�Ɨ���w���/��K�]�nI�7)��;�۫��������Kٱ��iJ$h)���Ҡ>fE {ٓ@{�/�2fnI��A��N��	�1�:�J�1o���;�ɣ�&N�j3^��ݥ@f8�D�8�C�&"b��&fw�ݚ�Fk���Ձ���;�n�):)(JPNK2+\�:>�"7{�'{� f7h]�B�����B*�NJ!����{/m�w!�M�;{y�m;�㓞lt�%�.���t몋��cj�n�cw����!�O|���G���N2!�*��ww���Q:� �0�W9
�L�La�P�R�z�O���s��:�}����X�6�8T���S��� {�dV�G}3��Bv�� �fl�i�L�	8ےX�=�`wsn���UR[���76?S�tԦ�wRw(z� ?}��> {�h�����F�Li�4q)HR��ױR�nIÌ�v��=��;絜��,ݵz%���L�5�nn�%|c���gwe����_���3�� �5y�H�J���!`��r)�@<֡�m���:8������PNKr����m�̜3�e%B E*g<�s��$�ݖu���pEJ���qX{���z��@����%�_t��rMI�ҧ�ʰ;�4�=UKs}>.ؠ>��T�d��݃���@�	u�����Kħ9۞�r��Y^WBy(�d�Ls�%N;K�8Jl>6��o�Kr���B�1��䩩���$���,�7]����XܚXw6X�G���5)�H�4H��6��m�s]�7(n���f����7���M,;�,�Ū��������V�Є��T��0�HD��������z��<���"�58) ���r��mB�� ;���l>��κ^#O�\;�4�9G���Y����qb]�ɷty�q�-��1k�~m��Q� =��@<�g}�DG��րn��/rN�Q��8���u`ori`�l�7��w�s��a�QK�i�:Nj,�| ͫ}Fm =ͨ@lef�J���6
�6�,�͖�������V�{6�X�<���dR]UݠQ���� m� fk�JB0	9��"�����L檺@ݔ�O�t�*u��E�)��j�v���۰�0]8;$�u��Od�]v�vX�#J��.5˶Kq;[�7h�l��g����X�m���[���',Mm�4	�r��۝�[;���MvӖ�[c�h�zEw)]��{Q�����n��c�!�m�k�]���6�݋.��]��9z4.�hK/g͎�*U;�G��r�,�A������{�|��n;��8�0�u;��Z�˞�pO^�����sv�:T��ܩƥ1��4H��ͺ�m� fk��5�r�%E;	�7%XܚX{�,{Y���ٔ��.�w�A2�'P��̔ �~� �5�?G�9����@d1�)q<(x"IO���I�K�;���Ԩ��~���2!��L�����`}��V�&��͖�Vl�?w}��"�O��*�*M�T;A��ۅ8�I�&��q��B�s��q���|>��bb�������`��`|�f��ͺ�2�[�ڢ��6�6�,s]�����}��!!K��@y�� �����`М㎢$m�,��؀�֡�>��Ҁ���t\�򠉘r�34ܚ/;��|ފ �se��՛,�5��M����L�ב@ssFf��~}�>�e*7v��)��M�(bMԦ2D�gt�'�u���1�����n���]��:�q�7��] �v�F�@{P�s���uI�Lp�������~��3{� :u� �v�ݧU1/뿈�T�32�f��ٔ�^E&d��jK�j����)�"P��`T�d�/X��&��H�r���ѠO���ަ>��$�����}�P��iӌ���X~�qy�� o� <�v�xڄ�Ct�`��D@B�1@w�@o(�[��;;�Ձ����՚����)'L��6��oCTu��<1�[ιz�γ�n9S��Ks��㍻u4D'8�R1�,{Y�����X����s��},�z�un1�F�)��@<mB���ӯ� s}h�k���W3����6�$��`yf��]��ɓ;�k6h��T�|Pk$H�MND���`�͖�wF��mLY��@�d�_"��߱��{�Q�4�"��`|�f��jw] ��ٶ�H���H�.�oN�Φ��\l�Z<;e��m�e����򺒧�j��N*D�ȤNKw6��s�� 7����OOu�oQRWiԤȣ�`j��`����Z�v�m��#k+�v����Ӧ���;�ZΥ�@7�B��L9n��	H���ʥ�E�;��]X�5�z���������jF�F�Q37t��ڄ��(u�@yԷJH��ME�HFD$$!R����4���4�4�@�&�Ԓ1i�iO��$$B2��@`�aa���"�Wβ�ɤCbT�@$#0��BA�d�����0�2�2C"h��;�F{.& ��'t���95�lʮ1�����0�gPӀ ;� ��R	��f09â��3�IF���d!0�:����!��0��¥ �2.�)�����%�p�b�@��>~���-W����.�85q�����6$g�Zi���tI�$��:����'2!��!��*f�@�.\���MqL���Ʀ_�	�Rc�cHJ�\�ё48a$c�d;%�q��S�M�?9ƃXIj��Y��[�}jߒl  � j�     $ �f�H��e�� 7,�* �����;���[C���B���nXIND�E[���i��7M������P���+/3�fs�^ڱrsd�[��(����\%�.��mO�h-L�7M�#�V�*�C���avn��V@�ろ$P!�J�l*�K��f�;5�$@���B�����F�v�[r:]�^\n��hW����e�n���;ˎ�r���k[[�Gd+��N�}�,L'l�vgE[cy[>ϴm[v���-�b�l��&�y�<�]H�q\��9��]m��-�k�nE�{�J�ܘF�����T@�d	��-��&C�9�n]�2r
�nT��m�ՒO(�<���p]��;aT��s�!0�f�Pl�bKlI�n��j��pY��'[��L�o��2��$�S��g�j�{q{r���&��x.�a�wm��%:Ɍ���4lmֳ�Vx7gth-���Z�������M��؉��ݔ!��.��`�@��Y(�"���I���J E�g��x0^�ln�>�^\PsqaQ�^G��۵��qv�I.� {V�燌�	�C�tv㝍��Źt�1��m�z�g&��B%vIp�,�ܹ�4�/]J��'ocg��Zt��t�= S�(���4ZP:j�P&��� >���G5UO�i
�����u�^�3�q�Z6M<���b�<�jMaz�"�Q�&yk�\:�W"Sb��96���N�܆ʱ���l��S���4��Wwej7��겓�An��Ɯlg=.�lX�z��RB�=���Ap�;�R�!ԭQ�t�iX6u4��y�Sd�N��9�lYƧS�nѤN�����pkf�"��m�l-�	7a�%nx�}j,�#�]\���c; ��&��ٹřM@;u�4�J����V`�e�*�%\jj�쬶��+�;;gb�<��Ы)s`5A~������=�:�dʦ��]��t��:8��:�/x��P�U�DR�P��@dH�  5��C�N |�L��a�:/�����h�hݶ�2dR�s0q(�^���b�x�c�`��f\y$���ù��W��+��ָۍtB<L��)!�w`t��-�ͦ�)���x�����K��a�v	�%�E���-N��>� ��u��b,�=.�����on�v�G<��v���#66�
I�����m nG.�������p;���\�WFC`�&���뿝�ww�����q!:������xn<�ڻ;��X'�ɸ�oMm��=��ӳ�l�hK-Uq�=�� n�h:�뾏���r� =H�$H�MN%!`fl���ԷHm�@=�b4��\�54Uܓd݈:�����l@n����=mRڄ�J�����,��� 9����:�� nK�&���R�*G*��ɥ��W7}~>�k�vwv���x����E�TĤ���X�����c��wí�v�xCJ�[����jsQB�SL�T�'�n�x�>ַ]��ݺ�s���{^�XU�}#II�����o���4�H�� %����|�&d�(�#v����w������N���M	)��ݺ����:���)�E;
�5Q��s&�f�,���`wwn��m#Y�*jq)3f��^�}����T]�������O���l�O�S���\q�ݮ���nފ��p�
����;�����X��_C�E�̥@e�����fΔo�n��N*C��N'��ݺ�72i`fl���Z�w���i�e6��mJx�J�72t�.�p��I�&O���TZ�Y2f��=FFE�fR�=윉�)ދ���*�A�>��p�ή��6� �ɔwV���w�f]�dQ0�S)�$@yӧHm�@7Z��틤�$��������㮍�ժ����ƫQ�Fv���s��k���,63ηm��g��>?>Cn!�s�\\\c8�4��bX�'=�l�n%�bX��{��Kı;�k�A�<2����e}=�ᓌ�d�,�+�s[/6N���{�7���{�����}t���@H�&"X���~�Mı,K������Kı9�{f�p�,K��Ş��ͥ1rۜ�&�X�%���^�Mı,K�g��4��c�
P2���S/�N2q������_X�%��ú�ͅ����ܗ8�s4��bX�'�ϱ�i7ı,N{�٤�Kı=���I��%��f�=��DM���뜚Mı,K���w�/j��?=ߛ�oq���~��4��bX�'��zi7ı,N����n%�bX�{>Ǳ��Kı;���}�tD�;Jt��n���y�"��%�����v���8K�����m\�3v�-�q�I��%�b{�צ�q,K��}�M&�X�%����{E�Kı9�{f�q,K��;��8���-��q2g�Mı,K���4���X�&"X���c�4��bX�'~��I��%�b{�צ�qVı,O�s���J\������&�q,K��ٽ�4��bX�'=�l�n%��a��������Kı=�߶i7ı,N��mx�IL�J~{�7���{�������&�X�%��w^�Mı,K���i7İ?E9�W߱��KıY�W���$�S3���'8���;�M&�X�%�ᏽ��Ɠ�%�bs�o�cI��%�bs���&�X�%����ib�'���;~�379��<;v$��9Z��y��֜��S��%R�D� �E��uN2t�pu]I�ۅ٧%����F�ìl��vp1��5���m�*�ء��S٘�<ڞA;aW,�Jpf5�.n�hi�{�>�Ş��a�:������ݛ�5�q�q��\���/��x��Gnh�g���h��h
�tJ���ğ��G�nrƚm� tZ�]�wn��{EӐ�GoK&�L�嘞�^�,GN�xx�^��27+x�h�������ͥ1r˜Χ�X�%�����I��%�b}���Mı,K���h�Kı=���I��%�bp�;�L�\���K�c4��bX�'ޙﮓq,K���Mı,K��4��bX�'{�l�n'񊘊q��T<�Μ�!� ���_�d�X���߮�q,K��;�M&�X�X�'{�l�n%�bX�zg��Mĳ��R9KOh���Bm�P��W���(�%��w^�Mı,K���i7ı,O�3�]&�X�*%��g޺O�R9H�#����F�D�&H�HR+Ḗ%�bw���&�X�%��;5��I�Kı9���4��bX�'�Ͻt��bX�'�Ty�E���Ks�{uó�[��{h��ua���&�{a�'�-dֻ{F:���ש9znδ��w�{��X�';3��I��%�b}�k�I��%�b}���B���%�b}��f�q.��ow߿~'�ĺIL�������"X�'��4���CQI�A[@�/:8�Ȝ�b{Y�.�q,K����Mı,K����_�r��G+7K�JR	6�j��4��bX�'9���7ı,O��l�n%�%�b|s>��n%�bX�w���n%�bX����,�&fm)����7I��%�b}��f�q,K�����I��%�b}���I��%�bs����q,K��箽3arb�c9-�1�I��%�bp�}��KıQ��צ�q,K��3�]&�X�%��;�Mı,K��g��L��)���lk׶�.��d3�-�;i�oku�A`��n�0:u{p���&>{�7���{���w^�Mı,K�Ͻt��bX�'��i7ı,NϽt��bX�r��h���I6�(p�W�)�r�Ns>��n*%�b}��f�q,K�����I��%�b}���I��%�b{��7�`��Iq3�L��7I��%�b}��f�q,K�����I��0"SB��(8T#V�n��� a��	D�3BAp�P��D騖'��~�Mı,K��]&�X�%����s�L�4Ͳ����M&�X�
��Þ����bX�'��4��bX�'9�z�7ı,O��l�n%�bX��u��6F�hr*���|r��G)��ߋ�}ı,Ns>��n%�bX�w�٤�Kı8s�ޓq,K��;�$���Al������c�1���M�x��p��ͯg9�lY���cO���������;\P���s��'�,K��s���n%�bX�w�٤�Kı8s�ޓq,K���צ�q,Kļ���g�f�Ҙ�-�st��bX�'��i7�I�=즠�	�{�M!"�'�w�MD�K��箽3arb�c9-��M&�X�%�Þ����bX�'��4��bX�'9�z�7ı,O��l�n%�bX��u��|g,���an3��K���b'=���Mı,K����I��%�b}��f�q,K�{Ԑ	# �P��E5�M�>�O�R9H�#�硾hq6�
/��X�%��g޺Mı,K���4��bX�'�3�]&�X�%��{�M&�X�%���?~��91�&1�K���s���r���g�ܽl�W�ѹ٧v�OC��|n���CGi�_�ߩ��bX���l�n%�bX�pϽt��bX�'��4�},K�Ͽ]+ᓌ�d�.������u.�^eRn%�bX�pϽt��bX�'��4��bX�'9���7ı,O��l������oq������.�S5=Y�Mı,K��^�Mı,K��}t��bX�'��i7ı,O�g�W���#��R9]�//��dMG	q���Kı9���I��%�b}��f�q,K���}��K�,O��zi7ı,K�N�{9���ns���Kı>�}�I��%�b}�>��n%�bX�w���n%�bX��{��Kı=�h�ǌ��8�sY�v�sD�6�n�Ȫ+%�\�`�$z��j�k!��d\�[m,.�x��8JI��d�l�H�ພ�t��b�;���(n7&J_]�����fvf�=7l>�ɤds��PA��]]�z�֞�'�=�#�:.��V�r�4"�|͞���)���:K�F�m���h^^g�p�e���j�k��<n�������=gnsݻww�����>��ܻ�����kq�nv�._,����/od����\kK^w\w
�n.G5�M��w�{��2X��߮�q,K���צ�q,K��3�]�_�b%�bs���I��%�b{��������8)�f�7ı,O��zi7ı,Ns=��n%�bX�w�٤�Kı>�z�>rf�e'li���D�D Lfi7ı,N�>�t��bX�'��i7���LD�L��t��bX�'=�~�Mı,K�w��pZ\��Ř31�f�7ı,O��l�n%�bX�pϽt��bX�'��4��bX�'9���7ı,O`����Jg�m�fnri7ı,O�g޺Mı,K�罿�I�Kı;����n%�bX�w�٤�Kı/y!}>���c���L��.z��=={u�v�M���Kz62v=V��%3S�=ߙ,K���צ�q,K��9�cI��%�b}��f�q,K���}����oq������8�m���f�=ۉbX�'1��Mè�T��D�-�0Q
Kp�
��D1q�V
Ĉ�F�i\���`�@[�'s�l�n%�bX��z�7ı,O��zi7��"X��O_ş�3�aL\�8�q��Kı9�~٤�Kı>�z�7��19�k��n%�bX��}�Mı,K��=��\����Knq�I��%��
"s��~�Mı,K���M&�X�%��s�Ɠq,K�����&�X�%��wX���r��fc33��&�X�%��{�M&�X�%��s�Ɠq,K�����&�X�%����I��%�b~���>�s�p���]n9�Ȗ�nG�d��d�=ѷ�ʩu�jݶ\y�=��������nd5�m��=�Ȗ%�bw��i7ı,O��l�n%�bX�pϽt��bX�'��4��r��G+��}#��H'�PM�|7ı,O��l�n%�bX�pϽt��bX�'��4��bX�'1��M�T,K��{ٹĦq�f�pff�&�q,K�����4��bX�'��4��cף���$Lb� �p�0�Y&J��9a��L �+��f��8H�0Bg������:��a�55������Q�I�-#$�"O��s�eWX�9�,W!Q�	�7�bj�a,&SI��ÀA� EXVԕO� ��GLR�7Q����*i	��CF�`�CY!��	���1�ɼ��F��e�]���^�'���x=D �&t��V��J�ʁT:�N(A@�\�� *�𫇢�a�3X&�X�%����4��bX�'y��fL��pc9�q1���g8�n%�bX�w���n%�bX��;�i7ı,O��l�n%�`�؟s3�Ɠq,K����.ɓ9��.n.pc8��n%�bX��;�i7ı,O��l�n%�bX�s3�Ɠq,K���צ�q,K���߿~33�ns�ֺG/�3�l��8-�rs�vc[���u�Q�q�+�G�A�N�r\M?��X�%��{��&�X�%��3=�i7ı,O��zh7ı,Nc��4��bX�'�3�{��1q1����&�q,K�����4���8���'=�~�Mı,K��cI��%�b}��f�q,K�ﻬ\K��.,��&q���Kı>�u��Kı9�w��n%���b}��f�q,K��&}��Kı;���b�be��A�	�)��'9�!(d��S/�X�%��{��&�X�%��L��I��%�1s�W���-��w9ߦ�q,K��ݾ�i�g9���e�3�&�X�%��{�Mı,K��f�~�O�X�%��{_��q,K��9�cI��%�bs��mŦ��⦊�F��%oGأ��=����ݸ�N.�G��c�6��D�:=h�����,K��&}��Kı>�u��Kı9�w��n%�bX�w�٤���oq��������e�TZ��q,K���צ�p��1Ľ�gI��%�bs���I��%�bs�>��n'�D\T�K��dɜ�c781�fi7ı,K���t��bX�'��i7��C1�����7ı,N{��4��bX�%䝷�'�nf1K��8�s�&�X�b}��f�q,K��&}��Kı>�u��Kı/9�gI��%�b|�>�q��4�"��|r��G)��{�I��%�a������%�bX�����7ı,O��l�n%�bX�aA^
�CJъ��5�3���s`����:��MK�w�&#�����3[���� �b���6�+�9k������m��ֹ�dk�;v;���xdv��e2;��C;�됍�lc�*lqin��dzۛG(���]ɦ1q�ŧm�f�8��qX̶��tq���{87�V�;\Rdvtk<%�{�J s���vY��0�۷D��td�5�.u�b�3Lg8?(�T�>Uξ/�P��
X��ӧ�l�d7]qϵ���ou�v^�{�.\9�����ݸM6;t���Kı=����n%�bX��ﳤ�Kı9��f�q,K���}�|��R9H�#��OR�b�DҀ�ɤ�Kı/9�gI��%�bs���&�X�%����I��%�b}�k�I��%�b}��o4���nfs&Lیg:Mı,K��i7ı,O�g޺Mı���צ�q,Kļ�}�&�X�%���=se3��4�I���n%�g�9�_�]&�X�%������Kı/9�gI��%�bs���&�X�%��d��d�33���fs���st��bX�'���4��bX�!y��:Mı,K��i7ı,O�g޺Mı,K�1=freq:��7:���n����ή{��lQ�q��q2Wm�$���N�U����>{�7��bX��ﳤ�Kı;��f�q,KĿp�����>���%����맿7���{��?�}�w�S��Z�&�X�%��w�4��1�
��^i����O�X���t��bX�'y���7ı,K�w��n%��{���{�}�3��Ѥn�����x�,K�{:Mı,K��}t��c��������7ı,O���O�R9H�#����NRup�T��K�ȋ?w^�t��bX�%�}�:Mı,K��i7ı,K�{:Mı,K����1l�n1��.fn1���Kı/9�gI��%�b{���&�X�%�~��gI��%��-��ze���N2q��=$�/1#�*+q��6vs84�.ֶݷ������i��A�:����>��zҩ#��}����<X�'��l�n%�bX���t��bX�'����? 3蘉bX�����7ı,O`��~����i�[�$�ri7ı,K�{:M���1������n%�bX�����7ı,Os�٤�Oʡ1,Ow%���mM5j��{�7���{����_O��ı,K��t��c,	�R�!�%�������l�n%�bX��;�:Mı,K�w؛v���$أ��{��7�{ݻ��{�~Γq,K���~٤�Kı/�=��7ı,Os=��n%�bX��o�>����8K����{��7��=��f�q,K��p����Kı=���I��%�b^s�Γq,K�w�����~���쮣�֊��v����n8ۣg7�����ns�H���V�\��sfqq�i�Kı/:~��&�X�%��g��Mı,K��t��bX�'��l�n%�bX��u,�qsH\��fs)��I��%�b{�ﮓp�(�1,K���t��bX�'��_��q,KĿp����Oʸ���'_�����`Rش,|�~oq����{�~Γq,K��;�M&�X��"b%�O߳��Kı?w>�t��bX�e�{Z�&&yy��.�4�ᓌ��bb'����q,Kļ���t��bX�'����7İ:���\@��"H�#h<p��Pj���"T2ר�G�Dǳ�gI��%�bs{�\��9�in�ɤ�Kı/�=��7ı,?*��u��I�Kı/{���n%�bX��u��Kı>���)�&r�F�]ѩ��Oj�;nz9��?��=s����;nݝ�ju�����=ߩ�,K�s��I��%�b^s�Γq,K��;�M&�X�%��3=�i7�r���o��	RA�Q�H���ʱ,K��t��bX�'��zi7ı,O���cI��%�b{�ﮓq�r��G)`h��="iRjQ�_+�,K��;�M&�X�%��3=�i7��QH�����~�Mı,K�oM2�d�'8��I�}�O*�T��3I��%�b}��{Mı,K��}t��bX�%�;��7İ?�vo�S/�N2q�����:H�	�g�&f3�&�X�%��g��Mı,K�\w���'�,K���k��n%�bX�s3�Ɠq,KĠ�I}��{������O�ݬ�U]ˑJE�u#i�Zv����M\�D��	��4�:�c�V��D�K��ͣ���ZC;���N#"1^U��Wo[�7N,1�7n����8��6�;�5��;�f�x$f�n���6_o�������rW�KCuVn��"�6���<��V'�=p�nG'g� �q[nwX�Nn%F/lX��\�6LX�F/;�&l���{���w~�����UY�&GK6��ȹ��r�;ַ;��;���78�뗕��=��/C�� �K�K�-8��N2~���cq,K��;�M&�X�%��3=�h?�g�1ı?w>�t��bX�'���I�g��s&Lیg:Mı,K��4���D�b&"X��g���n%�bX���~�Mı,K��t��bX�'pN��KI��4���1��&�X�%��3=�i7ı,Os=��n%�bX��ﳤ�Kı=���I�����ow��q��`�f�M=1�7ı,Os=��n%�bX��ﳤ�Kı=���I��%�؟pϼ����G)�r�Ox�r�mD�pR]&�X�%�y��:Mı,K��4��bX�'�3�]&�X�%��g�W���#��R9K1h�ĨƔ����]������:��73`]{;���p��b�i�g�T!�n$���{��7������I��%�b}�>��n%�bX��{�Mı,K��t��bX�=����}���R�%o����7���{��z�7����uQ,L�ޓq,KĽ�}�&�X�%��w^�M��$��N2���"D'��Ď��f�7ı,O����7ı,K�w��n%���b{�צ�q,K���}��Kı9�x�Ŗb�\b���ی�7ĳ���Lw���&�X�%������Kı>�z�7İ? LD��~�I��%�bs��o��inq�2d͸�s��Kı=���I��%�b}�>��n%�bX��}�&�X�%�y��:Mı,K� s������v�9�S��i�5��s���ę��>�����0��n�<W�{�����\���vI�fi>�bX�':g���Kı=��zMı,K��tB�H׳}9VW(+������q�$�G#��В	"w�w)���bX��ﳤ�Kı=���I��%�b}��{M���{��7�����}��-��RmW��bX�%���t��bX�'��zi7�ʿEH�����nCE����g��&�X�%��3�]&�X�4�R��y�zDҤ9JI|��R9HK��4��bX�'��ﱤ�Kı=���I��%��@H�����ޚe���N2q��OC��"bb\���i7ı,O���cI��%�a�c�����%�bX�����7ı,O��zi7ı,N㽞3��.
g�i�v�ƽ���#�W`ܥ�ηy���Zϳ�<���c�vƤ��{Cg�������{��'9���7ı,K�;��7ı,O��zi7ı,O���cI��%9H�k�W�E�q_+㔎U�b_��gI���bX�'���4��bX�'��ﱤ�Kı9���I��3%�N2���LD��bT��x��t��bX�';�_��q,K�����4��bX�'9���7ı,K�;��7ı,N����iq�����&�X� �X�s3�Ɠq,K��3�]&�X�%�y��:Mı,���DJ����2o�����W�)�r���=���E$�#��Ɠq,K��3�]&�X�%�y��:Mı,K�{^�Mı,K�d݊e���N2q��P�%L;�A2�<�����ch�r�8�p�k��z�nںع獗�k\�j���|�~oq����s��t��bX�'���4��bX�'������$S蘉bX��}��7�N2q��h�:e��9�a�f�|1bX�'���4��bX�'������Kı9���I��%�b_��gI��7���{���_C��k���j��w�Kı>�g}�&�X�%��g��MıD,K���:Mı,K�{^�Mı,K��.i�30g��q��Kı9���I��%�b_��gI��%�b}�k�I��%�b}̛�|��R9H�#��}K��P��qK�f�7ı,K�;��7ı,O��zi7ı,O���cI��%�bs�ﮓq,K��ؖH��"p�;R�Ph�B ť(I$"�f$RX�� &�Q�ʬ$! F��-�	�2e��'���Ơ��FR#�2��7��0�v�)(�H�#�饈C	������M"�p��~h4R/��0g�1Ar
� ��� `0�7��6TA�� � sl�M�\AS �W\��CH�.a�	p��`8����5�	�f�0�L�l(Dr����8`H��iSi��(m�!�����PiPr�pL@ٷ�czXȥۥ(}X�a�I�dx�2�eL�m"��aC��ba�0a�c�Au$�t��>JJ�T���2��	6<�3332 � -� �� �-��[�#�m���m�R������YA�C��s-[�ѝ8�YC�"\R��E��;W(�N;\�N{kԈ��k�3�NجSF��"��< ���@�r�s���=�i3�vo3�#�3���;D4�9U��
X�!vC���@[J�1F\��#�T�T%�Zn�tT���L�Y^��E�6-˪�.qc'Sr�띌ǯ\d�&��w��0K��p\U�<��ㅌ�M�d�o�mmv����;�VNՒϮ��q���r�D5��فi����gK�s��i�Ki��� ;tv왑�>�G[\���{�eq�:x�ֲ�3j�/�v���>k�υ���o\��Iq�s��֧�mA��v�5#�����QPz�h�@����÷m�S��Q@bɴ̻�GUY̵�����L�OOM�˲����A�y@�һp;-��m)�t9�+h�uO��l�v�^֟.�s����t+��ɶr�B�1��yq�gh����fg��kZ�I؜�<=Uӊ]����vA�st����rs�9����"6��"Ƈf�:vgigF��x��삻1Hn:��@�3��ڄ�D�Ú�vvej!��nZ��V9۱�ᐏ�u�e�Va�6�Yl��W�Yr��&+`'H�V�m�  ��M�`����2O8f�5m�*��<v����� J��*����\`�����_>|�x��74���Mg4�>Я!�V�pq�l�/+T�f,����uZA2�wvP9֫=����S���3��z�ˡ�\�ݗu��A�f�����.��6�5�&Ik�d{T�M��5�*��T�*���^m�eAd6 ْ싶�M�h���mx��W�oe���1��ط,��l7���		�������ᶱ�ӳ��ئ��@R�(]��T���@^�5G��*ki0��\t�Ԑ�	����8��1������dF4(��S���a���� /D@r��ʕ�Wr�TW>��n�E$�@T�Jm
���╎�6Y�����(�Kq&tL�Kaؐ1��c�t޺
�nГ;m%�$fET�n��M�Վ���Ŏ<gУ�m��Z$��S��۱7�������m�k��b�[�X��F�\�ήz"�6xwf��-뉧K��jK��=��sn�'$i%�q��Nƅl����b�4���a[w/<$���rĺ䰦R^�̗�}�=	�D:�D2�LA+�y`�s�g>n��獹}l�W�ѹ�F����_���M�z������w���oq�������n%�bX�s3�Ɠq,K��3�]&�X�%�~�}�&�X�%��I;���I¢M�&�W�)�r���C}�&�X�%��g��Mı,K���:Mı,K�{�4��� 1�{�^�t.���e�?=ߛ�oq��s��I��%�b_��gI��?� �"b';���&�X�%���{�4����oq����};SvE�|Mı,K��{:Mı,K�{�4��bX�'9��cI��%�'9���7ı,K�;/�{9���c%��3�&�X�%��=�Mı,K��ﱤ�Kı9���I��%�b_��4�ᓌ�d�-��ؒT���w^������0>\�X|���۰qb�h�G������p)ն��Λ�{�7���{����m�cI��%�bs�ﮓq,KĿs�Γq,K�����&�X�%��z�6H�@I
a<�1L�8��N2�g��M�?��]�
�~��/O��MD�.=���7ı,O߻�f�q,K��3;�i7�8����}~���w.�p$L|�~oq���b^w���7ı,O��l�n%�bX��g}�&�X�%��g��Mı,�������䣒n��%_=ߛ�oq?�C9�߾4��bX�'1;���n%�bX��{��K�� �D����/�N2q��� ��.:x�K�A394��bX�'؜ﳤ�Kı9���I��%�b_��gI��%�b}�{f�q,K��=���6�q�[�2�u;��1��Ȣ���=]{s[c�S��f:62lmӦ"�	Q��ߓ�g��u��g��Mı,K��{:Mı,K�{�4���LD�,N�w߳��K=�����~����+�dY�G�w��,K���:M�� ��LD�9�߶i7ı,Kþ��&�X�%��g����C�����p���/:	D��I��%�bs��l�n%�bX���t��cP�D��A�抪l�>�����I��%�b^�����Kı>}�b�̓%���&LL�&�q,K,K���:Mı,K��}t��bX�%���t��bX�'���i77���{�����kɘ9�����bX�'9���7ı,?�;��t�D�,K���f�q,Kļ9�gI��%�bs�����K�!q2�:�U���6p�����;z=�p]���Enɗ����/�|MƋ�\	=ߛ�oq���s�Γq,K�����&�X�%�xs�Γq,K��3�]&�X�%����7N8SQʁ"nI|��R9H�#����i7��LD�/;=�:Mı,K����&�X�%�~罝&�X�%��I;���9sn131s�I��%�b_�;��7ı,K�w��n%�)bX��{��n%�bX�s�٤�K7��������2��ٯ����"X�%�;��7ı,K�=��7ı,O��l�n%�`\G�����Ļ�g���Kı;��b칸�n1�\c8���t��bX�%�=��7ı,UC�{�4��l��g��$�;��@�f�$�N��$T$T�%!��A���㱮��l�nv7q�5�n4/:�8����P��(��@{P�s�:@�� <�h��Z��JI�)�ʰ5f��*���˼�(ۻ4z�s333;��#�Мhq&9�����>��gꪪ�^��Ձ�t�;�SZ�)BR�jnf�@m�������,�fƩ�5�$��6���d̛"�l|�N��^M���ou�~��o� 9&��N���1-T�U��<�z��r�=s�g�n�����[�q�]��n9z��ݸ��ܽ�-p����K٧Ns����\�י2!�u�Żofr.�N�m�v�ms����"�%�j���nN��[C��Ǆ�ۆ7R�s�ɧ��ìq;��k�f�ڵk��P������7�\���<�'/]3��nѭv�=�`��6���v�� ���I���=���u�;�߇�?����'=bX�b{���B{Y�S����n�r�^U�\x��-��F����@c�b ��h�� 6@��jH�`�#���ɥ�r��ꪦh��ޚs��o�y��^�P<���q&�q8X}��wv�����vw&��V%�z�hT����fR�-��"��\�A�ܙ3D_oM���U�)&�d��`b�f�����]�7P����(��&jJ�%F{s8M��'�.<�u�p���n�Z��Ssc�x��lB��h��8��`wri`n;@n6������[�Bˉ.%�Լ�@e��K�l͉�&K�7��T�W�;3&�ۓcT� �r�I3Wv��v��F�G艖���;_]����I%'"�$�a��^y[�`6� �]�<ݱ �l�������&�Pw8P��'�͟����`j�f� ��0KeF�EPN;y�nV�˜�ûmO�O����t2Wm����X���q��q8X�6Xn�,]��`fd��+��z�lT	ݠ<ݱ �#] 7v؀k��JxV�$Ԍ��!`j�f�3&��9ʆ� 슍 � ��)�0AV��JE)3�>I�%�K̛$�ߦ�۹���,0`���vfM,{�,�f����V������BR%$�E �k��jr5�wm�{{���-e�e�g�n�l�FzTU9u۶�s6�ݽ��w3�{nqv;hi�2=r1[8��@y�� �#] 7v������-���"L�;�)!�J��+Y$�#n�@�ր�mB��7WWv�`�#����K ����ݺ�5ef�4�v������p��*��'}�٠=���{W�@��
D$�@�('��ֽ5$�>���^q6�	I`}��V���`fd��7�����ʨ=K��j4�t�]C��D��8�n��d��7oSLi��qָ�(%��*@$Ԍ���|�V���4��l�>�۫waH��C��t���b y��m�@9��K���#w�ɰ)ԈD����,پ��jr5�wm�=�u2TՁUuvM��͵9��Z�|��},@n��B�e1:�RU�������P�v��6����G�w��ZU)P!/{�}�3����9ɚem�z���d�����c;cîd��+�<�i�fNw%h��ۥk"K�H,���`�Z�!�e'iCWf3��/C�hr�nĭ���ƚG�B�l �����	�74�]�":�Ӝ�Iʩ��t\I˭���|��wk�wd����c'�z3c�nWO��8.E���Lv�^N����b�������Lk�&,����8N��6��]R�3f&1�"[u[أ��y-��Y�(���O�t�wǙ�Gmۛ�Q�pJGm��u#�ǿ��<�hcjr5�X�*&�&��J��&�P�v��6� �#] 3�5X}��S��ڤH�9,��t�s�����P�v��2�왚���)�ʰ��畾vc�+ ���.���=��u#86%N78�mk����j9�Pޡ�]�&��M�=s�� p�cy�ރz9:�������.۞��H���]X3T 6r6l��(k�u2TL��L̄33@}�*�3|�d�$&	�� ��V �� �p��p��ݝ�5$�q�� ����9T���T(P��6A�N��@fV�@5��� wtJGm�rԎ��^j��l�>��,]��`en�NRnD7�w(�@{� �#] 3+\��X*Z�64���aB�a��&��Nl��wv \,��C�\v���͙S��5v��;bg#] 3+\�=v�����z�t ��$,]��`w�5Xۛ,��K1�k���E8�8��� �se�:��>���
$!�\��8@p�a��LwB��c�c��$�h`��l.;�`̑��!!	��I����i'�I��0�� N��z8J&���C������rmS�к�����S��5v�l��.t&F��!J!ݙ �,@�S�T����/Óc��J	�ȳ}����Ռ`�77�
�#s}ڙ�S}r���x3�d�?�� $GG0��k���>�4�2g9M�I8)��b��CC�:R8xh��Z�C����lIa`��	�Ӏ�+�8*�4"��"d`&�t&2���".�/E� dxcOUr	�G`�Q��^c�k:��n�s]���i�)ԈD���8�<�}���gJ���(5&I'��נ=�;0�RF������4�1v�]�޼�`nl�>�k6GE%(!1S�:�vy�z.�m\<D9ۇ�x�ݖ��k]��[*HpN&���p�1v�]�޼�`nl�+��s�Ł����q��v]E� 3+\�=v��;bg#]_�#k=䭊'r"8�R; �����4�1v�]����`�ҧ���� �NK�������vWs]��F���C�ংP1�0+'f�d�ޝ��ho-���	�%A7bg#] 2s] =v��;b�������]�u��t���k�H䳜�)�c-�;{mk>�8�1�ŹݍgOS��M̕uu�6u� =v��;g}�s������N�E)BjF��l�2w={��{Y�@y�y��;�ܝ�w#�1��)$�;��Ձ������ ����t`���'Pi�â""z�Rg_R y��w�9��@{�	H� rԎ���k���h��J���Rd0����w{�����Y"��<;bHΘ�h/I����t==(q/,g�5�-3��x���cv2']�4��kO�<�qge��p1c���mu�;w7eѓ�� \�r���Î��g���7Y����? ��7l�٥���{���=��M�.����Ț���Y��=8����Y��ۊ�LYw/G����a'=v ŋ�kv�����4�rG���Z������w󻻽�����~k�{u���g;^�+V"��n����.�����ś�����{�Ħ�F����������mB�F�@d�@�ҧ���� ���ݺ��T��k6({͊ �/&�S$�yh�Z5���S#�`j��;����>��`}�۫1�-$g�A�N;��� y���?DK��Ԁm�*@��*R�ԍ�`nl�>��Ձ�������[n�C)�n��R�.��=�7�۬q�ɻr�������-=�烣1��Q9�&��I`}�۫k5�]�v����tc[
�)	��MI9~9�hO�����D�#��G����Ԁ3�Z�ڄ�HKbR8�H�u#�:����͖�ݺ�1v�]���Vڈn4�J8�R4���� 6r5�'5� �i�*z8�\R�"rXwv���k��?���ؠ��hI$���lI*H����W�
�m�Ƭ�rs�x���C�v�;8�C�M��� ."��'B�)���Y[�`d�@z��v���]��A_I��vWs]�}�����4�1v�]��F��S@RuJP������MI7�s٩�t`m� ~��`Dx��2 8����4���`}����"N8�*)%��;bg#] 2s] =v���S��q���8X�Y����پ�����Xwf���OQ��$��#�������o`�����qé��#�L�=�8(JGJ4G�G`uw5�ۛ,��Kk5���B��i���H��@z��v��F�@d�]!]�ZT��QP)Q�9,秋k5�]�v����Ҷq�IЂ8H����F�@d�@z��}�zFH��1H	�(�!X���"��o?jjI�1;;�f !�e�aD����P��}�>����(L�כ��q<<)�vxׁ��yw�:s��;N޸��p�.�s[&9φr���TJR7���Xwf�.�k�r�A�7�����QH��&��I`}ݚX�Y����k��6_�_��<�����N"��A��V�P^E̙������Ҁ�Bw����D�%H��� �se��viaꥯ+|����@n4�AG%��� ��h��o.<��Ԁ��u@��	 L��d�C�F)"I��� �+r�mh��ʫ�JWn��*�<i�8�q{:��1X�Is�hF�g�8����L&ͬ���=���v�b���:�DqQN��p]G�8��m��=��˰����|�|ƥ]�u!���Ob��k��'���4�u:lu[�k*�^9�\�H�ht�՝�B��ؔ�e�]�E��x3���*�m�B�q\m�cq��Wn�3�c%��Qؠq<��W���ǝ��gh��!��鮇�*�[��q�lAnv7x2V�7�[k.P��GlH5��nd�`b�f�����>��`}�6q�IЂ8Jd��1v�]���� ��h��/�#tq�t}J�*H�t�1g���͖W8�n���Օ�vz���)�ED�5#����@f�P����HN�H=j�p��!�#���f�X���y^���������`~�Uy�z5Qz�`�mlG��d:�&�u���ݍ�n�(��r���mR�*�>4�)	�$r�W���n������f�X뤳D�qĳ������q�&�;�k@�����B$G�X �!��4 �d��$��5��(f�*���6Р7$rprH������;�۪9�3���ؠ<�� ���uC��	�����@fkP���n��n�9���G�=I:G	LRU����v��N7H�j͉r��j&k�vkO�8�q�h��h�h�#�pq����]���9v5�}���:��y;>�g�����Ԁ�����B'!�@nS�L�o�	BjG#�:����6����n����`}���R�F�C#�@{ה��Y�G�3bnfvV��C!� aO�. w�P�sw߱�'�w�;�����N"��A�*���n�Ӎ�'����ބ�Dˎ��ģQ8IR;���`uwu��mՁ���v�����/JQ�)'$Go7[��=��������b�:+�גz8������e)9*I(M)@տ�;�ͺ�:�[���wu�}�c)�Ҋ�J�(� 35�_��M���@d�u 2q�@w
�2���$���������[�N7H�j�c�.��b���x�Q1A��ɹ��;�����=��TMs*X~
�(&Z�@2�*���&L�w�%w���]"�%SwWt������B'!�@fSs`wrRTQ�����(��NQB���ep�뷶�أ�v��*sY���Xf��奒����cj9�2��N6��68�ӈ�'������S'r�7^���ؠ=��U��d�[��jr�4�QԎ��~�:����v����n�6��)9$���MIzfd���m*�����ϼ���k)�iE@�Q�`w��Vk+�[��3#I��\P�&I�33��EW�("��dEV��*��U�  ����A_��"��(�b�E��DXP�0DX �b�E��B$Q "DX �`�E�!E��EB"A`�`1DX0DX�b0DX!E�$Q
� �E���`�DX��DX�DX�bQ)E�AP�QDXAbEb$P�DXAdP!E�E� T DX�*�"E`��DX*�T �$D��
P��DXE���T �P�DX�T �A`����"��pEW���*�AUj"��U�  ���U�"��@A_���H ��� ����PVI��`�u� �v` �����^���    
       4$�  � �-�  � ��  �D@	{�J�$TѕP)*$ �!*%PRT�QUT���HR��P[j�(U
Q��@*���     a�� �P
������^�M4�gE40N�0�wX�x 0	9{u����p[�}7�}����a�  �pro0|ך���=�r76�';�{�;�;��C\ڜ�=��N�t� �yғ�4`44m��X�-�'�u�ö9����6����|�s��{:���%�� <�o �Ǡs�\ W6N�z��g�_oZ���O�u��޳����ַv�|Y}�(��|�9q�����p |<��� @� sŇ^����$>��px�{�y�+�}��A�oO!���g��s�>�F�|O�na� �'��s���m��ٟ �a��`rw2��-�}���v>#u��u�� ���>���� ^��c-���u�C�� �=(}�����9{M��툾��]g���À �vOw�>��ml��ϥ��,�����C{�w ُ�\���7�� ��@   PQl}�֙R_ �އ�-:�{��t�Ǡ�G��\���M� Y��ΰS��x(w�y�J� 
wY�  )wp:QK�t��{��z^t��u� D
� �4�pt'Oe4۸�S�70 ��Δ
9�S�  ��қjRT� 4 ���T�S&  '�T�I���T @���EOڒ��@ i��I'��UC#��E�)$&@4<Sy\������V��s?�?�ZI%R�9��_�B�*�?�U�""*��
����*���PX�������%1�R�Y��e2��C�H)�*i� 0�F%@`�0da�4�� �6 N!�B�%����2�>9�ˡ�6J�.U�V|\����`�q��BՄd���϶l���3��f<XY�ɠ�� �6In����/M�F�F9HP�%~Zd�	��x*��JHCCY�X�. � ��2����.X�D��!H`%���c��� �
��e��vCF40a:%�_r6l��p��9��@�������r�e�����\k3���
��8����(E �D"p����1�R�dHX��C A��F�9�}�w��DƵ�]��;��(� �
�pH�Q��X6B2I!"�!dI%��d�X�#F�Xaa,�@�&y���YCD�5�JVR��D�0�>��_m��BF��\YS�؄NI+��ѹ	��}��4�@��"�J�c�W0ѓ�%1"�(���
Iq5��_���a�ą�r�$3���8�6gf��jks���ɷpɇS�b��)�i
�H��*J��lhFԸΚgA��S��8CYL3�/DP6��x/B$H2H$&�d#C	
B�p�nK�`щRd��j8	v�,�
�������P�D,% BH2@Jh�+��[af����D!��)�I��/1�����w���BF�N�т�0h�	�I�7���ۢ�HA(P܄H]�1!���,�4H�22�
`�Ð�v�!X[���\BM���F0�#P㵋L(wٸ��i�^zB�}�W��zXW-I1���gZ>����;��E>tB�_�k��mJ��.��Ą(�������X��"� 5�y��qd1��7Nh�&�dF,��l���#$	$a�Ɯ�Ѽ�N��e)��P���ri�$�E�*�A�HK��Ē"�k��Fm�jsY�)��#p�n�ְ�&ͱ�!dM�J��،�T�_���A�$�Ѩ��sD8�HXYh!Y��9&K�@�Hb��B8R@�Ŷ�3&�*p�B$P�3s��s��9�J��.P��+5��Xd��uO��q��wlxD+�WVLc�ֈc2˖�I�8��>��JO����0�Ė���I�+ȟa��du�)�A�@��6`�saXSD`i�$�p�#H0�e�P�0d X0D�)�Hi
�ă9��N�� ����)-�:F'Ƙ�F�k���F��6©!0�ZB�_}� ҄��f$IRO��>��8���%�(F�T�[4�sZn�bp�
I+��HU�u�9ᢨB�"F
b���@�i	X3
�i��͆l�7�3�L�����cL1�����K3�b�{Ϸ�$&1����^K�ı���`@��y��f:�l�HlK��A�őA`Mk{8p6D��'e����^�&Q`��@L0X,R�@�HB,1��KA�D
$"��Hš�*�>���l�ڽq�?}���M�T����$b�RB.>ņZcḂH��i�4>��.�c:sd�ƒadp��X�0B,$$# a�H�
�$H�WE+��<#\H9�MR����0��&��^h����h��HP�V��ae ��\4�+��Jx�*|�+��d4m��cB���2�i$6h�k:���8�`���q�Ipe%B9�H\d��3��Rl�.9XP!B$![!C�Xa��(�VB[�k��ܡ�9�`M�L|d������1����\E�4t[��Ln��%X�I��o���d+-��:�H[b�9����S�Nl�
a�X�s �+�����Ѽ�X�>�7�����1��C�	@�HX�"%�t͹f���
`ΥK��m�%�����;&Q�Ș����K�.w�$��hɢe��.
��P5��t��$!����)G+�o�*�(\9u�����t��.�>��^gp�&�FBI1�o���01�2�.�]sVcl�qS:Fyd0�4$(c7X���XӳT�
�]�b���V�8a�˟��e�)����eΌl��B��B3'Bxf��[�Xt lwK	3�e��C�3n-��ѐ�v$�D"E0RU�pĤ��.0LsY�LwRh։��0�Rl��B9����7�1>?���\�%��Y���I��X��b�Ŕ)���x�8!L��.]��B�����%���J�K�Rb�&#�$
�� 
T	�(��d���Q�Cw:�1�"Tq����@�B��E"2B��J&Ȭ�:M��[C���L�u[����D��dѽ'��ˊI�h�	�I�se�_���,�gӄ��o\�p8k�\�>I��I $�O����K����HR`�5�}~66����[��7�c�mapQ�p�7�Kf-s~�u��~�k	s7�u�>9+�Ζ��;q�/h�)�����}�_�l�J��V��n���}��4 ~�7��e1ș���F�]���L��`��.sl��}���G���e## H�1`FHF#�,�L#)"G	�$�b�����bSS30`��>�1�|˩	s#�%��b���;ɸ�F	@�Q>%`I�m"Z�Y��,���
B�!�):#�s�lD"@���F�Wp���$bB�bG�h)0Ē�#\G8����I��?n[����aX�9 a\F� @�
C	��1�����	r��>B$��i��>v��_w��}���??!��)����i�J�(dMD���Tj��J��!�|l���۪��FBB�
�]�Y�;!��F��*b��e��F5"�Y!H[�d��5L�%��C�R��-HR���B��In	!h�s����тH0�Q�@*E&2`&.O��y*�*B�����#�i\�]�$�nJ����9���*YE����}>��=���7i���cx���ϭ�\B̤)�%��rm�!��;c����Hۣ&�A3��|��0�!#��_l�����K�d�&51��9HQ�d�*@Ԯ!%�n1��
B�ӳ,�δ0�сȶ������2Fh%�.��K��9%Mm%n�.e%ѐ�$Y�\�!pe��F�.w3��Y�r}�����}�����Vc,�@��V�]��!HY��Fs]&>�Fc$��4k:��Ʒ�׹�t���)��AR�gV���ۼ�����/�+�Z��ӡ�b�_o���ڣ�EPs(�s>u��	�
+)��	�c�HζT�Ra+�I83R�2B�r��͚~�HR�#}]j�!	�%�iӆF�s��F�X;k��K��[�\|nSTq����~�R}B���^0���.8g��]c;IZ*��~��O�x\�4��9wʻԛ�rh�%�rt8���?�[��?�<m�@"���a2:��>�m��y�F���3�e0&�WXd5
�έ�s>&I�8���W�m>Wlny���6�	�R@�7���d�\s ���6VR��#q��ƾvk䔗"Ÿεi�]f������Ԥc�1�V.M\�_���>�������!A RѺ"M��+	��a���5]�!`Z$�p@'Ы[s����[hj���$�B�K�w�4�������!JU���K��A��� Ƥ��|�a���d�X�A3vo��N`����,�!×��dJ�:BB�b��H� "�IL>����$ D4�0�M`�GR!
s��BBCL۴�##%�ey��HSֵ��B84�a��#B1�3�.�0S=��aN�0�)��L42�,�K�N�0l��wY�~0e�H5^13�L����U˧�.��ۮ�̦�xVbT���8�$�3�7G�$a����g3�W�M�����N�S�G7�A�H[��b�Z��HT�oD�VK��!a�k�0�k�pD�6��5�*Bo::���d��
T�I���,L�I,R��m^�a�u��Аb����X֘Ί|�L�ѹLA�艞��X`H1bĉ$ B4UG-.�Rp[�p��|֙�(�d���)��0�P���J�N2j8�(`cLe(II
Q���&����^6�lgDi���^������>o�  l  �    -�8                                  m�@�                    I $                                  m�      ��  ��    [�     :p��ڶm:I*�sU�u�x�n��Cb�JTGQ j�P �kj(��2�Ji�&��9��&�X�z��3��]⃴m63�I=,�	�wz�㱂lj:��M�"ʂ�l�����We�q�c�Y�)%r)��kj��0u�2��F.y[�3m[<�����&�nQ�MTy�omT<����s�'�@mu� 6�6��۴��a��%���m�[BM�� !m��Mm�@��-b4�WU*�nWn����U1CU�\쪭Ĩ**�uUm�M����p��6ؐ �mH �` �[[kn$8���Ӏ��it��M)���X��ڡ�= jGm��ݶ��,�+I��m[Rvٖ����ɶ�����>K��ې[Cm���jٶ�H  p�^�m�-�l� ��V]��b�F�V�]��1U�"j����@T������|��n�6�Ŧ�n��tu�Ͷt��D�d�� 6�Ӷ]7`� l�$�-�-�[D��m��XBܛn]b����i������UgNÜ:A�R�m�`���l�Y2@ᶓ;��]��� P�,誕�iU�V��l��PÔU}U^��	"u��gMݶ sm�idn ��lK&�1.]jY�l�py���њͶ�u�Wf�.4�[\��;O<�ɜ�;\/3�����"�b7@i�t�K$�N��m��$�Gq����Vt�ca�] �1�&��6a[WL��a6�b�"�uO$�-�aX�[UJ�A�@K�v�V�G��m�M��nL O%ĳF5�V
�3��4Q�n�^Z����ܑ+Ϥ�m��3�6������
WpS�.(�R�^;g�9�Z7�y�:{)�v��c�F�����	`}��ג�.홌'E�T�X
�X#������ú�,WHl5T�].��e����b�l��2�*V�3�!��C�!��
���@ְ��K/ ��d�ݥ|���xOT���6��Ekj:�6� 6�mF�t�I�@[��L��v���E�P*��&  (
��T�R �qz� m�Cm��$ %�.g�l�K�I�t�G8��W
�{5U��u���n�,��ʛ��&;N�e1���V[��ZW7�mb�y��;�Kvn�����V�Um"� ݢ�������d�1���
�@5�I��q�n�*�m\��:tU���k��u�-�6q�l[Ie 6�	�ԃ[:1�v� Z��e�S�)��u��] ��[[gS��F�� �
W���iV����  �qI*A��)U\�.�5*��[-UJ�����V0:
U�q��l��Q�uR�@K�������@%e�w*�[UMک��65+ u;v�Ҽ�;-UP
^�&��-��ͻcn��
�U��!����J��P�V��l�byx�<�����j�kR`  �5ð3k�N�.�	yi��/=d�j�hZ�gB�� ���Z۶$7*��F�;5\u��\�P [cy��-�?_|Y~��UR����q��j_Zm�kr�rb��X�msj�e��Ŵ*��R�˽v(�m��vUZ��}��KvZ�z�/��|�WgeWj��Y���l���8�<�Svb�]��ʃh�N4��ӆK�-�n��쫱��S�`j��sa�_o��U��*]�vmv
nҼKǲ�wI��A�i:�*k�i�I�jŭ������1v��j�)���	e<�NC�p�W%��T�s�^�o�����of�hM�oyk�յ9�˴.݇�s���{�2b{e2Uúm��QR��4qī���Bz�j����0/;Y�k��[0\hn����Uv��m(<�Vy2hն�)��[R��VQr���]�k,���UU*q��@]m#n!&`����W�Z��������.�g��2�mζ�D�&��/^�[F��[Am� ;k�k'`�A���d��glն��7e�f��[b�2	A�� I��L�5sJ���6[�HIm[\ [@�[^�U[��R쫅��VYZ�����-mU�1�ʫ�+UV�m�I 8[N�٫I��`$�m���	Um�� 	bռ�Nbk�`����K� -� -���,�m�տ9����m��UWT/,ݗd�e���UJ�m@Ep�-l�U]�kcK�I+`s 3���l6�j�櫋n�I߯�>'Y�b@   �q� ����ٕ`���U�U����T<�7G��U��[�״� V�Z�n���I`x�
ڀ�ͳ�l�{�mRI�N�0	��m��I��r��Uv6��u��"�Nٖ���k��(��2���yj�n�c��\;�^~i:m�(�^�ض��[+�"�cg� Ճ� r�smȓ�v�$��4s8�a�13v�9h��G^��k�ڔ�G\k+�8�������ᑚ�^xwemTv�<�Mtn����7]�d��ys��4IEt�-�$�λV��J�UC��n��:4&xV��;AW��X�@�۰ݳi0H mf���h�H6mٖ��3��UUR���* +���)��`�l&T��V�t��,qH�VS�3:��B�e�8�3R��Zm�sm�D�Ĝ�ZݕeZ�2ݔ/��u�6Ă�(�D� ��]b^�U8\=�(�J���`�,��zP;e��-s`��[wH�riڭ�45���X*W�m�v�.��n�ձpMUl��9T�jj��8`6R� 8h���loZ�jUtT�R�*ԯl� 6�(��`� *�P8��"@b�n��mmA�����ݺ�,��nįWU��4���U�U6�X [v��ԗ�f�>���0qU�[R�|P��*���UUV���y�IW �֤Ą�]���T�A�%�vUX
)G%[��4]k�oP lnm�9�U-�ܑ������R�U~����j 6)WNp��P'D��쎛'AͶm��h�6͡��F�Z�P���]�@��������`I�1[mm� lհڶ���֐��8�Y�J�l��6� ���`qmu��j�ӱ������$ I'knm&���i�5�$�b�U�YV��U���7SP*�76�f�����A��u�����ۢ�Hl�Hv��-�e�h�d6 h �`��[v�n`n��p!rѭ+�\�T�ڕ�̠1.�h�� ᰺;i�[u�E�a���� �oYj�^Z���H�U�Y�dk����u��>� m m�@H�m�n�hSg:U���Rc"n��R�r󍴺s!�T��<*ҭUK̭UT��Z��34��m�� ��[T�t���6��U*��R�j�&�6�^�t���Rg  m���p  vܴ��p ��-JF�ѩVT�[ ,�h�P$�m� ���m� ���7:�Zf�9҄�@6��m	�m� -�)[kW4��4���R,q�]V�c3�}�v�x1Z��J��jd�2��� �"M��]�l)V�	� 0S��	�m�	� ��-���8UʵT���
Pxؕ6���� f�t�$�lv��Lo@PmJ�T�T�����YZ���+�0l5Tt�@���:�\�92tpmY�j� 6�6�f����Ӂ� �T��U.�2��F�۶El�� kC�՗v�P&��� ���m��m���k��o���RZ�q/;���`�v����.��I��L��ջ�@Uue�P�U���i�l []�;m�m���[A� �`��qrj݆�� l�С�6��@Bv����U��X4�f��F��D���0��bM��v�@7�D�GRl	-\F骢��gp��-��7]$�4�`�` ��6�mj�n�@���A����6���T)�9t۰E  t�-et����\�-UWU]UlR��WJKʵ.I�h  mכ-�\ �vZ ���  �im�h-��h��Y�( �6Á��6T���8 6춀]��eZWej��m�m� 6�m�� I�����������q�dP����8͖���  �	  HFKnݲڶ� ,kGl�6�R�m��  [@l  h�8ەB�[�8Bۓ6m����> *k�&�i�aM����y��Z��Ъ�+�	�l"Z	m� �]a�d� m&��U�!5*�m<���&t��p^�"�	�Mz=�
kp9Ŵ�6�bڦ뛥	�&�ԧe.�UIZ�C["Lmtm[-��*�r���>NNNNNs�����9?rh�?*�U����S ���R( $�aP7� ���(.���vB*�����1@ڊ�xH�� D�� ̙�{�&�X� �*�
��| }�x!PL��)�AA5YDZ�#�G`��2X���X�0=H� 8" 1���ʡ�h��<@8�:FA0�<C�C�M��<z�U���9�S� uMs� <*�=6#�Γ�z :���H�+�0�|.A"���r��PJ�'��.U�+�W�)�
A�<uE�0D�	��qQ!���P���!h.@:��뀜^���T:��DҎ� �Q���AQ\aq��j)��> :'�Aڮ��E�"��D�4 lx��[R��WL�ȝ�@:����b|�P��'ʂuE8"4U:���Ȃh� ���DE>z�Ӌz��$��5�A$!� ��"ā �!B��H�dEc��| ah @rDp`�u0�E�
E~8�D���l\,H��Q�@�EdH@"ńA��B�I�@`@*�'��N���H �?�E���#�H �H�rV ��x
�����N�+ �#	�P$P&�9�0D�@��� "�M	�v(l��t;T��0�� ��:����
�D�@a���)D�@�Z�R�`���ޞ��K�~�V��m�      q�   Ҷ      VÒ�jBj�d.�p^.�f��N+v��A<�s��y��OnNjGpaWt�N`#��N���m6m�Vң���	-uUЮ��M̪i��i,�<Xѻ��c�m�M�v̦s�	,S�.�����1�n�,=�(lH��V*�9u�nN�n=���q]&RW4��)�ڴq�m��6��t�m�H��L�B躌q3��3^ҽ.�v��p�i��كc��rYQ���	� ��)�ڀ�8���;JL��S�һqf��}p�0�7X��e[Z�n8m�s�3`�0t�ښ�����*�E:�x�N�����_&�$1.���e;v���Q1�!��vUY'��q�$��D.�8v0�-�%��[lѱ�m�ڌKl�`\�u�`�ܛ6]&�68z��/n��G�l���q��@���b�2��i��Nsb���S�
�u��p8u,J��5�I�7lu�z�{i�\��C�pP�
��vtZ0���
1�ظ�P ��kk�ΌBD�pl�69���kN�-یx��{H-�q�<X�q�Q�m��Y7�v)��<Vݷ/Bc!Zh&�^��e�vz�-l!���������p[�T9�7n�N�<�WJ�����u6����-C2ݛ�ۃXd�{_5��tq��y�R�#׷4͡�a�ل�v�V�N���ZUٌ>\�E�[U@���d���u����yU�i�V�"�; �[c"�/<$/Ss#�h]��ۑJ�r����Fc�vt��"��b��ܖgk�e�sr�&��P��(��M�&քn�E�`pfv!Q�r.ьT��2��6��{&췭Χuf9�ebA���*�m&�i��4��tf���˰��q�]�Gf���0'!�h��T�:lԆ�M\���f���4 -PV��s����f�6�N��6���1�q�a��tʣ��QpԒ
�a�H�AM�t��+���&ES�ʧ�: �t!��*d@����L�9�s�� ݵ�2�t	vv3h�+y-� �.ց���s��u��]\�ɖ�K�����nn�P8�k��cq��<�f�{;���֎����������7m���Y�g������BAc�%�N|�q��IH�lfL�J)��%�)�n�4X��,�5x��>�r=I���\� ���`��5��cr(u��N���AJ;5�۬bS�&-0�,��}��7�3��û�x)m�����`�ۺ��O�_5���(�	"}���j	 �K�\���1ı>���&�X�%�x_J☾%���g%MD�,K��;t����"b%�ُz�5ı,O��oI��%�bs��*j%�bX�c���%2]�ݢ����^B���ۄ�Kı7��zMı,K���SQ,K��3��&�X�%�y�� �6(j��<:S�:S�Ͽ~�I��%�bs��*j%�bX��yۤ�Kı91��&�X�%��rK�{���p�/���B����t�MD�,K��;t��bX�'&;ۄ�Kı7��zMı,K�N���M�)mهs��ó�-q`��"�h]�[sd-#�SX=��[�R7d���%�bs��n�q,K���{p��bX�&���I��%�bs���'�����/'�}{�f[q��p�I��%�brc��MC�9����J� GQ7����&�X�%��otT�Kı9��I��%�g'{и�fR�`ɹ<���/!}�{t��bX�';{���X�%��g��Mı,K���j%�bS�����l�s|���N��D�otT�<�q,N�=��n%�bX����Q,K��s��&�X�%�~/e$���-e�c9*j%�bX��yۤ�Kı91��&�X�%��罺Mı,K���SQ,KN�����>�l.�=DVGgg+�ay۳���ݹ�.g�̂'���0+b1E����3v�D�,K���j%�bX��{ۤ�Kı9��5ı,Ns<��n%�bX���;�,&s�LbY1s��&�X�%��罺Mı,K���SQ,K��3��&�X�%�Ɏ��5ȸ���'��'��c77�f��Mı,K���SQ,K��9��I��%Ga��a��`(� ��C��h������nQ,K��s��&�Yҝ)��wُ��nPSsT�<:S���>�q��Kı91��&�X�%��s��&�X�%����T�K^B�{��=�ff:�g�U�r{y�ı91��&�X�%��睺Mı,K��쩨�%�bss��n%�/!y?Nu��jLBo2R��s�5=��J��tv ��`X೹K�ɏY1�������1�q���Kı>�{��Kı9۞ʚ�bX�'1�;�&�X�%�Ɏ��5ı,N��C�ܘ��$�$��n�q,K��otT�<���LD�;�{��n%�bX����Q,K����n�q,K����L�me�c9*j%�bX��yۤ�Kı91��&�X�Xb&"}���I��%�bw��*j%�bX�o�v��A�E��'�����/'���j%�bX��{ۤ�Kı9��5İ>� b�t'�g��z�5���n%�bX��k:ǔ���a�M���/!y��s��&�X�%���詨�%�bs��n�q,K���{p��bX�'�t�Oo�=�6�I��m�S/k4SAَ�Wo=̨�tl(GE
�#����I�f��O�X�%��_h���%�bs��n�q,K���{p����%����]&�X�%�xzb���qn3�3��7*j%�bX���s��Kı91��&�X�%��罺Mı,K��쩨�%�bo���s&s��6��|����������ܞ^B�,M�=��n%�bX���eMD�,K��t��bX�';�f)��Kd���1�q���K�"�D�>����Kı;�J��bX�%�9����G)UȰ	���,V����;$��=UUJI��_�������8���t�I�>�y�UEr�UUv0X0r`]��֒�)6�X�0[{5���8�<��k�u���q\�h����Mװ��^يn����<u�d��e74v6�{4o\ODq���w�|<7������Z��O[�kq��Mۇ��1�=��v��3��������a���ǎ;&t��Ы�"%'VƘU4\n��l�p>[�A�v"<�C���{������v<`��f�]l���v�I��c��g�8���v�=)^�b�6�n�q E�Z�z<v�X�Ixd�XWe�����]��v�X�Ixd�X������Bm�vRWn��>RK�;�e`�ǀwnE�M�	X2���ݻ������}X$��;�"�>RK��Aۻ���5n�wc�7nE�|���vG�U�qM�e�~c���AwB�P(I�;h�a^X�n/�V�)<Y<ᇩvN�Ls�7M�Wv���o�$�y`)%��ez�� $�x�<�:Hi�wn3u$��{�4�dC�zR�*��|��@���5�RI�{�ԓ��{t�AR��|����e`�ǀn܋ �I/ �v���r���+M���URRO<e�� �I/ �ɕ�uv]�ؓbwV˻��wnE�{��z�g�����5ݒ�+j�6�`��2�z;i�=�Z&�m��7A�e�U��5�R�K��<��w��ݓ+ 7v<�r,n���wi2���ݻ�;�eg���� �~��>RK�>EB(;wv����5n�w{�I9�w�S:���#Z5�M���6�֣��'c��v�X�6�]��m�v�X�Ixdp�ݏ �R"��hHcL�����$��8`�ǀn܋ ����\x�C ˦&K��P�Te�n?ǖhO< ml�s�W�����J�������_O 7v<�r,�$�Q�"BWr�\HV� ����Ȱ�Ȱ�p�:�.��J�;��;�v�ݹ�nE�wc� w� vB����vR��X����X�?��xyʢ�P"uEx�}����'9�	����⦮��;�e`�W�����,�܋ �{v���Nݻt+�CF�Q0V+s\��<��p�#N1�Q�;K�si۫�N��|���c�;�"�>�Ȱ�2�����Wm�Uj�+m��"�>�Ȱ�2����	5"*�Ƅ�4ʻJ��>�Ȱ�2����ۑ`wDT��v�H�V��&V w��r,�܋ �v��I\��[u�uwe�����~��;$��3��NU즣m�퍶��gM���7M�����m�� �*�3ն
2�G|�LZ�\�'v0+���Ȓ����ݺw����b�V؍`\]9�����p�Ԝ%ڷt��qX� sC�D��n�.H�JK�`٘�N&*�ڹ�F;v�n��Pugmr��:��ȼ��	Q����pA ��˴�jț&���5�,LWc�uc(�vu��L�e���2mPO(gh)�&��JNHG\L�v��ב���6Ӻ�9�J<���,q98���]�k�dM+v]����׾Xݹ�0�� �
��;���J�m`v�Xd�XWv^�r,��D�lv�|��v��&V�ݗ��%%�� �߼��J�+�e�e���[���/ ݹ�nE�vI��}�d�N�m����E�x�Ȱ�r,�L���/ ��aE�5\KV	�m3Bf��4�m����Ji���2ʠ�֬#m�3��5�ܠ��v�Xd�XWv_�\�W9�	/�Xv�Rʵm��5m`�ec�T�C��Ċ�T�O��}����"�>�ȰGh���*�"۬ �v<v�Xݹ�&V�خ'bV6]��v��r,�܋ �+ ;ݏ 6B����vR��Xݹ�V���� ݞx�Ȱs��N���k��p]F.�Z�!��q-I4��Ɂ
i��Ձ�SpJ�+��H����_�������ۑ`v�X�%H��էe���[� �v<v�Xݹ�&V{����g���M�Uj�+m�_���r,6��s�U[TU2�#he:�*�M��;�t���v;���	�)94&�X�$<=�D��sTq��$�	r DJ)M�0fI'> DS�A(��G:&�`d����"�\�D��	>3�!���oY��M�+���c		I�.1�Fu:�bߓ� Q�c.�$�﮴ˡ4I!��R�8��z���|�2� ��RWqK6���.�C�F�3�x&�5�l7u�!p�Cjp:�	�H���A�Wx��g9�f@O�� �.�M
|�+�M�֢��k֢�S�BA�� @��j*o�މ�f�� ���A����;�����}��A�lll{���7�-�s3b�f�A�ll��z�A�llly�k�B��`�`�`�y��:w�@\A����B��`�`�`�Ξ��]���,�ę��Ѓ� � � � ��צ�������t �666=�}�pA�A�A�A�����������ħ�Lg71�!������Χ�AӤIݫ~6���7c�
"SKy��K��^)u��￿��;�"�>�ȿs�<�`���4%e��v���;�"�UUq#�~��6y���c�s�T�o�W�>wm+�����;��,�0����Ȱ��N�T�uj��0�����ԙ<!�<`Y�0С����N �Ȧ�7ެ �;^%��N��|f w����#���wo�Xv�`}�ݰ�]���JYiP��c0i��Al Y[5"��2ʮ�6e�8;WA�X��/����"�7�"�;�� ;6<�JP��hH��U�V����0�c�7nE�okR�K*ҷV ����Lf vlx��`ۑ`���	\��pBl�͏ ��,{r,�Lf�أM	+M �v�o ��,�S_��}�c0�c�>⪯�ww޲~  �wm{toNIF�07Qƶv�2�:ݫ��5.J_]��}���J�ʝ��ұZv��v8�.�m�]���u���z�,� n˓X�\�<� !����7A��
]����6�n�'�[�%���+P'�ޡz��8�^yNEJ1��T��k5�dRJ��0\<X�h��A�}��Q��V:A���l7%�O{�ӺN�t���ͭ��pl�0��l[��Х�Ѹ�M.�Y�3Zi�+-�+
�f<Qݻ�V+M��}/|��#xٱ�^ŀ}�
&��6�����XV�� vlx�ذ�Ȱ�J�WM�����i���c�6^Ň�RSo�X��7�}�d�N�7MU�|t���l�� �܋ �Ɍ�͏ �航�)��v���oob�=ʪ���{�|�x�ذ�.�Ww��ݨ�P���&��5 0Xh("�;y<�Y�з7
.�.l����H��_&�36��￿x�;��/b��9���s�����<�����&�R�S���ﯚt�s�!���7��c~��s���&3?r�����٪~_�$�4ݶ�?~�v�,?QʤvOc0�<�v>NڻV*�ف�����=��	ݏ ��`Q/c�M�uuj�X�ٌ�	ݏ �܋ ��� �ʪ�z�KIG��Zm[V���^�Fɜ�]��=D�`+5�0�B�95����)�l��-���g���wnE�N�ŀ}ݘ��&z�V��e�|tշ�/�X�ذ���6<{��U�Z)��m�k �{�y�fj?����A. ��a$�'�M�gb}&����'�c����DT��i[�]�M����`͏ ���l�� �j�EE+�R\�m��c�=�ճ�~:�_�,w�����t�齟v�Xz�l�vv�]>܇nrR&�nCk��@g�ٶD�7!n�'���e�$�4�m�����l�� �ى쓾P=�﯀ޓ�<Z��\Ze���g�ܮU������߽��v8g�Uĉ�
=f&:�mS��V��='��&Ǉ�����~0z� o7J�m�;t_��r�/zy��?�9۩>9E��T����P�PG����g�����{�ϱ�[�I��������s�s��=��� �c�?-��U�._��t*T��"�]���F����6�/F�<���Xe�8��W	�O5-"��\��~���|�vc0M��\��wc�OD�ʴ�,Av6�	ݘ����\�U�~��� ����$��=\�:�DH~&R�Zm��O<���r�/z���`.˸'I+M �wi����.���s� �ٌ��ʮs�W.�~����Ο��m+�"��%�X�W�{߾��I?~��:�o��F��D����=ߛ�'�f� i�[n����%�p��$ig2E�(C[�J�3�)!GJ��������=����h2[���x�p��Rb�P#;SiB�;q<���WS�Ն�vݖ�CU)P�\�k����j7c�9��=ێv��rVs�9S����ŷ47nN� �d��-�N.��v8Ơ8���ea��]�|�ۛIث"�q�u�Ϫ��7�5!᠎Xl���3sn���s������>���� lj��)����h+4b�a�郴�TMϫt㧨����;w�|1��j�]Z�׀�{�H��&O�w���o߯������j��77)�H��*������z��N��`�r�[�&Z��Cm�wfV%Ȱ	�1�$� ��VhH���۬U/y�� ���`�<�ɕ�l�EBʵv���i��N��`�<����$����qP�ww�Ti�g��n��`���f=�r��P�mF+�X�)Y��.�-ĸ��x��߯�}ݙX�"�'vc0�e�����L����u$���tC�0	Z�@��;�M��D�淍�`n�f I#���H+�����ZN���X�~��&��a��${���;��V�
�]6��իm`{������{� ��2�?W+�s��g�� =����e-pf�����߯�~���^��ݮ��������, �۵J�Q��V�v6��Ϟ����F���XK��		'�'8a�0���y���䩮y���$���	.E�n�qz��@{���;���R�+{9Y�~�o��ww�6=��� ~����7d��q#g��R��H���X�w�$x_*�|�U�D�/�آ�D�"E�)����}��}�w�R"Q��ԢՔ�C�k�O{� ����6\� ݎ��>]�pN��wh��m��e`���I�~X�����~�v�ܦE�Vٖ`�Jp[L��CL ql�24$�.��n���s�꽂QIЩ]��;�"�7c���#�|�O{+ �»��WM�uuj�v;� ;�<vL��r,�$�E��ؓ��E�۶�Oy��ea���~��o߯�{��~����~飇F���m�{�O{��7��,v;�t�eS� ���-DJ�����;���g�Ie�"�k���0ˑ`��U�����] ��~x�p�&�wIQv�� d����{v��ѝ��m����Y�o,.�	j�˰�m��'�оKU���7+�{ߝ�X�#�7c���W9�	���`��y"���E�)YI�k 7dy��*���ѩ'=��jI�;�ۯ �9w�~����;��x��V�z��W9Il�^X$��:�-#|Wx�䔸�MI�AȂ����5$�f���Ns�Τ�!�U{߿|jI��'�n4#4[��'������'O�$���~��O{���o��f��0�ʤ81t#1��� M)�1�Hv`	��Τnϔ�r�P�׮3��1�0��qX�/E�6'#��Wc�&W�45�̧�nWdb�a%;���-�E	��!�;_3bd� kc�h'�r�&�B$�a6`���U�@��#�<!�I�1��(���A`���2 F81 �@ �i�'.r�	.��sd�2��m�@Wp9I/0��āB2O��ʲ`o���`bB$B�0m#����:��l	��P>��w�#�ti	>Q1�&F�`�~{�?���sm�      ��   t��     հ��[��
���۷ny��f�hgi��Eձ��ç���79i,��V�+��@41M`Q!�e2�S,R�^�3E)��;�)\�;����k�y,�@�E�8��X�6�(��)�V�/�WT�fa��?�=��#NΫ%�A�#Kc,F&$��Jd 7��C!41�X&՚`F�iteƈ��im�rf�R�$�<nj��XPI�Ii`C�,UN��N-�&ښJ��0�9��L�@�!�0�6�=��g��؝jW���p�M,ihK��j�˩��y�v%�wn2�tB�v���<�]�I0:�4��)�4������,˃ �W&�%��,�[L4e;jU���d5�:s�Pڭ��#��-�(GJ-�F�� !6�H�m�h��+v�f���kg<y��A�ٹ�,�],y�l��wb�D�Z	`��˂R猦�aڛ5T*����S*��g��f�mYp㧔��^������Jb����e��\�v\� D«b�-���&��
��&�N�Ս�����ɧ���������sn����b^�B���	��as�a�]��"s��`5�l#���(76����r�)���C��,�!;���T�4\�j�]�q�Vډ�(d�s�8&5)RJ��&��v�1P�iaQ�h�lS7�����/N����U�儯kmMV�8�^v�+v��a;u��!�$O'm:���ḭJ���h@�[�Z�U��v�9������RyJGM/m[n���lR���\�69;n8d�+ ��R�4�j�v1������$�.��Ѣt護�k�E���墫x��r�3�i�Q��kK,��V��aΐm�:@���w-skm����1��"�j�j�BuN�
N-]�T�;mV�u�����İc�5���Uj��z"����C�^�(sV��v�k�.�^!�nh��t��h�8��r�iO����!D�?�J&H�D<
)��DO"#�0$=��>���� � ��J�ѱq��gA8Ml�N�md���B�ݧa�s���yܗm�'-ٳ�Z����4�0����؈�Gc��)�|�CKbCMm+����K�:&�a��`Mj12�M3�dݢ���XT3Xg��޶#�����lX�������[�W���z�V�V�ٲ�g���0h����̵��ζ-�T�-�̤�{�rs����I�=��5���m4ūMo[d��Tp;���S�����B�l5����6c��ؓ��E�-�� ~��� ݓ+ �nE�s���k� ݉��ݎ�M
�&��7d���W?r��f���`ߚ����窹I�yREhH���m���� �Ƣ����F��I�e`��,��ӵav�X�UR��^X�<��2�=ʮqv?y`Ez��J��$�'i� ��x�����������wcQ`��JU���:��M�M���2�Aj�%x�5�kj���G5��%L]x���X��	�V�݅Zm['���ݍE�����9����������Z��r[�K��jI�c���&QR�#���H�9�ȞEwO���������s��$��+����L.�]��l�^X����r�)<�`��, ���+vZv�e����Kd��$��}�"����+�$�￾_��>�=Y��s̪��8`�9����y�, ��xa#�g��L)t�wp�X��8v��V4�0��4�v3 �T��%'����,�����[�m�>���nƢ������W�Wl=���`z�ʅ�j�;Uuv[X�j,�9I��Oy��>ۑg��\�5�_�R��BL�V'i� ���l��Sg�P�`+���޺�w�������o����n_�I$��K���~0������X�UWs޶�򇛫I�W`��� ��L	�n�Q|�y�#��v���n��t��q�]N{�V�E��\�O�ݶ����g�]�p<Ĝ��_!�yb���]���}o���ǀl��+���, �x���ӱ�[���X�����D������nƢ�r�č�2��wI�
�&��'��`mȰ�W8��k� 6O<߾�@��1lT�s����NI7߼��5$�f���O���R~�"$"֍X	 DB.��HXP$䨪t��*��w�ԓ�~/�/�Uf��x���~� �?I:I���Ϡ{ߟ� �c��^݊�]�Ui�a�'� "]�޺Yt��?r}�01�v9��%Lt�:)��y
�տ�}��n���*���<ז�}w�5Jۻ��M�o ݎ����r��y�0	��~X��y��5W�<�ZMڻ�J�0�{+ �Ƣ��\�H�<�	<�`�A�n���WV�����R��^X�<����Wg��`�<�ӱ�[���X�����������'=���I>�s{u$����g�������ԗ�  m��6l&ixp�҂-�h����nvg�m��t��3�+�~F~��b۶���x�j"�f+��ۧfä��	��c'4v�m�k:y�>�M�t�n�:�e� ��X��bZ49���m�ƺ��%g�:��/�S��D�N�@X�lu-�7m���5s�v.���A��3�p����.��Qz��Q��*Yh�9c�^�r{<�$9ϧ���Ǝ��H��i�8bӋ��w3K��ib�KRŭ��ڒ�G!��$�%�|��մ�]+��I�����+ ݍE���y���RE,��M��v��&VݍE�ݏ ݎ�H��^T,�N�����v�`<ז wv<=Ĥ��v{�X{g%X�WR��i;M`z�-�� ����܋Զ{��}w�5J�ݠ�M�o ݎ�r�������t	��~X�����P�{�E�א��E0���4بb��as5�c�M!�`nk*�;��L7ŘF4�l����ݍE�ݏܯ�I�� �p�yj���q�ի���j,�������w�=���I>�s�&���������t�?w����GtL��=�� ݎz�Iv_���k� ��⫧M��һ|hm���)=�0���ݍE����Wꪫ���x�ߒ��Yi"�k���0��X�l�//��'� �0إت�̫ht�ҫTk��]v �J�C_�_�9zu�0���[s����ޜ�K)'M����5mt{��V�dp�+���v_��	��!�����.qsu$��ƿ��Eb{������_�� ݍE��*����}w�5J�ݢ.3q�jI�{>��o��n�%r��iQ*�R*�J��Q~v�{��r�FL�^X��<��7V����b���r��\��~��$�^X�9��O�'�L{�����{�$�q�S9��WV���7cQ`���R�<�{���܋ �U�F�v�v���+.�^%!c��5��k�lh���ơY���2[ltc@A���v�N��J��_ l�x��}�"��Ur�A'�� ���V���:J�[m�#�{�\�����'��'ל�5� ���N{߭-��-��s[m�0�����8a�URZ����~0�DJRN�����j���r����ԓ���5$�{��ID@�ڈ�vq(���5�z�I�=,,���1w�t&[0��x��}�"�7`�<�t��7���XYa�f��e�1hCv��8����^t�-4�2�.n)J���/��Zخ��
�Vջ����0��X�=�s���j�(y����ue�U�f�܋=UIx~0d��7c�~�9�'�����`~��c�:�i������ ;��*�����~��	ͭ%�;
�V�Xف�s����{� �nE�w`�}�qU�m7N����x�#�=\����/���������<�@��������������s��!�kj�[3)�p���NxN�-��7.S��;�X)÷-�Pfm���#�	z��F����s(6;p�t�ݬJ�u�U��wZN�*B�Qj,��E8�N�x4��й�Lg^���v�i̼h�mܗ3��F��ţ1�p�F�N �Z#&z3���!w0Éj��a�K[�i��-X�*��6�8��fs:�h:�ox�1���3n	Jd��3lv88Vu��;�ە��y��,����_�w��CK9������������� ;6?r�_ $��6$z��������b�xv�RA��� =�ߞ�מ����z�HN�Qw|WBe� 7�� 7dx~�W�}��6x~0�긓T���
�M�o�\�����׀w`���U���w?{��"������:N��&[o ��/ �r��x� o�� n��B�t];WuWn��c;�'f��b���!4��mDyѴ��D1����S�C���Wn��j, ���vG�W9��[�^ {����;h*��[M`fǛʨW*�ī��V.$XqT��)S�L�G��{�^�׀w`ឪ�+�����cLn�+��I��	=�Wd�?s��s�W+�ʻ������<�ؕ%��J�k��X��xv5 N��=��*��'��`�H�#*��wuuv1[��� �r�U\^�y���V�w�)��?�,-��[�"�ce�mה�p�
N{|�t�c�^%+쓤�^�S���Cmt�����y��e`n��U�r������7����~����BiR�x�X[���j, ����~�Iݱ������V����� �}���I�;�۩����Q�Xw��\�O��T�~����-��:11R&���A�$"���\*f�N�gʽ�v��L�H�#�	@�������������%4.0�g����`H�D����H}Q7,2�,M��7��7�8tgɢH0#	���(O���3�g(D�O�SdU(+�G#�e��T�*M�.����O�#�L�ez"U *�W��� 	�!�b` z?!�eN�S�}��:�w�����~��u�Ơ솅���$�z{����I��E�/ 6�l�G4&R���������ӽ��~W�yI��&Ƣ�?W�]�VR�&�*�՞D���h�hZ'������b	5�0��w�;�]�dlV2����=����"ݗ�}���Ur�Ur��`~��<}��RX��t���v�u�E�/ �� 'dx�eg���8����2�t��+w�zy�, ���������W*���߲��߿^;�H�MDw�t'w7RyK}�{:�{���I;y��Rl4A ��T�{��uu$����4���]&+o �L�ܪ��z��漰:�ܗx�K�;}vz�+n��:�N7nոӪd�Vͳ�f���[i�� �6H�u����Iʣ|c53CL4�f}���b��oy�^���{�s�ǐ7�[}�{g��~;-�hx#k�n�����w�/�I)w%�$��O��J\�f{���r����?G%�-aDO} ����j�o9����A�1�{>�ն߻�_]�н��-���n]����Ӝ�����k�K�����$�ي/�I)w%�$�߾�@��X��\��@;��o����_���c�1�m��;�{��~H���taeT�a0������_�|�a��K�S�2����͜�6p����Z�z!yy]�6�,�4&p�8��1�(b��ɓ�f�%�ܰc���ҭf��iVh�f��g�	`ܰ�6NŰ���е�	fH�K���	eI��\;�x�C�g����dc�壗�h��#:[�0)�&.�c��^�2�KWV4�D��;%��ݛ�m�Y��,t�f#c�l���N���r5�h��֓+�B�Y�,@�dN�ۭ��>��|��m���[vs-�������hx\�m�ڴ\��?�x��������y���=ǀ��axw��'��wo����&�?���~�c����=���m���M�b�t����$�d�|�R��X���s�6�z��}��o��x �O�X�M(�>�$�떱$���!��%.�]�K�����������Ƈ�6�6�L��_wL��$����]��K�g��I)z� ���ò�3ͥ�Ml.r�'����{����ջ��Y%�&!zcg-aK��������y���=��v��o����_�i�֬`g�r��۾s]��\�8����gA] 1� <�y��k>�ն�w�^�ݶ�o����}�Iv�T�����r�$���d>�z��w��I%�3��$�F�JX�v�.�&�bK��7���%��I%�^��)ʸ�%�I%�Ζ@��!��J��������y�I)z�I%��d>�$���JX�6���l�غ�e�%B��,':��=����TD�5��T�M�],Ј�z vL���%/\��$�ݬ�������� >ߎ�ch��ih��@;�{�%��d>�$��˼I%��C�˻G�Y�:���2�����?_} ��wՠ��4T[@
�5V �-������O9���zov����< �~){�T�U�f��
]�Ē_n�>�$�떱%�]�J�Ǿ�_�i��ݳŪ����y���%��r�羳�]�g��I)w��J������4?�Xd41,hM4cr���7m�gGm�烴;�Y��6�Ґ���M.��c�gz�R��1$�۵��䒗{.�U~�+���^�����%���%��-ݫL���{<���ܜ�c�������g��I){2�I%�yT�B�v���v5��%.�]�I-��}��r��w~��5� �w����@?�|n���],Љ����G�g>���7�m��~�&�������p��/ELMg��5m����]XSJ�p��}(t��k� ��NWg�^]�Iy\��	%���I.�ܺ�w��n`҇8�;+�Sz�%����D��%CB��X��� NI/��e�c�n�٫�$�g�y}�IE{�I-��~�s���㿼�� �;�'�UKuZO}{q��k��3���{_��m����.�����z{��$�ӑP��?�i����U�x�K��~>�$�.e,I%��E��%�}�x }�����45�S��7�@�#�{>�um��{S�{��\s���S�Ͻ������ǳ��2��s/��~ي/�I/���II=�}�Iv\�X��� H@`������wK	�:H�ڪ���P��6^:f���˵u�c {l�T�9�gi�<�݇]'8B������d�a��N"7n��*�۫����;]�a�ї"8*tc����[nwY���ԍ�n8Hn˸Q�*�3��;��Nx�3��ic�`��7��h�Z��K�"\p���ҽ#Hrt�s�)o%k��ign�B��%���yxI�a^�.ڪK��	'I=�������lK��;Z��ɁK�ԌbMH�v/�����8�.�is���$��W�<�؅�v������oIn����$�\�X�K혢��긣-��],Љ�x }���{��m��߼�����?���x �O�1�h�\4���ww�x {�o�����x }���{��Rnڶ#�4�ۥ�$��d>�$�\��$-ݟW�$�\��sw���/��w�Oƪ�굅.o��}�{���}�g��}��x {�o����}�`.ua��2����P�:Y��9�h@�"�s��m���ۉ�Z�4fm\�������@>��<����ʪ�w���~��$��=j�֪���Nge���W���=�Y-�N4! A��H�H�]��k�]�ݶ��q�[m�9ݛ����iᲄ��E ~��ߒKn�ĽWw$����%<ߒĒ_w��;����s}��ݼ >���=��C�߻���@?�t�[��Y�;x }���{��^���wç��}������N͂S�c�4��W{
x;%m�v��6�� vy���|�	�Q�f5�IL�} �uz �������� }�}��~����ф�P� ���t�����x }���{����� ;��N��J�k	qsw�m�1��f��s�5<�U�"���:��s�'��o���}�]�6��Z|�kܥ$�Հw�~0�5��y`g�R�˫�k���0�p�;5���ذ�>�-�>>ړ�0�(�f�<����9��.��g��������b�qg-�9���Q�8��u�ՃM���y`��`�p�>�� ��ڤ'��)I;M`��`�p�>�� �֢�>��
wi�AWJ�m`�p�>��ܤ�ѯ,K�XTZ\ZMիM
�0?�7�{^��s���ԓ���5%2�Q*�-
�B*U�Ujʀ�y2���W1��� >�.�&�i�v�U�l�;5���\�U����_@���`�� �AmؒE�A�An��;制�v|�y�k-�$n��pVknHMi�@@�����6:V��"ݗ�w�� ���9���5��O*�h��%|�i��>�p��UU���*�����`�k��"ݗ���"l��U����m�X�ـ{|�`�j,?s��%�'� ����%.�i(��J�.�i6`~��ݘy`Rz��0?s�T��g�}�U	?Z�vR.���5n��>�p�>�� ��7�RM��hP*�%�䁳z��G9&����e��AO����B*F(B1!���C_a�*�1�<�[���Nl�i`�Mu��Ap� BK���#��Yz�|�Ő��&�1��!7�$$FE��p�b�YX�Rc$�C8U��,Nq�Qƴ���\�dI��ښrH�'y$RBY���a�\�5%�,�_���&�&6��+�Jh�D�BO���jwB�0ǆ��3;�~�m��9�@      '    �      6Ͱ�m-�J�ݔ�뮭̕��g0qms��b�3s��Izj���n���۶�!�m�7N��:��+��kj���	�q�iT��qj��lmN3�-��l�l��^x�	�x �Й��i��l	����j����w�Y�����#z*<����u�1Ә��f�l��͊�n=
+]��
8c�J�D���DTi�7lhʯ9�⎻%g��
Ê���\��@=%���H<!MmP���Su�=��8w ����'=#;���m�nۜ��&p����Q�mR�x}���y�`������u/<T�u!/.�**�V!B�� b�M7	�A�ɞ�%�JH�j�̭�Om�^��̞0[�nU=����v�1>#xvz{f��ɷ!�G4��8ǎ�:5�p<b��7A�9�=p��gڳ�*KrS�Z��9�+�t�����p�Pn<��, �:�s�ԗ99�㝻�,s���=-�gQ�j����ݑ���5J�m;��w ]Mcfфuk��xݣF��+m�ƍ��0V�M�2XM@Z�v�8���a�<I�8n�э�-G�W�u��W��n;\U9��t;ʁ��UP���^[�C�g%D��v�^k\j�n��q�dv�pLI�D�o1a�Qb������R*C���p�u�`��\�]J�T�ޱ���I����5i1����B��WF�V'!:}�熸�f齺�v�T�
X�#���Q�5���#띮V�nGv9�P:�Z�'VɵGG��Ȋj�.���@n�J�j^��6�vJ��X�@m\vm8�,zJ���p�V
%5mj�SkD�.�I���6�.�7pm{XCsM���,����i�Ʀ�(�\�{Dlv�UQ�[A\�nC`%@t�/�s&�Up��5��t�D�l���H&:e�)*�S�ʪ��g9��1��J��K�"�����`C�H�A��_�I�����T>(�Ө6������������%� ��s����-]Eh�ң��5mq�����.6�h��h�&pu��I�����<vZ��m@ɛTa�
P6ZĖC\�sŚ��crb(��u�!�Ƃ1�#�KK�i"��ؓc2�+!��T���[\x]�z����DqŞ\�k��ՎM�4��ֺ��''q�%��]+�V:�5.�p��l��+I��I��%8�x��ȷu�SK`S��M\`������%�m4�&@��ÇqJ��_2v�֓KCn��~0�p�;��_�s�^������߆�n0�S�>}��<��E���c�~�s���~U���M:N�*�m�����wc�>�p�>�� 'u�m	+M`y)'����}#��l����'�Yn�n��|M���c��wZ� 7v<��ګ�\�Sv�C��K��)�$6�ѭY�q�:�p<���xe�8��-ڥYj�����~���E���W+��?�m)Iy]��X]X4ـwu��9�V��W�}�g���'��`H៪�7�%P���N�Н�����v8a�����?�ז�nF�);j��WHo�9���x�;�?{���9UII<�^P��M�X�wwm��L���V����	'��c��D�%�v����#��.ۧ�g/i�ٰ��Ϟ�L��86��9�c)��i�v�U�l�;�dX���v8~���Uv�~����y�X[tU��$+�ݏ?r�Uʤ������Y~�W
쇋-�M���M�RO���jI���5(��Q`mW/��b��, �����T����Smr�v��\�?U^�����{�w�`�ǀ}��J�[J	�*���j�`��,ܥ$���&V���;+����#
���\`��/lC9��V�i�2�,\��(���® ㆕��ݏ ��� �I��w�Ȱ��t����,6��c���+ �u�`�e��^P��N�+��� ����E����O^���H��Se4�;`��۬W8�f�����ﱩ&��{5'�T�\4l�T�H��%�D����Y!�L!��Q	��������DTVӥWJ��`�e�v8`I2��Y�s�[�Wt�/Tm��,�;�:�c�b�#��՝�;���3���GK���"��5w�;�~0��X{�� ջ/ ��I��"�k�+�`I2��U\H݌���s�E'� ����'m*�Uv>X]X5n��Y�v^�c���+ ���-!��]�k ջ/ ��� �I��w�Ȱ��twr���`�m��c���+ �u�`�{�I0 ��� @�ð[1�>� �4�m�嶁�<	#����I�l��NW�8d����8�u���f.��
% &�tt�������	�gnr��wX]��G:��#fN�����ڭ�`C3%0L�m�y�qx�.9���cgq�5���W/
�v��"4p���S�;0ݴ�2�t6���M�t���VE�����+������:�+��j���ΓN��6/|�VU�U�%�PR=�v�g�5�ƹУ��n�q�9 �����#\�Q�l���L���E���c� }%��1�I�j����"�r��H$�xw����s�\��ձ�m$�ҺT��cX$��>�põT�dt��u�`w�����j큟k� �u� �u�`�ǀovZ��V[���|�]� �G��E���c����o����xS&LD����(ۨ��ڈXҟ��$� �v5<�27�`9�.����>v3� 7v<�ɕ��������()֐����v5��e��Q*��.;��o��f��}�ȳܤ�[����]ݢ�Pۼ��e`H�w�Ȱ[��n�t$��X�wwv� �G��E�jݗ�}�2��.��:N�*�m�{�� ջ/ ��e`H�M��J�;S4[1J��£�,�l����7���uɂ5+�íl�Ir�K`���ˣ��xݓ+ �G�U|�v3� ;���L��V��?���y��KO�}|`��X��y�s���U]���j�ee�H����X���{����>��J(R�"�P@0ĨD�	Z�AG(����s��x�}��N�U��J�|���i��W��� $�xݓ+ �G���R��w�t;�� ���W;���������E�H\�)bb����=��q3���<!�.�c���3����ujj��)��4
l��l��]�?���x�8`�/UU|��y��/�:B��e!��ݺ�>��?Us�H݌��	'��d��Wꪫ��߮��Ʃ�I�V�� ����wc�>�p�>��-���wf�h@�j�[��{�Τ�罣RM���ԚS��`��"1A�/�Z���j�I>��:2ݕnؒT�M��܋ ����߾�t	<�� 7v<���`�;-㐰��¹TL�������\K(5���`�T�&�RV�ۡr���V��{�v^�nE�N�U��J�|��`�f��8`�e��Ȱ�p���9\H��P!���n���ul�"�׀w�"��w�~0�3� ��E�.�]ݢ�Pۼ���{�U\�)rz������ڶ��>�"�=\�'�ˠy{߯ �nE�D�!(�DbD�A�cQ ���{��zw�{��~�� UT�b�
h�Y�ݵ&t�u�xt�WC���Q��0��.aq+e�+�����[�ms���ӣz9�ϛl��V��z������qB0Ŷ��5�2BX���ƹ��x|�b�a����&�St��b�ys˵<{.�T�G]��l+Ʈ��15#5ī+.�3VR���FS>��m8x0��q:��A�f[����vC��N�wY�K?���[�6\��2�M�+��le�;+���6�{q]�p<����Z�Ӷ
�[g���E�jݗ�w��~�}�� %lJ�vƇI�RUwcX��y�#v��w�~0�2, ޭ�2ӫv���i��;ۑ`H���[��	ݖ�j�%��񤭬�0�ʏ ջ/ �ob�'m*�P�v>Yh����ݕջ/ �nE�|�K�'H��U�б�]_t�<���M����g�n�����c��.lZx�U�4�M�e����]7�����Ȱ��x�ʏ ��.�Z�V�)*xԓc����Ѐq8�t����.�� ��ջ/?UU$B���Uv>��v��=���j<�v^�nE�o.��wv�:Um�x��G�un��;ۑ`{�K�=��	[��cE�|T"��:�e��r�U���/��y`{*<�\�پ��W^t�m�m�k����@�|�n*g��p�[�iJ�f	?뼮�MY���Z���w�� �nE���UU|�T���=i��p�|i&��܋?$��<T����QZ��]���,m`{*< ��xNrr�s��WGU��9D�"0$D��bƉF�}��mD6A���)�h�H�&�
�3fUU(:�$�@�ŀA�����0c E� �)
FƤb�"@�
A����PmM$u 9k��H`c)���������ʄ*��#ā2�n%X�]�n#�Lљ���nH� T!@�U��$��P#c	%�P�!A��H���P��#B!R��J@�i+(B�KHP��%��. k"PA#4�	Md[�!���E���b�dS�c:�������^ �]f
l�@6��8��Q>*���\���@W
8��k�@�l8�M�`�EN����U���e���`v�Xv�j��m[k����x���<�۞X�r, ����5wK��b�M$RT�k �nE�{��W}����� ݽ� �/��ksu�ڲ&v����,0]v)��\�oG������m���ҠN����7m(̰�p��Tx��_�A�s� =����V�]�`�ն`wn<�\�H���n���6G�ʤ�T�R������]�x������8`{*< ޭ��iջbwwI�ف��.�>�ԓ��}5$�}ùԝM��X�#��"1ډ�k�/oy��	ݖ�j�ۦRv�dp��j<dp�>�Xꪯ^�]��_�a��В�.�DLe�eg����g�� ����呙����I_-m�iv�����=������ ��e`#���ڤ�V��;��dp�r�������	�?��G�ܪ��[��i_���J��0ｕ�l�~��q#vW�=�� 7v���ب�۶��� ;ݨ����+�r�\��������Ά�v�۰Uj�0�ڏ ���g���=�';��jI�5�ؼ�x�QirDB	h#������g�ߟ���  �n�.�i�ѧ�83O��ݸ4<�m-�Z�-��D�e��7Mː�2�����˶Sj�����Ō�&�! �ʻrj����#��n�$v�;v�V9�ۃ i��T�k-�3+Vd؁뱯<�6,0u[Y����T��{u4l0W�7m�lH��s����im�[B�1����X]-6(KUq����Gt�g{:3��I���[�[���Ms++�%n���0�5�;\�3zݓ8�T�f�GF0yk���r�˻&��P��o@���{{�8~���y�6_�-:n�n��4�0�{�8`�ڏ ���Us���wt����سm<qz�ĥ����� �����r���?v��Q�Jv:��6`~��s�wey�<�`v�,�0��I�;�����xv8`���ʭ�������������o�u؄�	wfJ��r얖���Ј�&6%t Ksm4�&@���HR�)����M$RL�f�c��0�ڏ�*����~0Ik�tm������ԓ��=��9(m��ҡ�:	���V�M{��ԓ��}5$���f l���ݫ���Uݶ`{��0�W����7�~0V�*]պ�B.��R{<`�{+ �����< ��<Yi��6��*i� ��e`���x�vW��0I��K1�*Z�0�]�+(dUg�]��4�it>2����Pۚ��i�a�Xdp��j<v8`wfV�Q�)t��VU��m���E�n���ŀvG����"������-�'���0uڮp�ܢ����j%�9��{5$�19�jI��.���.1���f��g�}�� ��%�~�R�{��{ּ'El ���l�>�� �Usc=��	'��������:O~��{����)�p�<b�&��P���Go5�jn�
DS\D����[�v�۰Uwm�z�߯ �ٕ�wc��+�J"���Qj�� �ٕ�wnE�}�� ��%�۱U����;�T��`�ذ�8a�K��z��~0���T^&�����k ���K�;���qV�y�F2D�.�����X1IHJ-����c<@��XƳ�&�Q�P�v:��6`m\� ���{ݎ����o��\T:����f��e�ݮB��Հ�42��#M0��EZ���R)V��t,�� �}�����Xv8{��|����X���HUu�!����;��`��}�r,����y��:~P����Ѕ4�۰�=��0�W���� ���, �9���۰Uj�0��E�wc�ݽ� �� ���t�5O���m`��wob�;�� �j�X*���'q�;�8��q$:�}��UUUPݵ�&�:$�uc^X�wa��k'&vι����u�:�^C=p#vH��Ef䋹o4��j��k�(F0�u��k�X]5�fU8��=��p�X�p����|EQrt�M���i�P�p���n��9�m<��s��������[؄���b�:��=��㮴���B�x1eqv��ՙ�a"	�dˋ
�%6��Y\��^Nsߧ9'�{���/��l��1<s���pr�.�{Q����8�@ڻ �k<��oZ�0��wum�n�SM�}~��;�� �j�Xv8`��J��n���o�I��wc���Ȱ�p�;��g��8�D�վX�`�f�W�,�0�9Ķ\��6y��>�j����t,����wI?o��������0�p�>ڹ��.�%WR�"���v�,�0��E�wc��}������h�TfV8�8LǛoV����̹�Jn��ZR��[v�����nƭ��wn���~0��E�wc�ݽ� 6NGCe�wv�%V�� �j�Y9\�eW;ʯ���l���>��Xv8`��@�顪|TZ�m`��wob���[�?e_����-7wVڦ�4ف��,}�� �j�X�v8`�(]+���+��$��;#���Ȱ��wob�;��
.�a�����c�-�t!&C�]g��=�[�w�3�c3�5k�`Ja��l�cS ���{� ݎ�`�� �h�!K�7|WB�m`�� ���8`J���]u,B)+.ـn�=��}��S@�6i�% Ȉl�T�-b�Qд��~�Je0GjP�s�э~��{���$�{���v��X�T�{<`�_���p�7ob�����j�J�[f�e8`�S߾�t	/ߖݎ������Mb�TŴQРj�Ƿf�3��5{z�V�\�8����u�(6<TX�ـwc���ŀwc�������	�x��wum�n�SM�{{~�8������?v8g�\�$z��¥x7W�v锓k ��� ��N~�s�Kg���s� 7B������	6`wi� ����Ł�9W�n����Gʂ]w��jI��!z��"�;�fݎݽ� ����8`*�T�Z���\����aa�GK�iڙp&��KvS�uEQ�9�GK���R��l����� ���}ݧUs����?��I��$�QI+v���=�>�)��;�� ���g�s���~t�.��%V�� ��~0�p�>��Xv8`��t�5O��[0�p�>��Xv8`~�W�s����� ==����WVڦ�4ـ}�ذ�p�>�ӆ���f��%@:�� Cp
(J���"�f$0XŁK��s�qx"�8iIk?d��]0�9�`������M�8��ih�@�44��1"�aQ1�Fe��:
Ȑ��A�!3�	H&Upf@��$X @bHs�q���c 0��7ǩ�BBL��tB�� nrGb�*�>�D!�ζ�e�L�(8{�b�NHB0#!�1M���d!BHM�9"���� @��B�'���"+7hŶ���e&�@�uۈB�R,#��la~���n�)�1�s@&DjD��/�g>�d��=X)�(}&SB8�O��a�pƟaM �L�^51�N���>���ڐ�      @   �      ��E�J��J�T�$n�zdu�Q^zwkh:M�.�I(JC� 㚸=�M���s+nJU��c1L�P�,����� �;,9�����i@�kB��j,�"(��X�`��Ț�p�ODq�+K�Ѹu��)�Z���Ga�&��[��ǯ�cp��n*�CJ��DH�+-Y���Zβ+�sAč���ss��g�[]Daxx��#�Û��uq�!��؋$�kH� ˹Y���ȳvC�QJ�V��x8w];�9�����=72�J��1rgP�ɵ�cH�6N��pV�m�<!U�k��]\�uS&K�u�Mi;qA.Y�Xl�*��IeG՚9�4��S�UH���x�t^kuFӸUKm���d!oP+%� �Gcu-�e��p-���Mҭ�-'jC�85��sY�h8��G ���A`��%W<�q�v���.U�s���A�9��r��	�rl�Z��ۂ�v�&'h$���.�=t/��6bh��9�0Es�H)����wI�$��m��y�q�ۚʽ�N�;����G��{lpB�c��
K�`i�7Xs��\�ѴԵ��HF�h��u�$��DKI����>檆É�wKMW���ݕͺn| .hǢ	��7����6�����ewF�F-�C�;�]3<�pVqꇜ�EƓd�.ԮU A�e\`i��ˢ	@ZR ��D��KX�s������É�{s�j+Riڇ]6��(^��FEk�C��T6{s�L�:*.*˳T�P���7\��%�c4c�n[�e�v����gPJ�jʙ�X+Y��f�mGNM���WmWN��HCP�ń\�c����u٫geg@���M�;+O�v��f�E]�iUV2I�s�ђ�]]&wn%x(���Nkѳ�Uy�����4�DaVRƥ`��/\^��	mlʹ�Q�X x��&D�½@������TZ)��U��D�DE"���C`#��T�=C�<�ܓ��v� 6�[kFDոX���l�n�c��:�4��25��n$�Y�Kb�J>xH�ku���p���N[�]g�2��җa�&�K1����h�Wn�f�J� `�.�%�k\�!#����-��R	���*"*�L���S��^�1ڤ)ٜ&� ��<N��D��\�.��l�ݭC�f��Hܶ���ӻ�O$D�hyG-KP@�a��mG�%�m[:=��8�%�ڈ��e�S^kHf��6x�S�}#��v�0�p�s�۞X Q+���ӷtZl�>�ӆݎݽ� ���8��$!�]�ӺE�wV�g����ݎ��p�:���AwiJB)+.ف����vg�g����8`���qRhCaE$�l�;�� ��Nv8`?����?�>��[�l��E�2��%�ZX�faP3�3�MdB3�ϒ�f�s.�����ّ�NӺJ�[g�we?v8`v�/����?�-]6��Qb�sRO���k�$~`ƪ�a���W*��nj�>��}ݧ�I��m][j��T�fݹ�wc��v�0�p�%HAR���|bM��0����;���Jl�Q{Ԯ��:v�M��ee`�U����&�� ����T��
�WwB�顺�Sjg:P�#�4c�+���'5�)Y�!a֡�����yB�_1�)��������7��wc��*���z��[R�U�ݯS��J˶`�p�;�� �l���3�+��/ʓ@*
)[���I9�g�RM��4jk���� �	�")Lk��{5$�;��H'.�7I�wIU�l���s����� ��� ���U���U�~����G���aj��Ӭ�0�`��}6VV�6ZH���:t��P\���k�ȦSVz�����\8�܀1��f	=�ҕ�˫n�M�7t��π���0����\��?�C�
�n���6��p�W*�\�G}=YX�?��,�U\�$����*N�tӺ-6`��e`��oob�;�� �jIRb�t��"�[t� ��{{.��s��ԟ
�j� ��{�)^�Uv]���)+.ـoob�;�� �l���0�l���]�RvswM/*�oX'b�x�6�vݭ�t��vy���|�P�v�&�!��)$ݵ�wc��d���=U�s��<�{��N����]�Vـ}�++?W+������s� ���\�) �IK�ն��O��j����������Kg������ �v������wJ�l��qM�� ��� �l���\����z�<�w���+��'l�;�� �l���5$���Τ���^8W	"��w~��VΕ;n�wQ�L��C���9�'J�u�\c\�i��w��,�A��e�� �2��mm�\R��T�m3v�,��˭���t�6_ ��i��ۙ��ϒ���&�]d�L���8�(X��n�\bX @���>x>�/e�c���L��K�k���[:x��ݖN��"m��y���`�
]�[��]���M�dÓ��Qړ����LDo&2ׇ��|������ �ڌI�:i��d�GK��[{�߫+ �ɕ�ݏ����6y��=(�J�=eӧt��mӬ�&V ov<�0����:�[t�]]��H���� ��ݎz�T�}=YX�{+ $ۊ�@��E�i� ����YXvL�r��vg� ��<�ӧi�t�vն`vJ��?��=��7c�wc���UV���ZW��{;O̄Mq:�ۮ��4�(V��j�ŀͬZ�i�&�+`�S��t��6{�X{�v8~�s��z��vW��n�ջ��L�dԓ﹞�aTSPA	HJ�;�Ur�UT���`ݕ��wd��%M"E�M���Rv��0�%ea��[=�v?���'T1�P�f��YXvL�{�v8`h�T�V��;�]+n�`�2�r�����<�`M���}���*	zص�QU�B����-�Aq���{v��v�<��6XQ���44b���Y��\0�p�>�++ �ɕ�mĆCMRI���3�Ď�z����V�� �*��;NӦ˶���I7�tѩ'��tjd�"��H� ��R`�M����Ϧ��� %n҈�lT�����`~�W�{��&�� ��鲲��ؒM�][�n�5n��`��}6VVݓ+ ;6�U�*�1�6��q	۲t���2��e�LT���h�<���N�TK<b�ꨒ�>����}�++ �ɕ�w��wlQ)IRuE[g�0�%ef׫��'�遻��z?��D�4'��N�I�N���e`�`ۑ`vJ��:�[����.l����MI��;�o�ԓ����RM��4jN�NU$F��yUyX&�H`$4�E$�l�;�"�>�++ �ɕ�ou� �U�W+�{|1��G3,�����kISms�pN�=Hn��X�L�V�[hmCk��Y��˝Fh�4�]{�e`�2��~�s����� z���Z�	�|T[WN��p�7��wnE�}6VV w�Q$�e��Lw`պ�7u� �܋ �I*��p�%n�U��t��c)ݳ�c����z� ���I�0�/%�J��*�8'm`)%^ݓ+ ���r,���RZ
6�m��t�m�B�=l6�^�,�f����q[
YiX�fB��L���]	M\�YA��1Ƿm<�l'`c6���Z.y!y��.�u��dw8j@�ݍQp�e 5�R�	C�W��3m&; Ĥ ٩�6��h���LSZ�f����4�V�ٳ���s��&t���.-]�ݹ�������	J��,s���2���3rI�����T�+��c��� C,�%� ��,�ZgMl�y��#���c�����`�t�n� ��e`��wnE�\��v�W�~��"��˲��"�e�Xw\0�Ȱ��� �ɕ����{����	;
I� �~��>RJ�=\��Ws߿e`�������:V���v�m`)%^ݓ+ ݽ� �܋ %M�j�&��Qv����2�߹^�{������>RJ��{h;��^kv�pD����Yַ�b�0fRE�0GD�mg�س@Un.�n��ذ�Ȱ��� �ɕ�J� �6�Rv�յ�wnE�r��R��  )U��	�	 Q���
�S��6��`�n��1�'��hԓ��"�ܮRF�K��h�ꊶ�	�XW���&V�%%�,e�� ��Jy��m)�2��{?wt�￿O ����wnE�|�J����J�.�U�P�-��;��`ۑ`-�� �ɕ�~����͋��Fc*9c����G���x��1q�g��w�=Z�H)�9��w.g�������E��������W�wd��;��`�
t�+v�WL�i����W�wd��;��`ۑg���$�J^E�`���E�n� ��e`�ذU�l�J�:C'$#6h,340!���G���� �E�@ΒT�7���0�`��L����\e6�"��m�`�X�`� RCa����L��!n�p��B��������> ɼJ$C)�[E�*XL� �R��I�#�r4�be�L.$"Q��\$2k�)���-5�/Ѓ	� �*�e ��`������0hАI1�02!�t�QN�#����A
�jT0��|� W�r�U]��'�CB��aS���c\��n��/ ;ݨ$ݲ��Un�5n���Xv�X����*��{��=^��X�O�ۦSV�ݹ��(�;�e`�ذ�	�
.�|�Nݴ�q.��t��n.zNxM�߁�Ԗ�yu��v�u�	H�k�E'TU�pN�����vL��{�9\�����QR�]ݺ.�ˤݺ0�Y�UT������}��0���*�VJ��e�Xv�,�r,?s�Ivy��g���v��N�P�I"�X��[���?Q�w{��], �B,@�X	\�}:�l�:N��C��]��X�� �9U_��߿v�����;�"�;���C���R�Z�HK0���V����h��D���`�vH�����26�u�t`�2���Xv�X�� ;ݩB����j����ݽ�?r��잿ߖ���Q�wd���\���G�<�U���R�t�j��6_���9F�s�Il����<��A%]���V��;k �c�`�2���Xv�X�*J�˻�E�Yt��Fݓ+x9���rNw�ԓ|�zMI8�TX�h��H
U\�@���'q��9�l0 �N�mY�ݺ�\�����anї[cl�����9mM�\�ߗ۝�~��9�3�igm���e����e�	�(nձ����<��1<����s�%-!������F-\��Z�z�b��1�q��ۡH�T.�\R����OFn��Z�j�Hպc*B����u��c��G�؜����iy�
��6�gFj�;��<�:y'�'�~lY����nX��gp^,�s���I������������Ч;,И,��!Le��{��p��X������V zJ�C@*
)$[k ��ŀ}��0�L��{ l��Iҷhul�����}��0�L�=Il��zy��	SiDZ�	�|TXۣ��\���}X˞X��w�1�;�(VՕj�V�V� ��ŀM��&6L�-����]/��b%��Z`\�<(��l\�w/�6�A�v��2�%g��G��q¶q�k �0�Ll�^��l��(���c\*�*�ـ}�`giw$A��O����o�5$��Ϧ����Hҥ2���wV]+m�6L�w\0��r���������0�k�%1��Y���ԞQO�=�o�����0�Ll�X7`����f68`l��2��`�%եD��۠m��'vy1�-��1���d����P�.��V�82��'$���Ɲ�ݡ��.Ӷπ���0	�e`�p�\�W>A��� '�Q�]�Bj�հ�&ɕ��s�ĉ#�zy��>����N�~�;`�����U�ܑچn2jI�{?����s٩�� ��C���oړRO{�ѩ'y��f�K�a�;'��wK��|���}� �&V��ݣP��5­��M��L�+�����G� ���?���v%�lk�$��-L9�)FjQ���y悔���Xa�<zM��2�E�YvZm�@��߲��p�&��&�]RE��P�-��7u�?r�U����?{��`���lp��\�A�O5C@*-�E$�ـzy��>�`aꪤ�<�`\����ح�]2�;l����߿t0�����Z�i��m�Z UhT�F�oɄ�{��sRIߎ��͕�|T[V� �0ܪ��/����}$��>Gv�E\,��:v�-'j���WR�q`���i,H����ې2�r
j	?K|kWm'E����>K�X��}$��&�nĨ��5EۦSV�68`I00	�� ����R�1�m�Bl�>�``c��ʪ��w�~������5Q/�t]՗e�l0	�� ��lp����}�|��tYIZ^�"˶`�p�=U���}���߰0	�� ��wi�wo?��f�?pp���t6:��ێ�kL�!8�vծ��z65����I��d�	�"�U�7���2��ifQKR�	G�k.�;ZZ�}U��cn�$���z���v�\�\�lb��O:�C�΢�i�d�����ݜ�����]���PI�L����E)�+��h��ak"-�^�	�R��%��p�K�4���Ou�r�^������{��|ܻ�^�iG]�J"r㝙';�Ξ �;�s7��6�Jh�� e%Ia.aE$�m@>�����L�?W+��W�6\��	�W�tX��]16�X�&z��s������O_�,�r, �[Q%v�I�|TX�ݎv�,�r,� ;ݨ�v�-�ݠi� ��ŀwc��Ɂ���� �����bt�n�M[Xv8`l��p�;��`umت��`�MB�3b,�,� ����w��w�'�ְT�,�Y�ke�5t��Eo7l� ����0��_��A���{�E^W�;t]�����7c�J�j��s��\�Հ}��}�`g�+��F�*貒���(E�l�$��wc��T�}�``<�`{�����n�)*V���Kg���{�v8`{�R9�x��4�WLM�f�� ��v�,�0r����(Y��wWZ�\��Փ����{m��A�⒃k6��XZG ��'�$���۲4lz�i��?�v�,�>��M��ڂCt�e7hl�7oF�צ&�F68g���RG�*W���Nʱ^n������&����M�W( � )�XZ0,��{��j��,-[IEI�QV�ƒ����F$p�7ob��\����ʪ������_ ��=�����6�Ui�~�~������/����x�f# �c�T�\;~��Q̝�Yܮpn�Z���^3�Ϯ�0�lȠ��ƍ��6f�Xk)Lf�m��`I/ �l�`I�����I
�RT���E$��ʪ�q#���`����n�ş��T�o��V/&��LN��;��F$�X��XRM���}�V�ѱ�U���N����{f���;�'o{�jO�#�(da���ͮW9O��Ȍ ��@Lt�[)ݢ�n�[�����}$��$�+o��chk؂�S B�&%�7v�vLM��t�d�eh�ˠ��U� n�rp���ٷLe�0���}$��$�+��~�9�?�{�������o�*6)�.w�}$�`I��ou� �Ixe.�v�webwl�$�+ ���Uʫ�/{׀o��`�[t���)�(B�l�7��E$���� 'v;��$��AIS��)%�M�f���s٩'>�{5$�P4p_�lE2�@��D�F"F�O�w*j!��0��Aq�)���6��}r!����E�F��d�6�S\[ӢL3b�,���	�����@���P��]���A�R4A�9���Đ:MS�E7�6�&E���q� Fy�+M�ā5��sL�4-Te*� ��o �,a�А@ִL�	"$���)XĊ��z�q�����@��$˸���N(a��aS���p.U.0�
��U0�Ck���h�T�B4Hؐ���1"�SX�"��������[RͶ      	    ��     j�rA��0Bj�R卻-�����0Oe�������:〴��͂@5�ab.r�voR�;@�5j6ܪ��Par �+ �y諫�ؚMn��9\j��6 �At��퇣��@to���wݬ&�ms�T��T{[5ղ�a3O&�L�d��N7g��z��m�����QΣ�ۮ�)��-n�<��tE:�vj��-��ю#d���۱��]�f�t=�g\�vPCM�g`ɲ�v9��I��v��M�،�\�!�s�v�]Lv1��֎JN����&�iV퉶����N�T R���		hU�'6&i�),��T4=Y���nU�ă�f�Ѭ���Ru��Kخ�F 4}�۾���;X�q�;����a���ϕ�1gD��s9˝�/7a��8F����9Ø�-��9.6E��������٤�A4�*�-[�@��ì���4�$Bv�v�.
�h�k}�Ѵ?Z�\�<���60��\/Wg�&-��1�����7\�3Ok9�t<r��ِi�tv�쾲uѹ�Ce�9ݵ���L	a�N(J�jݙ��.���۝�F�*XVl9ͱ���k
m����]�����)q����tiг���7�i���,��ncBm\u����� V�.��`�����Z�h�h�x�V���2:��:j���	�e���/-��:�˶��Tt��A؉�K��7����e�����2N4v�4�x�͑�"�,5¯/��a��a;P�pn��ճ/&e`GkY麗x�)Y�&��9ĩV�TV��&�#۰'M�z�g��jWe���t;tf��V��mSfF1[/\[��y�I|`�f���t��[#�]T�R�LB�*<e��F\VcG���<�U���ȁSα�l�
K���3�0uU+u<+�W.��Ԫ���꺮�Y�:\��n���0�m���{�y\��u?(�ʂa_�6ʆ��tDv�����'<>�'���!'F�����j�U!�vX��e�]�#	�&! L����Y���Txxyu%��@�v��sK&�������M�6�ݬO[��s�H�>l'�Q���n�����m8a�-�&��
�e!iƘ���f��0"b�6�Tg9P����`�G\ �mYsV�M�k㉗m�t�] �FS욺��RV��l=����z��t��2���������Ǜ����]\[k�Ŗk,�Rw����f��j�N��{��WJ�bi:T��۸��I0�`I/ ��*,M]45O��f$p�7u� ��X�8g�T�M�<�b�����Cl�$��%Ȱ��*��}�� ���`i+���T]�c.ـIr,�0	#��qM�� �ļ�U�)���V��������c�Ir,lwj�M���@n���I�F�Ŷ��3�鶓�<�a\���1��]���ݥ�.e�$p�7��Ir,����q\,�%���s�g�_M��^U��W+g���ߖ���0	#�~�+��y�0BJ��RT� ���X�\0	#��� ���](�N�1;����������~���0�`~����}�x�ﰇ��FǬ0��G{�RK�>��n�ݡ�oҙ���h���d�#���ƹ��l�p��aƞ�n+-���Y�}Mc�4K�U��`I/ �k����]�����`�z~���6R:����߻��t��H��{�~0�g�<��/*Un�m�4+w�w���$�J�+�U%9����!�H�5��:���{���6]^
�����-ݳ����M�����r,Wkn��wd�YB�f��?�z��~��$��ع��m����j�x���u�q���p�Ȑvʹ�3 ��8���$]�� N�*��U�g�{��,�܋ �8`�`g5+��Q4�*bj�Xݹ~�RG��� ݏ�%Ȱ	]�(�&[��U���$�{�~�s���~��;��, ���;l�]�Cl�;�p�$��nE��Õ��.Q\\�W
��}�`�����cT]�S�l�$��W9��y}�9HK���4��bX�'9�zi7ĳ����{�[.��}h-C�41�x�Bݠ��1 �����۴��5a��Z㛱�湶�7I��%�b}���I��%�b{�צ�q,K��;�M&�X�%��g޺Mı,K�'i��.d�,���9�Mı,K���4���H�&"X���i7ı,O߳���n%�bX�s>��n
�%�bw;���'�1	e��f�q,K���Mı,K�Ͻt��c�P�"b'��߮�q,K�����M&�X�%:_}�z	hV8��as<���N��b{����q,K��s�]&�X�%��{^�Mı,K���i7ı�}�v�M��A�h�O9=���/�Ͻt��bX� �����Kı9�{f�q,K����]&�X�{��W{�z��￹?@  !�-l>�l��h��Ku�v��!9��L9���`&M�2��tv�
/���e�+h��	�*з3k[Ss8ڌ�t��÷&�q<�؇]ۑ	;n��D��y���6�]�°M��ёj^�u��5�W�����lv��4�ɗ0��U٬���N��b��T��&&nL�ԻF�lf�Vt�\��ˠ���t4ڿ?}���<�Ϛk����(��Q�hk	��捭�ĕ+a���45�%�f�-����i���s���Kı9����n%�bX����I��%�b{����q,K��s�]&�X�%�{ǯ���Lc6f���s4��bX�'=�l�n����b~��߮�q,K������n%�bX�����O�����'�{���T%و�g�>)ҝ)������Kı;���I��%�b{�צ�q,K���Mı,K��q�	�b�2y���/!y�޿�&�X�%��{^�Mı,K���i7İ? Aq��~�t��bX�t�����ͫ`65�|���N��b{�צ�q,K���Mı,K�ｍ&�X�%��{^�Mı,Jt���b�q���K�A׫�aP����6�v�c�%DrM�̅.x=+ŏ<�s��ˋ��&�X�%��w^�Mı,K�ｍ&�X�%��w^�Mı,K���4��bX�%�}�I�,�&s.-�&3���Kı=����n�0:���'��zi7ı,O��zi7ı,N����n%�bX��{n&�� �4r��Oo!y�^N��7ı,O{���n%��!��������Kı?c����n%�bX�=�߅L�#�j��O�Jt���=����n%�bX��u��Kı=�{��n%�bX��u��Kı/>�y��i�Smb-���^B���>��n%�bX~AH���߱��%�bX���~�Mı,K���4��bX�t�����|�U�JYc,ݴx��d�c��k�����1$ ݻQpm���ͺ��s����3���Kı=�{��n%�bX����Kı=�k�@n%�bX��}��O����b~����Ը�)���6cƓq,K��k��n%�bX�����Kı9���I��%�b{����Kı>�;O`���3�I1���fi7ı,O{���n%�bX��}��K��2�����V6 H��0j�P��~@ ��M��?~��&�X�%�����I��%�bs/eqf/�LBYf1���K�,Ns>��n%�bX�ǽ�i7ı,Ns���n%�`~���~�鮟��N��~��e+��tvn�q,K��=�cI��%�bs�צ�q,K����Mı,K�Ͻ|���N��N����5��r�%Z�1+���й��e�u:�q�r�	��F�7�x������_6+	Pr��Oo!y�^O��禓q,K����Mı,K�Ͻt��bX�'��{Mı,K�z���0I���<���N��N���4���#���bw����7ı,O����4��bX�'9�zi7ı,a���?;2���&g���B�����}��Kı=�{��n%�X�'9�zi7ı,O{�٤�Kı����&��c��
y���/!���@�O����4��bX�'{�_��q,K����Mı,y+"O�h�����_��]&�[�^B������0�[��9=��K��=�M&�X�%��{�4��bX�'9�z�7ı,Oc��4��N��N����~��ślk��J]�=�˚ A�����y�H�[,8��۞=)���&evcW'�?�Jt�Jt������4��bX�'9�z�7ı,Oc��4��bX�'9�zi7ı,Nc��$��11	e��M&�X�%��g޺Mı,K����&�X�%��{^�Mı,K���i7��*b%�~��z�1�U�پt�t�Jt�O�����n%�bX����Kı=�{f�q,K��3�]&�X�%�{�v�K/��T����^B���{^�Mı,K���i7ı,Ns>��n%�`~b'����Mı,Jt�=���˒��fr�t�t�Jt�=�{f�q,K��3�]&�X�%��{�Ɠq,K��=�M&�X�%�P��&D�aS����?c9�s�m� 6�[ne!�5͠�"yڍ�	�$lmn�-�nL���{X�ѬvEi˳Q�v���(r����i�x��2XMG6RdX�|��y}���̔r�(���Iuf�Ҙ��%L�N�Qnܞ���{m���Hg�@�4��8肣	4fR�Wqt�ݎ1��W��-rSA�&��J!D���4�I��BLD3�����q�?�9����`.��X
���f�u��ƒ7R`�l�@��������ۛVk������:X�'?g���Kı=�{zMı,K���4��bX�'��l�n%�g!y?w��M�ǃ�.���^B�=�{zM��G1��k��n%�bX��~��I��%�bs����q,Jt�K��o�mb�����ҝ(�'9�zi7ı,Ow�٤�Kı9���I��%�b{�����bX�t��>�f�ɚ:����Ο��D�=�{f�q,K��3�]&�X�%�����n%�`~������Mı,K��})�\O�f!,��ɤ�Kı9���I��%�b{�����bX�'=�zi7ı,Ow�٤�K�)��?��{���{A�\�쫝���g�# ��!l�۹��|䍇���v�v���~N�:O~����t	����١$BA�;ܦ�z%�bs����q,Kļ��\��,�I&1�gI��%�bs�צ�p��b �B��R H
�X�1P� ��� y>8
'�ݻ��K{�4��bX�'��z�7ı,Oc��4���1��{�O�w91��-1�g3I��%�b~���4��bX�'9�z�7ı,Oc��4��bX�'9�zi7ı,K�=}.r[��3�Xf�&�q,K��3�]&�X�%��{�Ɠq,K��=�M&�X��b'�߿|i7ı,O���S|"���U�t�t�Jt�Ow���鸖%�`�צ�q,K����Mı,K�Ͻt��bX�'q��bY��汔��`�A����tP瞺w�o��}k �F,�s��4�
��M���.��>�bX�'{�_��q,K����Mı,K�Ͻt��bX�'��{���N��N�ޟo�h|��`��ɤ�Kı=�{f�q,K��3�]&�X�%��{�Ɠq,K��=�M&�X�%��p���.'��BYqs�I��%�bs����q,Kļ｝&�X�7ݺA9�a ��X]� ���>L� H���J�(�1(�Z�D`v9C���a��%��bD" B��*$S�	��}�g��`S�6.�9L&H,h粄���~�|;��B8���ЇGD��
�ѱO��Y���6�P���CkЋ���@�"O�g�u�;�Ak��@�O����2 E"��b,m&$B��C��"K�/�8I'!B$&�}j�a8L��&2���e�tl٠�U�>�o8N�S�ҩ����CX&�0"E����3�|�*�A7o*h"E�U>P'��	��*�ʡ:�C��Wh��b:B#�!�gDМ
)�h uE\�y�5�j��C���DM&�X�%����4��bX�%���=j�v���|���N���1�}�����Kı;���4��bX�';�l�n%�`~b'{�߮�q,KΗ����(A�3A�쯝>)ҝ,Ns���n%�bX�;�l�n%�bX��}��Kı/{�gI��%�N��K}1�Ѱ��S2�[E1<F�������l����L��tc�����au�2�7��n%�bX����I��%�bw����q,KĽ｝��LD�,N�Ͽ]&�X�%�u���9-�l��,&q�I��%�bw����q,KĽ｝&�X�%��g��Mı,K���i7�LD�K��~�0|�W<���å:S�:_}����,K���]&�X�%��{�4��bX�'y�z�7ı,K�Ζ��a,Q#�Ο��N����t�ı,N{�٤�Kı;���I��%��s�4�!! `)W ���o�{��t��bX�'ޞ�Hi~Lġ���Ο��N������I��%�by�z�7ı,K����n%�bX��u��Kı��������(�Q͙�k�q(��Q�ݳxA��6�����p�+3Fكh�1	e��M��,K��s���n%�bX������Kı9���A�},K��~٤�Kı/�~��f���]��Oo!y�^C�����~#���bw���i7ı,N���f�q,K��3�]&�~1�;��V<�ћQ U���^B������I��%�bs���&�X�%��g޺Mı,K���t��bX�'��}ߘv2G�j��>)ҟ�w�����Mı,K����I��%�b^w�Γq,K�9���I��%:S�������\�]H��:|:S���3�]&�X�%�y�{:Mı,K���4��bX�';�l�n%�bX�7��5"7;'�~�s��&s�� �%M777m��%�i�e��[�p�(s=Vޭ�'Ô��۷^�vBw=�6�e�@}l;tv��l/EF�F��{k�q�kPuƶʇ']]�����YcȽ���su��%��G3�ͦX�\:6��ir{s���Ǳu�F��[�]"�\���jv�]u4��x�����ۚ�����}a6kC<!lkRa뫪U��̲s�999�lM�4cv(q����ь�)e�m��f�щ$�{�ͨ�'m ]H�V�c<\)�Oא���/!����n%�bX����Kı9�{f�q,K��3�]&�X�%�}��-�̰�(����O�Jt�Jt�=�M&�6%�bs���&�X�%��g޺Mı,K��t���qS)��������f%�\�t�t�Jt�;�߶i7ı,Ns>��n%��������:Mı,K����I��%�b{�֘��'��K,�ri7ı,Nc��4��bX�%�}��7ı,N{>��n%�b����4��b[�^C�߷�R�Y[��w���B�X�%�}��7ı,N{>��n%�bX�ｳI��%�bw����K�)���>�����΀l��Բ�h˂�ۮ,��ԫ��u7�2��.�6�#�c��s��I��%�bs����q,K��}�Mı,K�ｍ&�X�%��w�Ɠq,K���zIn�&pc0�L\g7I��%�bs���&����U:�e��iP�D�%��}����Kı;�{��n%�bX��}��Kı/����̗���1�d�n%�bX��}�i7ı,Nc��4��bX�'=�z�7ı,Nw�٤�Kı9��Jc�3�i�����3�&�X�%��w�Ɠq,K���]&�X�%����4��bX�'q�{Mı,K�ӥ��s���fa�1��I��%�bs����q,K�9�{f�q,K��;�cI��%�bs����Kı?
����1JL]�?F2�X�P�0�Ķ.�*�ˊn`��ͅ�
*���iIF4������~t�ı,N���Mı,K�ｍ&�X�%��w�Ɠq,K���]&�X�%��N��.1<\�Yf3�I��%�bw����Kı9����n%�bX��}��Kı9�{f�q���k�^O�z�,���gx��bX�'1�{Mı,K�Ͻt��c��$Q�����!�#F �8��E¡TQٸ�D׿wf�q,K�����4��bX�r���1�MY����Oo!y�T��]&�X�%����4��bX�'{�z�7ı,Nc��4��bX�'�{�Kv`���0���n%�bX�ｳI��%�a�H���߮��%�bw��Mı,K��}t��c�^Oߞ���.3�b�Ml�xC�<��bb���w:� �Ӹ�#k['icϬ6ÜL����M&�X�%���޺Mı,K�ｍ&�X�%��g޺Mı,K���i7ı,O���K�n̖��˜��7I��%�bs����Kı9���I��%�bs���&�X�%���޺M�,Kľ�l���rR���3&1�i7ı,N{>��n%�bX�ｳI��%�bw����q,K��;�cI��%�bsݖzK�1��L�L�f�7ı,Nw�٤�Kı;���I��%�bs����K��CTO�."`�m@V�ECb ;� �^b&1��t��bX�'q��S���sYe��M&�X�%��羺Mı,K�D�}��4�D�,K�����n%�bX����Kı? '����%c$#�&n�n�+6��K���թ�8�n�L�;7�޲�t`m�m=L���K��=��4��bX�'�Ͻt��bX�';�zh?�&"X�'��~�M�)ҝ)�����c�����:|�bX�'��z�7ı,Nw���n%�bX��{��Kı9����l���צ:S�����-��n��7I��%�bw߿l�n%�bX��{��K1;�~��&�X�%������7ı,K�>}1���9���!���Mı,K��}t��bX�'1�{Mı,K�Ͻt��bX����~���Kı9�����7fKL\e�qs���Kı9����n%�bX���z�7ı,Nw�٤�Kı=���I��%�bg��h�am��K�  ���;v�n&#�G�EԆҐ�:�y��	��Q���-��}��;\E����<�>;j�K^W�z˻,��WQŇ�qۥ.��{#Y���m��;�hQ	C�����40]G���5��u�[��K�P�k���yB��69������.~nћ\���Yl8f��3���.2�e�41h�G!lyG�l�I��I�{��=����1qym�e��ͱ4��h@v�-Њ�݃��f��q�*]sQ@H�!�6��y?^B�����Ͽ]&�X�%���^�Mı,K��}t�'�1ı;�~��&�X�%��~����Qq]P��'�����"s���&�X�%��羺Mı,K�ｍ&�X�%��g޺M�Kı=�Y�L\b���e�c94��bX�'����7ı,Nc��4��c�a��������7ı,N���Mı�^O����p3m��<����ı9����n%�bX��}��Kı9�{f�q,K��s�]&�X��N���}#8ح�Wy��ҝ,K�Ͻt��bX�*s���&�X�%��羺Mı,K�ｍ&�Y�^B�I>���L,�jƐp�4��6��A��¬�]a"=vx3�%vՁu��'�v���c0�I�c7i�Kı;�߶i7ı,Ow=��n%�bX��}�h?O�b%�b~�~�Mı,K����1�l�6�&g���B��������'��$�*<��PD�@2���M!"�P��>�b{��i7ı,O��]&�X�%����4��bX�r�v���9+��O9=���/!S�ｍ&�X�%��g޺MılK���i7ı,Ow=��n%�bY����[��,Q";Ο��N�'��z�7ı,Nw�٤�Kı=���I��%�bs����KħO�~���*�(8m��å:S�����4��bX�'����7ı,Nc��4��bX�'��z�7ı-���_?����)���8�V��<�<t�wk��8f�s!DK�J�c�9�#,�ɴ�%�bX���~�Mı,K�ｍ&�X�%��g޺Mı,K���i7ı,Nc�ǲg�.1��`�q���Kı9����n%�bX��}��Kı9�{f�q,K��s�]&�X�%�{�z2ɜg�6˜�Mı,K�Ͻt��bX�';�l�n%�p!�*���p��5q3����Kı9����n%�bX�;�'��.q�V��n�q,K��}�Mı,K��}t��bX�'1�{Mı,�1�u���å:S�:_�{�~6e�F���&�X�%��羺Mı,K�ｍ&�X�%��g޺Mı,K���4��bX�'�N�~���&2\�g3J���7gr�L��u�F�G���B۵Nrݘط(�4ά`c<\)�'�������{��i7ı,Os>��n%�bX�ｳI��%�b{�ﮓq,K�{���}�Ѱ�$Cgy��ҝ)҉�g޺M��G1��~٤�Kı?{>�t��bX�'1�{Mı,�N���)�/�U�Ppۛ�O�Jt�X�ｳI��%�b{�ﮓq,	D�N�߿cI��%�b~�~�Mı,K��}+��|LVYf3�I��%�������~�Mı,K�����n%�bX��}��K��h|�HAڗpA�@_��鷞�O:|:S�:S����ޕ��n�1�9�n�q,K��;�cI��%�b{�����bX�';�l�n%�bX��{��Kı<c��-%�3���rj�]�wj9���6:�a�Y�v�\�v[l\Q�vHǈ9��Wy��ҝ)҉�{��n%�bX�ｳI��%�b{�ﮃ�>���%��{��i7ı,Oǽ$�wm�s�����t��bX�';�l�n%�bX��{��Kı9����n%�bX�{�ޓq? �'Jt�����l�r��F�y��ҝ)ŉ�g߮�q,K��;�cI��%�b}�{zMı,K���i7ı���o�M3��
y���/!y,N�>��n%�bX�{�ޓq,K���Mı,�=�{��n%�/!y>������`��'���bX�{�ޓq,K���~��$D���)�$�s��n��I�(����
���TW�(*��`TV��*��U��
���P_�� `�E `E `TP��(,E�,P�Q"@�AP�1B0B0DXD0BD@�P�D�BE`�B!T BT �@�@1B0BP�B1DX�P�DXP�@T!@DP���
���P_�����U��
��TW���*��U��
��E@U�*���P_�P_�����)��L!� nx��8,�������_���0<��6 >��VI�@�      R��@ pi.�� x�<Ҕ�g,(((^�9aOe����>��R��U(��p �Ƽ���#���k){�RyiR���Ԣ�+���79׊(�D�(��#X����S��)E,RJ(�}� <�(�33풊#�h�����L�J$Q2�$��� �ƼQELcEQ2�)s4tƲ��#MIR��($T	@�����JSjOP4Ơ ��  � 	*U� L   Ѧ!7���R��M� i��4�Ob�R��(h A�@4 M"�S"��O2��"4�� 2 �D �4���{B4��f�Ojz���~o�3�Bֈ(�J��/�TEA?䂠����'��29�H(�aPB@��b(��9�"�"���=��������mqϏ����-k[w��kn�o |E]�� � _1� @�F� +P � � ��� a�3 wwQ����� r���n   �h+UY� (����2 Aʰ���Q�� 8@ 	� R��j�� � r�X�   ���{�`2VF P 08�UUP �A��    �@  2p80�9 �   (��f���T ⌍�  r�ظo�[Z�#1x�?H��.���&\�]>��z��v�����f���bcZC9]�l�f��4mthM�6s��;���hax���{``7����9�gi���Ï��*Q@�`0%�����5�Zh5�FSN�h��2a�@�A	i�!���1��T	�ض�5�V1wy�T*h6���oޝ;u�����4�����H&N����)F��5
�b�fU�3Z��4j:�$�
b�`:*��r�wy��m
�H�0F)&�1�YWS��$"Ʉ�
,�	
����HIz�7w�f�M�%2�:�4�+/&��n���0d����(��BΤe�9����y��6;gKpRpBTYؑ#΀��.w��:h%�K$���	z����L!2�.M[�	5r�1f�h�0F��34�� �y0]A�1Ɍh�µ�]��(��!B D����&��gd3����q��//Crg"fA�� "D��� `���"@�P� �!�iK�(Z�R� �D�a�Q-.�=Ӛ���;n���x+G1�pc��^ݳ��8�6����GR�+kS&isv��m��[Z�3իq��>3[�����{n=��s*��W�◱q�sk��s���[�8�9�v�80*�]7%�Fm9uVR��gl{v���<�^Ş�{;J<s���b2tn۷s�T�<Z8�m���ܗ�E�u 	�8Q�m�<v�6f���h�8JRv#I��_�R㎁��j<\{h�ܜ3�n;����}�7��O��O�҉ǉ��ǻpV'}��ڮVJ���
  `6                                                                             6                                                                             �                                                                            ��                                                                            `                                  uK�R1$��$�� �񭪩W�j��)V��@� �]�( 
�h
X�j����/����J�UU�Ul�r��PI&f $��f`Z��@j����U�cH$� �@.�]�VԼ��,S	�Ӯ��M�IyL]���#0  Ne��
�����f`�� Ik� UU�N�2��Q^j��Z���KQ\���`�*�eRr�.C��;jj���Q��5������^٭�TI�.�5TF��t[�]UU.�:�����d$o[@�5U�)�@@�  fVڪ�sS�,R�U[USѓ��΁$��ZzW���vx��;k:狃���hԴd�   I�9ja�5.읝�#+hvX��ں�a��UU^�U��%�R�R�XF�la��EÝ�:�0c�m���U�і��c֮
��H��D�	'n��t^��]{v�V�4�b���������j�0�3�fݻ\��7\m��B�s�-�u�vb��\�]��������*�J�I�k�Rm��������^��i�]�>��}>|�Co�o�yyn
�)ζ�8�z��nz�����c��=^�uء�i��mW	��k;��;��i���هQbڕ���G��P�mv-�d�6�G�ю.�b�\��8�}����E =��͈���B(�=>@p��� L�7 bQT�eJ�+-��
�*b�EE�Ԃ� V���
�q(���W�#��EP
�`T-�0Kl*�$� D" ����Ͷ��� �ۀ ��v� Km��Z[m�!kKm��-im�ԅ�-�ڐ�����)�{�� v8�� l��� l��� l�� l�� l�  c��� l�� l�� l c�0l c�1� �� ��  ��U��-[j�ն�)m�KZ���m�j(���V�m��m�����il��m����<��|{���XP2	� &P6�m�e�|C �t�V;��ҦG�UC�ur�B��2��d� !��uBA �ʊ؅� �)�6�;b�Q2��&��2�Ŵ�w�����<�@��M���՗v��ڗwj]ݩWv��ڗv�ܫ�r��ʽ�Ar�����������UQUUUUUUUr����� ��]]�wv��ڗwjz��5�U^�Uw�^��֪Us�������;�wwx�x.���{������Ù�\�y��$��F�DG���+��b�[6�1GA0�0ie2�
eL1��Ht�����              I               $�              I               $�      �!J����1Ύ����DB�Y[�u��ׄ2+m�h��6�b�;5�n-Y�#el �=J����OV�v-�v*��zNR������F{3jϱ���m7-��v㓵�7lU7++�؎Wi�4n�mq�$��1�"f�@����1�u�s~�  	$  	$  	$  	#UVn�0K[tcD�r;�X���ݹ�������.������軗wE�/�I�������֋N��w1�����7xh!OZS��������R�~����s�U�<�  �B.\���\emٽ������^!,�c �ٍ׽Ҷ��.��K.���%�n�+����yW�O<o��o� �a��;�<;�IfDd�\^�3+*���y����[X�	<V�l�Js���qߪ�w��w���  �*e�ä3� �*���*sp��̮3j���P���̾��.�oH�{ߜ�����M��9�  ��c/ �̘]K���|s~�$�c�&S�E�2�(*yװS�칼�X��3�:UU��D�y�֩\A{�            
����q�#��O=�y�j�cv#s�ǚ����:�$����7� ���E�bT�D�󔃬�;�nT�2��P�u��V�u�v\��H:�;�:�B<�w�s(<�9�<��T��g�$�����:� �}�.��yu���U����s��  ��Ux�,�b��K�+H=�mZ��:�5��U]��e�q*�7�W��H7���.��Ș���<� �t#ٞj�V��"1H<�	���x��^1�r�u�H< 'ת��U�U\�M� 2Ȅ�K�e�XėXAַh;�7����A����IYA�iQ��r�q���,D�A�б��<���7������y�N@M�ND�{}!.�{�A�V���:� �=�@ p�b�Q��4�oUZ��]D���j�{3�U���9H;� ���zR�H=�:�:�vU�w�AΩy�N��y�W0N���s(=��:��w�k�r�Z�o�Uk�<�� ��n7ɥ��f����0'N���(%7kX�^Py�W����֯e�U �t������R��cW���DDr�u�Bn+ٮn��Dġ�@I��s�           ��vS;Rڢ��p�ړ��Ƙ`��$��c�y?'ΫU��  2����I�� 󴃌��{ww{�.a79T������P$���}�����Q��j�q��11h;�8��|��� �x�,�A�){���u�ח��s�� �/!&/$�A��Q}��(DNr�s�x�t]�P{ �5y�A��n3��8��S0�̫;�򊋽���뽵3}��;�j���~�  ��+t\��RH�wԾ�o�}��;�nҧ��ꪵ�S��2�DL�ə��������ֵ�j&fgM��q��{��`�uפN,�$�b2A`A���y'�����{���s�|�z��_W��@�y }P�|����=|J�K��ЪļVN{ ����!��Y�y��/(-�gvV��r���~��  L�0����4*��
�3�W����"��"�|�r�U�U��_EL�V��`��S0Dj>��=&*�����Њ���؊��*�t
��g�e̢�Ȋ����w��#�&���ל��j�{��c���>�  üD;���K�v��ݏq�;�/uUτ�����fU{Ӕ�^lN�#=�y�^�����y��ׯk�c�            S.c"Y�OK��s�[��n9�^�Ԍ�/*�j�\s|� ,Q:�	�w��wzGnfEb� �[�۾f`۶�������ŏ���fa���M�G���w+���{����9��y��� Ea�x�b �5��Vg��wp����%[���g��0��z�o�׻{w��v�ob o}˺"""" �IS%^Z�"�g�����v�7���:�ۼܗz�����>32 q 3y� ӽ��=���3�vn�{����Z{�kU�W��� ̋�	<�n��Gb���	�����9��Y�K���;�6�+�F����0�#�6�����������_{�>��^?O@ K�\��<a�C��̍�����w?u���׹��Q��^�ĔG�vh��f����z߯E��0ӌ�o툈���           �]�.��<ۿT�m��1p6�ϱ�����Yzh�b�U@ �˅��/#���=���_������;�v��)�;��{���-f�U��]���3{ﱉ|��j�^��� �C%�3�]��w�~�|�G1�qs�U��z3Š�M��=x�����y��s�꼹~���/�~��� �s ��
"�.6g/�z�|�ݼ}u�R��m[0FCK33 ��=^�H���?~�|�ew�����s�߾�  c!�"D:N�]�L% �U�^����'+*3U��Ux��;�2�̇�|	|��Y��@�s��S�n��z�p30�興��
�awRL%��w;��S����qq:50 
�52��ެ��禳  0���I7l��ꭗ��s~.p}� �r��5�+�Ig߉�x1
f^f" DDDL�̈�����������;�+�$ �FW7�����0�R�������AH�
���ovV�%u�����ˬ�����                                                         ���          \���E셐(^����J��jN#Q�l�3�-�P僈�ç�6N9�VےL8.�Hqn���s��.,��ݹSL1KN1���Y�@>f�l�lt��ngj�^�6ڊ��uk��ܢv8�R���`G:m)�T���_D�&E:>R�_{��Mj�V�7�            z�y�e�x�s1ߗ�t��R}�s�;l���-˻ɟ�I  30�̍�y�Sϝ����?��`K��S ��T �{��K2���A�S�`2�&v���{���f_9��js�rO|�  !�9q�i�	OS�}�ff_��y���NO	������;�s&��D�B��>�^��� 4�L���y]w  ��S���M�d�U���H{ʬU��I���0�՞��(���;�_I}�u��?�"""" 3
�����"��w��j����y��Y�(m���x�|�U[��2�~�����3?���Yp('���s��y�  &D���֪�V������fa;�tQj�0xY��N����@�U�/.�3+��M51�}m�$�w;�֫�����   ?�l        jR]�el;Y�۝p����:z���2\�*W�Uej��o` \�<C�O鈉;�L�z�x�����g����C�k(!�Q��P\[�m���󗙞s�V���}���  �1^k�D��Vm>��7r�.lg�|K3ٻ�g�k���TX���`d���ϼ���Wg�>����~�2}� 0"AN����C�w�������r�3"d7uMf�$|�<m���40�7���`�6���� �ꧣ��W���w7� �d�-Ir*�#1�2@qs�X
�o���.;�����߬@���|�8����+��]~�}����<�?� 	$E�_��Q��=�$��S�^�
���s�Y3 ����wo^��Y����f��z�uU_O��       �    ��B�I$Kc0���&�K���KsB��&d�j�����  �"^2�� ��$�|M_Κ]��	{�n&{zh�u)�B�<_�E��,۳W��֫\��  ����̳�:���c��|�32-��80}W\�~<�vQ��/I�|	s��x��u����]��sZ�rg������ $�2H����UL�w�:�{U�_�o�ZVy���W}y��_{Ǿ33� �b �<�����}�߾����{��/"�G{��#�58�%�U5�CܢySSȇ�:���(zu^u��=��?p�٪�Ȉ�� r2�2챒�7�ous��g�(�ox�V��9�H<�@B�6eVWWn��z|��a, hf�3�o����=������ 	��(.<Y��1����5Z�ڝ�S�=�����35b�f�%�n��C����_�           ��|�rm
���5��к�7�7�hT�1��	ְ]���T  �tf!WS/�������(�q]�N��чB���kv��N���7fK�Z_��Us��|�  fa���)i�¬���<�\߿U���i�fb��,����������v����*y�/U��_w� �I-ɇ�	�
&��uN����=��닃[>f5`3
��ɟh.�vf�Fsw�����{�� a�e��U���yX��/�.#7n�u���ي��(�A��n&��4�0���.g��b=  �E�$�I��̯<����2w�x��v����.pL��ר��u���eL����P�3?3? ĳC����"�!�b��;��+�p            U$I� �m�x.ą�	좹ucx��;}������T 2$�鑑x�������т�U�ҙ΋�3"��㪫�<<���6��wϿUϹ�9�w���8  ď �d��� �N�
���^�<����O�n�>�#f��1��ﺊ/}9�W����{yW����<��� SK���'��C�=ջԕ*�]\Sܭ����K�af��?4߼��dG��B�k?��EZl��|��Mv��1ٙ��w� �f"^(���Ȭ�xqG�-��A�_n�����MDI��~-v�Ғ �"an�qi��ڌ-�0�!���Y�bl�f�v��w��� 
��1�^F"�d�p�ZV'3u�C�1I��tHz��S�Q[�Z���e!/�$鮐4�ȁT�ۅdiD����B�����
 E�&K �-��v����q�݊`Q`,KC00�{vp��m�$Y�(��E�b��"���Q�����2�*�YW���6                                                                     ܬ�I&j8ۢ@�Tx A�P���j���q�^[;�r�[h��\�;׮�W�Ԧ::��Au�@qrE(��m����%��pr�vks;T�˗�� ui:�W=m��;v��y���3Z��r�Ȇ�-m�]��>��	��
��.&b�j�2�A }����<�Ѡ}�M��|E���������1�c�1�           1"�]�Y������Lh�����dVfR� ��.a�?�yx��Co��i��;�"bwJ1#u4���'���5��E���M�x�H��k#�������C��U�e]��U��΀ $K�qf!$������hu&�B�a9�le�>O�Ë������0�{E�과���	��1R]�"�
�v�(hM�9�/7_}��yu��ˮo�` �Yؐ��Q!&�$�2���x�����(��<l�3�P@p�YH|�<dHf���YO��	�Fb^���:/��]Y+/~eKח[�k~�π G���B.��!da�4�!�\I�By*���pĄ�E:s�8�#q$b�E�k���������C�a�a��3x{o��'��$E!��� x��  .�.���"�&�u�͛-X��Ns�tho&�F��s�눲�������t�4�4F�(�3tT(k"%5�E�|q!�0���D@            Ud-�u�J{=m�v	kN9�y����z�M}�-�3La%�������뗗�1z핔�!�*�|�m�x�8��������"���l<p��o�y7���k�^޹u���$�������.&����M��-)g���0,��;icd�����j!gzsę�����k�deW/�)Z��9y���s� �*�����8���53�	�x��]��a� ��bLD���|Qp�!�8��#>~>H��~qv�}���8_y_]e��.��3�  #!�x*	x�v�f$&�`�Gl�dn� �-%�狃DIj�6�ۧ/��@9u�w����0Q�0p�O]�9<�����g�o� ,Z�/��/#15�7y���|b��D��S�Zg�bp�F��C1Շ�(�g!��(�T_�H�L�a�(������U�j��^���j��      $�     WQR����-V��3�i�<5v:��T���̋�ir  �Ru�^"N6�i�*�y��O�
���ff!b�6yɸ�B����A.EE��:��J�0�-d)�]�~_/^1|�k�{�� $�r�I�	<di�BH�H�"�ܔ]���M�����Ӛ���@7��"E�pEJY��.a��"͑T�nw�x�����U�O~��5�ו_���  �(�xI� ��u�v�(�/~��7SZu;Y�v�:o"9g)�)�'�AE`A������n�n��뻹�������s�������o��vw�7������C���RVB�,`V����1"�;��++Ӄ*g4��0ƴ�T0�+�!r7c��0VD��H�+`�
X�E�"���z��O\�F�.����l-�܍�lF"�ꖿ&M�j��
|��o|�{p94q	�v[�`8��:݃���ܘH�����7��`��턠���`h`P(P���`PB��
B�(P�!�����
40&�@�B� P� ������*`}JQ\�A6��Ǿ�����VL���7SV?,��@�k��)6R@]� 3
\�Z�dY���+��#�Tc� ݿ0�1��C������CȾ	���8�S���U&�C�tX��L�_[,�|	y��F���p  ��\�\�@���p�$�DLÌ:�0��V!��MG���Q@�aaEZ_����ⴋ�6�Y�.g�.a����ERo��>}��           H����{P�����͓'lHq�\GX�A6�.��p� p�KU�C$U�Z=�9��s>M��d�4ET��HE��p/#15�� �Md*��K��$�&Q#���$aH���0�`�� 	�Ɍ�f�I���y�_���=�|!̎�ʆ�4��6��=����!G�:5܈���<���F�;Y�N]����E�e[=� �)��r*�%g+�s^]{mD(砝�&�ƈF�!v���P��}y���8�3�RN�DBj#�I����߹����<�����  �ȃ�TAa��%���v˭�\O-GI�ե��:k<j�YYV�FFb�/P�-���0�����r�ow��̮s5�y�� �2%��L�Bx���k!�v�+ʞJ� +B%5P��ޮ+�&��0��(��E�BO���vk��Z���MQN>�f`�_���           UUS �Kă��!T�/A���[��P���nm�  fd]�dR�v��Y�i
���u�Qs�	sCu5�����.��DU&�&�7wp����f���l<b䔝������M���숈� 	X�).-rE�es����ח���B�.o�j?m0{-�����������8ա7U ��FbSaI���]��z�o�R��V�U\��� ����%����מ�;���)C�xj*FzBw]��1�S��C��i�	r4�tw��#�)��l�Qj��ƹ�y~^����{�>� y�� �p�D�t�j!�]�������|Zl"�e�fC*7�T=ఈ(�*A?�ä�^!����CF�7���H�z�׾�S^]I��  ��AxB"
$�] �/dIFe7ug22��hN�;��Jw��*e���ݕ\
y�t��j\��9h]�&	����*�By���-(5���,-�QU  �翿�����X�P ��]��z�78�Z֍M��Z׋�-�F���� �4�FE(���hrL3'���#��V��&s����Ih�r;`V �b�,0h�����K�֦iz��@                                                                  
���������j�9�,Q�&�U��][S�N\���]ƫ��mV�c�g���b{\�	nnep�r�4����<��R�i:4F�)ڹ-��\"7�r����1�@V��gcc7m�]V�^5L]n@�`޲���]Y|̀�b�UVv�\��+U��W��U
��             ��Z;P��b�gCn�|8�>o2%ZB�Y+-\�UZo` �@�"�Au|���Z����
��D�u�ӽ��R4����d��R�j"�i�0��g&Fw5����ۯ.}� L*f.�˧x%ц�D�j"ޝ����x���ff @�g��<eV@.��4�hQeY��f���KQ3��hJ������+<�M���  BH������'�	���Fh_��"��BxP�ȇ@z�����h�#�����a�0���	�m7(l�t�W�+"�aj�����W7^޷u��.����_�3�I  �Iᓼ(�S��8d�XA"�)��K����0 �#�Y
|�	t�t�k"�- �٨��YT��w� �E:Ye^fJ���/|���뗮u�� ̈]�;��x.dNk�r�!�"���P�l�d`�M�=������ݗjC�@.��"�5�[Y����D927qڈW��W���~���             �l���.���:�Iǩ:�n�nM�q��UUUUVH�v	ol��Im>5K���JF�"G!}Έ�B�N�E�HxM�Iz/��8��e-N��{w2����eWn�������߿z  �[%$I�)is<��[����.��pK��+u�ރ
+�8��Qٸc���������#�d=s�%�BKQ��5����I���w_{�|�W>�� fC2	b�.�wSy�]n�ɟ{;�J;���-�����0(��,���f3��;��5�C���j�k�'�R�u7�\�.k�W̯����� X�:�'��^�jk#N�D<��%�Y�@YI�oh�����U�v|Zx�YPa��bi�G8���3�~�H��&�^:y{�5��;8  �$�Q.�eG�.a�Т��0fqv��~�tdo&�Cu5��1��@$�8GR�Ȓ����S���m#�5�qS!(Mg��l"���yZ�W�U��@             ��K����1�r���X{N��.f���7�� 2dH�qe)�HҦ�{�Q�t�r�v�DBl"�7t��^�CI��"�����Ql��z#^ߋ�F�#u5BҞ⪪���G��������jIkz��K��+��Hff�C�
,�Hy��J�ْ�
Rs}cw���M��	���)�;�7�U�6p���}��  	�a%&^.�GpXE��,���v�.S[�Tw�{��n��5��|���I�`�39��9���fff[��p����%��p��yO�ʯ�ϐz���fBC�uGy7��OU�.Sx��vÇ=�pGn� ڇ#�ǯDDDDDEU�)'b�"�l�������]�JM��ъ�:l�#u@"�f�P�DJl�� �Vqi���#��`��k�u�]ʆ�.�Ɨ�����؈�� �¯2��aw/}�o\���v���:N�Q���6R-[0fb&{���\FzP&��=�ГdQk"*.�{�!#I���_v�pm�             *�7L�)+�*�;^�-rٗ�S���qp���P  %�&%���e���)������(���N0�8
##8���$�:�v����)Ԏ��B��C��^I�_���k˯7���s�	$�2(2jLʍ����yu��K�3��>�
.�Q����)�q�H���%#H�%�"yU�E����E�=��{�[�����_^�u��x  ��K���9P4��e����s�b$`?0`E����4�3u�$�I���]�{�xC��|��z�M��v�8�ܖ��v���v�{�v����߀ L�$�H�)�7]�5˯}�yu��IA�A�!U��ha� ��>M:y&�q}���\��Ij#�@���31�on�I/2t����GS1  L�y�����2*�J�����Y�@����7SYi�WE]5�J�|���M����Ģ`�-"-�8��[e"����i;�a	�ӡ����@            U]����H�/#����S�n�:��A�Ϥ'�~Wʪ 2FeȬ��.����>���~��3,������l��+!"�=��*"F�6T�>�C���v��p�]��7I��Ak#��2"""" 1j�*�j
���>������(�;_wJF���dw!��3�+�) �F2�>(Yn��;�A�4����xמ�r��׾ySS�{�� 
E�2d�0�����2��9u��7�Rl��fJ"�*��]M����]hI�g��	;��Z���	���aH�8�J����럹� fB�%��^ �w��F�3�I�j�B27SU!�#e�+��FGH�.�Ş��/"�#��\W!���0�~Ɂ�#�ڄ�l>�;���z  ]��%�&dU�č��#�
.^y�]5�4D0j
h���-df�En��9e�<!�u��U�ɞ7�ވ2��H��޴��� �$�� �߽��]�o��{��{�K���rt�B�Zv`+�p�H42I	�:+()�s	U%kR�F
#*�
�)Gr⊖؉�B�`�ҖJ*,�fnmؘ�CD��6                                    ��6                               UW�Z�@���e��+	"i2KI]u�ړ+��:�eڪڳ��H��:�6Ү���BW�;�m���Ӯ5��ns37Y�)���7b�%�8IƟ[�[6�[cN.���|�h�o>,��7]q�{[`J�,�c*�(��)|��M�B�:����־�:             r��˪e�q!����GTw��  �$���ċ����I�8�L�mߋ�C�I���>����Y��U&�Bȳ;������i ���������AJ��*��y�� 2�#v]�"usu����3UHi���$Y����6��+~�#������RE���PӖ∃�x��Om�u#�I���ڳ,޴��Ij��yur*�]{Y��W�^�Y�;C�#ux1���!0f3��
�V�u	#���X�x��Ϸ�\�Z��	���7Ek!�5��V���π �I2E��I[���5R�����Pو]��C��6���F�j._����MW@.�2�> p����*ċ�qF� f!��� K�̢�h*�ؚ�s����.�=u�%���_��Jk�3ʲ�P�Ka(i�B�{ӴG�w'"��ie��3����Zl�s��bo���X 9舀            ���Yz·{$���r�n'�q��g�����d���Ɵ�UUUU�Wd�&n�}{���� ���]�+��5�?�1Unϴ���X~ 6{_s^'�혃���>{�i�(�6E:b���4�7J:�ڭ��π 2"ٙ�eȼ��<C�f=�"OuՔbF��<���<~ �O��"�N!�����2�x��]�r,��و����N�`�2�9~޿z�  
�K�c-D���k	-X�ן��z�o!��.{A.&N!��<'�B�rk��K���S�9�E&�V�P���g���Ŷ�5�Ǡ 
"�cwRE���,�7i�+8������A��8�k�x�nk���5��h��8�fl�n��D����	�?�t��T��=ƿ���@ 	1D�̻��DU�Q#Hsbi�8��J̓!5��G�GEm�D��q��ii-o|S�l�&SY��Yf<�#S.3����mWkZ�{��          UUUUU��c$
��Z�Z�W�.�m�m0�O>*�i� e2I��W3^X�\GrY�7��7y�1-d*����k�*X<n8���%�ij#u5PXz��/.k��o;tϥy]y߻�  $�E�u���ev���g>��Z�{�f��7SH���Q������^q7] �Bmai���dB��b$w�����~��<�g�� s���B)���1��\ݦ���]F�n��C�ः����u�J|"!��&I$0�$w߾���}��}���y�@�P�<Q�(�G�X@�GP��aD�0 ���6�<�fjS`a���я�\t�UM=��MUn4�`��ϋ�{��BN��=��� ��]��"֋ɜ���F�k��T��k�*P㒅�{��
$n��XIj���wNوQl�>�� �n���p.��-Dn�v���uUUUT�Yg	������qxv��8���m����eu�-�����	�p��
,m
���.v7f^c�^���}�ɪ�U/U]��             Y.&H]��mם)9M�CO[;l��VWզ̀ rR�e�!;�b ���γU�
��3��zlQ����]X-,>a���&ݻ����� ,�F�J�]�ߛ��Ysz^
��@`�O{ngk�	y��̸{��)�}ڬT��
���ݏ�g�x  ˆ"�p�ɑWW=�ɛެkPC���ݪޗyC2b>�`Y�3$`�l��Y1��6kj+K��߻�<�O�  2�-iy�"
H=骼�r�������"�^�4��Q�Ҏ��+��g���0fk������bW�+�Z�I���  �	��x
�A�xdH���W�����;�5���fVa�
�x��U�S�o�}�o���*�kZֲ���{�x             .*ap٭����bq۶�D��lĚ��S"򫼪��UMUJs8  e܌��r�y
�c���rM��!A��5�Ye���]ђR+0dOy�ny��<����7��� ��)<'w�\�Nf�ԙ�،��?z ř����qw�����E�zߴ$��;�|�O~�]�����{���  &D�XU�W�y}�y;Ͼww��������2�ހ@f��튧N�ê����;��w������  B�H�
 �{�z�Gz�p�U�*7���0��g1T�VHb|ϻŀ� �,Ny���w��}� 
d�� �]�3/�����" #�0�ݫ����|j�f��4� f���1ް�+��'<���
�_R���$�� (�|߭,iW�P�������kA�O�`�'մAEL�Q9�L�ZD`$U�Ph�(�"��, � D@EMDJX�/9�XH��)�`�"����$d�A�"@�S�.#��E���q���*��"Z(@ ��`� �!�F��o����{IAP>���#�&j�w���޼������mD?�#Ƞ�P1��D�@? �iEw�`����� A�}�#�� �=ח��B�����tC�@s��}g� A��u�'�D�pDC�'Oq���1>��@>�E�!���"��J���������?JO�R*���PD��3�1��>��O� �$PPb(��2( � �A ��"��wƏ��#�i
W����8�D4���U�_�\9���PT��ߜ��4B�b��~�o�Ѐ����F
F#!$���Kd�D�X"$������Q)��0R@P $$1$" ���� ��PTQb��H�b$R�������1�B0B !�	$��Ȅ�$R��|m@"0� �Pw���^ep�&c�����H�>�� �P�`�����~���?xO�I��|!�9�����C������� ������?�>����G���gĽ!F��W����}&�~$���ϗ�~'ݏ��"����������2~����s�����&�/�"���>�E�~����O�����Q���8H/�Xi�R("�	�$!����3� �(P���H�Y��&`��*��":4���n���!��}�٥@EP|��B���PC����/����ꀪ������y�q�0�O��O���{�b|�� ����>�����?(�����TP�>��=���|��O������L!b!��҂3��{I���:�^=�:�žS%ɿ��@E{L>����S����pװ�U�T>�z��D�}�O�#�=�y � ����/ޜ��Lc�� �(|OgV}�P��j��gp�z��_�{�@:�br�w$S�	��