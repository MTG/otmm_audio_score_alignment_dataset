BZh91AY&SY7�@^�߀pp��b� ����ak �	  P �    T � ���� �4( �
k*����( ���B
�E
BP
    (  D�U �UP(
D�JT�
U"��%"@   � J��   3�z���K������ԬzR��R�yr���8�]9:S�ܥ�{d�8 �R���@p�0�>�N-�{�� � ; >�:��i��@  ��	   c JD�wݶ���x�;ۼ[�Z��ޕ{rb�Nﻮ�u�U�wkOx� }}�w���<X� �7�uť]�@�ﯖr�m{o6�Z�����V� �k�n���;�6�����W���@D  � 
f� ��Zۖ�+�o/S�W}o�jp�gJd޲��|]�˥z��u9� >�ﾙr}޹��<� >��k׮�=�^x>�G{�N[�s������=�^��� �j��9μy�����/7� }@$*UP@   ��j���)˧M�k��}�u}�.:� �����r�Zw��YT�o{R� 2}z�y�xi��y��O]�R����}�w��<w&�����Y�8 wS�u��wT�&W��OK����*
  (P%� ���;�����d���ۖ� �9;�q۷���:��x��;� ����es3�    �}��{8�U� C�T��ٗ���ޙ� wJs�T����i��/'��      D�"jm�R�&&� ?P�R�4   @D��T�      تT�IH � �� EO�
&ڪUP4@�4i�R%Id��4)�4!z�&�ȟ���g��������}{���U_��7�TUU�"����UU�����$�U[�L�UU��I�����g�Uo�%����u������~l���˾����?����9׏V�S�˭�q�5�I���s�����ۂ&*�O:����ִ�kYμ�{��<�F����4��u�m����_sO��g�s��W1�[��ͯ���.h����[��j�Zߝ����g#:�[��
�s��^jb�٣AdF�qk�iM����+N��u����n�&�=Ѱ#F:MFj���w���O���]F����Iw9�'����v{�4^k7λNxBfa���E����Q���m�|5��;��g����l�}ș�v�s|��TO��3M�x�m�i@"��|���:M�ܰ�d�.9�G�:��J�V!��k*^��|�����Re���c9i �t�c1�f�E��j��Χ�{�)L��ĳ16N��二$�BbrW��>A�j����f��6�堪<�p6g�<�;��yى:�% ��	巃�ǁ����&z���9�y����te)�l��g(4�`�� I����F��f���9ӫ5��f1��Av�3E�$�!;���t�5KN�e�y�:�og}��ц�#I�P�9	`EEbe$c��bb�3�kBS����8!��#K�G��|����� �MG0�E]�ְ�e�Q���Ewa�X^{��#���2Д%	HH�'!i�"i���BP��Y�k5&�A�KI�rr�\�,8a���w�0�"2L#1q�MZd��`I�Lã�G=�~:������Y��<�w(����|� ��h���z9���g#�u�wV���Z��T��V�Z;彑��%�o�pv5����u��M�O.�g7�Zl����A�a>�Q�j0ӗ��k�p����Ԕ��nHfY$��K�r���q���Ύ�ι�5�]��p��S�o=�7�te�i3V�ݎ�;�6u�t��~o(��@a��%$P���#�Ώvp�ضWDh׽r��ۏ?��r���,3�=5���fO0�CKW�n`��ڸv�n���hU�;�w�n�3�'�wk�7��u�u`��`�0�$���.܃&3�$�,����:My��h�2�=��S�QTFL�Bw���s���A�Mf����%�2�2%�c&A%�14[1*2�9:5b��oif�ۮ��ѽ�:�ѫxtS��<,3[�Fn)��KK���	Ѥ�֭[籮���`N1�O4��p�tw�ηÁ)W]��q�1(JM�C�ds��-�oGVy���=t6�0ӭ�N�2,�# �\r0���<ֵ�V�N:�Za�J�*��&N壷�����N14NC�����I�r;<���G�kwF��}fx�xgX�''4s�9�<��E�a�]�h󣑇{L�Ώ���G���"�փFsy�ǝ���F��m��xg�a��g=߆�.q�|v����U��:��0�}u��+��ua��j��on`�&���7	C��20�N�K̎��I��5�f����h�5�f�I�ƫ5��FZ��MK�F�0�Idg�Ca��G	�'iL�P�"aBL���3,C!)1ʌ�"���1�Y�dDk���60�pg ��L��!BE�M	BR��f	BR��6ٙ�������)�NfFHS������,�5M����-g\�i�k"����y�0"��`Υ�-m#Z��Y�� �x��:�3��0�,�0����{�w;��7�����\�3y�zمט{���r�2[ys���pah&hK(�H���[��g:�:�u���a���h�͚δ{�}Z����͑�)<�<·�7���Pf��g(�1�['A�5��asz�7�k����,�
y��������tZ�R�ۂ�,MH�u�j!=�c�N�K�0ud�a������<����$4��˷ڱ��{���>�3�[�]ʻ�ԇ2�<�ya�����y�ML<Pۑs��?��I
k������F��P�;l��Y�c�rgu��~��!���I�.>kid8@�$M	D1��$������`�S@LL$bXC�X�.Cîl�OV!�t�t����	�X&�`w&�C��ĲLJ�N��w�.����M�K�!(�)��F����$����C��[��u��a������Y�0$#;}6N߳���90���bf'��>��8��L�{�y���8j�f�F�`��:�]��
)� ˲Նgӷ�3[�5e�偁��^t�4�M.yj�mBPh�1�Ajȭj�sM����ݭD`kY��E��Tf�����r�Z�P`x���F�t<1q���Z\rqrf{�S���!��|�����'Z05�f������1�kN1��kW���:�j��?����7}�ۜy�H��.$����������6�ܴ�����Vs�:��zMA�l
��a�{m�Fp4x����7��Q���2M1�t`Anb0�;�{���u��5��<[���wZ���/<[�I/��}��g���u�{׺�=�u�hò���=�(�Fs������]磧R��i�u���#�a��	'^:�֋O�kf�9����L߇�d�0�� �����ora��1%�74��f�j踦l��ƹ���]��@{:\�tu&'���Y�vh��x�(�駹��Ͷ���9�͵��s�]uv�tF�4j\�p�k|�˚���r�N�	��%��{����h�R���t��+���.�d�U	BrՉ����-�?LSg�<o��i�ؚ���r�{�3���s�z�E��D�l����w��`�h]-	[�p�ĥ�S$30�=���P�A�Fs���|.��.��a��q��٨;�^�h#{�i
�P08���/z���.0���&Z���#T��@��~ixz�Sh��(g˙�X�xg2s��v��1��q�lf,��H�Yg]��5�1<�	���q���o��6�S�E��I�7�y�4�d��<�ߵ�;�ї]w�3����4�;��^�3�p<�����������1#�4u��<���[�YfuCG�Oy�X�2~1�ہ���ɝ�?t����,Ɇ �z��;��Vuzw�,%�Ȁ�G ��̖(0r\r�5N�Z6BPd���C����J#P�'4&�%	�0J�	�w�9��14�1��˿;�u�#�nӽ�l�ўz'���m�yٝ�¼C@E�T�S1�գF�(J��z�k�8e�s��r�٤�cC�rq7!�����^�j����>Y5�m��0�4�6�ݎjjxj�Q���Y�܍y��!��Өp2�\�l�\r�2d&�43iq�i��z������}���L�6�c�m�{�Lg&�\3-�7S��+V6YIao��̂5�ݑ�ф�%3��F���]3�ve�n�ᮍ�̻�kEQ�Q�z�����Sם����w��Xh�X{��U�3tg}`hr0	���j]i�A�;�M��;�;��u9M�fy�cћ�5��f+���zd`n0ܚ��k�:}�_9x��pjʌI�6nM;&��]پu����MIA@d㢈�y�~]�`]�j3�1�!���	���qw��EY�fV{y�9ˮ��8���w����3LŘy9�Dn�ǻq{�t���a�asG��g3=�;�湛��-%���	A�#{�*�5�e�<I��ݓ�[=狖�"A��s�M���zk-���Rj�7�w�y	�x�b���9	�O-����\O`����ƌ=#_pXkS|(�-��u�|�՚�����o�<�v.0~{�=��z�sϗl��-�ӹ'��A#?s�E���=Yq�ۻ�<�	�*M�f�(J2ӳ���v��i��a����Ͷ�Z&�9���RT�C�f����[��L�3���mG�gb#[ �3VWwKS]��|��-	�'q���o�M]�u�Ik��#Ԝ�>����jo�a�=;���ν7�}���S��[�ÙZӆ:�]>f���R.�}��ϰ����y�#��O&DVs7ֵ�7S��t�PC�J^܄�CP��o�g}���h�����S��X�1��%9��~|��-��0��v��ټ�H����fs���xfZ������ɂ��=��7����'\���LD�l0��0�ٮa�ٴ(��yuվO[�5w6ky	Ӓc����Q��ךx��ݹ�}�ו��4��;>��Zi����0��<�ΰ���=�ӿ3�'[�:�zzf���=ˆw׆����%	X�F-�����0{	�{M&��8	�`SnLMF�w	���Z�&�u��Ow�����u	BPh#X��[��f����78�ˎC�d�r�F�hk��|���ȗ�wgh��g�a�����;��(J=��y����J���7�o=7���=:��s��y�g�hw!��*�<L������6�o��i�p4�Ltw&Df�������|��J�2����ʌ0ѳ.0�'d;C9���;4s�7à��%��G{�<�3��e�f;�4�t���hx��{�xxx���n�4yf<Ma�M�4H������n��v����{��gf�ׁ�*BZƓ!(M�k 4d�9C��������� �Ot`DgN.��y�):�6L�;�z��'p���=޷᫣lo[�Z���Ay���!奵�q�K�P�˷wlݚ��ތ������^y�z^k3М�&Rd�R`Z��[k�}�L>����m�����r�_�|3������as��qr���a$�"ǂ}Q��y�͎;����=��}j~{h�h��ǋ%����~b��ڛ6�1��������﻿_���_UUUT��U�m�H��      7m� �l ?X> ��+bk0Ͷ$ $8p 	��Y[e���R֒�\�j:f�%M�;	L`	� >����H7m�m�lm�Ž%n�i0  @h ����۶� ��� R�����^���9PU����U`���j��H֍�i0�� �f�h�a�� 
U��j���ӱ+���b��y�)-u��į&7a�t��/m��`ŗ��*�]��#��ٴ�$��"xl�J��לI�9٪��j�:���[�(��Z��
�L�uJ��^��әXv뀤0�]v�,�[�-�h��I:n�Z�:'_Y��%�n�:��!�8Η��ӈͤ夒Zi0.�k  %6u�� ݻm� �ؕMm �*�UN��YP6����9��ﭿ|l֣�C����7Y!P*�y��Q���*˷NZ��1TFL�*�,�DF⪗�e�.�Ļ�Unդ��3�J��]\�,����#R��a%���N0c�n�W;m�V.�x��lqezʵtq�M�ڐ��	���}���S�]:*�e`A���������P.����U��/!KI4��S'"aϱ�*�][vSX�8U��H�^��CvԜm�Uz��o���	�b�#m�}zK~�`���Tw$�R���]�mH�RF��4��Rݴ�-�`C�,v.q�`�4n9z&�A6&4⃍����g��M���<��qi��a�{`�q���W!��F$&��Z�NJ�@KO;<���
 ��s �����m*� �;l	��Z�G�7U[��c-���^���N �W�.�K���j��Ԭj�b�r�Gd:ݵ�(OUM���GlKK�6�P�1�����%�F�t�[��>  n�m(p�T�-zU��T.� v��(�jQ�m���Hl��V�"�g[C�� ݶ86Sa�l�0kΜ��p	q  �k�[q��6�ֱ��m,I�l�@.�-�A�͇�$��`*�IjW*��5�   6� ��� pIz�i����m�[$���l��b9t�� p   p��l��t�Sa ��� �X���*�J�J�r�N[q��l���f@��H�{L�    �[bZ,�I[n�Zt�#X��m����.-Ӏ��@ �m�$  ��T�V�j�]�X*U��@�m��7��֐�8   u�2l\\��m�)G눻�}[��6�    np۷6�h )��`�M��`;��@��   �$ m�� d6��( ���-�� ��ci68��l��j��IB��b�J�U)x	T�:�  vٶͶ  m��}��   �H l 6�u$��b�� m����`ii�3m���  ��] m�]5��:�   ����� 	   k� �I���n��  � H��  $h� m���j�m  [@      .J �]+ZKj�� $ mm��m�n��  ��cZ�'M�  i��� I$��`    m�m���i�^�  ��u�7d� ��5�amm� -n� -� �� ����6À   ��-���l v��6Ͱ   [@  �k: H  �@�0�ޜ[p	 :���H�Kw� -�v�G-��h�7W*ҭp�\���Εˀh H� �Ԁ �[d��J�HM@P
�]Q plm��86� �8�mH@�s��	��      	�鬘� ���ɶv��%�z�cU6  lx�t�ζ���}   6��MoP[��R]Wsl��{k��X�%���@m �a��� m�` ���j(  l�Jn�� p�3VÆ�� �릶�h�tĒ��� $m8�.�� �7l%��k���ۛ�n���:I6Zv��@    m��J �zO�[S�h   �ݰ ����] �.�   �m�    �`��b��6K�)m5�Ҷ(�l�[D�l8y���B��66��ڬd������S��cV�� ['KvP �]fmh�m��HKin�8 �断��i�ڸ�6�-�Z���G-P��m�u��`��n�r�:Ҝ7E <�1;�k4m4�p=��V��	 9��N0�r����ݓ����N�Qq.1��nq�!Amubh�[SoGNU���Ie�+ek��t�O�z�]2�L9g7r4����t{m�QQ�b�8�.̝Ō����G�q����%\<�4����ga2��`pa�Q�Y3������h���UG���`�
�𭧜�z�j��sV�94�N�S���=I��+�(�iV��b�vyrD��;�n4����g���'�l��v%:��Ų�9.�/T9Un.7N1�U-Tn�T'R�\A��!%���v���&�y�V].�	��'siΖ뮣`��\rSJ�U���|w�m�&���Z^-���VC�7U��Sl׭Ü[b�5�aN��j�k�k�ӵt��qv�n6�ޠpZ�EH�s�l�[�׷k �
�۴��y/C�-�m�Ŵh�m����-�m6`,7���m� *�u�n�5��5U�K�no\�r
� &�d�I�i�k)��΍cY� -,���hkm��  6�N�t��i�O^�l�]6Zl����n�i�^D�'N�a���jv�6�@ �vY�:v㭮��rUS֪uK�R�@;m���� ��#���܃U��d鶒�D	�z�ݲ�Z�j�� "@,mU�92�FJ�,�*UUKn����m����`�am��rT^2�s�ݞ��zZ���Rtuv�������1� ����j����+*��)-O[�%:@�yM��U�;��j܊��\��t��}[�A'�^X(�7 V����s$�&�[�v�q;ƻ��/�'����f�`���㟷�+&պ�6�v�WK��NՍv���Y^�<=��e7\)H�L�;Y.��m��f����	:@��[�lܥ�  y�bަ�WQ�l9eX6i���e�u�6����m�M���[Rμ�L6����@�uT݀��
 m�ԉ�-���i��m�o+ p�:A5��.ـ�òm���6��[x��P�4�.̡1�:Im N  l8lݖ�lт@�`  �9���8�ki�m�6ض�m�t�`K(�E��l�kn��nv���F��lmm�6ٶ�m� [d  )��  z�k  m���>�
��h
�@j�U���[@��mm�-�(�@4��u@.�յM���n��������`  �l-�t��րm�Al���&� 8H�l�l   |��vݭ�6Y(  ��;i�rIl����@��ӥq��[j�4I@kՁ�����$i:��zX��ɉX�U��P9�y���3Wg$�hZ�=�U�V�(v�d��؁�����z궐' �K�͖����KUJ�V9�l� 8څ �4�x$�[m��Cj�[�*�)���vC�����*�D6�V��RZ�"A�N���l8�Ҷ�#�\�-��Ts@S�[AmqͺM"�.����6� m h�#��u�X�/U*���+@UP��k,�� ,7;i&�1�	�	8�6�nm��Ԁж��ö͉�!,� H�]�ŴH-���@�� 9����5�,�EJ�U��T%Z����ݶ�Dj-6�`   (�K%�q�-�꺕eZU�uΚ��ЖP��6�j@;]T�U�//N�ܵ[l�����.mņkn�P�ۮ�2�
6]V�^83��XwDx)�w*��Ӕv������s��eyC��K���s�]n��1��Zf��Ԙpm&�ޭ�v�@9�-�}O���l -�9���6���Һ�HWJ��vk�ًn�m��Nڶm��mXc%��8-��WZ UW �Yy��8 �e��I�T� ����������j�(t��?��w�]��`]�m���B��Ŏ� ���H�R��X%.�`��m� $i �E۱ �\k;l�F6�H�U[@SƨUۗ�j�q#�m��Ym�`8���@L�M��h�v�6�ܶ�-��H�� a���������j�`-�m���[T *�[�jK]� I: &�;`R�9�*g8���3�Nq.�uV��Ӭ78� .�R.6�3�ZG�$�^�$   �j k���I[��*�n|JC���˫�E��u�T��ܗ���#f�w6gfu��āĀ    �M��� �$   m���      ��	 p�H�f� m�� �[@M� m�q�lm��-��mfպd��;���{����ߛ{�
��[�@�������?�������Q��G��?�~B�i]
�J�rD	{Gg �ؐ���H�*m��B))�x��:P9��8΄B&��YF`Y%Y �p��h�h=���dR%4��`����+�}v�H��v���b;'�O�g��pU�T$�A$���;x�:�����h��z&��{S�Bv����WB
��!�~(��DӤ]'�Q䁀��N�G}��j	��.�\�v�> /�=��>"�%"D��b�R���(�`  &�I:g��C��*�ҡ� �"�@� ‧�קX�8
��BH>���s��6�\E{�` 1ۚI<�ïu�|�����@j
=Ҁx�mC:@����U_���k�����?�����(�ǧ�Z@ �i��P�U����R�BX�CL	JR��&8)��f��.1����1 d
DU"Ф�0�,+Jҭ!K@�4- N(�AJ
QJ�H����2@�a�����w��}��ۖ�p$m�ts�Zl"\h�����IUj5��8N�`�mA�ʐh���<�zg�9��n#g�_n]�5�C�;�374�V�Tl��#<�H\���nNl����.�&E6�ŋ�m���z�\�;lq��x8�9z����x���-����<�b�;I���-����2/<X��q�� �82�Uur�;S��$�[����!M*��МV9Vڽq��k=�eB�������#*�v6�.��
�'�d���L�.J�6�iю���{isf  �˚:�����%P��E� H ���5�R� UPUU		e^�T
�ݭX�F�HU�6)�5R�@-.���*�ʵT����յ\�9�` =�0��c�n��Q)DT�=&�t��RV��M�d�YC;	97T�d��6�oW:�J��M��Jp������T�'CD�M,�D�Y��Qm�/2�B�/�ɀl�d�q;�^�=�b�[��<.��ɜs�[s]k���W��ƺ�kl9x���Й�{�5�z��r;[�/uџ���qP'n�[�[�p���X�6��v�p#�n����Hؠ��P���q�hʙ<�#W�m��lxFvF-�냖 �	����n�@Β�M[h8+]��li�>;���vv:�c�I¸�&�Bۥ�� V�� y���{m�j^-Ҕ��p/m�W�Q�9�@��UP�<h8�L�M) �R��E[�T�Y����M�J���V����3�U�T��=��Z8�kOG;���K�7^n��Lp2�馵���F�#�\�t�j��T��	��3b���ۈM��d�6p�P�f�"	���;�F3�9Z^c+���!��Z��N:J��5R��9�;,*�L�%�(z&��ۤ��n-a��ѱ<�H)��\d@\U��u������mѝ��e��Ml��Nsrԙ���l��l [E�M�a�$�����7����.�{��� ��z����ꠞv$;�}A�H=��F{Sv�߯ў�9c�"��1�ڥ]'	XgyзS�a|a�v�t�@��;q{;&�8(�d���ZU9�kh�Q�+kն΍�q��D��۫��p�[����1ؔ�45n�`��Q���sr)+u�-��W1�[M�h�x���5�x6���z�=g���7�6i�.vy�y'cv.Ut#�MZ��Ġ�{M0�az-m�sX�[�޵`�	��h�3�ɕ�ۗc˜��9x{>��{�o�;��0vU|A�Q0���@f촁����5��g ���W�c��by�98﷙@s�tPv��wt����;L �)���w_ 7�l�����o3�n�1�r%0���| ߷��;����ަ�9��(ݞ gh�5!~nG�n����g ����5{u�:f��$֊IѲ7�2)�ql�6r�=�$��k�ˉ��*��t��4p�fcj`&FӒI�>�������:�����g >��68�G������<��s�N�$�3o��0<,���޹Q�{g �ޚp���Q�1�ɒɊ�{��3{��������-����ƢS&4�| �۳�}�M8�ۯ������o��I�)4n��wE ^�M owM ��w���������ѳ�ݓY�.`8v��mì�t[v���gs�W�f�0�i�a�sĤIHtV���vpۻ8�zi�=�3ͣd�#"X�� ;��p{�hݞ(��zL���U醈��B\DD� $���<P7�����F� �$�Q	�A1��0ճ_ �����}�'��
�Ӓp�� ջ��u}�| �ݜ ���ǒ8�mD18p[��_;��;������4l��yi�"�u��i���V6�ϖtsb�Wl�7��r�vӡ����Q������|�������>��N�w_ ����c�5c�Ɯ������~H��NU����|~��)��2Iy�98������B������PIM{��q!<	�� ջ��uo���}�|�}
"T�N��=�.U��Ͷ�i�!�c�|�}�����{�M8��| �%������c5�]���b ^e<�6�u�!��*���N��	�#cQAD/͸��ݜ��Ӏy{u�����Ord�	��F�3@nl�@s�tP����4��Z��J6��p/n����@��@^l�@f�L�2�O��dv	����y�7�P����������:�a���Lr!����zh͞(~��;���?�p5���aн9�����v]-m���4v�n��i�G�(v��<���X���$m:,�q�m�3%�  Tق睹HjL�"��v�WG/'B졦뽈��z�N�$��x��{Ob+�3A��nmU�(҆+7cTH�۳�����h���Y׳�NN�w��wFvgɗZ�'O��9��x����6n�n{O+g1��n.�W��������������ז�!^�S�ﾙt�pv�rv��f쐔�s�`�f<r0�N��l����@[�tPwt����D �R1Hp[���������8�zi�7q�<����<q��:��(��h͞(}�r;�ix�ڊ
!~nG�?~�̹�Wm���N�{��u}����=����MD���<P���wE wwM ���=��co���nJ��ᴉ(��k�b�`��Xa9�c��m�Y۴�QCГ]L(��bp�[_ ��u�wv\���?g�Π��S�{��ɒI���9���ʺ���\�;��@`>�f�iu�N��Eʯ���}�\���u��/	둬Q��n> n����@wGs��t��k;<�$���3@��7���g��	BO@������>��76�r28��w= ^wM owM��@gk����ɜt�k�9ӓ�����b����Ok��ld���رv܎�Ҙ�k�bb�/;��7���̍�5��(Ǻ(��ڊ���I�n��|���yn��~ݜ�OrLq���H����|����ʼ�}�\����)��/��| ߷g >��z���m(�"%�~��;��7���̍���6G?&H<#�_n� {wg ���\�w_ �>k���8ۃO+��66�7;'m��m��;f2���l�1U���5OAM��3�2,��ߟ���}���@k�tP��g��i�&	g�bbf�̍���Β�R� ���T�{B\@���R28��TP����4do=����xw��KH��_n� n�������� h���s��^g���޵�f�����r> n��g�?m}�j�_n��@��c�6(��`Ù^8F-&vu��n܁��l����9�wjε`J�%����rN������8Wۯ�����N }��E0R&آܽ���&w1�(���27��3�M��8��5 �qÀu}����8��k��4�^^�1��D<D� owM��@ot�@[�tP��`�l1㌉��RN��ڸ�Yj�/Z��n������lq(�Q-�g3v#�7�Rʊ��r��������'mO]h���N�� 03����Z��LU��h�Ӣ7a�TjV݀[�Lp���[���%\/i#��n�f��=��.�^��>�;[ö��j��a��&��i-&�B�u�m����"��Q�x㙺�]�]�8,�ʕ	4g7.��鍰n�9J�I5�+r&9���5��cE�����;�ww���?��Q5��[�-[R�nR����g����8��Λ5�`����ڱ��Z9�S�?n�I��h{�h��z�^}M=D"X�)�����vp�~��=�4�_nk��i�d��9 7���̍�7zx���5�_�x�K'�16�p{f�����ۻ8�nj�DLM������<P����4dw=���!�~��*����e�N�[���9��Yu��.�\���s��'�ʅ+t7+=��(|� ��2;�������9)N�գ��G1�ے> {wgD��P�BH�}[�1<��O>wE��a�zF�shF(��|�W ��Ӏ|��| �������c�E�##��{vq@c��P�t�ב�M�?�!�xx�$�v���=y������^�Sotq��x�1�?}����uFa����'2	���u��k�s�a;л�gI���Q�8���rJ}W����z�7����%���-�D���{���8��oW���7�d�2y"BX�y���"&���z�7��ߏS'kR�}�W�Mn�;��>�κ����u�M#�<�DV���E��a��mW�sxHlbz�f��&�h�!�$�iݖ����Y�د��]&��zX�u��Y#��v`�ZT4h_�`bIS@RA�cdX�WFh�4���#�bȾ�$�.��$���|<Dt�x�(o��A ǀ|�c�0�^���('�a+�߿w�)JR{�����R��<�5�o-�ֶeoV�[��)B�����)K߾�|R���~��ԥ�VW�߹�┥~��Z�k�޷�[�[��\�=JR��}���)K��{��JS߾���)=�Ϸ�=^�m�w�<������CL��:B'8�q�dU�6F�-�
��8£[������O��>ѣ�5�e�����)JO?{��R���}��)JR{ߟo�?"Gr�����]� 9�Ff	�LEJUS]�\�)��o�Ҕ������)K߾�|R���~��ԍ)����Z�3Y��v���┥'~y����JR����i;�߾��)J{���┠r�بR�QTL�(T��#�s�����┥'}����)O~�\R������b	��������)J|�-P樕K�5"J���@s��x�c�)@H~T1����Q�߾���}�j;��ɣ\�#�b4ء�is[g.C��rO��ǀ.��=a�n�5?}���Řַ�5���JR����8�)I�����R���� )JN���=JR�{ƺ�&F�"&�I�����ٶ��^�)O~��qJR�߾��R��6��#`�9�����ʝ�&����TY��z��>���8�)I��{��ZS߾���)=��~��)J}�U�V��ݽV�޷�)B�{�����R�����)JO~�߸�JR����┥'_}}���Elݢ��[�o�ԥ){��o�R�~��߿~��)J}���qJR��~��R�����N�ܫc��qV�+�gmv�����]l�m���I�Џ��ϛm�Ħ�dk��m>�v5�@l�g�H��BS�����l+��'�q��e��pn�,ɡD�V��Bz�i�h�v�����3a��q���%��˱�����V���Z4"�����:�!Ͱv���kc���5ƺܚY�(�XU�ݬX�[G��� �s���������>�,�.p�N�uk)δ�Gu���Ή�������.S9�r��\��t��Ƭs�z���)I��?~��)J^���┥'����C�JR����)<�߾�vk5���Z6a�����R�����iJO��߸=JR������)I��{��ZS��=��3f�o��f��o{┥'�����)O~�\R����=��ԥ){��o�R������o{�ff�lַ��k|�)O~�\R����=��ԥ){��o�R��w��pz��#t�ND�Lĳ��,Dĕ�0{�l��Kԥ��~��|R����߿pz��~�_}�R����=�Y��o5f��Z0ՙ�ud#�"��b�ts��2�b�����9��m���4��r"
I�ߺ~����m��);����)J}��8�\����~��)J{��fF~ts[7��f���JR�����Q�����2S\��g�)<�Ͼ��)J{�}����1JN��~���7h�{����JS����8�)I߾}��JS����)JN���=JR����u��5���{���z�qJR��|��/R�����k�R�����pz��;���qJR����S$�J����Q4���Y�@s����JRw�����R��߷��)JO}�߸�JR������f��5�VY�ݧRt9Y�vS<k]��L<Ogq0�e���wS�G���ǽ�{ݷ����~��sԥ)߿o�R��{��qz��<��=� 9�F�cݍPUTQ55"���=�R�}��)JR{�����R��=��qJR�߼��R��x}�����fo[*�[�o{8�)I�����JS��ߵ�)�p϶
�JԴL0da-L�BW1*�"�i5#� A�HID"�����w��R���T��0{���t4;$���r���ԥ)�{��┥'�y���)N���R����}��ԥ)���e���Z�Voz┥'�y���)N���R����>��ԥ)�{��┥~���B�k&8L@�m�(�A˭��c�jp��|7]y�vq�ے�H������ss���{�o�ԥ)߾�ÊR��w��qz��;�}�\R����=��ԥ)�0ɔ%*Z"�"QSQ�r���?��y�)N��~��)>��~��)Jw�p��)I�~��[�Y�ݭ�������JR�~{���)I��{��S�=���)>�Ͼ��)Jw�}�}�ov�7o[�f���{�'�y���)O<��R����>��ԥ�ʃs�?z
:y��:�|R���~>�ַkN��5�Y���=JR����8�)C�~}��JR����)>��~��)J~�=�?g�ճ[�z���n�q��3G���M��=W����.��:w��g9�޶f����޳[��)JO�{���JR����)>��~��)J{��p┥]�{�Vk�-�7��5�����R�����?d�'�����JS߿~��)JO{�︽Bҟy�ڵ��Y����e��{��)<��~��)Jy��p┍'�y��^�)K�~�|R�������+6V�j�7�z��=JR����8�)I�}��JS����(O�
Y'�����JS�u�3F�3Z���2����)JP���}��R��"!>k�ߵ�)JO}��R���}�)JRi|PBPaa }�T��$���H�i���k�b�tйq�v�n3�-W[<:����\�&8�m`��٫m�y����Z��J:Bn��ͽ������.���v6uY$r=�â������n�y�#p�S��Z�c��]�ꢌ��Gv.{:�lш\�#�{=*�3����UcFLe��qm��f�j��]X�e�����m�Ý#�m��HIye�p��V����~}���?o�?���;^��E��pv��ˮd�ڹ�J�܇[��Jy��v��t���hه����)O~׿��R��}�pz��<�߸qJR�����R��ϗ���IN<�E�߰?~�������)N���R����>��ԥ<���]� 9�F<p�4L�MH)��z��>��qJR�߼��R����ﳊR�����pz��#߬�Ϸ��Z͙[ռ����R� d�����/R�����qJR��>��R�����)JP�ߖ}k3_h�ov�l�k{��JS�u���)JO|�߸=JR�{��8�)I��}��JS�M}�����{.n�K����-�F�\����\����7��İב�zF��ȯ}VL������>��R�����)JRy��}�:��>�_}�R�����߭V�V�j�7�3{��)J}��p�'�㊎ fb�`%	ѧD�AF�D'�oI�����w��R���{�qJR��<��R�)��3M�־5oy��z��)JRw��}��R���}�qJ)=�Ͼ��)J_{��┥'�����Z���4k�oY��z��T��}�qJR��<��R����}�)H��ũW�g���1���<ļ�<L<���R����>��ԥ�}���'~���^�)O���g�)=���`���;e�#%�� �;���<v�g.�H��e;v9yD:�ՍE�o��;-��vg9���JS����);�Ͼ��)J}���8�JRw�}��R��~���|�7l�ޭ���|R����>���~	���_�g�)<��߸=JR��%5��{����w�I-1$�TMUS=JR�}���)JRw�����C Q�J pAU�l�/����JR�_��c�s��|��*fQ1ڪ�D���┥'~����)O�׿g�(|�Ͼ��)J}�{���)I׵�V�c[4Yoy���=JR��{���)C�}��JS��ߵ�)JN��߸=J[�����#��/�%�N-��6sȝ�Ϛ�]=��݂���-[m�L�9m��<��7��Z�k{┥�����)O��~��);��~��)J_y��┥'}��3�k�4k��[��JS��ߵ�)JN��߸=JR�y���)JW"�������� �d%:%L�MJ�����);��~��)J}�������;��߸�JR���k�R��{���[��c��kyk5��z��>���qJR��=��R����k�P��H���"+��&��߸=JR���3�f~7Y��[ռ�og�(z�߾��)@~P'������)I�}��ԥ)�����������������^y��ʃƹ���ە{
\a�{!a�fZ��C�������3\0��6kv��\�9��R��<��qJR�����R�����JP�ߍ�9g9�G�rJ�J��U�$SS�r)JN��߸=H�J}�p┥�����)O�Ͼ�������-g�͕����o�ԥ)����R�>���pz�JS����)JN���=JR�y��+N�־���-e��┿�2����R���u��┥'y���(_��\R���5_f���֬6h�7�s�ԥ)�{��┥�$|�����)O�}���(|�Ͼ��)J��q8�9Mg�j5� ��&9冡C�R;�K0
m�(%
��i���k֔r�����.-$�E)��,�L,@A$$,��$e6e1TA��e�d�v�T���$d���C("�(�1'�4u�h#{	އ�B�8��Ra9ALHV�dDVe.TA���F��3���2��?"k��%i�S�J��`�P�!�E4$�fi&t�i�(`�E�!�VUAQbab�P�aD��2��v:�e)�AX�8G���WXAP1��f�KIH��n��GNYY�e7
g6�����u�}�}���^�n�r�< -s��M/,X��
���e	Uj1�����)]��̅�1�5fs�r�n|�\���91�>-����v�^�{*f����m;]�0��*��W�n��/�v�Vv,��� n���c����n���]l�6�)�{kg��ӛ�O+�;�osm؝E��uuX�LU!���n���\!�"B�m]f��a��lж�i��ɦfdn���X��M�[N�ә�6f #bg[\h�nv��g�}�Ǟq T�	�'T�n՛c���lfK��Jf�V���%f�����#jY"T��ejv����z�� ګX%Z�^mT��PN�����(�[R���O���T��)�XԴi6��U�SV�JPU� �:p�6�و�q��r�:�r��T�G[���r��s�Ui]�꧞]�
gq�]��rL�\Yku�'��c[m�id�(iX%�N�sl��=^����l��.8�ф��&�w3��:&
r[��D�UϬ���I��ny�^��lm�n:����7�_8�;&8���a����\��x���s��p�:z��v�u�i�&{v�p�=�!��Rn3֔��oI� q�:�r��Wl����s��xMۮ9t�bxts۵���s��[d�-vGP�����G%��1�a�����-E睫��;h3&���]��=��������W��Q�ˤ�]A4蓲���TФ���i{-]E�uSh*
X *9�;+�O*�d�*��m�!�UΉ����m���V���v�\n9N��N��JEۭ98+dFk3:u�v��َ���*�m2I�����x��s�Oi�T,i�mG@q�ت���kM�A�-k�� �%�l�����:�ew�SXx�dvp��R��+�����Y���q�v.�gl�8�X����]����m ����I�qUI�w-<�V̑`ՠ��E:�n����| ����&cF�kZѳZ͖f��������z����OE](L��'�  �?؈����A��6߃�~^IMZ��܅9ۖMx���͋���޻���'/�h��Zj��ӥ��ݪ�nxX-�Q����	��'�i�(p<9ԷoT�fز���u��`'��:4�;�zֺ���c�9�� �&&N6�zqȸ�G�5���+gIQڋ/6yZ(
��^��Y�;4�t$S����1� )���K׫i&Ų��R癦�5=�X'B(?�u��Y�ֺݣj���6T���4Pd���3�(L��q�7��;v'u�����1��C����m�v����?��ԥ)���┥�y���@�#����9�ǎ*��Q��5k[��)Jy���-)C�}��JS����)JN���=B�)�$�'��%J����9���c�)Jw�}���'}����)O}�\?��Hd�'w�hό��FoY�[�o��9�R� ����qJR�����R������)H�P��}��So{�_���G�3]�i�������}��JE��w��)J<��=JR���}�)JRuߙ{�Ϸ����kyi;J͐ܦA	ԛ.�&z�ݖvN2��*u��`�ݟ���4��]��a��~2������)JP��}��R��>��p? B#���~���RW���bǉ��c�� 7޷��~����FV$�RZ@�B�2�>��r�;���|�\�����!��T��T
�UŁ�g�gjWg��x;zQ@ڕX����CQ<M�������}oz��\ �y��os��zu���J�)I�ˏ�݁�Ҋ �{���J�u�(����{=��U�piH�"NC�ځ��.g�l�i�փ%�܊���].3��{_ww������9�%!n ߽o:�������o3`��P�C8��y���%�����u�+�f��� �y]����jUg����y�7R��>d���9 �����ڸ\;�8"�D,�Ͼ�Uy�{��W^E��e���������"�b�?{��t�ݸ�>O���D/{zd8�bx��c�ԏ�w}�������odl�P�������@7&w��q�-v���R�L�Nکo$�.��]v�����k=�6��7㻻�+��U�t��j����Q@f.W`f�'�3y�������M`��d�����|�]���3������\��}��oy���ݺ���'�Nw�|���}v�:~���/m|�]���V�9��1HM
�z9�,�{q`yc����wX~�����-�A�@��~� ���Eg�H��r"
I��/Z��f�yb�V��hv����{~�J��q���:��hCg�]��8���ll\n�1����wwwr}������b"f(����)�[ʽ����`|�k���=���0�F)�@7q�t�G9Ȅ{^������~�vr#���n�Y����q98��y�1�QA�f��[������P�'wggy&ᮞ����7���(�5o+�>[��3��߃o��U��XӬ�A�$����~�v�8Ds��{= {�{`|���	�[ ��'0���VM�@csvn^קBdh�-Ʒb�w������)��i���:�Վv�)6�iYmc��H�F��zN��9U@l[r 휫�,y��M�5��*���FN\�=[m�Ƶ�l�;l�:�n'qՌ�w#Y���%�������\FN�Gj�q-ں�r�N
L��Kj�q۝�i�UVۢ��t�&H�r�K� �j������};r}�q;<����l���Kxò���ǰGkv�R�	L��ϳ?N<�$��F������> r�U`c�(��0�+�C�Dı1�����n��@�{k�}oz��_33 7}��Pj~r"q��s�c�(�9jWc{�����R�m(�$��L�!r>��>���ގO@v�V����(�/���KBT�M]�����\�<����ye�|��{�<�yjWmA�?4ƃ#;mm�#��tq�q�#C�$����q�z9��֯��Y�bbM��C"��[��/m|��{�:��N�ׂ�,X�#I�J���>^�=�9����G"*":9�vͭ:{��_�#��Ȅj�(�L�"J%T�3S�=��vٔ΄D����>[����*�%1dM'���C�~�����v���{� ~�;����ss&")�p�[��/m|��{�>׵p����`�j(�cNa�+����0��q��vm�Ϋm�c��w#���n���x��$����2'$�t��|��{�>׵s0�m�tz�Ƥ�I.9L� �R�<����-�m`b�s��@��8�SP�UB���+ϵ���]������2z@!���ok�{���{B�ͦ��!ć���7�ݍ�>��J���J(�kʚ1(F��:���>^������o��8�@�}������`S��&��ݗfӫs�V�}<Iv���M8�<.�v�J�AbǎF��5�@��������>jS�z�3R��$�lNw�{�j�~� ��o:���������qDD ���f���%�a�&$����`�M3y��J���\ ��I�Hb���8�7��~J(��v�rz������3���1�vr��v����,�!rE�����Ԣ���I�u�(�����?�Y�g��ps�d\�s�-��fȁvgVeK���; ��ٮ���n�������u���BUR���f���Sj��x��ٙ��n��kJ�ͳ���H�3#R������P�����wxG"9��ob��TĪ�"�V������P��������Ԣ��>jS`n�Lv(6b��m<m�������z��}J(͔���\����" ��p�&b"n�ގO@�3fl$�?}��W}���uV��J�@��̣��$��4�X�rXѝۍ�B��PwQ��kf�^Zct�ɍ]�2s0uu��`�Vŉ�c�m%�b.���ݔ[��J�y�L��g�W��ɳֱ;�쵬H��5��[����|���X6wE��ⶁ�A���^�v.����4Zˇ*����w:����ss��GZ��.�f*�8é���`6�]v�,�UnN�E��79c`�����.��wȮ��4�׬
\��g���d�'J�W��Ǯ)N{N�+~����c����)9(���U����}���DE��k��F� ��28��.���_?g�>����|�{=���V�7�j�fhv���&b��Ԯ���Q@�񙲓�/Z�h��� pB$�s���m}�n�E���E�o7�33>���1�[0�J�$LJ������������P�����(Z��4uŔ���,�{�v:����Xⴚv��2�@c�7����N�3~>߀1�(�35+�5��W�����z�yc�d��i�n>�oz��g���zȘ����H!d���G�7u�s�r����}uWy察�f~���[�$��bq�s����}�}e�ȎDA�DG9������v�1�Uʅ4
�����@���� �Jh�J�{��ͻ��k�s���dg�Zbfj� �Jh�f��u*�7zQ@f%H�;�9ԃ���H�m�R��Zնź�{����h�&n��ܝ/Y�#��������u�c�1�j�m����7zQ@f%Ho5�f�4�9y�r�B2�U�̦w�q#����]��w���F95L���l!R�1STt{w�X��t|�\]�$AI��:D�F���Q���o�Y�ԛތ��WWvj�r0�,C`�5�c�n�Q�A�������3K���jpg8o�n�a�7��mwλ70�≜#{�f&��T���F�E� �o�Ѕ!�f,�*���C�!�l]ho��8��MP^T0BT�i�:�#C�r58�P�7��ه�I�*���"}ء���v��TzD��C�AΔ�zb ~�{�]U�o�yߞ�M�m!�������>����{vS�w�^S�{�#�sLMC�4f�{�f�E�g%4�}XēH���2H���gG)v8����\³�;��r��9۳s��=v��x!�`�"&��P������փ��۰h��PT�B���D���3R,9)�75+�7�Q@	k��� ���Ii���,9)�35+���@�n�����`4Ḓ���B���"fh�J��P����f�~K�p�z��Cb���Ҋ l�R� �Jh�J���W���~;N�v��fl[;�;s��/>]6'�v�`r��Χm��.ہ��c.qq��i��������䢀�ԭ��P��X8�o�b��}����W`ot����H��u4�)����w^���7u+�7zQA�1*E�}�g ���H,q��q��;�3=�P�R,}J(�J����$E#Y��}���@��>���{�n�zq����&8�h��	�SS5ԶJ4kC����<�U���T�΋n�4p��D�V�ڳ�vݩ����lq��ݣ�h��
��AƀwE& M�ɯ<=t��hy1����p`�<�ӭ�009���N��!�ݷn�Z8c9��yG�ț��+U�{E��a�'ίd��z��(Պ�L\ols�]�z�.�ܳɗ=�M�u����:ۃE�]�S�J�f���36o>TF  �Y��9�.���Z���mcjWJ��.g���Vy�[�A��TA�J������3��:Ů������M������Q@f.�X�K"DǎdC��{�[ޟ�`yo(�1oR,~J)��X��"$bX"�����<���gYg��G�ݞ���n��I�$M�B�������X��Pڕ�f��Q@f�t,��nF�N>��/Z����}o:������:��r<L2G	\F��v2d����p\q�qm8x/<���87��X�H�Ɏ$(�x���o�oz�r�1*G��f�䦀��D��KDn���oVZ���3�~�4i���-"'�(������몽�=��Q�z���m��B)����n�,~J(��o������V��ʒdY	��9á������v�}�����*DAw�w���*B�d� ���/u+�7����ԋ嶾���4��N4�mC䐓lP�Q�^ӍGj��Iڇ��c�-V{=-���^�.�^���q����/���]H�>[k�g�=���@����<B��'�L����`�M��]������[�D(&��Iw�@>�g ��}�]Y���1m �z�z�ֽ�9W���t/\Ova��(�������z9=��"��x�Jh��D�D�l��M9ށ��N f~����t9)�7u+�#���NC:g&Fba�n�lp�:9���[]�I�Ƹ�l�ۧe��&-��SLN~��R5�8t�[y�1�(�75+������ ��� d�K�,�SSUV>��f���Ԯ�����|����[�U��x�y$Ic���35+�7�Q@��7�3R� �J��3*�"�5D��]��"=�L��J�9)��f��ϻ	]��	��xhwe�bbd��J����rS@fjW`k�(�/ ܁ᥡ�y������H����z�R�@/]=�ǐ�v ɻVu��fg�rs8��n5�Iq�s��޶h�J�}���U�˦!���9JJ���������s�"!��������n���s�s����T�J�L�<Lv?/��3U`�M�����ۉ��Y&R5���?~�Z�XjS@v�Wa����{��W�@|�u�����Lr"r>s���l�܈y��|9z���}�=ȅ�e._''���%ΰ�զL��P��I;��'��6뇶�=��lr�c��O�lۤ��(ݜ9�9�e�����+<CW*�tk��J�ż�շe$�ڴ&<��{cR�?�������c�n�=�N�۔yƕ4m�!K����4�X�^:����ν]�KԹ:
`)����.��Q�m�̎��x��[gnUNM��(� �m�Jhȍ�Ӌ���n����}����������Z��:��m! :Wt��K����HlSۃJ;�4Oq�u����g_.�y�1UI(�����{�`{'�����>�g �<���ɀ��'z��ox3R� �Jh�J�f��y��c��5��$| ��[΀}���޷��־߳n	P�#��	u�UV���Jh�J�}J(?�7�y���f�Xv�jBb���B����������P��M�n�4�:a�ص"�p�����q�dm=��qњ��Gn��0�`h������]���t���5`k�Q@'�Jlu)��f�o2�{v�kb�T���E*�QJit󒫆��מ�[3{�T)M��]��־~�>[�ZLE�c����9�y��{��͎%�;��y���~ȥW&T�IP�f��Ëُn�̝�����/7=�b�p	���
�������6�{��Y�=�{��w~w�&���z�9]�.3�f��;��^���`ӱm�9zwc��Hs����"�L;�/@��X��P����������4�/$�,�p�UV���7R�vz ���`�XT��XD,m��>���@������G���d�)�Q d�P�DB�|���o��꫽����ܪ�,o���Nw�~���@��X�S@f�W`�Լ�4�d��,#��}��a�[8�v��yz��=Y���f5�E0���mz -�c���9X�FSO[�S&���i�O�p��9PI0D��UUUV��wr��־ wv�t��T�S�o$jb��O@�َ�aq�vz�=��^n{�	1���%I
J�D*��=��_��l�"{7k�{1���Y<J	h�]�b"^��y�U�v�4or���:eBBZP?~C@���_�� �˿�i�1�8ƺ>s���k��\�c��,ݞ�_��l#�$�';�\�,�;�mX��씶}�����:�ۥ��Y��k�v�9j���W`k�Q@��y�u)�7VU\7����Nw�yz�������y�3v����G#���H=�m*���ȢRE�q��_��t޶p33��{�<�k�[�bfTB1�d�9�UX�S@f�+�5�(���%V��V(�c�ɋ�p��{�<�lP�%V�������������9"�C��`lҹ0D�hJ �p��q' ��8n]�4y���-�7�ɤ֬-Qc���D�I��eq��e�a��2��"b

F*�y���$*����jӴ�DĄ�D�����On�~+u�Z)A�r%�ơ�t��S�kY�r�j����q�4U;�+rҭ�]�1K��Xz]�ێq,��`� �q��Wm��u�츱QA�襋�W���.Ļ�v��d�nz�<��3����_4�+�u�l��'nuW巳���{l���#�ԗ-��h6�q��x�a :��X�oyy1Zλq���c��*�r�7flĻs!<�ô�,�eډ�o'O��Sm<���Z*,�T���%�4�TՍe�]뮭n�X
@I�v��6�%���k iz�kSj���V��8�WU�\��f�6�հ8��t+km;E�2l$-�\l��X-�mW�j%%�@T�ʙ�j�� �+��&A��V��55 v��5mT�J�+{l4Va���ٻ	L�R�Î�9\ԊnH��C\��hnT㝨ۗ��V8�vG�f�B6v��v�F6�N1��n��$�oP� ��J������<��஛�)�^!�ۤ��bt�^C����)��W�밺!�]��s��VX� ����[��Pꇳ�Χ�#X�ŢRr+%��n]�7��nl��m�����.�6���2'�]��1mɵu��]����c���v*�g���{*N2酙�{c�N-9,��<,sV�gɧtG���WP�\��ݞ������`��j����JZ�L�Fh�[l܎i�X!��m�a��]���ٲ  �U�dV����6uvu�2:m��B��7"u.IUꥀ+�MN����9�+����������Ʃ�u@J#���� 3gk�6�9l��ܼTy;q���p��:17US�4s� 8p��u���<ӝ'�Ԫ�(�ʲ	�oe[k������8"�8K��b�w6SWi�J
�p�Ӥ�;^����u6.�(Ñ؜"��T\��J;�)7�J1���4��i�T���P�]K���9q7�
c9���ҥd�3.���Ω��+@Wm�]U!0,@��K��9�>�>�n�����{�T<W�T�҈��PT= �edP�fӀ֯=�+�4f��v�T�J�ڻ#Dt;i�l���pºv�d�����t�3��c�ӓd���	Vt�Ts9P�ɳs��(�Ʒi��!���*r9G j��k)=bOfKs�0��3�����z�S�9Z�J:�v����r�!�M�uօ�GL��ʥ��5�e���>��);��<��6�!v�r O%��cf� ��h�Ηo�w��w��_�`��v݃&�9@�sŷ�dl֔���:㗶N�U%Ʈt �˙�\��~�d�F''([lP�%V��׼wr�x!;;�C@�2�}�U�n�4wr����v"" �歀D�TUQ5$�"���;��h��v��}�U���¼y��	�����ݽ�^J(�����S@n�N�Gh�#DԉL��^nz�������]�ͽ���b�	ԐLn%F��6�nح��N{d<��Wӗm��k����t�}��}�ˉF����wm�@����}�����,ݞ���u)JF�R**+��{����U36����N��v?r� ��y�/�&Y"&FLLr>����}J(���_R��7����@��8�7`k�Q@ܕX��P۷���H��/�1c��| ��-�tjQ@jI]���E{���/;h��q]�H�v��u��ɜ��Wl��'����s-Iv���svK�fr~3��}��R�;�]���E _rU`jO0b�!D����1��BF-{= �������y�NhS<J����<D݁��E��Y��{���oU'���_[{�>��o&9�����,�J,}J(���u�(}�0�Y[Y��s����k��m�@����v�m}}�U�J9���4��k���v�}���a-y�ӫ�n��������d<s$��p�11������yڸk���<�k�Ͻ�a��!c��"^f�u�(���R�sy_@���$�<u&,xӏ����@�Ԣ���W`k�Q@vo
A�	�h�U"VO{��~DDrNn�@o݁���������3�k���}�#��gw;`|��$�D�!R��T�O@��W`k�Q@��X��Pڠ3��� 5nK�Ѫ�A�^ld8���g�G��.�Gj��ٹ�P�U��Z�����(���R��y]����)?DF��	#�m���fbG���K�^m�����^�T�$jTR�y�&����}J(��v�� ��y�.�^L��d��ɉ�G��^��e���}}ܪ��Ԣ����,8<$��!ܝ�^����y�<�k���ށ�߷����N5�B(���W�un�nn�ї��tG6�d�'v��-�sh �Tr��6��6몕����U���+��Z��3�g��mp"��89�0�Q��{�Ny&�)�k�3�8�vN�s2�r\Vۺ&�qD+���=�ҫ���Ƕ���ۮq���f�v��W�um`1G3�v`���y�V�0D����[=s�d+[���?@o��Z�Ixnű�ڝۑg�x 9{Q2]Z���ںml�;rh�'/<�rx�1�ci9> ������_ �����޶p��\�ȡ��t|��@��Q@_w+�Ԧ�/��_�����HX��!�ő������޶p�ߒ>ݳ�yz��=��KA���I���@��X��P���\仸�RD
I����@��_ �����l��mm,P�♃fҜ��p� ���L��v��q�)ʛ��u?���ch�2)�DNs���@��_ ����޶p��y�/�>#FLL���/�����������o4�wJ� ���`|���b=�hI%HJf�K�57`����V>��r�������c�����wm�@�m��}��� ��~����Ȧ%�*��~J(��v����V���6������=S��-2�"d����ta݅[�^U����4��ݒ���� ��0;LD���]�o%4��U���>�2����i����l����r�n����g�}��w���j��&!�bjF��8���΁嶾�̂Ha	��!���(�( �%	�B%��f"_@�=�/����g >��I���'�(��UMU���Eky]�jJh>�;���X�#f;ILR&*J�$�O@��w`A�l�������>�QZJ��rzgH�ƫ���6]�"�&#j;9㊊ ɢA7�����M�d�w��� ��U`s�Q^�ky]���B��c���$�������;}�� ��s3��]�dd�&E1.��ʰ9�(�-o+�IM vo*�9t�"�!�ő��˷�{�[��U�~{�:�N2�0� �8�6���7�Spw��$�M�;�6�l.C�=��4�g�[�;�=��۷k���r�m�\[iw(��Y�Ga7[�x2�N���^f�b1"dnmͮ�&h�yU���Eky_�`�M }�kI�[Y��D�9��t-�����{�������S#&&9 �����l���y�<���;�v����N�?�r=�������@�����$���&�$�W@3�7�N9{�ڿ{�ߺ�Ͼ�|���BH������^����[V���nWu���]m{v���x<�WR��z!�/O'����\ml�6zsֈL �� j�%�-�������W����lT����ɝqK��oAt�cr��I��CBM���c����'q�=9�����3%�3f��i%z��L�p&��tʶ�r��"����6ٝ86�'r�ŉ3�����3<����w����w�k�M8�mq�*�i]��Nٷ/��p�U�td��c�cjwbγP�;�U�����UU���E ��]�jJk� ���n�1\��idn>}�{���n�t|�{`b��x�2\�J����iIހ]�8߶�t
�k�{���}M���"�������}�Հ�R�7R�?%����2�v���yrj����O�E��]���� ����T�$�� �	��<�H@�:"r�����K�'�ci����Z��~�r|,c�Ǒ���}�[ށV����o:[k����)�BC��b{�]U�{���¨D��R�p��o7�5g��f�*��_R�7[���$7Д�#y4�*UT��}V~J(<f�W`'䢀�]	��"Dx.��s������{�*�_�}��΁n�BM\�1�F�F��{�݁�͗�6�=��cs�7��������?�M�:�s4�F�Tu���@�v�6�ƞ�4�'7�XnӓE�.�$��R������@>����nw����v�q�����U��I)��bJ���P���	�(����Q���/0MUUUX	�(�3u+����}�n=�4}H[��?F��Ў�m��
�ג��A���@�.�`ш�����x┑ @~D���lv�I ���0e�ih���*�3]���m���� �ډ�6�v�i5���2�4��o6!�M�g%��0C�a�&�`]�2���i���Jc޵�o@�tu��8��v���/`Ƀ 4�4= ��G��x��6'o���K�A� Q�8�g-Ƴ|�\������Y[��#&&9��܁{ٻv��= �珶X���<�X�`�1���@�m| �뷝���}�{�<�yq���6�Ę���V�:��&���*k��[���Nrty fSi �ٓ�5#��]��]��w޷�������14H��
�W{��n{��s�fn݁���@>�v�[� L�"�7$K#q���]���E fw*��Q@w�'� �1��Ɯ�@�v� }���@�־Wi�$H���uϻ�>�>��$Ȉ��6�"��n�t
�k������]y��F�Q�PIQD��Sp�:`�p:�&�m�c�-�:z0`8Jd����n���$���d�99�|�����;�[ށu�\ ���΁���q
!�Y�e��J����3�U��]�s�	Dn��(��"I��\���3;�X	�(�/5+�;�<��3�	�%��"e�3yU����3R�@��\�x."�I�6G���9΀���wy]��z �IU����%�OCh���`(d�� ��҉�c� �Ȩ������������Φ��m�2��,q��g۷.W��x��8�� �]����n��m+q�[A�xu/0Gh� �Hp�J4�*e�#���uq�fg�����P*I��cl�%����vƛ�8.lz�cl�z�l������a�FI�aۑz��W�,��s����S�.�0bn3�-U'O9�ll��z�c���`�θ#�Mti|�&�g���wwy�`>�3�n��*�ۘ�m�0��g��m�ug��ڕK����m͝��;DDƀ�|��]	= ^$��O�G �e2�Om����]���o���|�Sݞ���n�~�٪�����D����΁V�����]���t���LD���'9Ά���=3݀�7= ��}�3��\x(�#&&9 ��������[y�*�_ ��JՉBI�%���͖.����le�B\��g��b��֌�Y��?�8�1)1���@�m| ���t���Z�{vq1�!B�lR�6�{�*����[D;J`�$I�o3x=��~Yf�?r�>�lt�"����:^��}��^���v�[eo��6�
*f�����{���^��}�c�׭|t�WSq��ƛks��ڨ3�U��R��R� ��8��3�uixs<���aLw<:�l�p�aM�c�9�s�`ݞf�\N�F�G�c3�U��R��R�?r� Y�(�!���I�rs��:^������U�_ �}�g@�U�5ǃq�FLLrb��Ԯ�Oܢ�o0�7�m��ޥ6^�����Z��JLm1�N�
�k�/�Xy��oٛ�XĢ6)D��J����|��u`lDF�n���۰N5�/�I,U2A�
����@�v�D1v97\�+��N��P�b�۷(&,������|�����;����ڸ��o:���6O�M�&y�z�R�trz ��U`-�����J��㘘�mcNw�]{W �o�΁|�\��{�>��y$y2A�irG�z���	�(�/�+��f��i౟��i�֓�t:��� �.P�QJ�`E�1���"( %�$b�q�q"���*i����p�33�Q�{��ޅrhXu8N�1��r-8�9hu��s�{�w����RR�53\��U=���`-����Ԯ�]�����6��o{�������ڝ��v����g�sm��3��:��:�����J{���v<LƝqL��/������~�S`'Ԣ���CW�9���rw�]{W �o�Հכ��y����#��[$(JU���X����̻6q��ߵ,�usx5����*���w}oz׵p���tl�xD�~bm˴�LPڕ����v�>�W 4B����U�����yo[�nĽ���9���n��ط�z��9��%��n0�LN�]8:ׅ��6B̻;2�ٜ��\gD���O/^y�m���/;g�7=k.��e��nP���J��m�c�T��iŝ���K>�]y|X�]O#�̎�؇���&�[�dqn��k�7mm��8r
B�*��G8�ŋ���h]\�0�Bm��h�q�uW��벟l#񛳉՝��(6�l�/]��g/��۞��'�hf�Qcb�X�dx�mcN{�}�j��n�t
�k����@��\�A��# �/@�ʬ��P�������w�f�(�53<��Wk����՛��/޷��ڸ�۷�}V(����b�T*&�zȅ�f���z��ُ�^����q\'1��N����f>�y���7v�1�H'���=�nJ�@�����-�ى�ftl��DЬp��,�ps�]�dθ���g�5�/��O�E{�]��9=yγq�I�M��T�'@�־}���1�6��(I�|�S`.R�&}>q�j�3S�/�n���Լ��Ձ�7g�f��K�*bT̨�5w��DBF�z���ڰ�s���c��8�s=�J��`�%P��@�g�Ձ�F�n�@����'�|y,h&bD�b��V<IF�v8¶�={F�NI�]���f���@������p�dq��Ȉ���N�W�|��{�.���|��g@7�bo.	��#%�"f(�J��.�O@c��>��m��\'1��9;�.���w�����>�B�x�à�\�P&�}j��hJB�(JS1���X&�X ����G&9ȹ)N���=�2%	
S�
ISS���9��x��Y�=����U�_ �ږ�U����|�Xy���盽�M���{Y��߿Ѷ�wUqb���Mej��Ԓb#Z�s�F#=�����i�1�f�Y�-@v��ɹ�8�w���U�_ �o������=�1\+��x6�Ɯ�@�v�w���<�=�rwW@��w{��$���$!1ǃ�"��+��t�j�~;������wڊ�brG�&\������O@^�W`'�Q@{��#�P��0�PL%�g���� �ՃyRL�b���p�J����|�S`-����l�s��Y)��v���B!s��0ÔR"�3&��<TQ7��5��-�s���G'�1�M��R��R�xhʁ<M_�,L��|�ݳ�U�_ �oz׵p��r�'�����l��P�������ܦ��l�� *f�Q35=��f���z����V^nz`�N%WN�s��ڸ�}�t
�k��}�]UѠ蓉�N���'_C�m��Jk��a�r0 �	�Xr3�Q��JLh�e*'0�"��E<��EYE֙L�� �DЫ�莶"kJR��]���B�E��s�6u�Z�]�u�@�;�� ��R�C�v�ѭh�5�d���C�EUJD�eIkD$���*fEwk���l�X�4,!%EBAA3IDN	��fyh�a+[��=����a�O=jMj9��0��%������L����&��4�] �7�^a����p�tg�:;��`F��݀T��I`��,B{�CZ"f�� �$�l۪�7cNy�k]fk-����q�d�+n��%�]t�k8x���
�h)x*`۶�CL6j�;Y�*3p�xGv{;�����������u��v�9�Ζڮ��.���xOY$�j�� ����u��K�k���x7I��gn��np�֊����v�׋� ��]rh��hwm�n��4�l�M����F��/�Ӵ�쁺守�5K�� �u�7Bj��[u��6�J��q<��� �]<����e��j�G���04��͐*����`U�U�U\�8�X� ��RZrβ�!��&�V����/Zi�V�<F�h�Y- �+zV�(.���G*���Z� b�SPm�%�dx
��+!5l� :kSX6�-�M%�ԫ���M(ԯZ��t����XZܔ��Y˺��GM$��i��YFX��Tj�"I��[zm����q�rm4-�m$�k������t�K5�gJj��cB����v�"8���X�YL���-:�I����u�;�V��S�Sxq��GJ\g�t��3�B�9��e�^�W�qn1�Y�Kh��Hrc�8��k�=�����ِ� ���4@e����b�u#vf�t�k{6��ܙ.7�e�1m�\q\Q+��Gm�[�]�j�pg�tn"]�b�������Eقk��4��#U�6X9���d�N���[o]������BPn�:��)�-���y,=���*� ԕE,��iJ�ue*��Ү�+j�VM�H�7f�`�jk�S��li��Q��Y���,;uǁ��ޭ*�^�` tC��r��9y9�;!S��$Hk��V��r>v�F�[��^U��ٞ0��ڃ�T� ��2�+r��eZI��<��%�9����l�9��z6��kM��ʁF�IWO0��f������v�ӎ�5�[y������}k=�7I¼$.�R�;E\l�I��կ]��]��p���fn�u�K�ŷ$�H i6\�JA��t��I�=@�
���Hq���0�d��8�����w{߯�~y��5�ǲ�r�]K�\ԙۮ9�7QU�1ٝI����筞k�����C�*�;m�rn����6�n�D�Ea�\m�����n�9�D1qX�r����/U�_n�m����JA&sKY��l���l����ݶ��]d��]�P��r��!���8���9�p=`5�;���Q�43�H@�u�o�ƶ�W��|u�3�m�;n���������<�YveiŶ`��\c�Nu�;<�Ɋ�2��ݭ!99أQLq�Q�*�]��U�_ ����G�5���x�Rj��ĕRT�{�̀�R��R�trz���.Hlyq�D)�r>����^��>[�U�_ ���,nc�3v���?o)��Q@_jW`oa�x���b`�\��:^����@�����ǉ�bR.��d��B�/h��Y�L�>_Jn�gg����A�;�gA��A�q�Ļ9:^���7v^nw��Z'�j�z��P!O�nAcn>���������׭|�wl�n��=�1\+$����cnv�O�E���l��(�J�p���Lq���p��l��k��[ށ�v� ]���RN%H��=�j�Ř�o�7~�l��c�6�q�����y�2�-�5�'q�`, �v��m���O�������l�-1@_jW`b������?y�����z���BД�f�I$���>r��������Q@_jW`o�2gx���C����l�n�Ù�2�H���	�>�]{����=��r���AT%ԕɄ������-��z�7n�k��@�g�Ձ�aSʂ[�X���w}oz^����l�n��7���F�Xf0Bm����&��\�qK�,��,�;h��^�u�O:�>*,��cnw�U�_ �o�΁V�|��{��h��o$����H����oc��������۰����`�Y�8�Q�.s�}�ڸw����q-��]�q����	��UATTC���ڕ�a'�3�yE�{7�o_�g+�j��J�,�!cs�9;�.�O@gF�trz�_��=̤��'�M��Ȭ�F95���kM{Ob�U��� �4�����\kp��3cyE���E}�]��R��y@UQ*
��$%M�{6Y�{�H��v�Y�=�Nc�>��
xR&UP�T�tg��������ٰ׵�7�LWb�`�17;�5z��>�M� ��]�#�����<ᤶ�QUQ��29#�+�΀z�}���j���o��Ɠl�T�&H�D��"�8Ř�Kgv�r:Hɲ��簯[�}���/B��ntl�f%i�j�-��*�"Xȴv�%�m���OT��Y�'v�Xʖ�jmm����qw�5��]����8mi�`�%�ͷ+�B���k���t����z[,�	�0ǁuv����Y0Wb���D�ʛs�EYL[y�k��w]S��%��7m=���|\[Qۥ��HV�g\Hb]=����N{i��qۄ�L�U�M�w�l��8�Q�q����_��=�W�|����^+��$&<mI4�%v>�?$��Oܢ��s`�J4B��D�L���5f���6�������{�=�E�&���Rfb�������ܕ�	�(�/}��6�����N�u�\wk��7=卺�6#�\�I΢f�e��)�'b��Y��p7\c��ϡ�&�nV{[æ^�.���LBa�Rqt��n�k��@�cn������iD�V�5��e���������0��]�ͭ��%6}��%v&�wU��D�1BH�����]��{�oz�Z��Wa�N
(�8ܩ�\������Ԣ����l�f��Ĥ2bNI�=���W�|�l����=��LJțA�0�����8;<��
h��H��b:���vۋtpU�.΁�B<K"X�7?6���@��_ �Z����ڕ��0�3Ë�2�I#�k�_@=v������k����6(���y8��������ul� �A �`�8�i<�r�=�{X�稨B����i��=���W�|�l�Wk��\+��hm9ށ�v���)�5�(�;�+�y:ND��s�R"j��D.���1�&e��s�#�[pC�\�7 7m4���>�o�.U`k�Q@_rW`v�O@,�P�g���2w8�9΁�v�w7m� �;W >����g�n%C�27#�rW`n�'���V>�g^�!c��Q�;�=�p�n�t}J(7�oq�7���i�W`-K&�m)�
D䋀{v�|�k���ށ�=��wjH*k
��p�5?4�L ��,X�Î}q���Б���$���]'M˛IɄ�85���Ns�|�k���ށ�<kyȎE�=��l�7��B�R�T91�%v�rz{����P�h�iȒM����ڸ���l}J(�J��N:�LĐ����"�p�ݳ�|�k�����{W �޹d���⌝�'9:�p�J��I��V{���@@��VZ���d����l�����j�y��0����nz��N"�)u�0j�@��Rd�	�jQ�1wT`#e�mI��!�¡��v�]���0UÓ�Ͼ������l�ݮ��y���R�.{��b�
!�6N�=Ht���X7;�ӳ����N�J=C��s��5
<[F.��BLti����읹2k� ��:^ƃ/\3���Y�������{��!����1�j�<1GG��}�q�/;��..���/;r��2O@�a5d���W��_����mt�x��s��|��{]39�lQ3\�H���1y�����y㮁����##]#a(��J�B�UUS�<�^Հy㮛�$�n݀�o����<�7�5�rrt�l����W�|�n��=iy����21(�|w���j���|��:����x[�#�x�15	yc�L���6�6�U�Er��v�i���:�1��	?I0M9ށ�־�l�Wk���ށ��^14�h��$|
��}��xg H��]��P愮��;�oz�Z��V�1<�/0M�L�U�j�4�%v>����t��a`Ҍɂr>���߬�vz��l�t��0M9m1�ށ�v� }��� ��:�7v�fn��蚚���)B��fT�J���pG2&��6��.Y��7��)�À�d�ҟ��NH��o�:�p��ށ�v�۶��6)#y���MU�j�4�%vl$���U�nʛlXF�B�ӓ�{�W���ã�L!������&���f���L�PDG[�f5kYYF�6��
9�S�1'��ˆ9#R{qp�5�.��wf��:�R��PԵ!�9h�0&���#���c���ep�;��.��1��9���fFPekDd��f8�cfi#����D4mN���k�qߠ=���*�}<CPҀa�	����j���o���<�4�"&��I�5r�]r�s����E� �i�b�H����t+��}���o���}�Rܨmcĸg��ȉ���z�9��]��m�U���g�DxD�GO"�j"w8�9΁�v�ﱻ�1y��Z����=�f&$6������MT�����$<���f��t�l��`Z��!d�ciN�����wW@<��l�tg����L(��U$P���R�~r!/={���\��|�@�PIa�"�S�*:��1x�=���^{�f�4F��G;'9�<���=���W�| �n�t�TY�c����Wdt�n����n�N܊n�&|{Vu�
mODB���{�W�| ��y�<���7�5�#Ē��C&j����f���կg�{ͻ��9ď8hޡQ)L)��T��@37w�O�؈�q,�ݻ�ݞ��b��'�B51N���@�_ �����k��m�@>��aq�&9�1@n���턞�7RU`k�Q@.��/�ij�CN<q�RDI����iz8h��z��r�����q6����O[�U���ӧ�x�wE�_�s�m�5��Ȩq��  ���9�I �6TWa��$��9�7N��E���[n�3�N���X�Xm�6��4;�nv4�mۆYfޓ5����n��e��
�{6�����+]�n���,�8�m�J1�zAV%�K�K'��h9���@�Ff�˭fgY�7�ݣ{���S���ε�����S#�qmṽ��pֳb�䪠�R�LUT�eD�Wl��] ����Wk�����veǊcM̄JF䋀�����|~���j���wn� 9���5�v)9΁�v�}m�@��_ /��t�2��6�T�HP�MOC�-ǻ���n�@~�mt+��}���B�D(�7;�9�(�������J�m@���l�*v�]���`�@P;�R�\��@��Vץ�ݭ!.�ԣ�!��5S���V'�z�7{��r" �"<¯��}U_���F�)���B�>��s�S�>t�� m�k��M��Wt��O���[ғ�%��2c�0NG�/���Wk���Kٵ������3&X*�T�LL�����s�	ν����uX�9��oz��ˏ�����9 /��tWk��oz�Z�w�Aq������rYe��>ki��kgѴ�����6�bγ!UӮK'W��o���(��W`s�Q@y*��e���R*B�Jjz�7w��r"���������w���F�F�5UP(��B�I3W`5����o�o7�A�9��1���&���`��&h"���j*"���+���"��g;��U��~��Uw�b)$ �0�*&�����B[�w�-{=������b�3.	UB��������5�(��W`s�Q@v�t
�椱
̉Ơ��S�%����W;7���s����e��=M�0���2c�0NG�/���^���m�@=v�߳պ
bf)"��7'z/7=؈����[��f����ۻ؈�BFF�ИJ�J�U
�j����w�玺lBO7v��vz盘H�UU5Q**j�����%����ݻ��\�t��U��y��u���΁}oBh�x�F��޶��s�Q@�*�\����w� � �۷n� �4�m��`��Nn�'�u�(&�)�WY�O��]��$��Frߏ������W%V����+�3���w�LQ<n!Ĥ\ ��y�>V��7���ݔ����\��&F�'q�Nr�>m�@�6�͎G9��u�@37w� �V¼��S9�rN�[{�32��y���G9	{wk�}�׳EB��reD�U��L�ř���ۻ]�m݁���Dr����0�8-�Z3���'��w�9��\��V�2�����z��d�gO��}���kgms��&ĩ�=�H����,e(��헙�!,d�bxͱ�5��m���k\s��uŌn���y4k���ufvGsk�y`u[���d���V6�VL���k�J��*����P�6����ƀJ1�n�W�v;m͘8�;�n�a�дGRX�k���������{���/� ��{yL��e�\ǣp�Z�-�b�[�ʡv�u�Y�f����Պs[�ߏ�?;`6�g�w���n��<ݔ
`����U*������u��"#�7v��i�<o�m��J&"�aRL<L��+�;�Q@�)j�IO �sr�����Т��@��N j��1%4jJ���\LK<<cq(���o:��p���we8��2ˍFH���7��iL�-/U��f��:�B���۱�:���M��Ӹ;\�G259��s��m|���n� 7�o:����4���	�r> �%w�L�3��33K��(���X&��y�r!#��=ق�%J�L�UUvJ~($�X�(�I]����(���r �m�@>����v�M���>�n�$L*���'�*&��1%4%���P$�~6����������V.��Ҁ���B\�!$q�/`ކv��{mu	��v��E��yJEHQR���{��`fe3��|��ָ��5�&H��s�_y�����1%4I+��r+�����!$\ ��΀}m�;��y��c��y����I-�r�P�WTc����C������-���n� ��g@7ՍV�7#h����W@m�v��9��`j�ݫ ��8�[E����1,�	�X�8`�غ�:Kb��wks�k��Dg@ݹ�䚟�X����)�*�l����.�{�=G��!�R!�p��V�n�����L��H��[ȑU4�I���{ڰn�t����)�*�l��phl�i@X�MO@xۻ3)��mՆ�ȏ�T�9�j=�~��U�{k��()�"Cm��n�p
��:�m|���P�'����bys5���a":7>0�<,�b;'m�s�౶Ӹ��"Ja24�8��E�*�l�-����؈�G�1���<��[BUSQ��G$��-�����kڸ[m� ���[�r(�	�r>v�v�rz?$���䢀��\���I����Iށ�{W �m��|���.�{�=Gr��&2C ��$\�$��΄��\��z9=mMl��3
��A�PD�M�A��ٽ1#�:6�4��M�:l]�!�.@�$��hXnA�]�XWVk�̨�Р�C������g�R��DV��諼��.�}1��,�9���g{9��zC � �kL#L,�W)%0�S�NV�������,��" 2���8f���ƶX����A��a�Y�F%1�h�f����c_u��������~/�mZ�\��HyżM.�g�l{3V\Ӫ瀩H��:
B4"Z2�z{�n�v�;�ܦi��6k��t��z����ɞ�x�`�W4j/��|@}!�˸��n��n�m����������1�θ8�n݇6�ֻ�=	�O��g+Y�;�<+��c:^���$�#a�{rmĆ����C#�Z�6��V�����[^I����,�S��鵺��CʕD�ݦy�5�ϱ&�gT�������8�l�T�s�`UV�J�����EI�` m���MN���N��6���lm�� �i�m�Gp�պۉ�8�&�-�6��X��Se��Ң\E j�d �K�&C�ڶkXH-�sF87lNqm,l��M����Je�(-.hm�����j�0��@�0孺�q*J����m+ʁ9y�U�nQ�eX���)�Pq4-ض�t\�$[C"J�ޢ��� �.�#J[�y�۞x��c6q��V*�3����6.<��g�\팼�mbzsˍ�+�k�0��������=Ps�zN�{�������l�1�c�<�)�Ll�+U���v5���HR4U'3d�m�c����[6��pO]o���Q�_\c��G�v��v�$����3�YM�]���;E��c����N�f��8N�t�m\:Ҭ�0D�ԭg��rg`��̩���}��z���c]Zev�@y5�kj����UV��-B��&�F�*�+R�r�b��؎�ùu�C�u��i�m��;gm8�'��U�v��vlc�ն��jPv�D�wk�kSH�\�UӨȲ�F�̵h�gnL`'�%��X#av��#8�gKp �K=cq�#T����Ĩ�:׎�v�x8�g���MGP�P*�D��{b젵��P��u��V���8qڎ�l������|v��	<���1m��.<]�u�յ����Sx��G��:ln��뮓-�];f@ [I�5�7]Z��H�����������W�'���=!����*��6���W�
y˫��^�-�l�n�ӭ�K��-���d�z�Hw��vz���tan��W�[=���m.ڝ+h rYZm <�T��`kh���YEV�X6�ev���&gbB�����G1W�=�ѐ�K���8��v���lP�ֱxT�����7ezv�`��n� yz8:.�g�t7J1��\�xcW-On�w3��&�8�����aEc\�e�z[j.sg��ߏ�;����ـ{y�A�j��ӳC�.��Ֆq�Z�n,ݷ&�\��?�����~��j�;�=��t��}Q(��P�\��ށ���Vݳ�g������7^ΩDҊ�QHR����\�]�x��~��@x�݀|�ci�B�
2E�*۶t��p�oz�ڸ��EdC��"'QSU6(I�˕������M���{���Sיuϰpg�������3�ֶP��1��ӛiݰ�=4�E*�mTT5J�ׯn�̜k�5���>r��ϲ��49���Iށ��N}��N�F����w٭�����8�@xۻ����v5TTITE
��S�ڰ>�mt���=�L��Plj��sX�W9��3>�j�w`{2��؈�ql�ݫ�莩��DҀ�D��m��ݔ�m�t����5�84�2cK�Q�Hh���m�x�������mǧ�:ٹ�A��E���<Cm��n�p
�����DD\Bz���-�*J�B�(���5����"#���-ݞ��wn���N��P�8�1N��rt�nz���[�Aʦ�����ڰ*�Zi��F�HLI�8�oz�ڸ[v΀}m�ﰺ�D��:�JU]��8�@�pmm=��=���.ݽ���#�'q�S�iƐ(��������]!Y�u�켷a�%��V۰�n�,����E�o��[g ߮��kڸ�X�I:�l��.�s�`�Mع]����5.U`rH\Bl�i@Yrp۷���� zݼ��l�z��h�qdX6�qv�rz ԹU�g%4����f�DZ��-C���,��N���Q50�!�f^�$��3��RJ�����jW��rbs!	"s�@d�㭭ݬ�j�u��s�D�#��1�D�H���2��"m�f��9)�5$��ގO@گ:��m\�6�)1'$�[����$c��������t��C*fAB��JM]���΁k3Y�H��� ���ށ�=��9�
D9���6�)�/����(�9.���N���5�w�rt�l���ށ��΁kَ��=Ȉ��P@	'T�����eb�ч=R(`�\Wk�S՞��0���WY8f���`��d,�e �e�mT�B�m��Z�z�#����3��Hu!ڌ`I9�ۣ���8��� ���4nز�㶒6%��)�/��;�sں4�=��ڻL8ز	�����s�*ك��;���E�����8�P����w/e�&�q��s���.�ju�X��u��~�6�m���溑z�4n6���G	�tZO���>9x4O>}�:JeP����)P(T���gۻvfS:��u`|�s���/{�l�B�M̩����m֝؈�!#��X�v��1��G8p)'d�
�*
&�t~K�IM{ܮ��O@fŁ#$��P�9:��p���@m�:Ȉ�m���i�$RF�(���p����)�ݷ� ���;�y�C*!��i�%ȫ�M���X�|��8n��pm�=�.3��e5V�)?$�G;�-�� ��y�m����z�.LH�5!�R	Hp}�U�y�b)S@nrW`$�j�"	�-5T�B���{`�]�ݛȎD%���@=����v@%)J��ӓ�}v��l� 7�o:V��=�Y^��D6ҍ���S�o"#�^���j{��>x���0s҆J�\l��d��8ܓ���Ź��z�֐vո)�H��ZB]�g�5l<�L���U����J��Q_;���J��*fP���]�{`j{��>m�����ݷ��VTՊcQe�"f(I+�;����{���5�vc�H2�B�K HHB@��	"q��:%�9�n�΁W���A*�k	���X�j��L�f7� �n��/n��`m�ɍ�� ) n���(�1$���R�3E�A��:����8[L�e�ڑ�pMj�:S�i���{��d���6�lq��X����t+k�[oz����΁n�04��R�P��]�ۻ�s��i���lWj��Ɏ6�DF�nN��Pw%V(I�I+�3��\�qUIL��
��]�9��{��1n������_E'�!�e�f 9�!s��r"�7��a���EE*�R*�iz��%$���������~��~�����[7���!8��[t�bR	�Ͳ=�16ݍ����	6���ȯ]�fr&Xx��1%vtrz �Ԫ��V��q,�ְ�S�k����\ ���l,nzͷw��s�����T�H�*M.�6�{`{%��>x�z�ڸ�MC��X�q���9΀{���cw`{'�lr9	<{���l�T	T��T���<n��OU�y�����tG"#�Ȏ\<���s��P�]S nq����f��:#�\q�ז�ݣIlΑZ�	:�]�F�*���e:�y�P3F��Wm�P\���)��������5��b	�L��s�8C��lޣk�d'��kUk�n:CHI
��]�k���[�n"Wr�U��s�#'�u�2ҍ�=��x{�U�n������z@x�xiϵ�-鵔`��7V�w~������{+^ŷ5��4��P,b��\ݮ�o(:"�]�OY����>*����>s���c}�y�������p�ĎH�x(�6��[o:�[8�oz��p|{J��DG&K	���IM�%vwJ(um����v<C�����p���ݔ���t���=�\X���Ҏc�s���\U�΀_m�n�
���Ds+������%*���.Qx�fp6�����'��Y���gr���]bA�d`��0#1�D��*���| �}��{wy�=��\ۦ��`��I��UM��9=c{�����7��HJ��'��n�a#rwTĮ$�T(EM.��wn��Kk�bm��<���kwE?(�MG'z�ڸ��΁����m�@>���Um&�Qj�z�mՁ��OU��wn�i㞀_g�+�ҙ""�,�IHcM

e�%�)oI�z�չ��N<5����i�t�f�!v.5ʨ�O{ڰ�k�cm݀��;h�ݫV(#gjQ!SH���5K�cm�@��|U�΁kڸ�5+�4��1F�zWk���t��{b��(JR���i��1ƈ���%2�	@BR��i�Ck1�Z�pGdGr'�:BL������T�V-���QcE1%��+�y���hP�	V���H�d�&�Vu�F�g���z�g�C�'"�����]�,K�\>4�d� ������"�*�"hh$�"��Zӭ!�dQBUC@Hi���ri�(J��*()���2̂� �ѕ�%,:L"(�� �頦 ���&��4DƮ��O���j�	�k�&��J@���es�q���9ސ�H������wh��&�����d�T�4�4S��4�l�h���LD皎�L4�de.��Y9�bq�S���f��tt����2���M�0&(Z� �gYlѾu�ф�{	H���)
B�k�w&�fk�f�{��	��;��{�h2C&��IҧqH�H)Ü10�:�w����r\
HJz�1O<�A$H���]=�����[EE:��u��G�z��0����󻮍�� �5�HA'xg[�@�B�H��ҍ�;B�8r7�yA�y��ҭ����mI�M�-�a2�L��z�[�Q�A�(x�bq���p����(kʼQTA|;P����~�ʸ�[{�=�Yq*��l�)MT�M�Vs�tm��؈���_ �Ԩ���x��|�����{w`4��@���X��5-�ԦYVC�d6���9�XN{Z��9�u��r�z�/�#-۳��,q�h�<L~6߯��݀��=�u�Ȉ��z�a�/��#�i���U����΁�q���ۻ؄���mВS0*EL�O@i��X��m��1<s�Ǩ���C�9�N���\���]U�o����,��?L,B��wj�����*T%D�A3T�����L�cn�9ƺ�s�1�.85V㸷4��t�sF�É4S��=E��㳻Yر�u�H�<��r�gR����֝�mՁ�8��{�v�'AF����$UJf��f7W�ȎG3e����vy�:��$L%c�$cŝ�''@�{W ����o���U����x���ȒY1b����Z�w���6���x�{�sa�87�ƚq9;�7���5m�t'�z�n�
�G9�Ȁ���p�f6�fVX?���������5�-��a���BY�!]�wZ�u�$:��҇�]�@i�4hK[b�,C\l�6Ht�Z�=n4�;85 8���]�*[=�.5����m�֭��㶗o/��n�G3� AK��8W9��Ƴ�uGc�3͞,�ς��K7X��¼k��0�
�f�Kb��-�a��ȗh��Qz74�vJ�����j{��^�w{������?0�������m���ll�\hb�܃/m���47hӴl/%�UT���ݫ�㞁�ۿ����]|f�Q1��!PU���'�z�n��tX۫؄�X�s�SQB�*&�5S�3wv��tX۫��|�����21���@�YN�m��y]��]���]�Ă����B�)"�m�tWk�m�����7|��)1��M�𘍫<p�m���"�\��ǵe��M��b��Ф�1����j�_ �m�@���V�g@/�ŉeG�$dŐnf�Ԓ�^������f����?+g@-�8�U���Ɵ�"i���@Jz��S`	%4���.F�I�jNE�5m�tݳ�z�{�-{W ��x�F9�H��Jrjl.S@o$��[	=��)�>�w���Ϗ�j��q=3�8;xn9;m������s��u�ڃ��]9�N������S[�*&��U|���˰�3�ycn����/���'��
9ށ}e(~IM�.�4�J��<�0�����R�X�z��WE��9���""!�ܞG9d�ݻs+N���! trH8�ŝ㏠m�wm�@�e8V����5cřŐrN��݁���!�z�[�z~̮����ɰq��:y
%f,� 8)�ն��b���g�'FGûc����ݫ:�
�)�4M1I;�<�k�[������oz�cm�����m8�V����]=�݁�N5�h��R��5�4�n���lٻ]=�݁�N5�ۯ�uya�9M����p���Uw����W�����I"�R �d�ڠ��~{�U�^��ٛ݌qț��kڸ[u�����cw`o""#��RE�����$�LԆĹl�c���r�u��%��n,ڥ�"�vs�,�L?4A
F���U��}���w����<����h誊����k����S@grW`gG'�;�s����"8�}�@�EP�3S�{�`}��t�Kvu����s�>��M*��X�9LRN���\�up�{_ ��{���������m8��s��t������(��k1�y������v]��7eh%���GQ�b�b�����j�vݶ��g�x;���z�\�re�g��B��*v�ݕ2;R� �zݝ���b-�Q��Q켣\�vu<�$���wn��I�:�z�{np͸�A�۰u��Tw\�zP�r�)l�:6�F�rj�$;��t��F/A����ӕ)����LtGY��v�&v�ju��n�[m	k�q��Η~��]��{���\{�\�p��]uÞPJm��V����AcC��v��"k�����{JQ%D�G�*�f������n�,�<���W�=��bl���ۏ�grW`k�(�9�tP��c�uJA1�3��@�ݯ�jۯ�u{���m�@�,K*��I)n> ��Eo��@v�W`gG'�p�v9"F��x��-������{W �����}�@\�&L�~pRlpYg�K\��N�u��
]���\���}���۵gIe�TȢ
�r�jl׻v�8�@����:��|�m����"i��:9=Cl�vif�3;��=>�E}m�@>�
�'������y��(}ފjJ����bt�e��?,riNq���|��ށ����y{u���y�O�4Lrcm�����ގO@k�tP�t��\P�g'��m8� ��8ێ�P�my:��nv's�e��879�j
Ø�������������������O&c�Д�G �����vpv��-���V�$�yǝ㏠�M �%vG��=�Drz�;�����l_�ŐnNn�ށ�ݯ�j���^����i�1'm�'z�v��ۯ�u{u��m��DDz1�3jjjf���D���!��rK\���d#��a�b�����T�����G$i��m������n���oz��\~��!21���Z��V�7]�$n�۰1�Ӡg�1t_,<�I�Ɖ�n>}m�@�� ����}�8���Z�pQ��M��(�;c���zhc������Ѩ&�&�I9����uW�ڹZ�#@�iHp��\ ｳ�[���}��UJ��&$��yڒ�.��)W��H�]�є��<��R��������yǓ�.�}�[m�@����h��@>y(�D�P
(�����"3i�Kk��ep����D�N&ێN�{e8��W ;������뛊�#�8"A��Z��������������v��~L��Js��[g [����x����}�O@���J#���D*���U_��������o9�n6 ��"�$QD3��" ����j;���UZ�>���������_�y�?�;�?������߬ߛ�9O��������������1��o{������������yAUW��򠪫G���������������PUU�����w�ӟ��o���c����?����s���/����e���?������͠�d
$��@@)�P
P�P�D��"�@)$�$�)2�L(�B�2�D�*$�L*
�0�K*$J�B��R�D��
$� P
P�D(��J2�J	
$(ʉB�
C*$�D��� *$"��J�*$ B�(�*$$���
@B� B�(�H,��)*$��
$����ʄ���HB�� �*@@�! �!�BB
� ��� ��2��� �HH)! $�0��2 �"� �@@(�@! ���@��� J�H���2H@@@@K!�$�@�H�H@I!)B�H��	(�H��@��� �!*�!((! B@�2��!*(�H HB
��
 BJ!�H@HL�H� �!HHL!+,$�	!,���@�
� J��H� H����(��B@ H�!"�!"2�!+!) B��) H�J0�"��!(HJ�� D!@L�� L!����P D*� �%U2@��%!	� �!�%� �& ��Rd
@�!V� H�b��)!d �Q%!T�I�	�	Q%%D�L�g����?���AUV?������=��<-�����UU������������C���k��*��������}3�*��?�U��:�T"*��o������������?�f���<?�f��뗟���w�ڠ��7�_������AUW���27��?��������1PUU�Ͽ������w��������2����=_����C9��?�9���*����xg��ٰ�T?�濗��3��}���TU��z��7�����U�����ߩ?埖����1AY&SYZ*�n@�ـpP��3'� at��  �  �(U(T � �S�  РR��
@/�(�E PB��U(PT�
P  � B���QTP��"@���� 	(H ����    XH 

  �@Y� �Ϧ��{Kż�sżmqgYp �W7^��oD�vշ'R�  �Tź�8� 1F�� �Q���e�wr��!��4{�D糞��ﻏ��|Y�m�=ڼ x  >"�R� P&a�(��,� #�h  � � 0  "  � �4� �  4�d bS�   �4�(� � f 
$ h1� P �
� $ �,`(� DAz���iy��J� -ONO{)ɮ���^��/' Ozz\m�r��� u�4�g��]� =�r{���e]�ڧ���n�/��y_mũ]�>]92rr���  ��H�
   L`�������m���#\�@ ���^��ew�׽��ʦ]�W ��!�o�zy;� �Y^�w���w��
����﷝<��^6.NO^�{���>��W�����{�}o�ө��
UEPP � �` y�=�_y�WNM]��OWk� (o{[q�m_!�����,�. t�O]=�x  {���^m�����)���e��r�.�}��@�)���ɪX���:�     ����T�@ 4 j~��y���   ���R���� "{JS5%   ���(��J� �@E�) �58��ߏ��?�?��o�f�}���Ͻ��"*���EDEW(���DEW�_�DU`  ����� i�XU���b�#pd�p0�\
�����!�H�F0� �1!� 		!0���c�cZtP��y	.�;^��/��ͼ��*Ef|f+����=J��{}�5R/�^Z��╡Sy��s�$�AJ���&!�.3�\�F&�pe�1̰���N��OQH �!HP���}ǘΦ�Xc)���C��Y1`0�XEIِ̻ގBq�>�Ӷ$'��>���lIp���, �Bbwz�ۇ��shBfP�E(&� X����(q��C��d.7�.3�����1 �)���RSшۣP��i��3�M��|� �p�IC64!HT�A���.a�1)��!B-���ap(�!B����;��SSM��@,R�-��#dBSl�*�H�P�
Ʀ6w�f�j��9.���)	�b˲�8A�$n�YV+-�L:���xX��/��F�\gF�kA3>&���ѭ^|K�	H��@��S	������+m�)���SD��K�M�l%¬B#F�f9���)�$ �}��8��s�^h��x<�#kohΫުV��a1���&s�I��ٓ�°hXH���e3^�.3���K/7��c�$��D+Ys�������.���T�A���X�`E����6�(�
hX�$p���+�2�3�.�M��+��X��U� P�Y�F����9)�cC{I���Y_o��޴������}���ѧ�2D$(B���+gZ�9�5J��	�0�eM)łU�SI!�c�̩
"�!$+�L)�aBT�T�KX�X��K�-:���Թ�ֳu/�ұ���
�sJ�H��%��2�3C���XHR�%)�#���S�鯶Rn�2�\1d�pi�G��a�C���	+�>p�qs�T�R	�BA$�"�$�H�IE�l���B��`@�H�`Bvs?}�JbC�@�Jʆ��W#�5�$>Ʃ�Ή����rA$a�N�2����p��y,�Xe1�ep�!dH\h�d�R�<���5��.��k���1A����O�����@�(�s�o9���	脄{�(��Gʞ[_|!���1}큓�;Z�dL7)�й~���-	6���3�3 kL3)YJ:2d @%J���%I�Seɣ38�^.�Ja#(@��D5�L�@+�k�d�^�t}��m�@��qXT�R5�a�����ЉY-��� BH8m��BS&c��&*cf4cf�g�:�b\Z=+D	�%kP�^k�Kz�2�f,�U>�m��'�yR>Y�^	5^�-2���|�V�}������-X_�)��,�.1󫹯�c�Z�_�ۃ�B,a!H����s'>�d56he��t]�y8ƛ3  E����4h�Hh�D�ѻ��M	�@��� @� )B�үo{m�O䨫�E,��:�I��p��K��BD�F,R��)"\2�W$�� H��T�YDB.L��3JC<��X@�bGA
D��X�o�p�חxTySB��ʅ��j�U�"�|��b̦LvbQ�4�%If���G�U�Y��[�|��Mt�˞�6,(8ι1/����C�+�<ad##�H� �-a���{�j�Z/>׬{���M3�b�b1)��~��k]z�J��Ņ�9���!�-�����~6�.3�˝�7[,��K���G-�,i.I�t��$!q��$1���p`�"@���.3��#!@��n
�$�#0`l�GZ`��.s		
\D�BK�}|Bw�A*)$jɣ�������!���[�&�q����L�"@�E���^"�*-x�/b������>0��6������y�>��׉�Ɲ�q���R�ꗏ�!S^���ƬL�[�q�w�f,�#BP�ILl6��-�D"��BY�������Hda�<L��
w�>�s��(�FS.>�>� �B�b�AdF��y�fh�4�&�X��A��~�LB96L	
���$#+`ՁF���aXP�	F>&�n}�:�ε����gSa,p, ��Els�|���
�6�¯1��U���\���>�U�uu-�j���p����!���$�Rbgd>>���6�	�ƍ�y~ߋ�r�?�ܾ�|+H���!�є 5�� �B$E�@�$ �*E"K0ġ#
�(Y ���q�W��2�.��[W˗�渵�rR������,Yb�B��5��{��ej�ߊσf~ܸ�7�C�����b$cN$)�A�0���.�4��c)s����%��8̙12J�.S&2Ja�f�!q�IL�����cB"g;���Y6b]�i4I���0_�6$c!F(Q��G
e�b\g�t�2hڑ��xI�m�&"��y�����5��!re`�bP�wzFB	����hHG�ԡ���]��*3v��^>~��U��b�=�H<�Λ�x�Eՙ�����jJdhb��.2SYߵ���}�$����o����C�i��H\ �a%�q�ϳ��ԯ�B�bB&tf����k���#�k�����iHZF���3FL��ή ������LT+�QB�{���i$y%X�ގ��4��B�%9���}�&��}��� @�^�\#�=�~������c<7���="�CUd!�d#@ Gr�Y#��I��6�.�M���x��0��D#"�h<����ތ��Z�0r���e#dzrH�`�D��;"� H��H�B�wzɢ%�b5H� RA�A$X�,BF��`�`L���.q�a��U���
ck��$!�%�T�%	�\�S+"HT�d�A�!���K�Z.r�� �$%�1&
B�*I
D)$R$Y2�4dٯ��]���z1a�B ��2%�E��> F-�" 0 W��Ϯ���NB�]�O�}�B\r1
�V@0�!G� t�5�\9�4B�d# �0n�;�5�a H$�R%FY[����	RNO�ɈYN�@i��+��M
�����J�A
I%1���.Ld���း� �F�=��A��,����)��e%�FP�&�K�����̌���!pI)+�!Lfb�[e�MЪ�6�]:�}Wږ����BD�$�#RHŉ"��R}B���f�rF+�-RR D�I FI	
ő,*�X�S�#M`�3�1��!R�L�
d%HV%�_���`�$HF@,a�$+&�!N��ꘟ�mt�-��C���/����9�3&L� P�d�,�2d�Ύ3���!��	��^�(=�y�-��|�2�y�4|����0K��'a!��2�䲁
Ka��c�P�Bc?g��o{���D���ư&����n�,0XI ��>hBY�Y�D!ZB75O/'�'_T�<�V<�I
��׮�o�<U��u�\�ԭ&�0����0�ܳ�n}ˍ��F\ꔵQ�յ{��	|��Z��E^?a)�1�������e<Y!B<!tF�1��gP�J`2I	.>Ʋ�����>�m��zHR�J�H?�CF�$�SXu�s렌~��
c�5�+�bc��BE�p�Lv���ƾ~��� �"H�I6#g�8��\g7(���oj��L��f}�W���G��B��$!����Ii0��
��+�#�#R���e�~�)L0�j	��o&3�ˍs�`Ō � �,h1�@� �0`D�I�R9�b���mX�T�yK�g�U����p+�����޿�����.�����{�bAVS��G�ZMU��yY��Ϯܳ_���v�7zᬖa P6�!��n9�q�+��0d�e0��F�2h#L9t@��HS��LC	��p�FHP�D.B5�@�	����i�:�	\$\d�`S�����||ˉ�HD�LF�`aXB$b�H�c��
��k��R�.�D%BT������>LZ��m,��3   ��  ���H    � ր �`	 h U��e������G�������I���jٶ[��S��tūsm�����Wvf�+1�t�ua�H�-�ŽV� HX�6��Y���$��ۋk�p:۶E�I'2�H9w�2��N
ݯ�����;=Umhs��  �V�l[z� 6���  � I#m�m�]��T���Ur�5R�� 8$�Z7�Y
ݪ�� --d��Z��a3�N�] J�գ/\p��u�:%t��j�-a�iV��.�U@�jA8�ae���-�L촒Kd�i#u�m�8�Ҁ-�H׫I�m� �gZ�6��%T	@n�PR�@l     ���4�3�q��'@      $  h-� 6�    l ��`m����]I�    ��X�f�pA��> ְ h��l��зe���At��j�T�����	m�4�U���6�k 6� pd��h��7qv�.ـ�ic ����   m�褵�����Z�5�fR�.�Q���*WC���nI�+�j���t6Ѥ�]�Yqn�QmP��R촫i��k&�im 'M�����j�t�ʁ1@9��)l�6ٴـ���.���j�V�U���kn(��]6*�@j�.4s�� ؐ���Yv�P��vP��'Zn���K5^\�jSSGmU*ҹ�(tmʚȶ��	�����*�[UW_.��K�=+��Vv�@6��2�ji*��M��3TT�Xku�)� m���  ����*�p�@*�PP\� �]�kjmp�I��� 8       $p  �r� l ��tY [\�[f[Ra��Ç�v�c��m�͛` ���kn�-����%���Wn�!ܲ��TU��U�8Y�G1�-Ƀ�1��7����9N��*�N�j��mɺ�vӈ�L89p�R���;�{q�Y�L�g�%q�ꫪ�H�rm�	��ƎT�R�E�q8+��Tr�u�q̃�GmI��PM=��nh�{#VIg�v�[^K��J�U���D믥��Ŵ��`e�f��;"zq 5�Yzh�Mn��ԫZ���u�B
]��1�%�V���
��P��&�c��Rn�v�`ء�	�55*����@5��4'c` �-�6�,�eK:m4�d�Hv�I�W�$)��J��.d���։ mp�If*�ж������ͮ8ƃ� ��6ٻv`A�˱͌*�iV������[���   �Z� %�\��^�)^emm���k��[aܙ"I2�n٭�u,��T�����`]6��m�-����k.����@4�a�l��v� 	���m�mmKFNY`H�-�-���U���YE�m� 6�H ��5�ۆ���@��@Tj�]�ؼ��v���mnPl N�Jm�]���׭m  �L�l $ƻ   H 8	��s�m�� ��K�{H�y��D�us' H[Ym�9v�-� [���l�    I"�   -��)6��K� 5�n��v�X,�m�     �m���8�,�׍�K'[%87E�� 6�� ���  ���  �ŵ�K`�m� �]e����@ � 	   �mm=i$�6� �vam�����-�	  I  m�������y;"�88om�$��$]` ��PL�ԯ5<�޷iV�� � ��  �m�am A�n�I6k�m�L�1A$�5�(6�G��[d���l��� x�l �Mki0�, �5�	   6�5���i�Ԁ  ��b@�   q,� �l [[l�6�6�zl$ _�����TÉ�mm@ 6��   �[o[ ��`m�$8m�   �g�:�]TmA�'ʡ5A��t m�$�p�`   �T�ٶ� 	:@զ[Fհt��   �$�UT���
\��.�B�kp ����o_d�D���j�  	�e�������������-��  	���$�8lm�  �m�[@��*jZ lh.M�#n�m%�z����I��%�`oY�@ �`�Y��Lm�8s�6���knm� ���l�ێ-��VV����� �U�  [u���b�l �� I�`��#��  Hz������S�`[m� H��� ��$��Z�m82[�����}�,�l��k��A��IC�ҵ#�AF�,L��Pe�-��0[m� ���V� 6ͳ�[��#� l�� -�'N �       e�����al�li7���m�@         h�c�nܶ����hKc�����g��Hp�4UꚂ��6-��kOn�61*�N���i+m�  �K(�Z��``*H��	�m5R�5�Wu�C�	�A �U`LP ԫ@s�޻c��;��m��$[BU�W�^� �z�Gݸ�,1�����X���B�Xݢ��GoAԵN�{jmIUJ�z�g�U�6�u5��� m�Y�'�y�zi�mm�̲6�y��u�^�j�6���P2<�M���*經���F��r�	�VQ�m�6��{'<v���p�kR���-�tY����C���ggIӮ��y5�]�s�Ħ[ɻs��ٸ[#����=� �h�&wt�p�p�h��cH�������pl��UTj��t��4���ݶt�J��ؤ�m��.�UqZ�֤�I#�6ٴ�e�V�i��*r��U��S���D�YF�ig(Qs��)K�G��+S�Ƌ�l�f�D�� � �l�mZ\�p[[lD�dNX�Tq�U[J���D�ʵm���e����E���6T�p�if�Kl�:n�g�V�HH&� = qκl 6���Wf�"C�M����N���m��`��^$n����t��tHl;.x�k[s���pm[q u����M�-$Q7@u�� ؍�9�p��c;bA���M�٬���(ޏ"<�T��
Uj����v��P�W�;T���W�=n.��;t���-��[�����a�B�!J�9�k(���5@[UJ�3��[����5��B�^��^(
�ٶ�HH��$Hڤ���;P�.Z��O�}�F������[T��Wo5]g-�n�R���P*���&�̶�l ��D�j6�\7]pU�[U*�;3���ﱹ�$����m����l ]6�m�  [@��   ėu�ۀ �-4��m���ֵ��m�$�i%��l�٭` I   �[ kV�mH�6� �M�.��� $��� [wj�&���l�8������mH��M�Z� $��:��nymk� ,ӛxf��]�c���[Kl�nY �a��v�h�k]-��h�C�5UK�( �Y��UUU*�J�<����M9&��jnٴ� v �m�M��=�d��lS]UO
�H�6K[�8���m����ds��-��Ѻ- h�֐��!�n��`p�Nu�d���P�@j������U�y�B�U��)@����'9m�8$ im�`�i!J�M�m��l����m�6��(�    2px5��@8 ��86��-�����E�� %1�]����B�r�;:�e�p9����m����d%�'9�Dr��` h�m�{^:����[[m2s  pm�X�m}t��[Fݰ��dl ��-����;m���:}��^Sm� C�m�α# �֜�� �`�HY���XfVګ��B6�]T� �1t��Z�&<nKr⸵��܌���֥�\-��B�6��@��g�9�M�@p�N����i /S����rI8� l�kaZ��9YZ��j��eeZ�˲q*�Y:a���']��z�n�Umuv��xr�+Xm�  �$���Ȑ�L t�fۀ�&�v�܅���M0��e�+�v�e@eZ��U���l\����B�ҭT�\���[$Ε����}��[V1j�Vwn9ҷ�U���hQ�]#Z�1�3�9���6SUO&��3���	6�;���a�f|����eU-�	�]��:�X��t���f�}����3�T�<�U�c$[����zܯ75@��htt֪�v,������Z]��!B��q%ɼ�Z�@4,�z����<S�b����N�N��{�
�^x��sUA�6�5�:�$p-��튎�P�ԇL�U��E�e���yZ�8��6�� Is�A��i&�! r�ж�H��� �`6�    ��8 �    �� 	)G��o�C���T T�]*�*�A<���*Ҹ@��Ċ�����0�R���Q\��t�DS
i2�O��*�P]�T���b�@M��Y�D��0��H0P"H�@H@��"łE � ��H���	�@�u�_� _�1` ��@�T�)۳�~�(@�t u:�C�Tt�?@>C�l,2�,H D����P�M!��AG�4��>��� �4*}��@"�)��h���ES�@ ��ٕDt�t-@ا6��SJ�@~؆]�� =G���`��P~�	��lX�!! �Q8(8_�P�#���T�p�qG� Ep��� �
*��0��T��P �! �����Ȣ|��
#����T4�A ŉ$D`EO��e�@�Q�Q$^���@��bD��H0bB*| �#�`��0`1 ���(ew�F!  ��)�E��(.�	� �Q2)��U]��T? )i�Q�"D�+�P��W�GU��X�&+�zN�ow{������p�v�Hݶ^��B2mO;��bm�x��!6tt�Ty�[��H��^�S� ��1΂`��ui�@��d��˦٥V���l�bI.��p-�jۀ�`ky�;,�\h1\N٘�m\���[(��6��-3��Jsh��;DL���Z(@�6@����q����[N�,�%�r�j_F�ӭ&&U� ���m�U	������ָm�
�n�yv�yt�&K�DZM�nj8�����0�6��{ϝ�� !(�ֵf6���駎�NcRRە�ݮDP;��[�Q�j��)v/!��s!��ݮ�0g�4��m��9�U����y�n�u�p�s@��5��l�v�]x�;.�9U*���@��i��@ܤ��
�UUr�����s%v��Pe�j^v�����F�]�;$Ys�r��(OP�l�f�E9i�-��X�n :;V̔����v7a5���v��Tf�m���5R�E i��R��Lh�WVR�w	�0yc`  �l����%��N�[���H���n��2*��-Kkm��Zm� ���e_EHIgIb�h��8<Â퓈�7�z��ps�.���h�\f��ZY��:wg;���Ob�\ܹ�6vV�@*����"���̣�g;��N�vmg��MYWo���k`�k��ղ�-� @��p�Ҍnπ˸���n��v��y�]��ul�8�gi���4�v��2� +�.L��î-�ؼ<=���V�*�;jj�ړ�t����P/l����R�W��6�N�GO:�E���n,��<�h�͓�M��'�gV7s6�\���]=�U$+��ٮt!*ti��=6�Vl��m��x��,2�$t�C��n�ͻE�Z*��]pJ���V�b���G>c��u�ױ�;J��#��7f���8��خ���@S8m�d����Nm�i��0���cy뮑ՑKu���8�	�Omڥ N����"sD�R���qO8���m��@���D��e >���S '�G��T>Z#� ���0o�[�t�M�GCθ�ʬ�"���嵉� ��aÁ6�KH��#�ct'U�c�����3���;�U����� ps���؝V�%��S�d^1�1���A:��m�;�=T�C��5�bƤ�!�K�v'�st]��������Cn�\�;B�ă�Pv�1������ϕ���\���O�5�l�)�e����{�������"8�^^��m�`��	���QC��8S�96||u����L���lޟ��mwN ��)��ǑH�����}V��U)�w�ՠu���6̙	�Ʉ�H��d�4��2�ҘIP�h�$�$�m�f��۹�u����Zu.�i���#�ؓbs4nـyֹ�7X�`��`
"]���>��M��N5�K:�[
G�<���]�Fy0%�Xw<�m���P[i{g�oS��7Yl�7���5�f��)DEe�b�B/2�Ѝ?���"NA���+c�����hԓ��=4k��iV2�(�D�C��v�i��dK�L�F�.]R<o�A?(���y��hW�h���������[�|$��H��#���_J`}�Q�l�0&�����{���~�y�P���S�̖�e�jx�b6�;��$�˱u��ɡI���y���/�7���0;di�6F�S��=�ʏXa1'�%mI�{e4��`�����Ŝ�d���4E]+�&j��0��X��>�	y"!(E �Ei�)b$"��j��s���s��f��>�N�y�&���z����h� �푦�a\QQY�b�B�̶�*4��ӣL����㿾������U����9���x�G�j�,��J݊:ݒM�N[�D�3Ux�� ��ti��:[{�4�;;9X��Q���������č�}X�=� �;f���R�e7s57k ��u�{v^,9(Je�_�� �]b���h���Z�����0;fA����	�%����V��	�^�ԥܟ�'�%mI�{cL��06�K`}�Q�oEiݣJ-V[7NG�R�,�a�vpVM��T���w6�m�*�Ξ��폤�06�K`v�`v��-�Ěw8�6��h����s@�m��<��hz�p���������v�:ϻ��ϫ �q�Ͷ�k"S#j1�����ߕ��@�߿4�ڝ-���i�r��e,�02�WYx0>�4��})���i��%43����_,jDH�l�������l{�yZ�U�]nR6��\�q�#@\G2�T.ki�q9ӳ]���V�nQÚ�W3�{/-!/��X�C�7	�:��@ն�^yy��.�9�Bjg\�R&#R�z���}ƨ���9���*{fxB�b��m멕�k��~��}ۮ�͎��]̢�k�GD���V[��K/F-�O�΍�@�8�b���Tz������υ��Ca��q���Z�N�m�al���vx��,<\�:"���a�gB�"O�N���@��.���M��M�W�'�b�~ra0R-�x���(��b�<��yֹ�7ƌ�Wp��$�m�L�;�w4;�4k�=��hZ)A3l�	&���{�y%[#�0;�����x�0;di�sۄCŎ8�iHh��h{�i��#L���Iw`���e��ƙ*QK���b�ԫ���ks�ۋ-p��79uG�o�)�R"cx`�^�S�X��X۶�P�(�_HoS��=���k>�IȚ�s4����3럒F1d��e�� �"H@/\���*[�������07z�� ����0�#RL�<��6_J`wq`v��r��+wT"�������P��[��gb�7��h^��/uz��,��&"�;��0;di���e���e�Dv�s7jӕ�"�5�����g����lqPs�6�l�pq��G �JLލ0>��`}/�07��	���a��4I�nf���M�����)�w�)�v{BōH��;����������2��/	,G�{��o�2�d�ª���+�"�)��Ր`v�i����}���K�X�����MHh�]��Қ��Z��S@��7��y�Uǈ9�f�7<�B��vV[��/E��&:�iF�E�9�b�F&���yzQ��������0;z4����E�*
.�j.j��Z�9B��[�ŀ=}��yzS~���_����"1Ʉ�H�	�~i���Ӳ���i�ܙ�cĒ�o$���M�Қ��S.X�����|��VD#���Wd��]�۶��B�[��6�����W��.�ňh�LrF�JM�Γ�mg�Wu觝��wC�V�����=�p�v0ĤBoR��M�컚�����t������L�����r�07{ ��� ��fA�����c��Ǒ���������M͙o,� �˦��(Uuw���2�Y�F���j��~!"O�4=����Ji'�s�5$���f���R1+���֝��\�l]{m� �i��Z�gd����8x���s)�!������rp�I�9�sO^��ĝb9�T�!,�VM���)7Z�˽�G��u[��� v�n-�q�^����Nq[c,� ��6�[�q���e�c&��[����Z �pΞ����sh�5����c�n>Y	;`��,�n�^����7��n�o9���m�ck7?��^�u���{��6�b���N�թ�6!�v�v�b�V���w�;�;cs��d\tnk��c@��g�`v�i��̃����Ka3"`�Q�ㆁ����<��h^��=��S@�ԥ��1���N��Ӳ�Q�oF��Ѐ�e�H��1Hh^��=���������XRꪈ2�*X���F��`}� ��vA��G���#�&2�ܭ�(�tP�z6��`���a��\�(-<)�z�����k.겋������Ӳ��������\�c!�d�щ��M���k�D�< ��Q�Y�M4�Ws@�zS@��.�%$�*���x0>��`wuF���`}�S@��M�Fd�xL#������0>��3j�fJ�UU[���c�b��6��<I.�*Z�K�{i�%풥�$��W��Ē�?}�*��c�Fң�p&����67Xi��.ا<�4v�<ss�vnp�������f�X� ?��ߏ<I/k�Z�K���Ē�r�RI\��3.2D6�C�K������U�x�V��$�����>�ٍ��`����7�&,�I�$�U�x�]Ϻ.����:F� ,� �U�R@�0f��"�dN���	q���&F��^s?�i������`}��2_�.B��8P�F"ΦlH,9��%�0`S8	�e2�I�ˌG�5���$q`$$� H'�����K�J߈�*�N�� D]敒��Yvo"�D4.�r`#��3�=�!^�ǉ�@��8
:>��"��� _�Ed��!�@:8�΋�E)�P�^g���Ē��E�$��"9E"�5�<�$���Z�K�{i�%겏R_f~����7z�><�$�Ǘ�b0���M91jI/=�$���=I%�q��Ē�wx� �;��Ͻ���������֝����G
�WQN�B\�8����Oub
��S�<�$�VQ�I/;��y�Iw;������i/z�Ǟ$����z��8��dNRIy�_3�>�m�_ۋRI{�~<�$�VQ�I/s�Ux,d&"$(�d��%���Ԓ^{�O<I/U�z�K����x�W�[�d��E �m�Z�KϹ����~��f5m�|����ۗ�AKL�(?�����m�����C�g&.K����~��f5m���O�}��9m�|��������Iy��l�ذqD`F8���m�L(&삌�=m\�ܸ����GJm��E������dRĒ^�S�3�K��ũ$����g��֒���z�KۄTM��4#j9�x�]��-���ن1�~�u��o/��[m�ܽٽ�TLa�q���$�M91jI/z�Ǟ$���=K����۽W�g�$���ũ$��܏������/������z�K�O��<I.�w������Ϗ<I/��4���~��2'�$��/��%��}���o��7�m��=�ն߱�2�p�ZKm�X�8�4�\!��ɹ��X6ٶ�4.ۑ�i	vyꃳ���vS�wB��Mr�.�sn��쪜qs�!e
���EVR�v7Z�k\��]�() �fx�gU#��9sn֝���ت����b�/q���ض�u��;��Z�v�kڱ�#2>͹��C���>R��pv|WI!��Vtmڭ�G��f�;�[i���D�\7?��w���ߝ��~[��#hL���w;Ne�����L��=7Y�@b�2�ˋ������w��0�f%��3�$���n-I%罴�Ē�YG�x�J�_y�x�__���Rol#M��RIy�m<�������z�J�_y�x�]��-I%r�j15�"x�!�%겏RIw�����m���Z�K޻��%�,9\Q�bɄ�Z���W��$���ũ$����x�^�(�$���X����<��Ng�$�s�Z�K�?g�|��Ԓ��Z�K��|�<I.�s�c�p�dg@�t����^v,Hu���/oX�a#�\��N3�v�՝`5m��5m�s]�ݶ��g���o>���(�b�k�RI[�oȋ�k�O�p�ĕ���e��p£�q�q�^����{�����y�߱����M=X9�H�b�RI^��3�K��-I%罴�Ē��E�$��z�Kđ�`�Q�5&y�K�Sw�NL�ϵ�}33�o$ə�z缼�$��%�L1�Q<#M�-I%罴�Ē�3�߼G�$�U���%��������������}r����uPX��5pnTN���|�Fy0%��M���o���p��N��Hm��rI_���Ԓ]�+�y�Iw9K�U7�[~�u��o.));|g�͔Y0n#RIw����~�٘�V��$��w��K�.�~�ʹ��D��b"e̷7�m�q�K�m�������H� r0�V�+cDdV0#1Bc��K�%� �$Tp@���S !�y~�}��F���O��<I%���d�����%������Ǟ$�}>�jI/}�g�$���l߅�$���i�D����S�<�$���5$�߳;�}�{�IZ��Ԓ^{v�x�_غ���}�	���v8s�q����t���.WnW�W�M��kb����̙���$�$y1'�I+~����y�g���n��<��}�o=�j�[R������d���F��L�Ē�wqo��?����w��M��{�?�f�������}����T������7!i�+q�LϷ������d�%
��Z��L̷]��$�e��ɦ\d�m���$����k۳V�yΞٽ�o9�躶�O Pbex�&�߾�ݶ�⒓�1��D,Y0n#RI{�e�<�$���Z�Kw]�ݶ���X����@���|c$���s24�D�	cG�Hz<����5�X�IC٥rK���F!O��<A1��Ԓ����$��ݧ�$��]F������y�I.����!��4�ũ$���<�$���5$���_3�K��ũ$�e�|#R@r�6��f�m�w=՚����;�{�Aq�k�Q�$����J��P�`�d�&$�-I�{/��%���Ԓ^{v�x���L���}f����`�ݹ�1m�1f����t][e�
��w�ߧ9e����.����٭�o�
�(P�A�����;��m��.e�s�nx�X{,�2�k;/��SӜ�)�L�y����ݼ7�cp��i��Q=S�%���AۭdU�����Wv��Gh���������K��zօ۰u�t��F���ז㊚�Mv:�\Z�>-';>Ÿ��s�t&ɬ�]-uc�&�jUn�۬]]]b5��*�ka�5�1�V�تt6v=iěH��T����˜�3�2�'U1y֮�g��f�+��uаs�+s�v#�X
�����q�^��m���w
?�<N[��{g��f|��3$��O���L�w�&���>���L�"x�!�%�wr�����t����y�gغ�ۿ�����~���U�����D�,�71jI.�{f�m�c��.��(���צ�m��=���n�L���v䤦n,3f2ov����u��um�����{��s=՚��1�����ĒV��!��QƵ$��ݧ�$�߳���1x�K�>�<�$�n�� ~?����?��OI�y�N�Q嗱���!�1�ښ)f��]���v��{��{�p���S�=�$�n-I%�q|�<I/[��I%�i���P���@�LI�ԓ���t"0H���#D��TH�(�0�B	(�E�\���޾0{^,�V��3�1(�I�����{e4��仯ۚ�s���R���Ԙ�j;�J'��u�,�jx�:��o|���)�M�؇��)�z�ho(���-���A����E��x��P�*�\e��/�8ݹ��n�ttI��l)�m���<�X�`���{.�ղ[��w�L�]T�Qf�Yv���-���A��Ѧ��4���OeQ�,�����og�RN}���� 9���&E
B�K�Y� r�V��f\ҺV��2����L��i��N���ޔ�<�Σ��<Y#ɉ9���V�T�l��ލ0;�-EXH�0S�%3��O]nC�sχ�\�91�@[�6�l�v�,q�l�.��m�N���{ ������%�&ʨ�L���I�#�<��7�H�~��=V�=�z��IO�L����)}���S�9~���߫ ����6M	�Yw4�IR�V�9)�k]x��cRM���jM���)'��w��s�K�	Ș��I�x�W�g�������x}� }�N���R	ʥn��Ō��mrQk��XY�;<9��i���7fLrْG�vX�ރ\j�\bg�m��o������/�=<���+�UҵS7r\V`�x��D)���׀zy�`{m��(��d�:�!=E�ڥ�kU�`�~��:[?/{�J�zύ��s@�ӊ,_���J,m�`~��/�BU���V���o����/m>���_fĚXԘ�I4�z�� ��\����7��x��� �l�͆�!Р�*�) # K)�$a��!XB��!	!�#!�Z:a��@�	�Ƌ�����%&��~� ����k�0BD���1�2�)Ȝ�!�`��*��@HVZFDDeD$͢��@f�Z%։
�I����	��ijMTtL���romw��Ҭ��YuB�PD�vBb�)�)`��q�o�w�������u]O+V��<��� �yY���eKq�+�������2-.�諪�ЅY��;�drVv�̹��Jө��vd��WK�U!l�R�T��-]Z�=)q �ʬE�5;sk�628̩�; �Hܰ��[[6�M�ܣְWB\��Ut���l�m�C �5��ʶ�Qj��;N�S*�:�!�[��W���~U�V�Ƴ�\�@m`�=�4�w]��r�����`�om7mεq�$y���V��ֶPU{��rbM���$.���s�1 ��m��oO^6��m$��W2E���u��n�8[�u�1��p���֢�:$�H�g*i�Fv,L�� 7:�k4^��n�O�Iw�jZ&��L5�;BMmv��K�+R�T���*�V��5��]��Y��W  [h�B��7ɬO���N8:؈�mZI�l�^Yf
�
������{T�[)��.�ȷ5=.� RG<���S��5��b�R2Li�Wm��j]��ewWJm�:6��A65|�}D��v�JNa�6�'T�*��U����s� HM5���]�9&�됹�]�%r]�O4�]�s�u[;����о4����r�慓=a`n��'b���[��\]��6v_�絮\Υ�c�l�\<Nnq��u��N�y۔�T��h%:�j�[ ��9KCĘ��\clZi�On���j�&.�*Wlj!8���`Jܲ�Nf�;�{`����sv��f�t������\��kY��]�����Ym�7;k=d��^m��\�]��� �#��	ej�JK�F�������vNm�cW�B�V�۪K����S�����A��)���E*Ȫ�U�+3Y�b�ql�-+I�;<3����Vr�̻`�u�#�]M7\���Ƌm�P-OBL�6��k�:�Q:v�A�l�P�A�8�����Q���8��7"�b�@T�(�sֵu:�E.Tl+u�� ���d��{��w{������ފ�_��-�D�h��M�C��qR��Q �D����{���O��u,�Ԝ�g�x��š���)-��<��$���mm6�`��ƙܜ�sqs�۵�>���&���[�u���ڲb��g�D��el��ۨe��cv�r��lS��lĠ*��h�&�����\����s�Mn�\C�i�N8莀�.N�<يWp�m����b��ϴm
����6�*���H���r�=����	��Gh������www{��{����;R��3-H@��6��Xyƍv�����[h���8��sO�G�{��S��7�x�!�������+4���� ����*(/�|�O",�UZ��˼�(��������}�}빿~�H��||Ґ1,�d���ϫ ��l���UϿb��׀{t�.]���.I&���)��q�=}� =�N�:J}[�X5�p�UʵS7r\V`��X(QM�_����<��h�c�,eci�)�&�h�nk;��o89�k��<�P�=���k����~�Z�"x�y1'3�9Z|����{��ʉ�G�I����nı,N���)]�6LR���9�n%�bX�c��4���
����Ȋ�� JEzAC�(���I�&�zi7ı,O{�٤�Kı/y���7�Pq,O��bcv�91�[qs��I��%�bs����Kı9��f�q,,K���gI��%�b}�{��n%�bX��m�f/�n&3f1��3I��%����w�4��bX�%���Γq,K������K��,AD�}��I��%�bw�W���pc2R�&1�I��%�b_����7ı,��{Mı,K�w^�Mı,K��i7ı�����ڳ.�c,��3�vv�m�[A�f�cVW<5��M<a�����w��/���e��)113���7ı,O��{Mı,K�w^�Mı,K��h?(�U>���%�y�O��n%����q� �eU$�Uu��!H�%��;�M&�
)bX�'y�l�n%�bX��:{Mı,K�{�Ɠp@,K��OjzfS82b��̳8��n%�bX��}�I��%�bs��i7ơ�4eXaL�"!"b'1��Mı,K���4��oq�����~���i끾�~oq�ʨ�EC9�x�t��bX�'1�߱��Kı>�u��K��AA,N��j!"�9��upٛ&)nn-���$D���SPIs=�OD�,K�﷤�Kı>�zz�7ı,O;u}!��I��&q���y��8:���a�.v�E�f�]l��n;q��������<ܙ&~�~oq�X�'���i7ı,Nw�ޓq,K��3��H	��%�b}����n%�bX��m�f/��`�l�0bc4��bX�'9�oI� %�bs����Kı>�=�i7ı,O��l�n%�bX��엳��pg�2Lc:Mı,K��O]&�X�%��9�cI���%��=�Mı,K�﷤�Kı:c�ޤ�ۊb�����n%�g�"�����i7ı,Nw��Mı,K�﷤�K��P\*FD�}���7ı,N��E�Hf���q3e��8�n%�bX�s�٤�Kİ�@�}��I�Kı;�j��Mı,K�{�Ɠq,K��Ӻ}�g2����%�%�R�[N�tx���\�1�җ;���	t����ݞ~�q=X�k�m���{��7����;�Mı,K��W�I��%�b}�w��*��bX�'��4��bX�'y�\S��38�Kq�I��%�b}����7 @,K��ﱤ�Kı>�u��Kı;��f�pı8s�������f[��c7I��%�b}�{��n%�bX�s���n%�)bX��}�I��%�b}���Mı,K���6����g�[��I��%���;�M&�X�%����4��bX�'��q,K�{�Ɠq,K���-�'�fn�3��9�Mı,K��i7ı,?�{ۿ���%�bs�~Ɠq,K���צ�q,KĊ�O�߻+U��v�.��{,K���5���H���N,�_ƃ@�@Q/g��a����]��9��2��n���:��=l#�]˳4�٨X� j���}�>�ۜ�n*��c[�r���O[��=��pd ��
7y��mۗ���w`�=n.� ��P����T�6ܻ�h9�����sq��$t��'n�w<�%�-[l]6A�n��R�E�3*7#s�������������X�fݴ�kgN����c9�cE�����r\s��չSv]y���x���|-t�`�L\d�n%�bX��]&�X�%��=�cI��%�b}���J;�bX�'{�l�n%�bX�1��[3f3���s���&�X�%��=�cI��%�b}���I��%�bw���&�X�%��{����,K����I�d�9��%�3�&�X�%��{�M&�X�%����4��`�bX�w���Mı,K�{�Ɠq,K���k�f���e��.34��bX)bw���&�X�%��{���Kı>�=�i7ıR���צ�q,K��3�`��%�3�d�4��bX�'��q,K��$�{��4�D�,K���M&�X�%��w�4��b]�7�������E3�����rLdDy$O�\tnN����g��.��t;E����}O�=LIsne������}ı,Nc��cI��%�b}���I��%�bs��� n%�bX�w���Mı,K���6n���gL�����{��7����~��M�
����(hȚ���'9�l�n%�bX��zz�7ı,O��{M��*C1��������͙�[��&�X�%�����&�X�%��s��I��bX�c��4��bX�'��4��bX�'1;%;�c38̘)�c4��bX��s��I��%�b}�{��n%�bX�w���n%�`��w�4��bX�'r�ҙ�����Y���Mı,K�s�Ɠq,K���צ�q,K��;�Mı,K�秮�q,K�鎽����6:�I ���oF8�kl��t��.���q?w��|�n�]�3��Kı>�u��Kı9��f�q,K�����7ı,O��{Mı,K��u��9�%�a��f�q,K��;�M��D�K�Ϗ�I��%�bs��Mı,K��^�M�ı9�����%�3�d�4��bX�'��O]&�X�%��9�cI��;G*��ю��+����צ�q,K��{�Mı,K�;�oaq�������L�&�X�*'�罍&�X�%��{�M&�X�%��w�4��bXb}����n%�bX����m-�.p\�[��gMı,K��^�Mı,Ky��f�q,K������n%�bX�c��4��bX�'{��y1�2�e��A�c1�w[���;n���>}`y [�p�3z�ci(������~oq��%��w�4��bX�'��q,K�����Mı,K��^�Mı,K��%;��g%�d�L�ɤ�Kı>�u=t���%�b}�{��n%�bX�w���n%�bX��}�I�������'Lv�!�&.m������n%�bX��~Ɠq,K���צ�q,�,Ns�٤�Kı>�u}t��bX�';٣ؒ�̆s��Kq�i7ı�>�u��Kı9��f�q,K������n%�`e0&C %��9�cI��%�b{�/�s���3a1&\fi7ı,Ns�٤�Kı>�u=t��bX�'��}�&�X�%��{�M&�X�%��������=�C�6��эq�Ɖxhg=#Ӥ�ۣY��7.�׵�F�x��w���~lK�d��sL��&��%�bs���t��bX�'�罍&�X�%��{�M��X�%��w�4��bX�'y���p�99t}����{��7����Ɠpı,O��zi7ı,Ns�٤�Kı>�u=t�������������6���I��ۉbX�'=�~�Mı,K��i7�A�,O��O]&�X�%��9�cI��%�b{ݖ��ٹ��fd�0b��i7ıP,Ns�٤�Kı>�u=t��bX�'�罍&�X�%��{�M&�X�%��N���n3��2`�I�d�n%�bX�w==t��bX�(��{��n%�bX�w���n%�bX��}�I��%�bh�Ϭ����*q\���ѸYr���R��ü��B��(��R����tdK�ӈӖ:��h�^�uz-��!.�U�vC`Ԅ�YNP.�z�z�8�b����9��^Y����V72���nj{e�9��&�ˆy�?���羴�8(㣪�Ovnл���`�0^л��cF3��R� �m�m���]d{f};&tn�'^Ӻp�#6�;-�����˾�֍��h���v,�k���u�N;fD�hv`�\�z�]���c7&).�ۂ�1�7I��%�bw��Mı,K��^�Mı,K��iq,K������n%�bI[�:�W5`��IUw��!I
H,O��zi7 ı;�{f�q,K��3��I��%�b^{�Γq?����b{��������si2L8�34��bX�'����&�X�%��g���q,�,K�w��n%�bX�{���o{��7�����������w��Ȗ%��'y���Mı,K���t��bX�'��4��bX�+�����Mı,K���v\��c3�3t��bX�%���7ı,��צ�q,K��}�Mı,K��O]&�X�%��wW��\ه�aLM��G���kk����ۺ���q�<ͷ[`
�-n���~oq�ı>�u��Kı;�{f�q,K��3��@��X�%�y��:M�q���������nl�/![�w�Kı;�{f�p�ޫ�:)��0Ib��B%$*i@�� =E�4�T�h��$�N(�bX����Mı,K��~Γq,K���צ�p@ı:{2Ӿ��r\fLY2Lc&�q,K������Kı/=�gI��?� �����{_��q,K��~٤�Kı8c��)��`��Ld��n%�bX��ﳤ�Kı>�u��Kı;�{f�q,K�;��z�7ı,Nw��ؒ���3��Y�g:Mı,K�w^�Mı,K��i7ı,N󺞺Mı,K��{:Mı,K�w�n1o�3�
���;9Lѳ��^1��V78��X�{7k�U;D������t�~Q$���c3I��%�bs���&�X�%��wS�I��%�b_��gBn%�bX�{���n%�bX�����i3�یg4�.2i7ı,N󺞺Mı,K��{:Mı,K�w^�Mı,K��i7�$1,Ow���sc��������n%�bX����:Mı,K�w^�Mı�p �O�t:��6)�f�i �;�*G�����S@�1`�&$ܦu�������@��y��a���
Z?_����|����eB�@�>ƌ1��(M �!!�`��d3$0`L�HB@��% Q��D�XhR?oDt�Q�  ��F0L$�@��$m4�h�ʀl�M���h�:D>�Pz�zT E:lE4
>dK��i7ı,Osھ�M�q���������ik�E_{�"X�%����M&�X�%��{�4��bX�';�c�I��%�b^{�Γ��#�#�#�_�K[_���4�7�%�bw���&�X�%���X��n%�bX��ﳤ�Kı>�u��Kı;�C�=��1#s�f�7��Ő6[\�VKY�w]��M��S<s�K��s�nS�Zc9��Is&)2\c&�q,K��{�z�7ı,K�w��n%�bX�{���~@�D�K��~٤�Kı:c��c�3e%0�777I��%�b^{�Γq,K���צ�q,K��}�Mı,K��q,KG��u0 �idD�I����#�!,O��zi7ı,N��٤�Kʄq=���Ɠq,KĽ����n%�bX����$��.$�&c�Mı,B��=�Mı,K��o���Kı/=�gI��%��Ă�Y�ν4��bX�'q���)����g82[��Mı,K��o���KİK����n%�bX�{���n%�bX�ｳI��%�b~S����d�y��ێ�6�n� e�G���nmc�/GX�n7d���p��s�y,@��'�w�,KĽ����n%�bX�s���n%�bX�ｳC��%�bs����ߛ�oq���~�?w���^���v��Mı,K�{^�Mı,K���i7ı,Ns���Mı,K��r�)!I
HO�3�SŖU�T�����Kı9�{f�q,K��;���K �,K����n%�bX�s���n%�bX���/o��s%Ė�%�2i7ĳ�\D�u���n%�bX����:Mı,K�{^�Mı,K���i7ı,N���c�ť�XLd��n%�bX��ﳤ�Kİ�����I�Kı9���Mı,K��O]&�X�%���v~�?g9&-�EZyU���:W��f��;�I��܎9�=t�@J�s�j�`z�(\n�����ΐі�)j��|���jrC��ї۩ф2�i�<Y�>mt�ya�5�K�uVҼ�㶽.���Nր�dx�9���ys��<d�;qAJ��ܷ!�q��y
y �ъx�K��=q�i�u��Kk�F�tl��c^�4�(=�{��{��s�w�{b['-Wg<{k����Z��睗r���f�Ɏ^�g�#��ˮ��Aպ;]����ı,K��k�4��bX�'=�l�n%�bX��zz�7ı,K����n%�bX����$����2L7��n%�bX����I�	bX�'9���Mı,K���t��bX�'���4���bX��{�|d�3�s����.2i7ı,Ns==t��bX�%�}��7����LD�k��n%�bX�����&�X�%��v���c2�\b�3t��bX�%�}��7ı,O��zi7ı,N{�٤�K���O]&�X�%��v{rb��q3�.e��1��7ı,O��zi7ı,W���i7ı,Ns==t��bX�%�}��7ı,N��-�J�PֆI�D݄�F�����>�{E�ꎩyo'4��b��E���<�o�ߑ,K���Mı,K��q,KĽ��� ��bX�'��4��bX�'Of[;q���LRd�1�I��%�bw����n���D۔�Wh���%�}����7ı,O~��4��bX�'}�l�n%�bX�1����9��,̷�n%�bX������Kı>�u��K�,N��٤�Kı9��oI��%�bs��=�fRd��&If3��7Ĳ����SPI�}�A$O��ܦ���y�{:Mı,K�<x�n6g�0���n%�bX�ｳI��%�bs��ޓq,Kļ｝&�X�%����M&�X�%��ƛa�6܍�뭜s3�7Q����n����iK�>�������F���~C��9���}ı,N������bX�%�;��7ı,O��zhWq,K�����&�X�%��v�fm�qs�fS�b�:Mı,K��t��bX�'��4��bX�'���i7ı,Nw���n(X�%��z{rC78��%̴��s�&�X�%��{�4��bX�'���i7�b��* Uв%��g��4��bX�%���t��bX�#��Mr��	�EUZ�_��$) �}�Mı,K�g��4��bX�%�}��7ı �;�{f�q,K��'�glǌb\I�L�ɤ�Kı=����7ı,K�w��n%�bX�罳I��%�b}�{f�q.��ow�������h6e��5��k*�c�3כd���p�=Hj�[�ם˜�y�)s�f���7ı,K�w��n%�bX�罳I��%�b}�{f��W蘉bX���O�I��%�bwޚ?bf��a2K.3�&�X�%��{�4��
X�%��=�Mı,K��q,Kļ｝&�X�%��<`�ۋ��&fq�I��%�bs���&�X�%��秮�q,ARı/;�gI��%�b{���&�X�����۱�s=8n�����K�=����n%�bX������Kı>�u��K��U."w���&�X�%��N�lű�2L�\b\�Mı,K���t��bX����4��bX�'{�l�n%�bX�s==t��bX�'N���$�s&�4�7 K]�q��Xm���v��b,�71���Md�N�w{����izT��c��bX�'��4��bX�';�l�n%�bX�w==t��D�KĽ����n%�bX��zK�LLC�.pLc��n%�bX�ｳI�~@�&"b%��g���Kı/}��t��bX�'��4���"�"b%��Oĳ����\I�L�ɤ�Kı9�x��&�X�%�y�{:Mı,K���4��bX�';�l�n%�bX����&0c�%3��&q��K�[��t��bX�'��i7ı,Nw�٤�K��E�Ng�����Kı=�O�f��a2K.3�&�X�%��{�Mı,K��~��}ı,Nc�����Kı/9�gI��%�bt2�i���}Ij��Mq<����$ �2�FGm�.��`�75��q���L�Vևb��)y�8��fxvْ��w��}:�=���hK� �1�i)+!���]W�b%6�x�
H���v�UՎ�3n�[���J����7�8��2IMķ�%��r�6��;t����s�i���F�i��8��e9��9+e!l���g��s���8{k�jk�/�wq��=����{���ߟ{�%�l��.� �!]���=k��^��u'l�%ݺ� �_�ww�:�7�-��I��M&�X�%��w��&�X�%�y��gI��%�b^s�Γq,K�罯M&�X�%��9�[�IL\ٜL�l�ɤ�Kı/;=��7lKļ罝&�X�%��{^�Mı,K���i7lK��{=�H�$̦1%�9Γq,Kļ罝&�X�%��{^�Mı,K��i7ı,K��{:Mı,K�������$�2�\�9�n%�`�bs�צ�q,K����Mı,K������K�� $1���gI��%�bs�����1?9͗8&1��i7ı,O{�٤�Kı9��{:Mı,K���t��bX�'=�zi7HRB��>>�U��pvQJժ�����1؁��Y.�n���%�<Xz�*�#x�w���ٸ�L[&f.2i7ı,Nc��Γq,Kľ�}�&�X�%��{^�ʉ�&"X�'����I��%�bt�o�������
L���:Mı,K���t���v�L��T�"X�'}�zi7ı,Ns�٤�Kı9��{:M�Kı=��XI��C9��..s�&�X�%��{^�Mı,K���i7��1;�_߳��Kı/�~��&�X�%���1f�s��2L��34��bY�Q���߿|i7ı,N�����7ı,K�w��n%�`~D��'~���x��{���?��춌$i��7}���bX�'1��gI��%�a�P�=�߳��%�bX�����&�X�%��w�4��bX�'9�[�[�s��b��e-u[��wc-���H�{g�qE�s���5�uu˴_x��Έ2[)�Km�s��Kı/}�gI��%�bs���&�X�%���^�Mı,K������Kı;�Ol����q��I��9�n%�bX����I���bX��u��Kı9��{:Mı,K��{:M�lK��ݒ��+��9���1��Mı,K��4��bX�%�g��&�X���HE��F@l�P�h���N� 1�'�.~��:Mı,K߻�Mı,�$/Q�3�\��h*B�n̅�
HS�/;;��7ı,K����n%�bX�{���n%�bX�{���n%�bX�1���`�Ŧi�S1�i7ı,K����n%�bX����M&�X�%����M&�X�%��tﱤ�x��{����������Ft��(���ٻ�6<�;+��i'N��V�u��}����	3s�g0�%�1��7ı,O��zi7ı,O��zi7ı,N�}��'�1ı/;���n%�bX��~?��昦1�e�1���Kı>�u��?1,OcǿcI��%�b^w߳��Kı>����Oܞ�{���?�����ã.�����%�bX�Ǐ~Ɠq,KĿs�Γq,lK�{�4��bX�'��4��bX�';�퐰�a�m3a)��I��%�-�~�}�&�X�%����Mı,K�w^�Mı,�!"9��� �b*���ȝ�M{Mı,K����L�3f1�i3��:Mı,K�{�4��bX��*�;���O�X�%�}����7ı,K�;��7ı,O����ߗ<����Y�G&r�S��\�{u��p�s�@�{a�O�����)��F��c&�q,K���צ�q,Kļ�����Kı/�ﳠ�Kı9�k�I��%�b}��-�ǋILɒ\�i7ı,K��{:M�[ı/�ﳤ�Kı9�k�I��%�b}���I���1S,K�;?~�s��2��6c9�n%�bX�����7ı,O��zi7����צ�q,Kļ�ﳤ�Kı;�w鶥���C���~oq�����~�^�Mı,K�w^�Mı,K�Γq,K�/��gI��%�bsǏ�͙��1�e�1���Kı=���I��%�bs��t��bX�%���t��bX�'���4��bX�'����@�P�����-	Fr�Il�,�˥����]hNSD$!	c!$!#$���E�c	�E�1�!�Z���	���AA�!�SD�H4����÷��A$C9�ReXzOw�ӫ�����C���{K���rB������B X.W�\+q�'	 Pfε�i6�m1Ė�&u�ă;��W �,v�ٴK��l֦�RL� ���`n��j�F<&֕��/J+�E@�g���.z��!����ܖ��(�k�13�y�cs[�=,P�퍶J2N�������v́���*�MR��6���Fz�]6�f�vt�@r�*��c�;���{v�Q[y8�lqs��s�6WgcG�;P�Xt�6�!�XgZ�\e|�J�8�eA�:�B%��!���Y{�]ӵ�dW[v��� �=u��Mv��o6�z�$�`�n<ܒ7 :vƃF����TQRd�v���Uyղ���L�*ԓ;�UM�h�(-�S;A�R����W\��2ԅ+��X�1W�t�n@h��s��'r����R�]T�n.̫*ҭ�L�8;D˸!nhKc�)�Z��T�I�ܼ�z���$5R�5g���:&*ͼ��g��6�ej�k�ݖF"����v嚘�e�ldn�3���Wm��r� ^���Ͱ l�ޒX��H�tX�2�qR܇"�s�m�{�kg�q�v�I͠جlm��q����r�Ɣ!�ܘz��ݼv�.�0Wuz����vڍI��bu��E��6Ჯ��K�cV���0"�9бئ�	Yl��@�<!�\L���;[�
�űۡW�A�tr��}I��6�Ux"��V�9k��N50!�����vM)��B�U��
�����5s�zBj�r��6z��۱/g;]%k��!�u)�l���q��ݎ	�h��OXA���m�d�ܓ�7`�%d�S�+����	�T���"����e쥲�Yyk��]�i2sM��2�4vn6\�$dw+;c0@��
lw�=�ݎ����u!���ʴbTR�8���9�\mb��<�˕6MGXì�.˴Yv��n��u\Is9u���%�]������LrC)��ʻ�`�8k8��9�ʆ" �@6)��U	�T�T �AG��� :��G(1��pA��Uz�c�ݿ�`��f9�����B���S2<k��͵ڬ����؃g�6�s���/T%����*t1��[���6rVݍO%��^I�T�U�S3��c�غ7��ͺ1���7:���)�Ϫ�{U�"r����H��$��D���z�Ӣ��(��L�sӬ�FFknj���r�6��0g�zn{<�F{@7F�e��kt�&���d5Lܰ���{ߞ�Oww���}|{<����i�q�vr�$n9Xx�����P�ɱu�F.�k~�}b;[8�Ɍ���}ı,O���gI��%�b^��Γq,K���צ�q,K���צ�q,K��{=�[1sIl�l���Mı,K���t��bX�'=�zi7ı,O��zi7ı,Nc��Γq?.*b%��ߧ��d��&q1�6�9Γq,K�����4��bX�'���4��bX�'1��gI��%�b^��Γq,K��ݒ�ǜ�ˌ�s4��bX�'���4��bX�'1��gI��%�b^��Γq,K�罯M&�X�%��'$��-��1d�.s4��bX�'1��gI��%�a�#�{߳��%�bX���_��q,K���צ�q,K������c���t��<�z��dN3���G>F�
^����Q�gK�s�hØ�
.s�&�X�%�{��:Mı,K���4��bX�'��4�A�D�KĽ���:Mı,Kݙ��3s����L���s��Kı9�k�I�`r��Ȧ]D�,N{���n%�bX���{:Mı,K���:Mı,KǏ���d�.2L��34��bX�'��4��bX�%�g��&�X6%�~�}�&�X�%��{^�Mı,K���������X���}����{��/;=��7ı,K�;��7ı,N{���n%�bX�s���n%�bX��g��LL�JS6Kfs�&�X�%�y�{:Mı,K���4��bX�';�zi7ı,K���:Mı.������{�v#� �su��Q�kd�\��{ ���{q�m����iӔ̈́�1��7ı,O��zi7ıRB���B��$)!I�} s����6�;�D6�6�4�S�?f$�׀�� ��f ��L˦�BU���V`�7���$�Ҵ?x�T$� HB]����fdl�0p�\Cu$�4�C�C�/���{���v�Дα��J|7Jf<��5$���h�M ���@:�4���4�o8�E�~qsɗ���u�ϴ��/R�us�v���\��li�	�na?F�u���� �٠{l��U�$d�"I�Ls��h��%2ϯ ��� om��ې�	��Ɓ"I�����h���{ų@�K�,!�D`M��tD(���0�|`�n�����#��NR�� �RA��N'�	���^Τ�礹1���$Cm�ޔ�x�h�f��\g~�����Ǎ���ír8�Z�w����K��i���FJ8��l�$�BBǍ�Hh�[4޳@��Mޔ�C���&8�b�+����~�7���;��zv[����o	�"��M)&���æv\�^ w>����93!j��E��Y��'�����`�]�~S���@��~��
D�qLs��<�� �����7|`=�`��[R����ĕrl����-��UR ����ݪZ]�g�^z)N�YIv�[Y��l.X�s�������tt��V�Ș��.�x`��+uc!�x<N�k@O�J�����j"^9��8���n�I�5�
�V�z����ҼG�.^wZͶm�5�rhȥ� %۰�]N��m�uu�ٽ��a�p�s�uc5���A�9��OE�hS���=��ww�ߓ����(2��<Oc�s<��nΡ�����m�����:�I��&�p�<�Z�������f��g(��=�� ��}�%$j1���I&��t��~H�;� �Ӟ� �k���G��k�J��8��R}?��_*������wJh#�v$,F	����U�	�~�����0%
ኘ�������f��t��m��<��@�[f1�?7$��4�	lَ7n{qkn=�s�٬q#qWZSC����d���k����<��-����U�[f����֛0����n[,րE@_�0��U�S�c.�ͻ�>ݶg�K�Q߫�+$�6��E1�I��= �l�<��:�M ����1Hd�,hm�����2���7|`ݳ �ղ� �c�$�MF7��@�S@�e4=|������%�	1Ɇ �9yss�C�l���s���M��C���K�w�F��2c�m��!�[e4=|��m��ҚG��6��,x�&n������$�d;�� ��� m�oٟ������I1ōbdz����I����N�$E�!�FD`D#!$!����ńF AdP��ԍ#�`Q�(�FIP �""�Y���h�x�@�^֛�`��`�&����^q�w>ŀ}:���S=�׀n\���Nӆ�z����uz{��<��4;��Yq�6���맭�Jcu����駳_���������	�9����1��������1���A�6F��K��]��,���]`�w��L��|`�ذ�Z���!���I�`)&�}�F�`M�%0	�c�"�U���6�ڐ�/[��_zh�I8�"�	"��T*$s�k�4
�A#��$��XLm��.���1�7�	�4���ES&��n�[nL���t���Ͱ�<��ηڄ�m�p��&�y�6
��������0&�R���f,i�4D�rh�S@����/�h�l߳?bG���k�&ӄ�x0:~��l�T�;����0=����D���V��X�}������فЧ_w� }U2).�xŔf^aL{�0&�A��#L	�!L��x���!z�/*�-b�.���9v��^:¤�+u+@g�����.���\a��-lM���A��tml"�1\�Gj:�����t/[K<��K�v\�X
%��v�r�[��;� m�-�U#Z(4yk�(	��#��I�v�b�㣣���dܕڵ�g�Ƕ����F�u�K��<�eV��y#Ѹ����<��I�K�:�:���ևb�n��#��Է�6qpg&t�ՠ2oy�܅�d��)���d�+�OA��v��/�k=��l��Fgt��!��D�$İRI�ޔ�7�������y���|T͉Im��!�w��h��Z��4�)�bG�ZKc�X�#i��?u��0�1�;�	:4�5QP�Vc��	9�����-빠__Qh=|�e9cDL�cwd�4��}
`�c����/�mv��Y�$�`7�6�E�h܇7����r����|'}�
44��~�s@�����f�{�4	�"E#1U"��yE^&��S���� h���X�ĉ��S dP�"��z��|`kx�ۮ�J?Ha�y#�Z��h�SO�?%��}��z��=���K$PĠ�����f�o {Mw��"e�׀w���9#M�6�4��$�X�� �����`	v��֮�#vܵ]t\|�G�iCc�#�lE��S�%�<t=;���o���`8.~�9���x�߯ ��ퟒ��C�����O��6�d�&�^�7���w_ov, �Z� ��u3C&˺)]WUy���0&��'�=��%7�C�Ì.�0�D0�V`ho&�w�j���2D�LR��1G��e��>?	��@ a�e,r��ƃQ¨H�L���t�D6�L��J�]i\�#˜`!Yc0�$F�QpL�y%�D�4,�$�I$`E�b�) X�V��`@R$�b��q3	�R�KCH@6ˀ~bX����B���bHB��hSV��D�hB�E��:J}&H�Q!��h�At`;ʮ:*��\�0"�0� @"�6�8 m0
�p ��4�EC~����/W�`�|�vɌ���)������SV`~��~����� ;�~� ��h[)�_]��bpK	�$�� n�w�~P�Ko��=�|`��}����?��?��0\7q̅�Fs��m����9{�����n�^ӛ\��K����ȀX����M�e4-��ݝf�ﴻ�d�"���M�e3�%
d|� 6�^ 7��=D�D!�H�o܆�o]� ���@-�4-��;BĮX$�4��`�L`$��drHI�"	j�J���tjI��N�nvLY@8�&�{m���h��h�u����\"k��ڍ<B[X^x��F�{j6��L��;�.�'Z�|������'�@��Mηs@=��}�h.v]m�"i�"Kp�7di�o1�}�c�2���Q+�߁�K�N$�� �_��ym���0;�4�7z"ꪖ`��������I�`v�i�䒪�O��{�������nI�yl���Ѧ�t���
_%�{��<��-�΅�\ �p�8S��;������Q��v�0���̭����[VKe;{y�q���@��I.ª=��Y ��yV�6��{�l.^� {&M��ٍV���+;6B7c��]%�W9xt�z�s�ݎt�<��J�;m�	��]�X��l�M�5������#ţ/�{�Ԩޭ�w�ӈ��(��L���e�F�׳���]���퐼�4=dRN�����7?绷w������<.Y It�=��`�<wgA�e�����a�ɱ��m�خ��Ҋ�f ��, ��� >z�}!��� �9��/�$��d�h�u���4-��;��h�ԫHu�����>�1����F�r�4��M~2&,h��ɡ�/~�~4���L�]-�wt�Qth�)b�L�FD�ym����4���<�S@-���SMJI'�7G��K�˵hZ�;v(���&�Kц.y��omp�X6D�I��x�4��4-����~����a$R'�#c�@;�w:�}2,K�B�A�O�j<��Ԓ�W�IP��0>ލ0�&h�j�LqIC�XH��=�S@�����h��h^�K�!��5U2UMف����9k����x��h�ĖV�Ȇ�� ә�r�%�����2ލ0>�S�q	�+���y��r��ݼ�� �h{5=Y[�G]���f{q�mۛ��`�d�ɐ`n�i���K`j��N�A�DLNM�e4z�h�-z�h.[�&,��Ʉ����0�&3�{�^�cd�0m���� l��'3@��k��cd�0$�������yW�T��wX �w�r�����;��`����<� �mI�? Ѷ���v��`6���o%㌼��fۮ����FaT���`l��4�;���-�h^�K�!�H6�&܆�m��r�l���2��*�fD4<Y�� ��f�w���e4�`mUR�e�T��f,�`�cd�07di��������y#�|$/Ѣ� B��`�B � 28-a �P!R1J,�"��
#	KmjJ�7�M�x��}��O��E�N'&����`�n�^��:DB���;����!�8�U�nbt��`�8�{��\丄���{v:u���$r��I>ŀ����w���0��D�p FD����l��٠l�΍9�Ut*�WB���������4�;���푂R"D�D`�@��M�z�h�z���@���C�n1bm�0'ti�j�1�+d�l�0)/)��dB)F�g{gg)�K:MU�Zҵ8
iF���[s&r4ղ��S[VQ�u�@���1�a-�q����ź����8�.�H5��Y@2��A�s�v�a��c�jG���m�۷N�M �l�75vj����
��:𱽕�:���v�L��*�#�Y-��T�/p�������L�lʈ����6oDv{5��as�M�=�r۠@�ι�T�-��w�k���ywI��،�ۛ=�X�b�]{A���Z'�غ�i�F$0X�ɑ@R�^�@��K`ṽw��j��-
�R��31��l������u�b���(������>��0S�0>��l�R4P���aqsV`t$�)��� 5s��>�z������"I�`��r�t�ղ[�dod�Ox��p�ږ��'�+��v�"�; 1n�v΋��WGX�;n95Ӗ۹kq�ܛY��z[�2��0]���%&)i�b"�=�e7?�?��˺c��-��Ȭ���w�m$!�h�Қ��f���נyl��޲�Ĭ����R��f��l���L�w��j������,��2I4��-��;ޔ�[��J!F�e.&�wrL\���#K�0�j�mk�0�Hlj�C�k�C�6�������bQcr? ��Ɓ�)���h+��e�tnaR	di�@�zS@;;��<W��<�S@;�E����	�4����{���6���A�% *&"��9�*���%L�ė��u4�)�{�]���/��,�M��S����=�|`�l�[�����H4�����-��>��~< �o�@�^�@�g*�'�1�����drW[nլFSk�:g��i�pÉW��a�y�#��7���!�w�)���h+��[)�{�(�VM�E��� 5n��ߢ!B��g��`���0�m��B�����(����pU�$�=V��-��<����4�ն�R%�X�@��M�릤��9��M*�-�!*%k��H�b���"�9��RNg�n��@�)�4�{�w4����mz�e4�\��j6��7+���5s[m��ng���wq��zt%��߾��s�5��&�)�9�,d�Lp�s< ��x����L���Lޔ�`�1QK(WAK31��N���L���L�u���K	�����@��M�׋�&F���=;�X�Bm��%U�4L�Uف�"w_|�����٠yl��y�,,�DІ��Nf�r��6I���0;�i�k�Hg�$!$���U��!L� ��ʡ Ġ;�*��b��l$"�N�32Fl��-Â�[�T)#�]cY����S��6I�H�#���1���� �p=��1Ѥ L+�&�H8��VL�!qA�0h9Ȑ$�-!�v�v_���|��	Ά�~��g$����܆�<T��>���k�83�$B$a�Y0��"XF�����%6��k玊�h��_�	 �0�B0�;!�;��N,�mѼi>R"� c4�,_���19(�=�,I]SLF{3���c�Zc�gs��,��'t�;��y{�������	  ���{;9.�D�G��Q�pG�O/E��TI�m��Ƈ�ղ�c ʭ�0��%��i�����$���iZ����l�m�[@l�׶iURm���f��� 9\��j�47h���nsT�;u�)ni˷KN;a�/T�S6�ۡ�D�l�e��0id�\Lv�rUT�Q�@�Ā�R�T��UW;��r��k�5�򱆮�t�nG�rd�{mۜ�na�'gl.[��m:�&���q�d�a尲g�h� ��mЫ�]������3`Н��d�5;\禗��ڭӞ.2XCc����t�>��)�>�!1�m$��_'L�ۛ�N�l�����L��u�]��M��Vj�[%$�b��L�:{)� ٪{�l�nYڡZU����j�ݥ��K���
� ��mSj�ڦG3��
���h�iZ���8�v:��Kt�5A�Ք���r�ݜ�i96*�o�-�6*�MhJ�WsOG;�U����(ZId4��pItں,{��v�r˳��88��V 9Vt^�Z��u*�KP�ޭm�4v�6�K��E�r��\t��6��m����lnz$�p�ۄr�ܚ@FKO�y�pv�ļ�λz����r��Z�ѭu<�(�iyx�p�zF�7n�`�.�����ڭr�^�f�Z�{4��(�X:�L�];ڶ�zN������:��A6���x�ҞˬtPZ��]'d��t�V�En��
�x�R[@����UI�j���Y�\櫤$:�UT�P�WbBt�*�u�[��Q�vw��u��,�ԛl�\���pɜ[r6ûg�s�gb�fh���P�D$r���[2�z�l���T�uE�[V�ҍ Kj���ˌ<],��ȓ�+mŸ�m�Y�vj�g�xU��ث[��n2i��z;E�bƍfy��F�A�^�T�Jq��� ��{Z:M�����4O)���6ؘ���ZE]ְr �d�~����;ۻ��������	���d*���׉�h9`���J�"�*���M����q�g&1-��Lbc>UD��c��W+*��vʵH������c�јؠ�-V<�ka�Bێ5�0Cqk[�6�l���;e�0tpJ� N� �k��Iy���pyH�<�l5v���r�.`�Z�X�ݝ!�\�E�a��8ң���s��{f��+ֱj��6xض�Q�p��ս%�<5�V��+ny� oL�ڸ+�;	A�gU�oe�PT"�(=�������o��������jx��:2,��e۳��0r��xx��fI�ϲ�Γ$Li�bŊ~�$�-�@��8��:_H������u����͉6��@�ڴz�h�l�z٠y�-����I`'�� �n���F�� �u�{kZ	�j���Yv���P��O�����6L�d�07���[Ak(WH)e�0�1��d&A�r�1�;������n֍�y^�!�ҏ8�`������:{E�ٹ���]���-�W��1�HWx��`�f j��>�;ﾚ���aC�"bB��m�{�]����/$`R��0	�cd�h�p�n�Q�a0R��� �L`l�I�`r�)r*��<X��̎M �l�=�S@�e4�����V��$����I�{lf�&�8����ͻ�9v�d~�@6Fx5�"����z�p��8�HKt�3���xڏnW�6�����6���`N�u�m�D/�<��uw�0X7�1BFә�x�:� ������`ot-]U�UZ�R.�f[ �wdK�#�P^��/|���^�sZ`mj�l	$fe�eUP+R��B��7�`���>�Z�@;���/��y�4l�0>�]-�l�wd��Ŗ�$���Nb�Ϯ؈6zA��0�����q��Fw/;�vs��ƌ����~W.��'I���	� ��җ;�,��O��H���~�٘���@��>4gW�v*���DQ��"5��Қ�S@�vuzm�@�;:���̉H�Ɠ��m��<]�-�I&0�%�	/I/W��#L���FLP��!�z�:� �٠y��h�M�rM<TQ4���:*1%g/BB���/�~� ���L�d�W\=��n��n���?�m����}��u��-������/[�F��c���&��[��[e4WgW��4�
R&DĄ'3@�e\�[ �&0>�`NW�J��IHh�ί@-�hu���Q=ݜ`Y)��*�V�ʔj��� �>��wu�zuk��G�r^�.N^W�kn�5��t��l��r��i�)Id���B���<�g	��u7��ң��O�v9ۑ�b⊪@�QT�:xT`�V���D�73��	���x��X�͜�ۣ�yp����t9;�/�Vq���'��u�V۴@8�=p����_6�.Ӧ��h�mb�P,OI(�h�Z��9ݩĔ���vtiZ��W��w�������FT�+;$ծ���6غ�Pӎ�`W�m��]g0-�}m�>P���U�I5�lv���I�`mr�lI1����k!#�D�,j9��S@�vuzm�@���=����LP�� ������c� ��z'����y�`���u�hu���S@�vuz�n�ف�%]�0>�`I2�]-�I&0?��w������.������ۭ�Ӌ=:X��tzE��$��w=�V���77��lV۶��d�j��wu�{h�X ���>��4y�$'����"JC@���[�rȣ��1"a\��%�⃣��푦I�`uq^�.b�85�2H���@�����_��\w�v*��	�I���`}�4�ޙ��'I��.��d�D�D�8�����?��K������x���	�#�����(�L��:�Ug���P��6ݧ��F���ٹц.y�M9��1BLnC@���h�٠ym��;����uM%��d���Eڼ�`$��F�� ��W�hڶ48�X$��<�w4���{52`G.F*Z&�'�:�G� J�)uC��ou�ډ�Z��lHBs4�)�{����l�<�j�=�p������ɉHh�]-�l�wF�� ����긂>D
�n{"���%٦�u�;:m%U��y����㌺��d�S�d����4���gK`j���!!�	2"8���n���] �:� ���7=�{5F�#8%�ǉ��d�t��L`}�4������C��8h.��= ��0>�`�<yy?/\����Ү���L�?�`�$z�hu��u��=]�^���Pi<M��Q��3�F���[t�`K��v�LoZ����q��p\k�S/o&�
$�Iɠy��h�S@�vuي��u��|�˪%L�լ�d\�[ �&0>�ʣ��I&�����dĤ4W/�@=��ηs@ܒ3��Mc��,�`$��#L�`mr�lqrUԔjI$�M���<u�`}\�[ �&0>�h���Yָ.['����Ԁ�rm�����=I�6�}����sklv6�&Ҿ��������9JJ�ۈ�n(��ڐ��C�����Ѧ�v/k���9�v�{oR=q�x�z�T���s�n�]��Ps���#�=��݈��Og�7��F�s;���*�C<��yȡ�:�z��K�9G>������K�c���+�[��.�ϩ:+��+��w����;����::{;e���2�pgF�S�zL���
�h,;M]W^��Ac���#K�ԙ�[���>�Z� <ۿ�IG�}ذ:��"��LPx'�gW�m��n�[�g(Q
&Ok鬪�%ڴL\������׀|�ŀkv�v�u�^�\X�1)�PK�������h�*����
~�DB�bCs4�S@��V�u�h���=��?յ��4��G#c���"�Jv�]E7���6G�\���.�9���83�G�p��X��v�I1�'F�$���Ԓ3�pk<�0��@:�4a Y0H+ )
 ���`ñN�SUuT��wD�H��#�@����/YM>�K��h�女s���-�D,pK��Sϳ���N =n��x���x!&�L���__U��Y�^빠yz�hN�+h��M5��U�ٞ^z8;GQ�.LXĜ&V��-��s������z���,1����@��s@����/�ՠwu�dx��0j	`U�0'ti����m�L��?���&�,,�ꉒJ�X��,m�L�'�R����V�#�� ��LK�*:`̇C�m�!c�&����hYXE),9��"�R�Y0BHH$,s�L@�k5r��S
 o�Ɇi�waQ0a(���
��z�T�eHC(?G"(�8����&�<@: `&���gRN�����cx���dcs4�p}����`r��}ϾX�I2��X�A�"�;��/u��<�ڴWQ�����)$I��0����%S�(��as�\Xⱅ6�۬�$�pN7 �q94�w4;���M�����߯ ��w�T�eT̪�eUM��>�x�򉓶�� <�^ �n��X�,jL1A������ �u���7ذ7ذ{\��Uj�^�B��L��	�`}�a��I�AE*3��5$��ȞcSY�'�{���g����;{�`mk�ez[����-Q�gi^H�m���Gk�=f�݌��z��2�W��a?<i��O�B6$!�hw]��n��)�^�M��$��(��]V���g�Jd����9�� ���x��qe��/�K0S8���V��Հ=�f�!B���ŀv�b�<��G:�$�
9�@�Қ�Ѧ�`}[%�"��C/(��W�R�����Ѧ�`}[%�'tf��X,M��vv���e͹͸�>��W��;p�snM�
k���%ò�u+V��$c���rn.��G��e�Nǂ��Bd�g�M�y���땫��S���9]ڮ�l�����6��r�rդ�gT5�7Hק��,�Y��5��͇Wa�I��/^���ݞ[� j�:0�e�SF�f���hŷZ��]zoP�ϖ�;fh����Jt����w����׾^.x8X�*�'���u��E�Ӭ�'u��N"������;�u���Qnݞ��1A��zu���z��s@�z�h��5���d��k䆁�^��ti��Ѧ����u��^*��U^[�����L���)�_xR�E���ٙ��w� �}� �v��׋ ��ܕIc��s4:�h��h�]��n��ج��
8D5��<Arf1����[)�;*�����2ONv�׭���+Qj�XY��F��`l�(��Cϯ�T��詫ݩ����MI>�;�[j���Ej�S�ix�d����0;�i���J�L���D�D���n��YM����빠Z큍H7�b�����$�/Å{�ߌ���X�^,ͼX��z��Ƀ����]��빠u���Қ�cW��1�V��E)m��Z�=���ܱ�o%N�p��fg��M�8����d�����N�0>��0:ti�7��aUT)lHCs4�)���?g�H���^}� �vٜ�Jd�]rU)]uv\��Mـy�� ׯ�D$���"D�a$aBB�HI#	!�� ����E�b!$�B��]u�`��}�$ɴK%)WHWWf(���,����49�Z��X��	?Loj$�hn�0��0����׋ �&�;�Hp�dgm=�5�{:�м��=���`��+�N7J��j8��O�m#�ݯPo����<��h^���Қ�׭ҹ�-Uڵ4U�ـ}��s�DBS'��������P�d�����]Z�TT���� �wb�>�x�ݶ`muZ���i��I3C�������I;���RM��ԝ��"��iN�aYL*#��8�I;�"��I	����)�yϪ�-�s@��h��l�Q���ى묧cc�#��H�k��p�<���v-ܼ��yݱ4cx���XLjC@�U�ym��<wJhsB�B��x�<?L̦�F�wF�ݐ`}�ҘQ�]Bx�$�m��<�Ҙt%3�O� ��ŀo�˜���Z�2��Uf&�du���#L?{������3@�}����px�ɍ�9�� �ϻ����`ݶ`$��$ � ��%�ni���H��bɛ�۳���F����a�ڭ����ђ]-R��q\`zv�m��{Q�,�l�	���ez��r�)e瀠8���UN���C��	��R�9�`ڷ�}��VYaҮ�@��q�/[�mʬV%X�oX�v��s�v����e�&!��Y0��t�JڒJKz�t�x�&u�Wm'Q���F�k ��M��J=]q�����t?m�br�r�m1i���������iP벯����B]�*4爻6e}7]�'eX��?~ŀ{��`ݶ"!}!���9��?7D�&�Rf��w7�߳�G[>4y���<�w4�)HbI'LX���`ovA��ܔ���i��Ѧ��Dcx���XLjC@��j�<��07{ ����)uQj�Z=�yL�F���`v�A��ܔ����_���B��I{j�9�u�����.�[m3�	u���li�;�4s�س*�w���0&�A����ۇSSq�$�D�4��7����I+&vA��F�{ �{�$�Q��|����MO�$r�gƁ�빠_zS@�zS@�z���D��Xcn�� ���}������_��dyI6����Қ{�������(��9�_5%�\�308��Z8���3���n��n��t=��������o�w�����0�8���~���0&ܔ��z5��	&,�vP���rHE�Ƥ4]��{ۚwV�od�y*�z����+T�Ђ�.��{�ѩ'y������X
8����}v��^�b���<I��� {���f �M��B���߼�����kqa�$�D���e4興]��?��ŀ=�f }�0M r���Ygd�m�m̵�s�S4�;�$�{<]���dv�l�:k󉘟I&ܔ��di�;���0;���Ƀ��ԋ@�����ؑ��nh��?Ss��!L��ՖU���UL�u�����w�	�%0>ލ0:�Kb@�i�JC@�ޔ�=��ԓ|�tjO"���"8�P��'�@���c���4Ϫ�&��m�L	ݐ`mw��,ʺ�x�89qWV�Z��*ت	�vx�����^x�:����f<YŠym�����7v������p)ّO��	<m����w�ՠy�)�^}V�����<�u���
D�(ԋ@�vA�:�S��L	�%0$�w{  �E�$r��h�]���L�do�Th1b)
�2��`M�)���u��T������&x�A0� ZM�7��*�Ҏ�tE�7�(a� �hgD`MZZMP�L`:,!�ST1��,�%�)"�����L\§�$c%Ns��X��.8pεIi6Ԅ�m�ɒ���+YJI�1�1L	4�xP��E	bFL��5ΐ�jJ��,���"d�cW�J+^��gw�s�'���8� 6�u�hM����r��x�yP�:W�k6�^yN�vjh��ZT+r�U��Z)w7i}�=V�������M��o0�5]�f 9*�UUP_�>$���R����S��=����T^�1��۳��.��.ru�:&�ۮ9Z[��b��M���~21�rV�m-�J��+َ  Yˀf�Z�#^Y�FֵT�9��v�N�4sA�^�gre�s�e�5�p��˖��{�Nym��vxs��qm�%;
�]mO`G�Y�VB�vNk�S^��t�=c�O6燞�j���ku�)���-�,[ɻ�{�n['^�:��z�˻��q�Wm�̯ck	5��I�.���'^���l )�9i�pr�P��]��+`�_�|���}[lB�ь����R�.�d��T�J�Ny3�(�ʮ�ig\A���][El+`�fA��V���d�(ݣq;���K�m��m�xӖ�	e���q��֪tC��ӈ�R��ny�n��N�(oDl �qS����ծj��qE�W�@8�3W#l<��UJ����ݥZ���T�L` ���Ӧ�u�#]'D�N+v��qV�1d��ې��X�h۰�968A�^-�9��C%��Ut5�f{n��^cF��&�P�#��u�3˳x�C k��`�ch{Sʁs��ң%s�������R�R��+T�w�OPu��;0��O<��u�๲�:'En'`�v���w֛\S9n;V�rʺ�9�:0n��1��R�=f�uE�ss�t�m��m�}{l<���Ss���^^�{M����s���lF"Yc�FU7l��!"�)ݵ�AW Jl�M ����4�6��p����u���e��V�����]UAղU�ҝ£�g�Zl\��]�TY^�=kHs���v�x*]�����R�Uf۵$�ʺBV\csm�r.3�C 70`�z捳ۥ[�d��،�jZ��
�f5��2H�I�ְv[��9�s����3���~:�m3�E'D�L*�ЛTu� ~\�>�"i��y_��g�#Y�$trI:5��66��u��1��Y���ݵ�Y�|�,c�|����&�����;�d㮄�ɵ���R�fy'�f�Z�ob�9�����d�����na�i ��A� � wX����`6��8�.�8���慜�[R�n��w7,=�ks�5��)6IJ�k��-u�v��5�\kE#s�������7~�xe�\��fU���:q�8\�����n�P<[�o %ƻ�OX�J2L�_�-���/>�@�n�֊X�LX��-��`k\��ŀ?Ss��&Mtq)�d��LnC@����:�V�}v����=愎�D��L��*����Z�S@����^�"�x��nM��Z�S@��� �����Q��D��!�6��{+r�uɩ7.w�-ٵ4W9�%�Z�#���L�Nd"KjE�{�)�yzS@<�f��Қ�Um쀈��䃘�f���sٯ�(A��@"� ZV�&�G�N�������
d�b�_k1LQ�,!4~�����4��<�S@��U��F�6�b.�`�l�7vـ|ݳ�B�>��3@���f$&��!Hh�)�}&A����wdu�`���TXn��Lnu��M=��Q^Ռ�>��g���.�u��<Xdb���FLY1��e4��X��:�_H=w� �I2wId�R�*��՘�or�P�dm�u���hb�"���cƚ�U�}����f��H��
"�zO�������\�c��IX���dN�0>�`v�A��*]���H<�q�h^��<��������)�u(�x�;�#MF��η�e^w`1���F�&��WZP���A��Ʀ9������;��h{Қ��4nuIfě@�j18�0;o�0>��0>��`}�`oAKb@�i�QŠy�Jh^��>ލ0;o�0;xF �0V��T�]ݘ>�`}ذ�k�
J!*%�,Un�d��ԓ|Ŗ��YU~�j�*��t�0;o�07o��<�)�r�yD�	�$cnHH�(�X�����mǛ��x��h8����q�<���2Ex�Q9�}V�ﯪ�<�)�y��9�UE$�"KjE�{ծs�D��w����7ծpmU��$���cNE�yzS@�{ká(�{O� ݧӀ}�%]U'h�6�)e����K`v�J`n�J`};!�uΩ,z�bj1(��;��h�ҘN�0>�`r^IIDe��r�Y%�ljp6�Ц7�g���YU�6xn��nV�j{i����:9�$�Ւ��ۍ1�HSq�gr�*�J:�<0��sk\��y�.^7@X���ݴ�EX�+��\H㌇�����j��{m�jy�F!���[�������r".�^S�;u�h��[����clUKҜx˝*�'f�i!"�4�A�f�?��q��r_;f�ѭ�K�@�ԧ��<�����)7n�X��7,���nw=�f�Gq�0�8	�������N�0>�`v�J`}�#(�장rR�sws�|�ٟ�D)��݋ {O��ﯪ߿~��G��o�ǋ&$�߿4���ݹ)���Uu!\�G��ډ9�z���]�@���DDN�w� s�t�]U�2��j�e�e07nJ`}; �ݑ�od>�?��5��iNRnش�rD� �tQ]�g��:½[^l���_g�t;��\YHVLA�=X���L�07di�����L��®��b�V�2�`n��^B�A����L�dIP�O�e
�ˬ�����v�=�%U����;�ۚ�E,H�b�LI%!�}�%0>��`n�i����P�n�Y&<J8�/Jhg���������<�ڴU��g��@�crW�LI��&2u��u���(<���=�ں:S�^�KT��^]׭Z�����F���`y��/Jh�4��Ȥ@���*�0;{ �ݾ���vA���� �B��6LY#Ib�8h����e���P�b�)A�)<�2D34�T*��w�4����UM�F�c�ӑh[)�yz�h�)��/�@��D�Y�&)������Қz���e4�۱����$��������U��c��8%��O��C�f�׆�T��#t�Q��	%RL�;�S@�_U�y]��$��s�X�&�.T�����ffn�}M�tL��|`ϱ`�`wCm܂ȇ�G���M�Ѧod�%07�T�]\˯Z�*��՘
"���,�0�78O��|
�Ĕ��2f~>���-ƒ��d�)�����v�A��rS���`rٞ�Y�yx��k���;+�=��6P�����8�]p*������vvB�k�6M��`�)�7��`M�zT����c���/�)�y�]�޻��������#m��x�0XYuf��ŀ7������`;��#4$�$�4l��m��v�Q��w� ���ʔJ���&j����f�.��>�v-�)�\y�V��&��n~���vx�˖Ѵ����GJ�b�����6sm��.V��-m�˭�i8��tb����٭�:p
:�{pq�#���=���K㍸,ӷ9'3k���^��v�ڞ��X��>����5OgW��\l�oj�nua�y��-ul���Unq��۩�ZYkv����¯Cѵ�����f��7,Am���a��X^W����q�_����k۞f��c/�Q�얰8}��)��\�lsv�/;a�m��n*$L�px�����S@�n�[l�:�M�G��Nƿ<x�bI�@�F��cI�`I2�uU�R5���&h���)�[n�m��ޅM�L1��MN�0;� ���L�&0$�v��J0�1��h�)�[�s@<��޻�痷�M4
cn~q~���;�s�����}�gp'eP���r�^��b2h���x�0X0n���d ��{� ���@��(�ČkQ�I�I7��:� �WK;�wF���3�@���ׅ2�H�bRG&�'F�ݐ`}:4�>�cN�+��2A�i��;�S@��w4+�hf.����{��|�,��d����kŀt/u�O�{_b�7vـ}�;��wxMΫC�^$5�b��)�m�[>���6��������Ɠr�v�f��rS푦wd?%�t�� ��O�< ��Z�۹�wvA��#L��L�R���!]VX+�yW�����d�/yg�Z,���>�X@���]@��N�h#	�(����R�x�����"�r(fB�$ �i�P�&4$�9pBB�x���t_� uoB$a�I	R��]� =�S]��I�v� w9K2������H$bBZ� bD���,����F��MI���pjPX1�F0���\HrqG�Z�,��]���K"eii��p�q@�攂�
9�vpK5��K��%��3���2|M�A�Ī	�1�]��ԹF�E�`�!v����#���+�iG���1CU �Ard \@ Af�22��J��� �w�3��M(dbR�e�M�� `�&����k��qC{"�,e��nQ�JJP`<6�G���R R*|���i��*B���bk2�����HFc��E� 3Y��U�P2)M�jG�2�� � h �ta!�W���]`���$��Z��y)��#L	�X*��g�������������7[Ł�3�+n�hqO��bxВ�)&hT���4���d�06uEi�5�AJ%�l���G�q��ZnS��V�۠���c��8���m�]{v��K��~u�X��0kx�"#�OwV����##&����4z���z�޷s~ďxx�}BbŘ�3Oߚ`}[%�7�i�����Iu"id�ɉH���x�W�{��I9�3٩0�"_B#�(���*����jI=���3���.s.�AY��ޑ��d�4���G�}�����	��his �~���wN���.�Il���=E%���u[];�	5�j&�H8�� ��@�Қ��_��ϱ`�1ӔQh-PR(*��5�9D(��ON�V ��,��f}8���dǍ	(���^�ףL��0:vA�ӊ�F*��.Ĝr=�]��zS@�Қ��z�Bb��ऄc�ә�w�)�Y��:[N�0)#�%�^]��Aŧ�c�nJ�ûNؒZ���K��V�j��%��8��m
��Y9j�U��י�ѩ�<E.��:�0b�JBLQ͛vj��E[Q��}q�|��қN�DمM�gv��v���*��Ɣ�`�ɮ� 8�k��8���ڊ�cq�ރ�n�%�QU�l�N_�=-�6m���U�JV�fȝ��/�vX�ꖻ�ٮ��179�����C��(�q�m�sL�Lb4t�`�,�0ⵃe��dI��ۢ�$���yrZܰ��c�ȓ����d�����x�W�[�s�<Azύ�b��4�)�p�<W��-빠w�)�[Қx9;�cr�8�z�`v�A�'dV�l��t�<QJD���{�Jh����^�o]����Z�Ɂ1���p�-�M�mz��4��:�� �<�fV�N۩� S�&pd_<��w6�՞N�i��M�Ɉ��"���I(���l��0;� ��rS�Y�738ķ�3�I;��_* A-YGfdnJ`M�)���]Y��S!Hh�S@��Z�ڴ�S@�=xqSr"($4�%0&ܔ��2	ݐ`oYEOL��LNE�_]�@/[4�)�^v����?��|ܘH�I#�Pv��Kyf�޻J�r�H�h��ٓUu'[�df1�ȌQ)�}~���/;V�}v�����Cx�JdRC@�Қ�j�/�ՠ^��w*-X� �����h�*�/�զ�3��CH�]��\���ԇ��Ɓ��SP3#i	%�"�/�ՠ^����/XU�u�)CIGؒqŠ^��ٟ�}n�x��|���9z,�<������VE(��MjDz7L��[�N��Zv�����r8�!Hh�S@�rS@��M���<��΢n5	� ���:,�l�0'L�wd�K�d���LS$4��/YM�Jh�Jh��`�B�#(U���I�`N�H������(X�	HL '�{�x�>c�<��+�Y�X�/0`N�H�	� ��2�I-����x�������2Hdk�3�80��]�mZy(�|�;�v�P#��Fv{!Ug�s�|`�ـ=v�P��n�4����IF7���h�A�;�	�d�I{�D�
��a�QB6$���>���^}V�d�w+� ��� �拆M���\�t����:�StYِ`N�ްY�SQ�LX��h�Jh� ��2	�Ҙw����UGT�~l,.�\�p\�;��7���ԅ9�6y������B��Wh�����Cu��{N�^�Dng*���D����j^M��ֹ��K���j��I���!k]<i�g��F��6;&v�=<;v��h0mU#h7V�۹�<�b{s���n^��]u�$�e���6�����v��f읛t��'n�xY�:��0����ì��������w���{��w��=��sߘv0�e��]F�s�K=�\u�=�HE�.�D�6�Ca��ˌ]n�n1cRHx��M���/>�@�T��^T��(��QG��`N����ِ`N�<���"S"���h�S@��M���:�����?7���-��l�0'L�u���t��ǉ�J4�p�/�S@�e4Ϫ�:�)�~��_90Ȉ'1����_m�y����L�F��َ��x����-�n;q(8Ōj�$ԇ�}~���h�S@��M�ۄ�E#Q��f���9ۭ�`E����V*+!|:oL�[0ݳ ���]R�2bœȴmR���h�M���VS&&L5 Ԇ�6dL�u����� �P�2��[)�^}V��U)�_l���w�D�?7����2)H�P�h;�D4͸W�k�1��}���65�8u�ō�<11H����}]�h�R���hl��{�Z�j0'�&�`oJ�0&̃��0'_J`HR��dx��i��_l���j���{Փ��`l�`vʬ�0I�<��&�4m��/>�@�U��/�ՠv{p���#��4�Ҙ�F�o�07�A��^I-���߷K��G��c!���s`��';��gf����z����'J��Om��~�Ob��\��l��\�X�̢��`��4��z�h��h������x��(��Q'��YM���ڥ4�h�U���1�H�����ednJ`��Kk֭Z��z�� ����V����A���ݖ��2~raH�j��/�ՠ^����h~��|�n~�4������G7K�pF�-����,v�g�������a ��6	(�i��>���@�e4Ϫ�:�)�w�) ���lIU�� ��3�)��>��M�?Ss�\��?ENo�4Ϫ�:�)�_]�@�e4=`��WL�v�^e07�d�%0:L�e�Zv4�X��5#JC@�]�@�IC��� ���{f��?(�
B��TDU�
"*��TDUj�"��E_�DU������P� �
�P`�D
�T`�@��
�Q*�T��H*E �@D �AE*H*P`�D��B
�E`�EP��*P �@Q�� ��P�� U��  �E �AD��H*�� `�A�R� �D
�@�� �DH**�R
�X***`�E *b�D������  �A
�T��"*X*X*
�A�� *P��@B*�TH*P
�TF
�UH*@ *R
�X�
�Q��DH*
�
�T��EX* `�DU �AD`* X* �A� *�� ����2
�
�H*"�H",`�F�*b*X*
���E �A"*@��R�P��
�U��@������@X*"*U`�AQ *H* H
�T*"�*R�`�@X
�@b*F
���DX*`*H�H
�@��A`�D`*"*`�D * **��T *��
���P*���E��H""Ȁ?�QU���"������Z����DU�QU�"�����"*��(����DEW�DU~DU�b��L��8y���ó � ���fO� ��� �3րz    � ���      ���  |��%A��D�T�T (  P  
 ���T�	"
 �HRIQ@�H HRJ	"   h 
 � � �����qg{r�z��{��\�C��ۛ_F��ӭ>�z{��zz��}�Je���^m����W�.�, :;��>�������i�n%���v�� u-v��NC�`u��  � E"@ (c  �4�u8zq۶�k�B�@.� �
e�e}��ﻯ�S׼{��� �U9o���5�}<��n9ҽ������ڧ}�z��=ԫ��� (��_q���Ϲז�MW[��>�o@�J(�U@� (9 9�_qjU��iш(� �� 0PR S��
����)J8:��Pt� �@ DJP)�0= `z" PDJD  $�@ &�h,f�P"hL@&�@  � 	D   ( )�Q�4��t�is�M:p>@o)X��ӼY���T��Ҝ �N��m�> Msڕc4�}� 9���}i{�u���z^�'��y��������Z��p�{���| <�$ �T  (
 ����{���Wk�+����s� 9���ζܝ}���{<��� '*o����k� ���Η�K��@Ωb�Y}��n�����{�� n��z�qjWs�w����I56�T�  �P��T�@  O��*3�F 2=��#jR�  S�	)J� h ���ʕ	� ��|��=���u����?�����w�\�s��H(��CY삈��D UO�ADU�"�����"�@T�/�H�������)/��d�\����>��띛?\�;!IS�$��s�!\!H�$�c @���̭�Hs9��6k��C.������V(B D�BH�B	\�qcT�HD!`T��4A�AĀ�H�!ȄR@��$�"�ьH@��ЁF#X��$��H�HRB5pe!%���L#�IL#Yt�����8�m�qol��v9�]m��ۍ��}�s��|���	��.�)�,�+~;���U�ݤ$?}�R��x��=V�{�
b��j�f��Ϊ�|��s��o��:*�nz��{����*��S6I�]w��Ҙ˚%�D�ˁ.i�3L`|�7a���zNg����L)�=Ӻwu��I�'K�;r�HH�a�DJ�����\�����wy������;������&�)�VUB�)J}���xMF[υ�%�D`F,R+��.��?8[���&�D�jq�R"Q#e$ɋ܅�\���}�2܇�u#1��@da�F �"�$`�� u�RH$ ��� ����1A�"�$������w���:��%����¨޹ЅOɢ��L���d���a2FB0Ѳ4čI$��k��å����|�OƵ��A������$aF#25��ᐌH��8wd#.�HB��\�L�1Ŭ>4N��$H<�D�Y~�t����5��6��
*B���R��x:O�����ޡ%�}f�B�Đ AK ��F�/�h5�X4! j#�Č
�aD�VS~���JԁjF6�!,!q��~��.�I �$���������)Z�F�H&����! YO��53���s�E�Io�ւ���� �1$>;�R��`D���X2 H!	V-R1ȑ%�Ɯ����lLf,�ۛ�&����S�!�P��Lt�
�(!E��JA�B���#L�]�k���r|k��2M}�t�J0�0��$LHE�RY7����vW.!�Q���#]0,� au.h+�@�3pi��B�K"C[�cp E�@ �! B%��Z�	,�����0d4d%�n]:&�cBB�f@��	r8h��h��əkl���9�wF���Y�0���4Lѹ����3k��H�f�wZ��B3/�ɭ|rL��k���?c��4c�`H�$`B,c$a�`$���p�ĐHN$�����ֶ5���$B���!q�y�����	 �$ۆϡ]
� n�-p"�!p
�S�v��Ш��c�S�A*���
80�֤�2���f�gd�7�w���C?޵� �޹͜�@�=d4�!XC��XB&:�$`��o��~; �M��t&i5
��a�!L�T�"V��r77�g�=����?�ň��/�y�� M}�V5�K~ P���0�5�B�(ke�P��n�	HSd&���k\��M�_���;�����tF�� Ml*iMˤ��%vhZ.�%����������!�F;�d	8J0�h���F7&��4˩�PP��(J�zޙ�L'`6-�Q۠�`A�?!#~��s5����A���-��`o�����D�	 !P�!bX I"���� �\ ����~!����W>��N�}��]5�VW/{K�E[��E��_ ��/7ܐ"B�E�$#1(��J��i!s[:~�]��Dj1�!��@a$Z�8o��yzW����?�]m'K�]�/WU;�H��������D�GAs\���B/�A�X��Ԃ�E�0!u��ޟ�F0��5�����zCT�t�	L�
`hd�9{��!A�C�Č(f��Ð�s[c��/TwL|έ[VU��GU����~��ȱ������d!��u�l,��4��E
#���$�{��,U0�"��Mw{�5pe�	pb�7*b��$,(F�d��BF۩���b@�E���,+��a B�Nw�p���z�S�x{^���Q�E�Eu�}Ҩ���/+�
ϊ��g�m��^UKu��L���Vi���ٮ�u����"H�, �b!L�:^���5����?0�klB�
H.ЅÝ����i!�*�F�B��Wi����9s����  D$@1"�2!���l�J�jH����k�����0���ѻIm�7��t���0i��*B�����s{���?p榋�ͧ0I5,)��$�$�"I\�?|}����gu��l#9ZY
��Bi�|���}Ο��c�H�F�B��X��$#�|������^h]ȱ�	�s4��?l:˿��D/��?}�z~6�:Ν�t���I$j��bDb�B�?�˟��%�H�$K��Ow]�ݟ��y�l�~�y����F5����gcIy�����U�F�I��������}u��߻����4l8B��E�V�]���>�vp�@��>F Eb�H�6 P ����p�3�ۆٙ�Ȱ�f�.t#bR�X��B?>���+��an>�����D��w�9���!�������A��\#\��3��H�%ō��߂�L5�ƈ~ЛH]��ѽ��:~z@�/{�q���a�� @`H`R�l�h�E6���n��<7�w6l��kхaLP�ė��I
۲�j�Se���Ԇ�N��\�2*���9���0�����2�3�����E![�f�L�Ο���0�b�i���.:�G~�>I��w��p!&�����,
����I4�$��q�����i��(� @�J����3�k\��>	��Cm+Jj~��~�����F���!�����d�q��x�&�4 RHԃ`�aO��K�o9-�)�!Z�P$�"H 00���R0H1H�V?s��/�B`Wip�F��S>��)���~�s9��s��7���	�kd	$���6�,&�M����8G����S'�w�ջ7�y�B�~?s�.�$?&�B5�Xe��Q������RNZc
�*�B"�_�Ӷ=Ϸ�6ٽ���a��a����G>�WC��>�?>w�|����]VZc$"�D�@��
#�1�!++,(i�
	���ZƆXV�(VK�"	P�[��w��!FǵG�*�#���U�����$�;b�����"~���Jd!��~�o�f��)����z~>n� C����ĪŃ  WU0�,�K�.��� S�VB��
a����_h��Z���9x����|����r��UU��ο���~�0��7�4dh�%᫮p�.����p&o�w�{&��R�Bu0�~;���t!B$�rn���7���?g.���Ő���?\�M�F���kl6�8ss]�>sZ~e��R�9���r�[���%p�FA"�Q���H9�LB
����(�+:���R�k������K��7�?L֦w�Nd)���J���̻�Ϥ֧�O�"�j�?a?�"ji�qi�%P�����.�r��bI@jn$��L�R�36� E�a��:�$s���J�c�"Ej���#$��,HA��H�c�JC>4I���e����A�B<4�$i��\8쐺ޓD�]\ǡvO�Ca
aBS�0��0v�Fkp%3	r.��,�����z�"������G�!H�$H0�4B���ko�i���F�$(��
*�
0$*�F�B��!�,�J9�sz�˲�p!��10�J�!"D��f��_�$�t���u������3;K�C��n!YVN�XW����)�P��(�4oa.�&���l2�	��]���a)��c(L��Syr4���A2���t@�a��4����¤�I�IL40���`�~5�RMD�L��៲#)�m��󟸘�j� @Ͳ�L2�JB���i E�6��/x8E� 8�R��lK$h�({�W.��>
UER�;�$�H� D�m��   �� ��B@  ��;<��}��i�Ш��"z��Z-�k�R� �`]T���pD y� �W�pm���6�*��W��މW)�jwDUmU���J��iGV�i�4h�V��dU��WMX6y(-����W�7�z*[�.�۔�p15�]�,��&�dm&�E�	�DVڦ���q*�RҭT�U q�<�Pn�6p�lkX   �        m�m�  Z�-�fݱB�8��̄�U*��UT�V^V�Ή��u����}��`^�2��m[��� �ꮝ���p۲@�ۀ��am ��5�1mh�'E�k�PI�,-�p    �h�}��`���²ʪҭUP
�Vʪ�P]�瀩`(L�4�r��q�P�2�JѦ��I�-��86� 8m�� ��$�*���UU^j��Z����- -�kխ�H�cjZ�m�@KM��.���N&�'���>[R�� lp*��t
��S؛l�u[ͷ^� ��J杧����^�N��˫�8��)��m8z�겹����<�,�:S�t&�r&yܽ)��M���'��2�U����l|y~;�uN�f��lqm#Z�ΓׯX��n���mk 8�� 
P[Cm�%�ܛ��K��U/-�u�R�)�qT���Wl�@�WJɉ)����! 6� m[ �ْ�N��pn� m��eė��` <�z����iRem���U]/n؅..j�$ۚ-��$u([E��V�%:���\v�U��kh8$�I�/Yc��\u����j���M��\����-ђ	�mƮj���B���̅��2%]N��غ���s��"��m�.q5mJX���]�	#g��2۽�9�$���j�!tVC�8kn���sM#&�����=�v���N
5��v�:pIf�J���h���-i�kU�'-<�VQ�v�(ݻi^ۓ�T��K7�V��Ճly�Rwf�Í
��iz��Y��ۤ�D�e�7Kg�Wvj�b��5N��[@���9@6����� �   -��/���M&�Q����]�0	 p�����ٳl[!�@HI��m&m�H	lr�[m��%��y�[vۭ�JGm-Ba���n���  �[���p  6��� ���6m���}���m�r�] "�C���n�ƚ��yZ^�[B@ֱa�m՚M����X���h �  �sm��[m�-�m[H$m����� �`m� �À6�m����l H�� ��� � ������&ݳ��Ծ���      �  	   �� � $ 6���Ͷ� �u�;V�f��Kh�]�E�m�I��p� �	���n     [m�č�l�����2m�.M��m�p �@6�q���I/6��� ��nH � 	کUT ��մKԵ�� �d-6 p� �N��; 	 �B�n     m�  mp  9b��IM�  ��[�� �@i�  6� �m�ֳm���    ��k����-�       �> ��5�n�m�m�mh m��� ��-���If;lH<$l��۶����}���<U�m�6�     �8#e��$�   �`�� 8�[D� �� p�`�m���"��ַs�$ӵ�b&���mp$$ � ��l�    6�I m����@����gh*t[T�m%�6�0   ��     -���  ��8[@:� HѷkV������u�$�   h      -��$�ݵ�Mn*��g�H#'l pp ��N��!��l� � ջ(   -� /;j  ��;UUU��mI�)�$  �N�$:@[:Iy[m�^m���f� � m�	��� m� 6طS�ŵ�n[mf��d8  �l 6� ݮ��o9��@   5���` H'mR�R�T���`4Y4�P �p/yzHէl�gKb�    ��  �bKh܂�ekA�� 𓄍�m���:˃ �۶� �I�Ͷ�5�[A��@�V�����j�g�m&��V�  ,��d�ݖ���i�2@h 	eu�m�"��%��
Z�j��yP-62��I"iX[`����F`H�N[D�mW�E�'C[�`���i��@$�d��äe/-][·,���$�Z�  
u�^	.v�5 ׁm��!v���"��<��ӰHC�g�`zl�UZ�@{iK3h8��`68 y]�v�[T�U��89�g�)E)�Y6���
d��m�mV�K�Oj8��;|���dPm��B��Q�]��'hFJ ���e���wR��Q���T��n�g�����\Zl9G��Iߟ-��R��'m۵-�V�m�k���`8���[y�����ְޒ�lHB�iXv�R�Y0-6ӯF8]9kk��	�.�WUJ��Wm���U��幞^�Be��VU���1�W-�����ER�W*�r���� ph&�����Ci7N��$	'I.�6�:�B�mٔ�T�ǅV������Ege]�U�Ij�n�m�zAm!��	ݦ̖�l��mjO���9�lU����w.�cp0nSkY�5v�6��I�����T�n{l2s����ʳօg�n���w9tKSV�.a�A���ۧlt���M�ؖ�媺�Umm��F��ɰ�;S��I���R�*�U�d.x-�e�V��B��]�$��T���[yե�Y@�M�n�LkM�9� 8m�    I�u�6�pm���&�]d�ȑ�m��m퍷Im�l)�6%Zݪ���mR�U հ8   hlmem5[GZnE	,�{�i�7kn݀� �Y��Z��۶�xq!6��4^�P�ۢ�v��$qm�p�I���-���\�a';v�e��n�@q :�m�ف��a�ɕ9���wgP<��յ����L;�3�6�v<�B��k���*���Rt�k� �UÛ�to`�Eѱ�Q���V�e�)VI�l,
A�;5QEvq�c+�iT8��e`��mWUP��U����O��;C�]\	�7����y�մ�ҭTkQ�C����J�Y���l�   �������V�W �Ul&+��Z�4+*ZΡ!�HK-��m�$� A� 6�  6��g-��� 9m ���p -��mv�V��c�v���U��TjD� Zl 6� I�m�G5��m&�h8�N��톨gp��J�UK�9iVW'e�V��y]�zV�Ʒ l$���v��`�Ͷ�m� ����Z��UU��v�6r+Um+gpgn..M���[A 9-H���V��.�s(v�d�%�6�sj�2   �v�Ͷ ��vm�m$6�̀r�(U�C�%��ۡ���ր	ٶ<�m�F���snBJ�=V�����m��+�iۭ` m��h [F�[@-��h 
X;6��M�Ѯo��_��u��xrtuq-��+u�Z���Χbs�kX�v��r�m�Բ�%�:�x�,�W�⭪x�� [\:;m����z&K��5l�@X�ï�>s��7
o\7��J�Q���m���Җ�ݖCg �J�m�&�ն�p�����ݶ�`	 �l����      �6ۖ�'E��[[[�� @H�   �`    4u�6Z �`l �$ p��  �m� .� �IJ ����4ۭ�36������D�Qms�ba�n�h5�Q�-uQ�ѣ��בu�I�@�@m�@��m�KF�@�l�+��kMٻ` [Ro�)�S.���]*�UU@L��6ؐkZ�I�E-�1�m m����X�j�%%�ສ���)Nr�P�IKO(m��$β��l���l���J H&��vj�c�@��U����f�j��8 [@ ���@k3YM��ˡ�[@     � �*2�ҭl��P׮�*�v�Zau�V�f�c���I�	yyj��܎���� h&��S�km�m���m��۶�0  $��ur�Η$F�u��*��v��d14F�m��q�MSR��ۦ�6V
���#��I�4�@ -���R�mݰh�ׯ;Yǧ۵ �ĲU*�pohjW�Umt���հ���mR��QUU;&٬����L�s��s��[@ '@ ��m�  M�-m�@  ,gF�-��EpPb�@`# "@ t�m�� �   l�-��-�Ze���L[��ZƵ��n�8m�   ?�* *��P�0EF��THQ��U_��#�B(
:;�*�(U_ȴ7TA(� QL��EN'"�J7�Tq���Sj�?-�&"�����sH,���F)�����(;�A�A���E��@���ۀ��"N��G{p8�^����
~[�	���ɨ���H	E� 
@����h�����A~����VE��x�*?w�p�a�r ��k�6�p
~@M"
�o����C>@a�^�� >E��O�>E���b�T ~,�!�/�	�_*�E6�0�T������S��H;O�)$���,T"��7� <��� G� � `t��%A�`"T�� �b�T�����"~ ���S+���1@��`$� @P�0��U�����;V���� ~`�������򗪊��buP�҈����hOƔS�?q�DQ_�|?�,�d�Z,T$E0@mF�b%�*�$��5bĊ5�R����������8,8�iƍR�6��iL��vR�eq� �p����:�*����`��  �[%�1��>�<�λ���u�������-����i�ª�����b�Eܳ��/2�m��V9�����.&��lݱ����t���<v�,O��6��S��i5�0Z�mj���^]��e�H 8�6�B:�xx�L��O;��
ƌ��&�
�.a���Cd���kQ�����]�t*�9Q"��es��<��H��jշ���2�� B[`�g6��m��E/q�{([��˫�V����ڛj�����g��� ��9{pJQ%�w)UT����jy%��`��]��UT��+0mu�ؕZ�j�ڹ�`�� ��y�l�Zl��GKe�^��#J�UJ��]���Z��6�rmmv�iW]M+1��������2�"�M�B�I�l��m�	�<W��a��`\���T &���k/r�H㖞�Nul�"�qI�v��8���G/jnG�-0�M=!�;1�f.Қu�6��δշ8���U��)oX�"m�,�S�1WKr8�<��mg'r��̙k�����[;�b7dӤ܂����aޱ�z�Z���V��69��G��b�u%ˍ@�	����չzeUi W�L��]W�r�ܖԀ���qdrY3����Ǔ�ɮ��󸠅�\�q͍��������;����g:rHUK���0s:3!T�-Y�az�&�p[�؃�C�8�'K��(W�'�e�Y�ڶxG�ZU"Z���Q{ b� 8��B��i��\�]���	�ʫ�0�z�*�R�l&��� K"�e��:H�ɖ��ѱ��۳\���Q��sd�;9����ʹYMTe�x�l�<i7EB����]����(�q�Cn�^�%�ʄ�r6�� 6g�:L;�u�&ɳ	����1��lە���-*�eP*��^U��xY�kWZ.�,�[�kE�9�A�p���@z���T_�ت��h'G�Z'�wH~E>4��w��q���ԥV�ڪ���$f甫���p�����m���v(��ÇyZ]ڲ��w-Eё\H�����f�[�8�c��V�8�L���]�aիi]����A5n��ڞn8����q��r� �6��T�d���-�����h��V7)@�����'%��ʛp�"�KD�2ض1�ӫ� ����P�73�zxm�����w^�z�7Ǔ��p�<�˞��˅QE�N�U�\�ȣ���z�-��3@^�����]f)LI�RJM��V1�`s�uX�mՁ������Ѷ�T�29#��$�s������e�=��#e'���� �V{�u`w2i`skv1� 隝6�7�#��@w=���@{�K@w8�����w}v���}�湜T�j-��C�U��\��v�|z�F���3��eb屳]�f��LJC�w^���{���sn��&�--PT�N$n��[j�B&b	&�3?Mp�=��g4�>�MJ��y��IԌR�����m�������1�.Z���o`�R��r��&�;�R�wvXz�f��`o�Ɋ�A&�9(m����=�h����qR�� ?W���U���ד���S��cX���4.֍�V,p�r��Pv}j*�p;<9N9�M��3����� :=�����u G@��Q���{�u`wri`qw4v�ݗ�H=��:l<�UqT.r�9m=V˸ʳ�333$$PG�Q@^���;��[�~�mՁ՚-JJ���858�.昀I�� :c��wusr�on��4,��� �M@w8���1�`n1V�u�iI
$���1$e,��7&Ӻ��'�Ms�@�b��	���g$	(�R��X�mՁչ���<��;�,n�V�E �R��r����f%#���X��X�;��jcv�!�NJj8�c�n�;�|�bbb�{q`b�ڰ��@���U�������;��s���%����ƨ��Q����fnI���knw
��3 ��@w8��6<s1 w�����}_W^y�h�	ʉ� u-��P^���-�jGK������i��$9Z3J6$�r���)������9�5� �we����XY��9Q�A�+��t@y㙈�M@w8��6�O[Q�� "H݁���`w��V~�K3�Ł�{��]�blRGI�J�Gaﾯ�噾�X��,c�n�;��`r�V�rJ�9�$�r��`���3t���qR��������c���ϭ#S���続p��-��W��Sgg��n[F�Y"{:���v{�nX8�HY��^w��[�L�jm,INWbTr	ne�ʬX6��re^ف2k�hn*���'��ܹ���9��[n�iڱ2p��f%�7[�H����T� ���L򡵮L� =q�+<Z2dh(r�4$�/�ԡ�e�IBM�ܛ��K(E����|����&hc%�x�;+�ܙ6j6����i��.t�����g�!6Q���%1�>��1 wI�� ;��#���MRdC#�7`uwu��H��]X��VsG`s5PGCOaMJY���� ;�K@zۗ���,�uQUT��*�\�.r,6fffn&�������@;�1��[��HF9��!`qfjvu���q`u�`l����F�HQR��i0�6�bU��֎k��n��-�盩�	x����D�I@R8>�=�`w��,��6""f&'�M�=�Hn(�6)B�H��6��}�?��+́$�xČ�Bq&+� ��:9��N.1wu߾H�{�֣�Dピ�q�Vy�y������6����T݊�M���4Ԋ�f"&%u��U��nՁ�㸰:��7qi-e)��+w]��qR�9�s�v��&V-��/v���7<�7Ai��:9�7<0����qhT����v$��eGM�RR�h$���sn�q�@{�˴ �M@ܼ2�˔��Hԕ`unk�9ܚ��gwe����XY��J��A�%�v;�iXu�Y335�D�O#�+�㸰:�k�7]e4��5�%5"V�݈� :c���=�h��ff^�oɱJ�G`w��Vu��ɩXwvX+��eDҡ�4H�% �[�K;��K�4rӅ�B�U����<��0�u��u�ۍʰ;�5X�MJ����`w��V�je�tF�t�CMH���i^�̤5��`f=��:�:����5RA2'"V.��ͺ�;�5X�MJ��M*:hoaIJm�7w�*@u�1��A��}I}J� �;��w��$�׷&fzI����ԕ`uwu�����7����v{�u`wv��P�%M�����#�Ɏ{Y����|���Χ���Wv��<�%��	�J��Vo�`uwu��mՁ���`n��il�J!@QH������������|���f5VVc��JM�P��;�ͺ�;�4�8��;w]��ե� �#��q�H�`��� �j��H	L��6�Gӎf�`��rO߾���?w�vnI�x����������;���tŸnu��n,q]��9y���\�� @.��Fݸʡ��;&�`�%�����ϟ>V�즜��GP+���M��*d�\�9�����4�/)�I�Z�"n�sƳ����3!���@�=�:�Fڮ�\�ui��f����g=����N����;SJ+�9�g[&�n��Z7f�ح����>|��.rGF�����C���iv�>\�C��7W���]�{����P�5��\qm��e:����뗛��y�{jR7fz���¶ԑ��j��d�D�}�,�6����`qfjv:V��齅%)���;��H��=m����w.�e5�Aӑ�*���`qfjv.��ͺ�:��i#�I������I�� :=�_hժ($����E"v.��f���3�|�,�N���)�CQAӔ�p�75�y�r�yoSge��úڂ�ճ�ĳ�� �n8䊚N�JRRI����Xu�X,ƫfbb&>@�nՁ�ե�¤�r�n7*���y�e*�����P�]� GY>���ܓ��{�{�u`f�B7HUDێ��x�w�b��H�� $w��@����	�I�1wu��mՁ���`qfjv0�c�S{PJSmQ$h� :㘀��/�L@~��}��M��z�ϊQ�(t��(dl`�����)z;M��w5�h�\"p���qX�.�k�;�?b�ܼ@;�1��Vh���b�RH����<���o�{�����:���X�(�@��HQH��w=�`w��Vr��QOﶪ��|�4md'\$@����D�H���W�����"��$b�5���5?~�p�S���KG��9���qLH�a���x� ?5��٤'ҏ��$b�Г3?]`�A7/	d-�b@�vLL%BF0�,%r$3$	������A��M���]"5U�P����ZJi8H
iU�ߓ�|��ʊ+P��Xǿ�^�p�ު+�/:5$�&feG�}�wU��=U`b�u��8���4�$ܒXyfo�Vc�+��[��U_}_}Iw=�`wƐ���(G)�f�m 9����@rj��H7��~��gC�u��ln
�뜚nn+לݮ��'�Xi�ۗ6���V]���GQ6� ��v�ݖ{�u꯿WXo�?��R��_�ک��� ���f=��3)�>��U~���U�G��IF�dNKw߮��ͫ6e.�{U`{����B��\F��a殺<�;����;�,Gk����'�~ֽ��rO����rT�PQ�2G�ř��_�����UT�~}w߮�.�^w�4܉�<��Zs��k����Mx9�\n��٠�wf�S~��j�P��i!E"| �o�`<�q`w��l��57����Q�8R��I�M�%���u~�H�{�`yf�v����ԑ�OR%(G)���X������637y`k{q`n�
��Q�M���|��~J�ś�`<�qa�+5ޖz�Ph�+�B���Ĭ:�,Lzc۾�t�~��7�5+>�ϊ+v��mRcdQ�:{WQR�ju\���P�B��
7@�Kk�]C���n-m�i6G˲�v�n�H<�U[�[{m�R)�v�A�T��{+cV�:Q�̶tg1�ev���:��n�,v�S(��Y��WP\tB�z�r'oEY�������ٰ�1��l��n�l�/
f�l��/�\Qƺ�6�h�y�b�B��O#tN�SW5�&�j�Tp�U��o0ɇ2B�p�x�ȁ�cvm�[v��ŗ���ۛ\��������[�ו��	E������[w�q�� i�ՀkZ�	�z�I�TiHX�۫�Gq�`b�y��M,�5k��b�RH�I��k��n����4�37n,���	J�$�$'����`w�4�;�۫�y��2�p�RO�j�N��wq��� =�e������1���"�a�2���ǵ��y�����u�� �]qk*K�ž�[_���}gmQ���9���q`}��VW[�LLϦ:�}���?~���\i!��H7�`s+��c�8��1ޝ_oj��|���wn�����l��(�I/̤ԌL�HZ\�1���*@yㅠ9�o�z�J6�"rX̚X��Ձ�y���RY���j�6S����p���"��?��~�7�[o������=�����Wj+v�YAw#�u���m���i�m�j��W���O���b�nF����3�߅`��;�4ؙ���6����7H*=�G9�
�\���_�ffR1�i`6����+4W��2��^��TEH��$�3�צ�}�vnTDz�$A��(b�Dq�`3Qh�ZQ�KM7��U�<(w��s�w$�{�Ձ�0�N%jSld����w}ʰ:����,6ecw����E�%LT�A�$���E`{�}�N��Ł��u`~�:�6*�:l�ȓ��IU]�.��u�-��;���CJ�����[�>��F4�[)ē"�����`w2i`fc�؉��u��X���
Ў*�UGs�s8��Ǧ&&���\X���|���D�L�A�j�U[!s��H�������<�Y�ꤎ�ޖk�+�MBk`�n(�	ʰ��K��E`��X�Ƭ:� ���S?%����|�o���ܒ�=3�VkSZ����������Z� <�4V諭�v
�M�CJHP�M���5(Y��Y�z��:���i��v'^ӫx&6#�c�t�UH��$��|��۫��E���ޖ|i=N%jRlc�X��/�1)t�V���ܬj�ǚ�+�$StB&���c��swyf�JX��{q`<�ʤ��(
�]�{�Z ��P�� ۊ�~�����=~�+4)��P�|A��"rX�ƬLLD�o~���Ǫ���,
^��%@" $@`��ov��w���=�-��i�
���.�Z���T �2�j����<7�8�`�S-�*:�aGk�Bx���i�S
&l���))��k��d>;�B�v����%=�v�g���ܻh�v�vr�h-�6]������]��=n��Ȳ��/�kѶ�%U.�vWh؜k�Y�lg���gJ�G���l9�-�l8{���svMdy�ѫ[���{~_���m����%��_�xl�s��Q��p`ksSO=	��΍҄vF�C�9N�#��g��Ձ������?���׾V/M3Ш��J�P��`|��U��1蘪����o����u~��� ��+kҢ$$
`��; �����V5f�DJM���;�����'��H�a<�*���,=3>����{{�`n�,�X�6ff&kwj���G�ģmJM�r+36����}ܛ��W��`wj�32�7M�:lnHv.t�"�Ě�O%��.n�����k�u���s�O�T�����!�!NI\����&�X�ƶg���$��8������!�9v�Iswg9��+�+*���}0ҡ� �B���Q"�{���:�Uݪ��]׿G�$�j��W�m�ܢ$�"'M�E$�K[�7i$�3y\��}_6��ݤ�]��9�����#�z����'�>�w�ܭ��}�IeSҪ�I/�|����LE>;�� ��}�ޱI\�a�����ʫI%�D�G3��3Kky�V�K3�����޸w�^�7㬮�� �eͻU���mp�˷\��n盩�	x��wz���6y��4��$�>$�]��9ĒǓZ��Y��������X�J�$�EkRDV���6䓜I,y5���m-��+�I,�<Ӵ�K��9Ē�F�p��9Cc5�eݶ߾��9�m�~�m���36(!�
l���׿�ߵ�[os���i$�sS�L�$I�$�q%�y��Ӵ�K���8�X�kV�����\�Io�JN�n�dC#�6�$����q$�d��I,��W8�]�5�i$����I�b���#�K�S��;*���EǱv��q��:�W��\u��K�b��"�mb��KM�����s�%ܓ[v�Iswg8�Kv5I�3jHԥR
A�I,��W8�]�5�i$�7vs�%�&��B��S��)"��Pܮq$��jN�I.n���m���$�����$�[��Ȝq��J)v������$���jն�����-�N��:
";?�}�|���]���Q"�
����I9Ēǜt�$��"c����Mo<�ZI%�{9Ē;YQ� �#tF��nnj6��7X���C��5n��<�:̆~�N��w�P����F��Kwo�8�]Y5'i$�7vz��֒׳�ZI-��0t��*aM���$�[��}���Iw���K^�5i$�2��=U�͵��Cv��t
�G$i�I%�{ӜI,y5�K�}�owo�8�Y�y�i$�ڂ�&�m2)O2��k9�o�����컶��{��9m���i�K�7��y�${Ѥ�H~�F�*�R5i$�3y\�I~���o���}I%����s���g��ݶ�:4Q5kD�H�	$Z�-!V�3"�pʫ�$(H�Q��	 B�+��%�n�W��.r8��m�⨚��"J(Q�!
D���Tf�.��0���l!! �$�*�"7�b�^!E��$�C�B(�$5��# F)(HH�"���]�I`A�V �� �"@$!��XB$̭��	!�0�d�BE`ĉ$HR1X��#��l��O4I#d`D���
��a�RH@��@	@�@�!�k�~$$4���b��bF+��w��~k�*�4���L��W����H�Waֵ�qA,Bu�3�څ��k�yZ�*���iT^^7b�^�H�u�ݮ˳�d  �ً��m��\ે6al\���UT65&�-��S�84�9�J�:�pu@�Gm��ݮ�n�t]���T[l�.���l��Vh -�cs�ٝ���s�9����;%�;{ ��.+q�e�Fݱև��b����\%��� (=ft\���Y���y�ԧ�8�o����Z��p�x�h�疪��b8�l�x��p���"V�� �Ƭml���вst�!� ]6�P�l��Ԅƅj�ݓ<.Z]�&����uWlˬ6%,5U (vl����ڃ�� �T� p6Ͷ}�)��qUJO=F�Px��C�j��h
{l�=��ݵ���  lٴ�͵m�b@[��L�~�>���k���w`.�6{���ڥj�>[���v
�ٕC��]�-1��e�� �A�im���=O+E�s���k�8��"�ڭ��;Ӈ2�h9�)�6���m�8�sA�u��
�k�]Lv�ltv�h��t�ܦ-��{)S��e����$�9q��Ѐ���b6c����A��3����v��xi�m82m�3{\6�ً�C�7!��;���l�J��q�ݳ\�T�O���%�Unm�ݛ�c(lu>Ok��רL������v�	��6��tm�r�����s�Y���T���؇��\�*����m@��ɘu�;	�|���
�i�ڜ�9:�Y�S!��&�=��nF��7;Q
���m���GYQ5<�Ƭ�`6�7���u�]C'�e�j}j�����7-֭�� ��T��b�kU�ӊ��2�n����T]6�Hm�<�m�C�6�^����f��7ir5Tkv1��z p�'P[s��@�����]�ԔSt�!4ԖY�.���܎����[iT�Dפ�-� 4k�:ƽD�+Z�hE�C�U�L?(�!�	�]�y�8�C�.�����(��z(�T�w�Wd@m�] �7/�v�s]��n4��[���ĺ�E�ۛOF�&�eԯ���9�,u������@��''F֞اd2�T���vF��I�E��yūt[�]};�����N�9�e�P���spF1mێK���2S�e�ݽ)�dL�卲���ٱ�J�@��:��j�\�P�TnW��h�ƺ�L[L;%�#��`H�PA�mF���{��{����?9������v���b��Q�'.&E!������7-g���+�s7���G���#��^�I~�v�K����Hǚ����6���r�Ē+��l�G�t�#N�Iswy\�����$G��)i$��~�s�%�sZw���YOux��1E��+�I#^�KI%�����勺��v�K���_�ꪮ���ǈ�[������������~����$�k�i�I-�{Ü��r�]������Ʌ�5�����q$��kN�I{ﾯ���{ݮ�$�{�-$�f�+�I,[ZՍFAIAq��דe�*$���</$i.�7he�:��9��.ٍo��{�k៚��lsl��-���r�o��u�����������[������� ���Eʖ��9m������9Ԣ�A �@HF Ս�Q_*�5o����In�杤�����}UUM�{Ѥ���(6�*�9�����\�Iw֝����m��W8�K^�;I$��5�b���	��^���y��Ӵ�Y�{��$���ʴ��=3<�ｑ��$G��Ģ��q�/�"HӴ�]��W8�^�����|I%��r�Ē�9�;I%����FEQ��'*y����6�{Nv2�V8c���>�s�%/;����{#�G�
y�
�����wٛ�����r�}��\����Ȓ�߿r�Ē���7WN$����r��If7�}��D�L�U,��UV�K7w㜶��}�f�
"9�o}�\�CXaH��nJ�K�&�$�ww��.������D5�^���ݶ����s���{4f�r�!LѓW5���o�"�ʊ���G�$��o��$�cG�$�v&b"8���I%�+l��W�F6�$�q$�_�um����v~�m�g�뙻m�����K~z��n��T������۳��6ֆ�#�:V�T�
������G��{�4�1;�)S����Kw��s�%דS�I%��ѳ�$�SګI$���R�1HԌR��s�%דSw����ig��W8�Z���I%����=_U6��b�Ȝq�暑7i$���+�I,o5�K�}_6�}�W8�X�y7i$���P�Aqp�������/LǦf#�w����[����[o��]�����M�w���C�}�����$�~?ܡĔc�61�݉%זϾB[39�z��I$�w�����[��YOkC��dQ:)A�6e3�M< %�/��K�`9)�ח2X�$}��w������TAM�]�Ic��ݤ��n�Ē��[�UUW�m7��_���Ӳ�)�*p�'i$����s�}UU�mw�ZHY��+�I.����U}U�6��-RN�Ԇ�6�$��$��|夒�n�������l�i�I,�{�|I%�lzSnR�ԎZK�W�����K='�v�K����^�����-$���4�~�Jqan�� �~��0c���{ǻ������/}��ݶ����9�mCN�~?�����-W�`C�̼ps�m�gF��I&4ȓ�h�����ѵZ�q$�`'�� �-H%�)�V�O r�r�	T-�M*���\;/�����|�<N�'����vrV�;��]�^jٻ�;��ݪ�
c�w�5�s�si�F�CɸEqۂ������\2�b����� d 5J�m�n+B6���9�h�����t&.�\ӳh�{���~t>DИv+h�*�r�X�^+�:��2)��h�������X����~|wEǞ5�R�$���_�HY��i$���6'���l�i�I.��h)�"qJ%(ܮq$��l��ww��$�vMm�HY���s��6�x��DlR�e)#��K=�r�Ē�ɭ�K�_4�}�W8�If�KI%���r|*�j8&����/}��=w���ov��>�>Xl�,�ߢ��3b��>`��q��37n������}�t���Ձ�٭Xǭ��������������X�͝���Zr��ڵ���un�����BuWHjSmBI\ ��K����|t�c���Xw���)Vљ�4B��Zܓ�{ݛ�� @.�;Ϲ��׷����DDG�*��ꢪ?A�F�b�NU���?5`fn�Y�H��K=�]X�j��dRΑ$j�������}����]{{J����F�2JR�nU�gse�ݑR�l�@7"��[.n��`Nj�\8'>�,1f���%�;E[�Bl��@�ҤIOQ#�C���Rl��=�]Xw8�X��l��oy`n��/��D�Q�4��`s�5����}��Ձ������Ձ����g�$��I3�O��lܓ�����Є��U:���QR�8Z�Jۼ���f^�f_s�a��Ձ��q`}��V���,��M�My
1�)��7sn�u��u�Ł՘���Ff�	TUok�&�w��btڵ�5���kr���tn�^K��
Ĥ�z���n���`7�����u����K�4��JTp>T��+s6��T��w���|�����J�>����~�\�$�L����`j��;w&�z��.��%`{���a��":jSlc��{�K�w~��~�u�w$�~��ɥ���e����y���N�DpLq���f˴�*@u�1#� ?�WT��(�ι�f��p�l�&մj�A׋��-n9�g��P���uMy���w����;���cj���q.��o�,��Vy�l�D��:��V����5^5)��$��3]���Ĥn�i`u�jVx�/�艙�l��Ѧ���!F9E7v��ߕ���4�و��Ku�Ł��� xꊨ|�I���"���W�R���+��]XY��׺�4֊Z�&�GΔ\�Vm�X1M�|�n���4����v���p_˹v���I�{y%(+��7;k�]*��5C��GNٔۜ6��7. ��6��-4��6H���m��-�w�nի��{ive��Ŏ"Z
vi���Tk�p���;)�0��q�c����L�]v�;N<�l8��Z1��cl�f6�!�mŻ6蝓�L�;��ǔη��rE�����3uW\����-�cYZA��Y�]����Kr�8��d�R�cU<�f�[��u��L;�����X��ʾ���=��G>�IS9*B�nV���;u���R�}U\A�{�V|i�r�N���\�X�j�"e#��R�7wn,�������&\ut�#�cN+���X�qg�&R�S�`n��1�:-B�0A ԉĬ=U�����Vq��V�����L�?}�8�\�G�Jm�I*��^j�=��UW�=��;��J��ݺ�?n�Κ�q�ܤ��m51`��u����|у����F�uG�Y�լ΍Ҋ6��Q
1�>nE�?~�+�٩X�q�3��=V�j����K�+5m՚�]�9����A���*�b�4\0�0�
!I�+����y���߶l��+�Ưf&"fRimRG+Z���֭ܓ��nI���n��?�,L�{վV?s�X]@�B\�\�s�.Ur,�XՀ�q��|iXl�LD���ܫ�4��&H69I�E"�7q�X3ͽK�7^�Xv��������c�\�<c�O�=x�Z����]q[���Nq5O)��=�{���þ/H�q�J��O%`nf�X��^���g�u`o�<�J|�H5"q+sŁ�k�[��>��J�1鈊�ލ�GI��q��I*��~����Ռ~�Nb��T!�,-k�1\���M��|*q ?i�d_�g-�.�m�n���8�p�	?PH���F�֐(ZG��df�F,HJH$�����~' em��փ�"�B��+\�4h%�bX�p� C$��\&0i�����I
�+)����V�r���$���v�'���Q� �
 
p�U��j�M(|�o�p /�O�!�%��T] �O��~�n��z����I��blr���X{���z��o�� =���avM�7�Mʰ9ݚ���g���ǾV�M,�z��hkɤ��J]�Y�ٸ�[�k�|7FNl�u�3�=˩�0��_�D0�F����E��������k�72i��︃��,Zx�
��*N{�����1� =Ҷ	�*@na��R4���(�;s&�:㌳ff&�ݸ�1cڰ1���TP���1)���5X��VWs]��1��L�ݻV郢�E
�G^�ᶀ�EH�s͂�4���}�߿~��Cا��$[F.`xHd"��47n0�n0v��9�5�i�
��|u\�8��W ś�`n��`s�_���������Lm����>NG`n��`}�����,���ԃ^�	����Vs��7wn��%�����������RߣJF��Xzf'��{݋��+�Ƭ��5`ut�6�Aq��Q�Vz�U����rN~�n���ٹ'E
D4��'�^ɗ~ڇ�(��΋���M?�#��5��ؖQ��n��^���e��e�k\���Z�;YNjM!����D���!�3�e�S+�.0	&��h��+i��;f8L�n	3����[�@쁻 ���ۑ�J���W6��X��a<����y�nь������Q��q���g���<�+��64���&��Z���<���2���~�����w{����o�9�^#i'*J���0��khx˧�F�uBV�7H��R	��7_9�n˜��"�h���`s�V76���^j�3wS���:JD��E`s�W���{q`fS�`gk��Hz3h�P�cdQ5"dV}���:����}�}����~Vo�~V2��Se6�T8���� :��@>�-�KA���?z��Q44z���7#�3�4�=��6/O��:�����5@�B�x�.�fܐ)���ӊ.rX9�7����l��M�q7�*����(��[�m�����>x�,���LD��>i`c�P�j�j�K�kSrNw��ދ�B1RDR��C� >U[�~�rO��Ł��M,Y����Q9������:�;��,ؘ��������;���70��t'(Lr�d$��+�}��=�Ӏw+cU�}�\11��u`n�2:Q�:RI`s�kU�s�����k��6X�z�*W^d�)J�х�eF1-�Gc�:�st%]�3�x�j���m6K��U)�lj�T�JF�������K����;�|ٙ��w+cU�ס
9��Ɓ�'RI,���ɥ�ν�V�����I�Q4:^�Sp
nG�'�w^��s�t�ܰ`�� c�!����:�|�s^���A8������R��M@u���rE�@f�j��Q��O��X7vX��x���M� =�IhQ�1V��GZ��l�nN7i�v�v�[d6���LXubݴ��X\�Z�Tz*H�5_6����u`fg`}�pק�1=�3��,n���%(Ӕ�!$vfM/�_U}I���`��X]�V6�Z��\B�&�p�9׵��9���UUURX�|�͞,���:WI�$�����bbf�偋Ձ��2��㈘���vj�;�6H�DSQ�ԒK����ٙ�x�O��oV����iw��ߦ�m��-k�ա#Y�SjΙz�f�ܴ��A������.���� ��|sg��ښX76~��Y�v���H�j	JJB��v���虉���o�`4��`gs��D�Ͼ���l�<�&Eq?��*�������b�� =Ҷ	2�/+*)#QG#���_RǛ�`g�x�9ݮ2��3陭��������Q�\�\��	#�;�4�?}U]�U����v���srO����"��9�њ֬�h^p�������*��~t���5L�9���X�b��1�`�y��Bq�r��Ω�k0�,�Z�����s����N`i��A��n��c!v-���9�@ra�i�g(��m�]��:�5on�e9-���lO9m�0�ǧ��n���B����ꖘ(;^vB�nn�y�BU��V.�pR��u�&M����/d4�wO{������ݟwڨ|�4&�g��ݶ�>x�}���xNnawVn��Nr%<�"�wy���%��lUs���{�9��������:�:��X]�m&��܄r&E`b��}�ґ�Ձ�������W���gZ�!M)M����|��f�;��`uwu��l�"87#�و�Y�zX���`uu�������O�_=����=�����r��R�!`{�T�_I��s�`�w]v�M	��te�;���E�\w7|q̆��=����É�۹X��w{:�|�h��Ǌc��1f�X]�Vz��zg����`~��~�7Q���9����e/��z(�*~D��}�vnI����ܓ������#<i��$�nRl�����,�N��)b�ڰ1cڰ>x�WJ��#�rG~��m��������`uw5�~��������o�~��l
ND�����:�=1��k�74�>�8j�߿��v�v��0+�L���7#B��f�.Y콬n���e��t�~{�M���D�$��b��7�4�9׵�����`f�m�1=�Q8'#�7�{�ܭ�V�{VWq��jN8�jP��iHX���5w5ت��3��B�
J�@� ѥ)EY�Q:9̽߳rN~�,�XE��Q����u����}O��z������,<��f�V�6�L�H���9����`~���o� �zV.�6��M���6P�G���N9X��#t���W�4@�
�z��d�T��謅�d�&ڔ�!$|�����^֫s]����`ssP���HR%K��ݧ_�c�F�������٥�����M�]2��(�n��1cڰ:���؈�L�Uc�<X���`s�A�m���cDq�{睊c��ܓ��צ���;w'Ő�.��u�TW��3v10boi&������,DDDG�&'�<�O}VWq�ͷ����ym�sD�9Kqbn�h��;Y�5�;K>N�9�qq quņgJL��)���ԅ�ν�V.�����W�}�͞,4��QGe0�#������DĤbǵ`w4�>�8j�3�UU$yV�ڧ�5�X�}Vٜe���K��5X[�X0d\6F�mJM��;�ɥ�ν�V���|������+cHD��9#��4��=�j���s� 
��M@���7�B��-d#K�����@��:L���"�!!��;>'�zE�@	"r�0�F$"��$���~shK{1N~�kF�QU�P����q�>-��͒8�q�X���n-U\��Cz{ �s[GI���I��=]"y�X�k�TUm�F�]�i3Ɲ�o:wm�d�]�h ����+V�x���*��xMZV	�̠[��9۳;��b��Ga���%������8]�	���[lݶ��m1�,n�ո%6 .�d�H��w;ky��=�*[:�{�[a�5��7W9=6[��� 9�-��m��=�S�x፸r��mػr�d�U��L��l{<Vr	s#jc��uW-ܗK����c�M\F�Ȳ���
{ 5���x���{h�� BE��t���6�ڹ%��Il�� ����I�b�#�{&v\�UR��ѡ;�wEC��@:K+.�-�*�WK��UTc���-�I�ҘX:�-O+UF������.��f����k� �.�\�F�m�n��-"I�&�r�I�[1����2��R�,p�6�iy"gm�ی���`A�X�Պ���W��t��ne��u/\@�GLէL3%�囤{D$̺Da��v�v��g�gx�qɖ�J,'�u[��y����F��R����e�s�c�8ƎѶ+) �pk���Vuʻc��ۚ�����=n%q��� �s8[\4<��n� �8y}Q�  �T��V-g���h� �.݊^�����o+m�Yu�0t���3aNxzS�R!��8���NǇn�h-��Oa�R�k�l�KF�2-UJ`vɞeUbUp��\4�t*$<�'S�2 K�Ɲk�L<���X�)���88����HrK=W`�nrY6�3[SrH>&��S�89�g���0�J�-O0UΊ�UU\�1 $6�U��A
������eN�����
0���@�&`m���w�fn�!�]���t���n��������*:{mS�L�I�ш��<�N��� ����Tu&�ʛ������lsv�g�JTi��j������5��調�����{����l"u>�b����/�S�=x�Ơ�O�u��w�������e���C�5)/8�Im��0#Э��a�x�5s�v�m�K$���T� ;]X�8����VJ��3ų F��:�c�˰
a�;-v͐�a�"Ns��YصGc���pF�0jwWF4��	њ��84�ps�� o$k�
�ñS�H���Q7�%���r��{!E��.S���mץM�g�����8��8]��0�3SVə3W	�m0.�\y�)�6���)����l��L<�R�MȔr&E���`uw5�̚X���`s�A֨Ȣ*(�u#����1 �� =�*Z ��W��Ѿ��hb^��r���X�<X���`��`w�5X�N�q�:j{E�\�1 zI���A��"�X�V�����S�n�<齯�����󡺰P��P�H�d�@��;P-�Ѷ7\]2u0�Nz�0��j��-�����>s-	�j�6�7�`w3��>t7^����{��7t�Vء#b�6BH��M.����|�}3vR7w� �w�M��>Ƅ��D���N8XKw]�swe����//{��������c@���"M�*�,�o�M��;��Xl��[��3UOJd��*(�u��ջ������7�� ���X��,�c���Ev��zsΝ:��IX�x�Ӌ���s�`�-p�L�j�7JY8.������q� ��aw7yq�0��L"c��{6��bX�%����֤ˆ]KtK�M�"X�%������?��DȖ%�����r%�bX������ND�,K��~�NE�,K���ɪk5�2d�K�kiȖ%�b_�����Kı=���iȖ;u 1Q�$vr'"f��M�"X�%��;�fӑ,x��{����>�M	�Z�{�7��`'���m9ı,O���6��bX�'����ND�,�dL����Ӈԏ�R>����W$lR��I�\�bX�'﻿M�"X�%��=�fӑ,KĿ�ﵴ�Kı=���iȖ%�b}���3'
\33S5��sL�Ig�+�����[Tn�1!a���qs����$��D�,;{�7���{����߿_�9ı,K���[ND�,K��{6��bX�'��~�ND�,K�z�L�əL���˚ͧ"X�%�w��Ӑ��DȖ'�fӑ,K��}���Kı<g���r%�bX����>����G������7���{��}��r%�bX��ﵴ�Kı<g���r%�bX����m9ı,O���L̹/��3Dn���r%�g�"g���m9ı,O�?���iȖ%�b_�����K���B#�iFT!! B#�b4����>�Mw��fӑ,Kľ���5ud�fj[�[��ӑ,K����iȖ%�b_�����Kı=���iȖ%�b_��kiȖ%�bǿ�Y��;<��!͹W;C��v����y�rs��'6X:����TpO�n�|�G,��}�O��X�%��{��6��bX�'���m9ı,O���6��bX�'�����~oq��������� �Бۦ�iȖ%�b{=�fӐ��L�bw����r%�bX��fӑ,K����w�p���#�G��x�lP��J55�fӑ,K���w��Kı<g���r%�bX�������bX�'���m9ı,O���۸z�[�֜�f�SiȖ%����k��ٴ�Kı/������bX�'����9ı,O���6��bX�'{�a.Hs&e3SW+.k6��bX�%���[ND�,K�?�����~�bX�'{��M�"X�%��=�fӑ,KĂ�ڞ=p�e��-��r�λ��u(���V�7i�u��ڮ6*sZ�[f�ݰȍSNK�֓��d�N���d	��� �<Ö�*�Kcm�k[!-[v�����	[dUv����0=�6;vѸk�n,��3{^8m�;:������yW��pr]�g]f(]^����l}�V�|q�7�Y:�/!�WF�9N���Hr-�td���N�A����iW��اl���0A��Ү���Ti�#�n<s&��\{t�i�:��m�f�D�����oq�ı?{��ӑ,K�����iȖ%�bx�wٰ���dKĿ{���r%�bX��2�I�j�5euu��"X�%���ߦӐ�B9"X��{�6��bX�%����ӑ,K����m9����oq������r�#�{�ı,O��6��bX�%���[ND��ű=��I�$�~�u�$D�������B���n	"z'��}�ND�,K�ﹴ�Kı>����r%�bX�3��m9ı,K��|�.�";t�|�~oq��������ͧ"X�%���ߦӑ,K���iȖ%�b~Ͻ��r%�bX�x���m�Y��nUp�.ݱ�5c�9��l���v�������\�1H'.�O%#���k绑,K�����iȖ%�bx�wٴ�Kı?g��m9ı,O{��ӑ,K���Ym�>����NeֳSiȖ%�bx�wٴ�>t�	��\A��D�K�~涜�bX�'�k��ND�,K﻿M�"+�2%������߆Uu"���~oq���������r%�bX�����Kı>����r%�bX��wٴ�Kı��
|�)�#���ԏ����2'����v��bX�'{��M�"X�%���}�ND�,K����ӑ,K����a�g�]f���5v��bX�'�w~�ND�,K���6��bX�%�����"X�%��k��ND�,x�￿~<�{}���a�u;c�C���۫ɺ��3�����U����&����5-�˭N'�%�bw�_��iȖ%�b_�{��r%�bX���ٴ�Kı>�w��Kı/��N�SZ�ֵ�ٙ���Kı/����r� #�2%�{���m9ı,N����ND�,K�k޻ND�ʙĽ���S�DGn������7���{�������Ȗ%�b}���iȖ>��(��F����U�b)��`1�z���	��D��]�"X�%������KǍ����ￜ��8�\៞���7��b}���iȖ%�bw�{�iȖ%�b_�����K��	�=��]�"Y�#�G՞�����#i�)�q���Rı>����Kı/����r%�bX�g���r%�bX�}��m9�q���;�}|���m��q�ӄ�p��ێL�hծ<�^�V.K��L*۬�qٗ2f�fj\��r%�bX�������bX�'���6��bX�'�w~�ND�,K�k޻ND�,K�}�\�Ժ�j���Y�kiȖ%�b}��i�ș��}���Kı=�]�"X�%�}�kiȖ%�b~�w0�d3Ʈ�VSY��m9ı,O���6��bX�'~�}v��bX�%�����"X�%��=�fӑ,Kľ���j&��Ĕ����ԏ��gչ{��Kı/��m9ı,O���6��bX�b�ʪԈ�����=6��bX�'��{SZ�ֵ�l�j�9ı,K��{[ND�,K�{�ͧ"X�%���ߦӑ,K���ߦӑ,K���t�g�[,�l�l\Ƿ'v3�E�i����F�I����5k�tg��%��wFB/F�߉��g�����iȖ%�b}�w��Kı;�w��Kı/��m9ı�{�W�ME ����㿫�ԏ�'�w~�ND�,K�w~�ND�,K����ӑ,K����iȖ%�#���	_�MILc��p���#���{�M�"X�%�w��ӑ,K�����iȖ%�b}���iȖ%�#��{Γg)�i��7"p���ԏ����{��[ND�,K����ͧ"X�%���ߦӑ,K�&D�����iR>�}Y��_�ʐQ���G$���X�%��=�fӑ,K�����iȖ%�bw�ߦӑ,KĿ�����Kı<�=<�̆[��Ve���Z+����-vWvz�+#c�D$[K
���9:���Aћ�]�Ncm��y��5&1���In��\��Y��[X��Ӊ���H��he�j��՜��ۖ9�Y�u�z�5�ˠ��[oN{s�[�f�bt쎱���i�$]۪����,(ダ��IyT��ą��!n��ї&��i鋐��
��jۅ�Vf�k� |�V	�7Na����5���rf�����0�:ci��e�m���f;
�r�n��t��=���7��,N���m9ı,N����r%�bX�������bX�%��{[ND�,x������k-�e��V�����{��'{��m9ı,K��{[ND�,K�����"X�%���ߦӑ,K��=,����5�ji���SiȖ%�b_�{��r%�bX����m9ı,O���6��bX�'{��m9ı�}J�7ġ:#��
����R>�%�{��ӑ,K�����ӑ,K��{�M�"X�%�}�kiȖ%�R>�n��B22F)I��r_���GԢX�w���r%�bX��w��Kı/����r%�bX����m9Ļ�ow���Qq�0Bv�6�۶!1]�&��]N�\��7�k';.���Lͪ��֜˚�M�"X�%���~�ND�,K�ｭ�"X�%�{��ӑ,K���ߦӑ,K����2p�2�L�L�j�ӑ,KĿ��ki�xD�:�C��m��K����ӑ,K���ߦӑ,K���ߦӑ,K����w�Z�Y]�k5�m9ı,K������bX�'�w�6��bX�'~��6��bX�%�����"X�%����)�����YK��kiȖ%�b}�}�iȖ%�bw���iȖ%�b_�{��r%�bX������R>�}H���{�r����(e�ND�,K�k��ND�,K����ӑ,KĿ��kiȖ%�b}�}�iȖ%�b#������f��&uCi{hq�s;�N�n�������-�S�����ݷ+.���j�x������s�dK����m9ı,K������Kı>����	�&D�,Ow���NF��#�GԼo�M�HHJTG$��pKı/�w��r%�bX�w���Kı;�w��Kı/����r%�bX��a��.�fK��C.k[ND�,K���6��bX�'~�}v��cQ5��0~���=���_��	NE� ��������T"y� �6�׃���" ��@��t�U08���%�J�*	�B�ԥB'�e�iH��Qe
��A ć4�mw� �IE�ؖ�&�H�� pO����Z��I)H6�
i� ���� @a#1B� �s�5�Ǝ�s��+�A:���?B,�9���kiȖ%�b^���ӑ,K���[K箥�5���kFӑ,K?�`dOw~��ND�,K����m9ı,K������bX�'��m9����ow��߯�9�3��=܉bX�%��{[ND�,K�9������ı,N���6��bX�'~�}v��bX�'��n'�2e�Y��ѫ�i^w<kZ\�t��ˁ7V�ռ�Q��]�:�#t\�M_=ߛ�oq���Ͽ�u��Kı>�}�iȖ%�bw�w�iȖ%�b_�����Kı>�w�*�1������7���{����xm9�V9"X���v��bX�%�����r%�bX����m9ı.�O�p��i`�����7���'~�}v��bX�%��{[ND�,K��}��"X�%��{�ND�,K����{jK�k![5�]�"X�%�w��ӑ,KĿ��kiȖ%�b}���ӑ,K�]j�����U��D�o��ND�,K�w�p3j�����{��7�������bX�'��m9ı,N���m9ı,K������bX�'�5�}��3MB<��Ֆ�I�B�qm<���^��6��bu�n�]N.ssZ�r%�bX�w���Kı;�w��Kı/����r%�bX����m9ı,O������5eִܹ�h�r%�bX����Kı/����r%�bX����m9ı,O��p�r'�S"X�����3'ɓ2f�fkY��ND�,K����m9ı,K������bX�'��m9ı,N�]��r%�bX���=�f�,5��љ��Z�ӑ,KĿ��kiȖ%�b}���ӑ,K��u�]�"X��J&+7���|L"a��m�QT���\�]\3Y�kiȖ%�b}���ӑ,K��>׽��O�,KĿ{��[ND�,K�����"X�%��ȋȡ R m�.A,QB��Qi&
# �����w����k��-���L�x�,3u+x���R;F;�B�\����cGW���4�۪^۔�VG��D�Z��; �^@��\��j� u���ҹK:!<���kȕ�'/�:ۅ�qmc��Z���ы�:��l�ۥ=@�K�M�s��[�j3MN�M\�"li ���˜e� �HGy
ځ��Yt�g����}���i�u�f]��_�߾��������t�Z���a^���5�
/lj�O��hk\D��]gJ��sY��噚>Nı,K���6��bX�%��{[ND�,K�������L�bX����m9ı,N�����a�ї5����Y��Kı/����r%�bX����m?��2%�bw����Kı=���m9ı,J}�}���$$%*#�K��}H���#�]��Zr%�bX�w���K�!�2'���ͧ"X�%�~������bX�'��{9t]�K��C.k[ND�,K���6��bX�'s��6��bX�%��{[ND�,K��}��"X�%���@��&*��]�������ow��}�ND�,K�ｭ�"X�%�{��ӑ,K�����"X�%����~������Ѹ�����N掇��Cr%��P�nn��q�Nrr/
]�rfr��Y��Kı/����r%�bX����m9ı,O��p�?DȖ%��￳iȖ%�b}��o�5��5-5tfa�ֵ��Kı/�w��r�ڠ��B)�j `�gtU���"X��ϸm9ı,O���6��bX�%��{[ND�,K�wy�2[��s&h�3Zֵ��Kı>�}�iȖ%�bw>�iȖ%�b_�����Kı/�w��r%�bX�ݾ���f�0�|�~oq���{۹������r%�bX��kiȖ%�b_�ﵴ�Kı>�}�iȖ%�b}��O�Z3Zѐ���Y��Kı/����r%�bX,s��ki�%�bX����m9ı,N���m9ı,O��;�.�y�*�K�r1n�f�F�u�%�����́���'���Wj���v�Y�k[ND�,K��}��"X�%��{�ND�,K��}�ND�,K�ｭ�"X�%��v�]F��蹐˚�ӑ,K�����"X�%����ͧ"X�%�w��ӑ,KĿ��kiȖ%�b~������I�ִܹ�h�r%�bX�ϻ��r%�bX��}�m9�zQ��7q/��5��Kı;�}�iȖ%�b{��pg�ܙ��S�������oq����m9ı,K������bX�'��m9ı,N���m9ı,O�z|�0O�t\-�~{�7���{��?�}��"X�%����ߍ��%�b{;���r%�bX����m9ı.�{�������aY�:ws�A؛���-���7c8�x�e���KU�i��%�&g�4MLֵ�q?D�,K����"X�%����ͧ"X�%��;�fӑ,KĿ��kiȖ%�b_v��u�u���kV\�3Fӑ,K��}�fӑ,K�����iȖ%�b_�ﵴ�Kı>�}�iȖ%�b}��x��Z3Z�Geֵ��Kı?g}��r%�bX����m9ı,O��p�r%�bX��w��r%�bX���珞kZ�F�K�kY��Kı/�w��r%�bX�w���Kı/~ﵴ�K���C���2YE��)Q� �HD�R���, *���"@���A(���DX�JF0Q)h��g?D�k��6��bX�'���=��.�k-�3!�5��"X�%��{�m9ı,K߻�m9ı,O��{6��bX�%���[ND�,K�W�?�������j]kWZ2�\�m*�����c��6X�E���'u��e  �F��֛�5�q?D�,K����ӑ,K�����iȖ%�b_�ﵰ�!�&D�,N����r%�bX��޿��Rh�[3Y3&����"X�%��;�fӑ,KĿ��kiȖ%�b}���ND�,K���[ND��S �'����2[Ls	rfi7�I�����$D����n	"D����ӑ,K�����~���7���{��~/97�K�5Vӑ,K����6��bX�%������bX�%��{[ND�,��}���7���{��>��~����0���bX�%������bX�%��{[ND�,K��}��"X�%��{�m9ı,N��l+"��OS��u��M)UDm��eZ�7lV�(�$�g�V�چfA�æt��M@7	����Ԥ�<���l�8�9�]�B�k�z˲q���V�`˻9��[HW*���'��Ͷ8�n�7n.lΥ��K,ݻ<��\�lq�Ok���Y�s<�9;�&	;X��cu��6������-r�gL�J4[5t�u���6q[�*�8��=�-���r�d'g��J��m.-�7]k2cX9K�C�u�ڶa�]�	��w�o�M����U��ؖ%�bw=�fӑ,KĿ��kiȖ%�b}���ӑ,KĽ���Ӈԏ�R>��j�u#��)P����"X�%�{��ӑ,K�����"X�%�{�}��"X�%��;�f����{��7����w�..����9ı,O��p�r%�bX��w��r%�bX����m9ı,K������R>�}]����U	�$�ӒU�"X�(@ș���[ND�,K����m9ı,K������bX�'��m9ı,O{��W�2�Y�ə5u�m9ı,O��{6��bX�%���[ND�,K���6��bX�%��K��}H���#��o�|n&�'�Ԕ׺�5�9�&V�ɞ�5�ńm��65P&	�fz���P��չ.T��~oq�������[ND�,K���6��bX�%������bX�'�｛ND�,K�m���68I$w�p���#�G���m9?'L��K�}����bX�'����ND�,K�w�ͧ'���{��>��~����0�|�~d�,K���[ND�,K�w�ͧ"X�%��;�fӑ,K�����'���{��?�N�v��Ϊ<��|�~g�B&Dȟk��ٴ�Kı?���ٴ�Kı>�}�iȖ%�b_w��ӑ,KĿO�}%�kY�th��ֵ�ND�,K��}v��bX�'��m9ı,K�w��r%�bX����m9ı,O��=�3��5�S����]8ܻn���+h�d�`�縙��a�v�y�� ��Z�����Q���oq���;�p�r%�bX��ﵴ�Kı?g}��r%�bX�����Kħ��yy��>P:$��q���R>�}V%���m9�,K�w�ͧ"X�%����ͧ"X�%��{�M�"X�%�߽�%s�-%����WZ�ӑ,K�����iȖ%�bw>�iȖ3��� A�S� @F@��mj����+�X���\���r%�bX��w�6��bX�'{�^j�k2��&�K��k6��bY��,��w�ٴ�Kı;�o�m9ı,O���6��bX�'�｛ND�,K����9C�c�㿫�ԏ�R>�ݿ�Ȗ%�a�@�����O�,K��=���ND�,K��}�ND�,K���|�����/7����/k�#�ri��Փ����6��J��M�#�Ƭ3\Ƶ6��bX�'�w~�ND�,K�w�ͧ"X�%����͏"X�%��{�M�"X�%�~�;�x�Z�Z�Ӆ��M�"X�%��;�fӐ�V9"X����6��bX�'}��M�"X�%���ߦӑ?�*dK�w���̺��4R\ֵ�ND�,K��fӑ,K���ߦӑ,[�����iȖ%�b~��ٴ�Kı=�����T�#��RGW�R>�}Y�~/���%�b~�w��Kı?g}��r%�`` ��]\#C�����m9ı,O���d�楔�֋�5��ND�,K��ߦӑ,K�����iȖ%�b_�ﵴ�Kı>�w��Kı<;iw�R�F�5�,��Sic�f 9�*��I�]�������m�
{�s���i��w���oq���｛ND�,K��}��"X�%��{�M�"X�%���ߦӑ,K���H�`TeP�$w�p���#�G�w��ӑ,K���ߦӑ,K�����iȖ%�b~��ٴ�Kı;�z�Bp�K�5&���m9ı,O���m9ı,O���6��c����>�fӑ,KĿ{���r%�w�������1��b��w���D�?w���r%�bX����m9ı,K������bX6'���6��bX�%��釋u���f��Ѵ�Kı?g}��r%�bX��ﵴ�Kı>�w��Kı=���iȖ%�ba�����%g�M>�����)��m�� �H��&}\6FH�I
��~��1�H2C��`�#!��1�'��t�<��C�~?1"F$�1! �BB����w��|�a�S"� BPg~��cC���'d)bdK��M�&�AĢ"�[��a H���IH��U{\�I	$����`�)�D��RF,!�@�@�:����U�$�r�`H2�b��4�E�>֤�E�9M�0�@
F�| ���I,�M �H�C�V�}�EHE'���$	J���~�u�[I�d9�/m���r���é�5�Iu�"ۭ�{��[�%n�0�m  u�H��]*#:�;b�ƅ�;"�LRn��_A�������nUV���vm���*Q�#��Q�iZ�m�C�\뜗0x6�������!���Z�H�V��m�ѣ�2ܴ;ɤ�-��e���u�Ë�=���.�nys���ݰ� U��L*kX���Zϝ=oem�[f#�k��p��u��꽀�ܼ�n�T��u(�T�:n�r6M�k�C�q�Ps�[Y�sT��aU#*�V��Ul�n�FV���Z�T�/ ;��*ȨX8�ଧ5��Yv�$m&�l�6�մP�]2� ��PN
�س�qUT��mZiKmP��oNں۩h��׭�MgE�` ^�lҷg-�u4*�tn��mg�`��KY��8vK/4*���P�=�H�� ;UT��2�0�]��
TTkgQ� l��;;��������Ѷ�×nprl�q�鵚kt�^ڌ7-X��5Mr���Ǡ�0vׇ�;Cx�zp�ac��H�n���s�������睸C66�8����r�cB�;h�˱�]�u�=/ ��'��j^MA\�nW.u�=��� ���mJ�J��:��k��*�Z�a;j�,Q9q��8]�v�X�b蓵��8r�if��ӼK�b�F�	��ϣ���[O�e���49�G�uA��	W����ch�@)�$;rE���dL-ڜHMC�ʆ�;m�e�4,�ʸ��Ìt��ZMm,�5��ў�y�66��v*]Oq���Bm�z�(mi.`S%U+* `(vݪ���P��C$�6+�lRk�:�nʙ��`�f˰�������uYT�3�v�:��XcdB�=�˺Ne�5�r�֙v�C]�U*����+#�6dJ���v�ڭ(s��z����+��ڰ*�l
�c�96��%l�:�˹c�U_;���;GA����8���|�G�P��6� O��O��@�(0D�C����9��Z�Tv�т�F� �KbN��l\��0�uέZ'�:�h�Ψ\a�1�W#X��5F��#��7'1)�a�آq���Z�ґ�mĶ`gr=�؍�M�h�0�0�$;�5n��IwG*�ͮ��η`�Ъ��.k��OD;H�cCh��Ub�@l������r��SF7LE�#b�oc�u�i�I��f@Lm�i`.��������ٹ�/1� 1���>p�v5x-�͸��j�{���d�t=\v�����7���x�����"X�%��{�M�"X�%������dK��=���ND�,x�����j�19�\�|�~oq���b}���iȖ%�b{�{�ӑ,K�����iȖ%�b_w��ӐlKG��yy��D�JM8�W�R�����"X�%��;�fӑ,��Dȗ����ӑ,K�ｿ��Kı=��✺�d�3Y3.��m9ĳ�BD�^��ͧ"X�%����m9ı,O���m9İlO}�p����Gԏ�V���A�PO�9B���r%�bX��ﵴ�Kı>�w��Kı=���iȖ%�b~��ٴ�Kı?�?۾�/��Y�˭R蠵�9ۢ��ד�klqfv�z�n�U�,�aca0�/�$�'Drs���#�Gԏ�}���ND�,K���M�"X�%��;�f��F~��,K��fӑ,K�q�����h+��l7|�~oq���?{���r�������K�﹛ND�,K�w�ͧ"X�%��{�ND�,K��w�E�Z���i�fkSiȖ%�b~��ٴ�Kı;�wٴ�Kı>�}�iȖ%�b~�w��Kı/���
fM\5th���k6��bX�'s��6��bX�'��m9ı,O�{~�ND�,K�w����7���{�����ﺪ��X����bX�'��m9ı,?�������~�bX�'�����r%�bX�f=����D�&1��{iU�B\E@q\�k�ZLZ$�I�K�)s�j<>�.�Zh㭆'����,j�F���7���{����o�m9ı,O��{6��bX�'��}��'�ı;�p�r%�gԏ���W����$i���\>�}J%��;�fӑ,K��>�iȖ%�b}���ӑ,K������K�R>���"qGN���BH����#�,O���6��bX�'��m9Ǌ.u�R(A��~U�{��~��o}�ND�,K��{6��bX�%�a\�ڒ�]Y�f�Y��K��BD����r%�bX�w��iȖ%�b~��ٴ�Kı>ϻ��r%��oq���sQ�r�-�����2X�'ｿM�"X�%��;�fӑ,K��>�iȖ%�b}���ӑ,��ow���~���y{6���;k8��.{��'kW��,�5����:wm���Ӹ�.�Y�E˭M�"X�%��;�fӑ)0���j�����>A��i`cڊ�5�BrG`uw5߾�ꤌݞ,秋�7]����9 ㉷)7��o`��M����_9�Izݥ�p���q���vi`qf�:��A���}T}U]�uA�����aND����,�vWs]��ɥ�ν�`r��:u���J�)A��ha]g��@�,��ĺ+vg[��wW���,�N)B�I����`w2i`s�uXY���E/�6mDF�;�����& :��@̻�k�SpJ��8���,�vy,Y�vn���[Q�rO�(�v��qՁ��2�f&!v��X�n�N
��S�9#�1w5�̚X[��,�vUtu��4����N�ڶ̴����D�a����Y�x�{�݋�l�7�q��v�a�°��/��
��U5\'b[k���:9���XE�`<��8 ���u�5>\ƒ���u�i�"4�n����	c�#C&�-�髇n�t�`_n54�7��j���Ҡn�[�X8X3մ�s��Rέ��U��Jp\�4MqjՇs�-����\.Իj������w{V>`M��XY+��\tZ�sKe1˥W\s���^��������6�8�H�m�M�$}7'��9�[���@wIy�����wj��sD�9�[���@s{���7<�&�6&�I������y���@s{�9��T^��iYy�^��|� 9�����n�����F�M�j�#�;�4@z㘀��1 ��ꪯ����yG�8+��.0��u�d��=��!=e�v���e�炜e�ҒPl\�b���~��Ɉ�s�� s�[Q�#r?�'Vn�T��|J�Ā� � nj����}��7$�vi`;���8:j)N�����:�;��,������x�1o�V]�Mq��'I�����f�XܚXY��]�v{��e��l	%&���G�@~����x	n~�7 =\ɔ��g˙�s�����a�z����8��BGg�[s�g����r�&Ss@�6��Ɉ�s�T��M��jd@8SnRL�;�����Fn����zx�8�u����q�ڢkY�'����9ߵٹ���"�H�� h�PH? ��"�(<����:�5�洵� �)�%9V3������j���:�;��,��cm�9ΐ�,,�v.�7 =�0&nnnN�#1Cp7Mm���7n��;r=.��ج�mV�[������.[n��*(�:�>�7� 9����[��B�o+tq�)7���۫�z��<�@;��VWqO���m�Ѱ$��rJ�;��<���r��T��.j��mT�7"p�����Vq�ͺ@�ꯙ�|���{��-.�@7J�ͫ��ݴ��7 =�`�������릮8�nP�$i�H��s�G����� ���psqٲ&:��R4r�~x�YӾ뀣�6���o�����ri`qf��}��}�ǾV��iy� ۈ�q�� <���rb��7 �-֓q��B�!�XY��c�Vs6���d��:w5�t�r�	�� <��@sqR��/�~���|P��C�N�RH��mՁ�������`s�uX_V<z8�u$Q��B��Q��7Cb��x�-�v�'($Ч/<���ۣv�g�v��Fa�wT� 9�K k�7�7?>|L٠����ew;5m)l5��l�A��\���틮�x��mksx�W����k{9 q�O�8��j�.�u�����ZB��`}��`7Zx���)+�(�=�t�T�e$�渰�Y�^�N-s����+���I��Y}�ww�{�=|;����;�⃮'vҮy���u���6ɘ�E��&�w1�@�m4�G�l	%&����O7Vݦ����~v�������P+䔕9m��`qf�9׺��mՁ����}_U|����&O�J�IBH��n�3ś����,^���o��-�ێ6����ͺ�;ܚX[��u�Q���ԍ7Q9N�i��\����� ����~�g��^^�M��gv��3v^t�i5���؞{�
��TpN^�*��6��nm�=rL@s�- ۊ��K@;�]:n��G*P���Y��9��[�2�&a�g�7�or���S�`|�u`qw4�����$�����VVI�\�nL@zK���>��wiUW9Ȱ��)�}�1?yU�՘���ͺ�7��t+�T�I�'��y�@u�1��y%�:I���������⮐��å�3ݸ7^I\�k� ݆L(ܶZ�T�_}�-��k�z��6?0;�� #qR�$��p��e�J[�m�����ͺ�9�uXך+�3]��5�'�(�iʉʰ;��V���N��}�ҕ�t�$�|Y��D�@�c��Z�YL(ibF$�h�t6m�FT� ��MD���!���2�#!2�0����!L�b�� ���I$cA�T$��c!��$7�nB�S�4䐐�6 UWh�|�(�\�.��x�|%WzD/Pz�"���V�GR����nI߾���9z[�X��M8����`o^h���v�mՇ�]��+ �<�y�U��R���b�Ɉ�T��Z�1�[Q�(�C�$�0��J�2����D��`��s3�sv);k�ם�4��zٲ�f.IW9ʰ31�X�mX'��Lǣ�{��`g���vG��Rm�*��=�~H���X��X��,�eB�|
b��bqXך+�7]��-��Ձ���`n榮�'�RHr�#��:���3��X�mXv&bf*"$��c>��>�=;}���R�R~�Q��S�`gs��=3����;��+�����O>^߽����Ьj�1¤�*e��ۦkM�3��\6G����7�*q�eNTR5�����XY��̚X�P�[N��܍S$����_�H��j��>i`w)�{2�i�B�S#N2T��"V-�������U}U�%���`f?xVr�p��"���wq���K@>{.�nL@s5jv9>�u��rJ�;�uX��z��b{�`fc��2>�%�D

���22�[T��4�U�C7�Ņ�j�ۛ��[=���8�ױ�p&��8���m�q�d�I، *4ـ��#ٱ�٩l���CuԻkZ��^��Fwa�J9;1kݡ�b퍱=��7b�A��,zݞ��h��s�לmL�똍��wm��V�.�=�������k!�@�OOI�m����-�?����+�Ơ�hz��N�A�����������wy~'̖'X��`�<S���k���8h�a	]m����ՙ���gs�dI�'��l���՛���d���=�`ff���'�RHr�$����vn*@s�-�U�#wv�y,N4�j%#�33n���V7&�`uf��j���!��NQ$,?���7U�׼�VV7Vw8��(!`m
A�$T�"�9�5��7]��ɥ��{����/�Ԥ���Tk@#����]�k���{)�DBj�{�������ӌ�(MH��՛�������Skfb~��$A��jVV8�\P����n�nkZ��>���7�ȮBP�13����Vo���ՍՁ�թێT"��ۑ���=�`s7����Kݫ���:����Es�UP���bbf=3Y��Ԭ�ޫ;�K��U�n��)��9D$ܴ[����$���v��߿�_'�eKP�yn�m��2�]r72�`rݤ�f�.-�w1�6؏�����~di���͞,��V7f�`uf��j���!��NQ���U����H��m+ݫ;���f&R5Ң�שR�i�2H�����:�u��u=R�	!2@ ���è��;j��g=�rN���nI>�����������}�[���=��Ձ�s]���c�8����D��
RY���	T�w�L�q 8�ߧ�����ă�B�z�gd��R�эlc��\��J��`�MX�u>E���3\��Y������w�L�q 8�${����`�s�ND�i8��ݎ�1	׼�7_4�1�5{3�kz5 (��	�)�#��zX�4�;�5X׻���i�M8�M�U�Xj�w���OU��M�c�SIT *�(oy�krI�om��;!���ʊB���`w^�v��,ܚXTuf�8))�jTI�c��1�'w �5�x->�賄8yř��V#'n�MI#�I��{��nl�7�4�3^j�;�-7)�N9�8�'M��r�d��_:�[�����nK{�K5�=UUU�[��G`b�y��n�l�$r�n8XǺ��ݎ����a���{=~,f����R9m��`f�����{����,�6��=�LDTC � b)Зل�$��2�i�QF��<��d�=z����f��d��n���(�ם(���ŉۖ;rH�c���LUAŨ���u�Y9wR�5��b{P������9���[�ۙvon����;��'aa3�sq��.:���{�|�>|��:a�=x��lj��c �(0ZC>GU
�۫����52K�u��eJ.�F��n��<GcfۅK�f� ��f�p��3Z�h�Il�ήÓn%�fb[����������;����QH�$£��܏ ����������=���7�ގ���P��i��ۉH���/�U�|����`o���՛��;�[e:zr'(�U��rZ̓q �Ih	�*@7�EI�h�I$NT$���{���uX��Vu� �߱h ���E8�vy%�'H����&�<.]�߼8]`fck�:h灁��S��^n�����Z�M��7N�LlC=="]���5ZG :c���n =nL@{��wj��q�i�%XY��)}��Urf&ap�V�VW[��w�1���`��E!Sq��v����Y��ܚXY��s6
H1&$I���,�v�M,��v���{g�݁��*�����mD�v�v���	2L����ﾪ��n^h1]4�{P�v�9'����c��ۢw.��mcn�㒝��	yyn3��U����䙈_I��a��#��u�9$�H9M)1�P\�v�*@w=� 㾗�o6̭��UX.�Vw8�BQ3*�UT���͜,u�`b�V��H:�j��wq ���`���3����N��rIM��,�M,�����n�|Sݫ;�e���eTS�p�G#�{O6��kg�uk\aOc�/nY��nb�J{��v���+��0y䙈[��������$I�G)&7�8�u�ܚXǚ�c�n���URG�P�ROȍF�n%#�76x�9�5XǺ݁ř��;�[��������HXǚ��6���f:��ى���b&6o^��k=䑺�JN�Vn�`qc��|�<r�al3ae�XK��һl�bI�tΝ�Vl�[.�_]O�ol'�T�8����Y���q��X����G�V�*�Ŏ6�Ñ%E�$��������{�`n?z;�3]�����?��0rRj7���q�nb�� #s�Ӧ*r$�JG`g^�vf�;�K�3]��ݷ%HP�)IB܍�nb�� =m�@>�7�}|���p4G%Ԥ$V�0#
�V4cw���~ m/XD������+D!&���������i!44�!�ا-�2��4#�̡Zڭ��aLՔR�-�P��� Ck��^�hCqA�VŤ]�jD���B��2BB$bH��!���JBĄ
��#��|P�p�H
:R	��S��$)e�]?��ܿj�0M;� z�Z�ۃ-�ݹ�t5���7��T�v��O-vz�I��`  x�����MK��k�<��a"���T2=&E���.��N�2���$�ڪ�4[&��%Xx�z��^:��9�&�ݪ�NPb6�/k�<��2J�p�e��a��{h�����ʦ3�ls��sɯV��͇�n��<!�k��ⷊt�[B�E�q���ZGPm�\jxϷhv�����@��XD4pV���&����2��GV��C�+�;v�j��j	�;*�ͪmR�R:ŝm3\�8��.�Uq�܀׀��ڮ�y�C^���-@���H��N��_�ʭ�@m��'��R��n�mf +Lئ^�Y+E�V�gWi�Iq@,���geO�|���@�:i{�n� 
�ꪔ�8L�;<�J�F��9�3J8GL��i[�������z��	E:*N���$����* �7F�{mv��*�s֐c[-���=�/l�d������.�۶|B������].1v݁z�(.��l�{۝ѷKc=�y�Dk���������l�ӗ�S�w'0��ͧX��L fw;�k&㴆��6�����ێ8�nH�m��v���mv�������m�k�@mՃ��d��m�Z�^n��)<�&ɊRZ�U�;���\�ӕmV��W[7M�n���P,�<�F$���`�Ϗi	�C�e�7\�m�Z�MoY�mmJH��m 4� *�s�v��iX�;!ݱ������V%�.�gSr�Vӧ>~*�W����:�<���Bڐ�B]<�. �ӥ�.6i9.�ѳ�,z.�cx�RV���m�"%���ڭ�p$Jkp�GI�,������UA�ǔ���p�(�)3�u��l& 4�\3�wc�M&��Rޝ��Z��� "��-2�*�����[UU������s��2��]uA<��Ƶ�%�a;l�<��� r�8�T�EJ��W���(Y�o{��߽��w��L8� �
 O*&�ۢ��
�  �:x���M �|��u�=�i���&R�:,��Rz�n��[$d�m��W�����%Z�JLm�+�g�eLVu�F��u[����Xۊ��ӝ�8�;MT�l�qP[]*����C+�;��s�o_Z��|p-뎞'h�q)�ء�yD�˝�N��ӥ��f9��WDۮmqsu�G[��f�FG� �
��I:�Az	-]�#zMۭȠ�H�*�$�U�Օʷ�M�r�%��r�l���惃|2��&�A��s�.����n�ӓF�dU��ʹ�����1 �$�@zۘ�9����I����HXY���ݎ����`gri���䎣�{Ѝ�I%'L��~�����1 ��o`�şj��"'QN9�ř�������ri`g^�v.�kC�IQD�	8�3�4�=����7������m�?��~�VC�����Aу\c�펂ܛ[��Ґ�3����j��i���7k���{�q��1 ��,��	5h�ȓn':�c�C��h�@�@ D1D�b#���\ߪ���`}��/b!#��n9I6Rp6�vVo���ɥ�����ν�����ƙ"m�%�U����k߼X�<X'�*��14���v���/H(I)���;װ@z㕈_I��`�l�ef^�vϝ��l٪ۊ��`�-�2#�u��ں�eg���v݆�	L�3/K��y
� �6ʰ>]n��q�1? �|��յ�Sm��@8�����~��������X��X&�W���8�G	RTQ)BNH�͞,�M,�WO��s؉��[zU���j��F���O+���Xn�<r��*b���ni`osX:N�B�"M�H�-�����@y㖀w&\��/K��p�X�c�@��>�����]����l	����*��K"�Ȼ��2���o[s8��Z\���wtT���D�mD�v�mՁ�y��ջ��8�5�qkj�ڔ��JNTrR���!�[s8��%n�M�)N87L�+V�����d���ٹ5�S��Q�-3[���պ*�I����(n����`H��9h	rCS�jVѻ�Kv���;��9Px�>ݘ����ޡ]{c���,��uJJ$JRI����u`q㖀�$1�nb��/�ۆ���RJ�9�5_��#������;w6����hv9m�E`j�Ҭ�c�6"bR�{q`u�i`6��*ARM��)�`qfk�7sn�fM,[�;�5R�&����ډ=��*@{��.9X�����������~��ꝅX�UY�*��jVr�ʑ/PuNn��<N��wi\L_S��n"#G��s�S!��3v{�{9�8�b�ݎ��H\�F6���w+���y�#;2m=;(5�'��u\L����9�6w@SӁ��e����L���|����p��td�LFF�z��\��x)5�	��e��X�]����̍���@�X���t��{������ǟ.ߜ����u���^�k�s{&�d#���o�>%+�-��U���v����G%x���,[�N���k�7sn�?�R�=���"�ԉ�������U���GV=���Ł�s����Hk4U�QH%JP8�`uf����V:�U��si����$�H�����@8�����b�W�W�}�|����܏�`��)%X��V�!�_9�T�ur�]^C7(�b.vm��O-v[˞-�N9�t�O�*7<����'d���s@���m�?d1��1 ㊐�� �e�m�4�M���pv1櫕_| �ͺ�:���[�;�5R���`�ۉs�`c�q`}��Y�1	5��Xt����-r���#�rJ�9�5X� <��@8���&mfi��+���9\V&�V�L�������V1�;��MM�NRt���T."� �.�iM�!{�'Q��r�UƮ׺sñb�ѹQ4�(n��<�`f��Xǚ�[�;��Z�Q�4�$�{hT���- �Hb��q�m��8��LRJ�9ܚX�tw?"`�V,Ep���j"	"&	���uV:�[��c�HwC)S�&�N-��`qw5���V�w6�X�yZj'Cl��Hyy[�_9��T��=��J����_��W��۝h�f5-�۰7kDӮ�ѭm;��v��J���{V����m ܊��@u�S?}U^�����;�~m�R18���*��ri{1)�cj��S�`f7q`|���t�J�����ν�V:�U����X�M,]�V��(N��RIJ�fbs�U��������XlF
fW�,"���P9��ߋ�'�ߏ\ɬ�����+�ͺ�9ܚXܛ�μ�`b�i�lB�Rl��t�I��3�Tv��\�î�iV�Ӓ+sǴ���X��-#��9)��V3&�w&�`sj�;�۫s5�MZ*p��G�ٶ���-��H7�_���'�y[j&4�M��I$Vu�ͺ�9�4�;ܛ��֪Dc��I@y�^�9���{sٶ���}UT��|����ܤIC�A9%X�q��_��:��X�w����{۽�������.�N�Y�Yj�RcUl���T#/��:P���j���<jF�	5�<Kc��1���bړ��Ol���T�W+۶ӭt[tK:w\���gs+���k]�v�w�Ϯݹy觚����-�]���$d��-h������&�VlN����8ұ�����K�ь��\��t�К�N�<W''9������]]�ꬮr�+�I9)��t�lb�T`�Ӽ���xb}�\F�ue�/8�;����m=9���%!`o^�Vs]��ͺ�9ܚX]�]�(lR�H�.��7 =$T���@z���4��sKڻ���@sqR�EH<p�,�v�խ܎�N@�S��l��x�hm�@sqRt�f^]�b��mIV1��ř���f�XݚX�W�U}ڕ�t�z�9HK��su.�gk��3۪-�]:ҎӵH��A�㴹�5�4�L��$�����]XǄ����9�T��KX���5n���~�����O�G�7��y�Ł��E`b��`��I'E �t��@zM��- �n*@qn���u*P�m1���E`b��`w3n�=�.���X��N�F�@lr�H�Y��Wٛ�W ��V:�E`n1bI:�L��GT2#�m1�����i֗���nx����.ٺw�cb�Π�QAJI8�;�۫��u`s�4^��5f�����ۓ�ڔ))��HG =��h|� ;�T���썈T�M�*��^h�]�w;Әi�w_�N��h�H"�,"� H�)�~៤�?�/�Ȑ$
VR�b,H�2]�����H,���$	$�Z� �c1��&d��$�@"	�B"��C� �G	��J$�0D$ �L�'���B4��P��`��<$�f��r$�B֒!�������!�21��ҡ��T1S���Ƶ�7�@ D/�!�>a�.F�����arDy�M��uZ\P��%�H����@p��D���qwpИ��hu�>S�L!�f�~��1 M?�TVҔ��"F�G��#Ǐ�^���6~L;�tmhh�Q��ȋ1P�;����5���s�7$���́��J�i4Sd�I$��y���q�X<w+�Ǣ�1ƨIr*+b�����m������p�u����4l�	ʉ��8:���N�;K �BW60���N�o\�ܧi��m[����NF����u`s�4Vc�^�꯸�3}u`u{��Q��J��5�Hv8Z�r��T���R��k��r��NP)���U��ͺ�9��V1����5S�F��+���@sqR��H<p�U_���$$D� �E�~D�o;�=���'�
9LrJ�9��V2���̬j��c��6f��TUB�Rkp>�i���g6�\㸹�<���z���aY�N���W�����?_߸�ecVs�����q`=�E󊐕EG�9�X��^��L�F7�}�]Xǚ+�RGv��%)����/v�Oʐ�*@yㅠ�- nk{$�q�)��a��{ܫ����䖀��\�2��+kn�w74/6�x�h<���T���*�꺯���GԱ֋[dPpRD�vn�=���ح�W\�9vKW7��#o13:rj�x^m�#�l�n�`��mմڛt�j.�RA���W �٤�yut9��c��#�n��3�ƹ�Y���=���U��c��[K�کCewaJk^���ur��Á���״�&E�ٵ�	[�2���6�1���o��㫝uJ�R�4��{:�e�힬�m��tl(AK�[Q�����{�c�r�v�-�Tl9p�Z�'Jλ#Axseۮz�盩�-����(�ʃM9@�p]:��`w3n��M?}\A�{�X�O&Q#r����ݴ7 ;�������~��#�yy[�}Q(�1�*�������d����re]fR۩*&�N1���^�;��V{�K7u"���"*I �vIhn*@w=��-9̬�Gpᴥ�'r�Ns��|�2�F��\g��+�7�uبK'sͳ�A,[~��R��x�hvIh=m�1E �����&��WO���?AEz9����.䟾ϻw$��ݺ�:�C]Jn�D��8%!`sh�_I�n*@w=�[u�@���//6��sK@z�L@sqR��ǚ+p�L	�!:I9#�;��,�q��1�`|���=32�!�W2�D�Eev!n[E��ۍ�vM��V���Ir��$l�U^�M79�� �����1�rb����tRv�m���i��`qfh�.�7 ;����w�Y��ه9\�V˭Ձ��qe���?LN����4O������>�}雒}��$�!�2������7 ;��@zۆ 8���s[od��QH' ���j�ٙ�7�|VnՁ��q`f��o�l�ڃ�e��\��.۪Ѯ��Zu�/Ot�l4pJ.ť�H3.�[p��Ɉn*@s�--�l7 �NP'�ś���f�Xǚ�,������T�%D��w���'�H�� =m��& 7��W$�E%89HrJ�;�5XY�fnI��{����
~����X��Ch�M���i�#�8�4v���|7�WqՁ�13������b� �� e�v.N�4lqqv�&���\=:��e:�(-�Mˣ:�A������ͺ�:����Wun�vt�BR�~	Q4�"�;��VWqՁ��eXv�W�130�kڪ�M�!"�NA�Vc�+�3Gg�K�=�`fﮬ��Z9%'���J��]����7j��c��;�ƬY��N��&�r�8��.���R�����*���UW�F]8S�Z�1�Yy�ow�;Z%*Q�{T�ߗ}�Y���J�']]W^�|�7��G���:Z@x�@��t`nY���(�����<�#�a�E�m'H;]��9'I�R��YI�#��Μ�5�����[��j
8�td��z��^�L@��m���Ӱ<�ƫgp܄�%�)K����-�GWZk#5��n��my��4<g6H{����������������w~��k�'�������^�d�;y��íڥ����-�a�s�c@Uw{�����T��{��b�=�"�9��\��	)��I8�X̚X��[��T��L�̱�eniy�nh���@y䖀��<�X���I6SdC$r��=�@sqR����9uue�+o.���m��H�@wc��u��}^���l��RT��$Nnz�N݌�#ZzN[ct�ZK���|"27sQ^�[�p���u*)���7_�+�y��]���3w�V/x^�R�i�+���s������RLvfg�qSu`w3n��M,Y��cR8FҔ	ǥ�=nL@sqR�� <����ؓ"MFF����;��u`w2i`sh�,�v7V�q�! �R�y�����7���rb���o���C�v�Lp�g�HC^����� �/oN�#�IuոV�������ʑ�W�י��sٖ���-��Hoa`nb�Te	��8��Ձ�{����7�@{�̴�]]]�e������X�۫��K3����&�`qf��m�C[P�H'��v9hsٖ�����9���.�5I�)LQ�`s�5�����;��`w��X30�T��*��*��m�l�X,��m�g��`��/W�d�RqN/t�T�7jI �(�k�ug����,����E`n�ؓ"MFF����; �f��Fc�+��°8���n�V�E �R�'$�;ך�x�h_I����rK��lun7���֬.� �se�����=���&"t]�U���(�φ�J�F�j����`�l�;�5X̚Ձ������o��)6�7��m�f&�-��a�uې�gN΢̕5M7�e,��M���1�(pi�D�| ��K��U��ɭ{�:��v��:l<�IN�,��w�H���VV���;��`un�I�)8ґDȜv3&�@zܘ��qR����e陻y�Y�f�Z��b��H�sǚ݁��bo��"�R�����;�lNe�]��\���`~��b&a_�Q_��EW��EV��*��"�����"��؊"��"
�����
�`**��
���",��H* �",��0 *�"Ȋ��"�� ** �",��)�"����EU��EW�(��DUx�*��"���Ȋ"���(����*��"����EW��"����e5��+� �� �s2}p3��%TРS*�M Ѡ�T�!E   4� R@h[�6j����"�
�*T�@I(�*�    $
P H �  �T
��QJ
�T�%P�IJ��J��   @ P  Pc �R�U/��=c�=kqn� ݵ.m�soV�E�s�X (}����}�{| ��&��rz�������8�T��|F��]z�jz��}�꩗�=ܯ6�MϷ_mo6�_ ��  � P +4{�*ͮZ��n�Z�MW[�UO�ЯzQc>���^��#U��� =}�p�2�X F���5� ���y����ɯ^�6UX�*� zou���uJ�ܾoO,��rj�x�  )@
 �q�4�}�ҹ5����\����/t�� 4��ws������i{��a�\@�>�Rͻi:};� ]^/9�}���� >��}2����x���+��o)_8 -����t���V�N�p �   �   +�� )�ӗ}5;������
R�)JR��R���)M���)��(,���,CG4���E)M�t���,������(� l�)K,����R�)c4���R�Z�t7)JR�iJQ�)JQ��(� ( 0  �P� �� cJR���)sP&���lz}x�3ו�n�9e�5ͥ�����`��������π  >��i{���Ҹ� =�˛}�\��N[ٽ�Ņ�} >�zK�.����r�ɩ���=7�S�&�Om)R�  E?�e3U)P  Ǫ�*�0�i�=��Hښ� �OД�Ҥ� �	�R�D 4x�?������p���vw��G�7��EQU�g4��
���QAU?������*���TU`(������p#HD�@ �$	 �ЍHBI����N���Д�hPÖ	C
f T�X�R0�J)J��g�,e1K���
C<�4�.7�4fy�%$dH���4���@�aS�e� ����!�b��u��ĨÈ�
|s ���2�1��^K���r�PCD)�����9F��r,�>��뽆�9������H�#d�S�
cw�� RD�"I3Mw%D� ��(d@b�s1�#��yF�L�?4�D�V�2�ɜ"I�EɒH�%�������2&��9�4?�߆�����T���������K�O�3צ����K�\��U=���Q��NL�[ιCO�x�����wL�ַ��Mf+a$L&F%��I&	��2�?P�!B[M\��Ǡ��N� �HK��6gp�^�.��`%YLo[/oN���ǝޗ��[�dx��2�K"��/�ӍK�>���7h&)A�A���Iq���9��s[����n�ʺ���[׮���^=ý�5��P�B��"A��3�.����3a�����D/�3[��L0��}��S��s��׬)�:ݚ�ޙ��]̝泞n!GuG�/��������ʢ�BR�мO۞t�!q���@HX%Ƹt�;����q�"l4 n@�Q�~���y�#NHC<�FX$H�r)��.l������!�|f��'&��L���K�	$`?0	�R�s����e�)^�1�u,~�;U���/�T�t�X��b`ֵ]Y�����L!��>0HB��1+��f6l�Ά�\Hr�bh?!?�|�rp'�'CBgӉ>@�K��\Hr�D�ɨBYD��4���I>I��>?Z�>b���}ƓJrdg>ʟ��	fRYt�º�aI.����j^\|3�V�cb��ƗQV:�e�Qf�<�j��FW�+rl�ƍˍ0�lN��$1���Tr!,&��d6F��
G�B�$	A�F�# �LA����$����!FP�\��h�n�!'\n1tF0+�JĒ�H}�:aoP�	�[�2�hѦ:�Yu�ϭ�k�U�V<ʢX��K��8�ϔ_D80b��V��� ��L2�ƍ��hu
���c?��\����^+�=k3�(���Ҷ-��}e�ɝi!G$l��Ñ6|��D$k����R��ɭ1\����9��3���`������!VG2&��f��d�y� ��@�+�# ��`Q�0�ɯ�I��p�F�0F��>`C/и��RM�}\�C����3�4"LL��Fp>-�9�j��j��~�o%�XL��=���C�]�0A���NZC}.~�w��95�k�l]@�iƙ$�4�jK�����h�@	(*��^S�ǲ|^9ꢯ�3+{��-�\G��Fg:I\�e&��b2��!��wz�����0 �H0�c��"�5z|K���'{��B�~��I�b�e IO���Hg�SE����Ыի�.�hA��N��d�`\�4K��4BS��1�CD��b1��4�7@��.L��Ҷ��i\�����{�tڝ]��>��! �~	s�_=#��3s�w�,�3�T��!{N��ʣ羫��mY��z��S$\����B�(g3~.���)��[	q3��HR)FU$�SZ�h�L��� �B��B��B	�|��oS��|��}���s�XR��B��8)	��}>�A
`����ha���ц2��F@X�H��!+��5�1(���ψ}v�E�q���]z�S��_w2���s3�^�E�"�:�Qx���d#��ۍMk��X�Ĝ���Ah+F ����y��|�t����#�	���US�@U]VW�-H��D��,����{�gF��
w[zSS�5$���
�!��J`I�l�cB7!	\���! ��o�XR:��%2JbP�YYt��F�C%�]������U�6�Sw������A��X!q�\>��y,6�*�JDbD�U�)�Fd��w���Da�8��C�aB5�HAL"��E�)c;�	�gP%4i�Ƶ60���5K�AO[_�\�I �%�O�b|���-���±�~��$�$��>���O�5�ʩƧ���Cm�k��f��,��E��]�%4"�9��T.vUs�ʷ��,����P��滸b\�3z���Ƹ
�7�|;۽>�Ik)��eɬh��v�E���~XO�gSF�SAR�B @�eaw��2�*p��N*�÷�j�bj$�5șa]b��,��5��%q"Ƭ��7�+�% L$�SK��H|�8�_��RP�\d1�u�Q	Ȅ�HMA4�GC�f����K۷�ᷘd��Z$�@���tˍs��l��0B @��F"���4�)��i�j��E�0��r�!��y���Z~��L$F'S��!L�"R5�Y̟}�v���p����:����|�HS!�"�A��շ����%�����3�,i���bG���ә�dlR�B�91H���pa�����'�w6}��n�\\�%2M!���f���韦�Y#'��~]w�Y�m�]~�#���|��rr���!��o	����~��r�0b�M�᭘�(l�4����JL��X��97���Σ�;y���ӎl�7��IL��87�&Ǉ>7�5�a3��=�0��a��0���%����v�D�8�D�"�b� A��`P�!R,	 �I���b1�#$�E$$ �h.1�˟���F)`�2YY$HI1
�B`aq�x]�ϴ��\EB�R2����S4���@�A��J$+�Y6	�M������^��*=��|��"�*誨H"Dd$		��/�λ2�i�͚��H@�b	$`�X�V�!"�(ń�`b�3�u�t%O�B�0`1�"���
Ʀu�5�s��s��Ƹ}
�g[��1��8�*ĥ7�}����p)�BHP˃4�����郠���!�D�qM�.t��&�c�yj;������O_�X��NW��q�T��"5�H�)K����&�������I�d�s�!���T،Z� ��9�;� d �&��K�\m��	Cex�)��B�	���[�ے��`X������"�@  Y�#I�����H��)## Yxc�p�22@���(F�,+�����ЅH��u�M���.&cB5!$2C䅆0bŃ$�0��ی�<H�4"�#B50E((Bgs�CΦ����`�d Dt��X�y Bk$Hr�fd�ә5���F��a|!�%�e�d���Ɛ� L��!�&�����ʦ������f����1� Q�$rO��a;>�>�tR���$�?]2c:xCY��:d�7���q�M}{��I�T�2b��"�����
�����bi�
1+����
��%p�K��L�[p��D�,a,&ZP���Q8��B"�1Fg9��!#��f	 O>�U��bpn\+ D��c����gS��y����l��!!,(Bcp��!����:��a	��B6P�	cLXW B�1��	YD�F%0ƎP�
aI4Į\e#d��FBHыB6LK����nX���T�������P諭��+��Yk���䆉q�s8e�q4�k�aL,
%��b1���ܟR�R6��s[����@8��~��ʑ��3�NH�3&KB�0��ڼ�Z�3|���BU��^�z�q�,�Sfp�b�3���8���Ed��M�ĉ� T"�D $ � Յ�Z�����#\,B�X�t�1�dY�	%�� $�X����H�.P���%2d!
`X� ��Ҍ�ǽ��Oյ�V�eo�����}�	V���wgI l�pP��!HX�R��
�:�7��82�R|0#�[����/�6`)��]�gf~~�1�I Db�j@���FH��Ą ��1LR��ܸ˨\e0f$h�`��ab�a0��%VP�$�!Hf4!d!L,
a�WHT�B Dp� r�N�E�s�~HN�

���v�g�x��75Ԭ�U�U�T~.�TU��G�|f��i'ox���JK�q��y~�}xa&S!)�!I���Q�k,�(����X}
�MG����`�q�4�0Fe����96�q��UOt�e|QB����x���nk���Fg�{U_��_�U�=�N�����	ߨ���3��v�m��m���           [@   䃀��o��`  m�       �[@  �` 	�Ѷ� k� m����    p �ִe���7cm��k�i�,
��T��N��[@p[�}��}����Z�Ry�MP;,�q�`N��m�I!$�l'D�Ҁ�ifI檺��$ܵ�c`[��su�I95t��YiÇ����j��!z�p�$��-[@�b@6�kh   	8��v��w�j�����Ue� � ��Ã�o�Yx����ΡB����wOD�u��[uRA��R��t�������L�f�J�U<��kjC����Z5T�d�j�e�Vj��` 6�����RklIb2#]m����   [@-��ô��n li�m �`�a!��m�-�v��5� �@�-`�j-��� l    $  m�M�q�V� R�5E��Ԅ�Y�`Ƌh$�iZ�i$�ld�!R�]M�2J�R�WP  l��ؐ�`i0F, mU�I���j�i,�m#m� �` �f H�m�q�M��p?e���PFy'�1��[��Umm!;HMƑr�v�յ�+:6T	S=rT��`��6@檕��A�`�,�M��+m����  -�m� 	  ��q5��+�iI�l� h��ᵴ���T��v�!�L$�Ơj����'MggN)��KjmB:U��*�vU��N1̣UUMn�,���I�oi6e\�5�V�UER瑍\���S�[%��m�NX�R�i�dld���ӆaf�Q���e�S�q!Vw����죸���<�k#��M��C��e^��قc��@/.ͺ�j�!R���~W���N�e[u"���M�����檪  gi���t��6�:�mt4��qN�Zx�0���Bv`@&�KIuF���U�ݨ���T�PYw$%[�����E*�VԮ��qN�0lKëg���:���(ݫk��c��J����ҹ�]٪�"�2K6=��J�dc��q��kk��Uզ�f�`�\��@��x�@�&ac$*�ڻq:*�Cj]*��&��bS��2�]m]�UV��E�hEk��jM9ĒI�ͬ�n��v��0�m�r�.ٺ(	� F��u���`�ڪ��Uv�
�.ݸ�ds�@�  � mkm�[@��WKi��=c��m �u�2iӑ`�!�k�nհpKZZ�v$m�Hm�z���n����)PA��ͳUT�*5@\�,jg���  [@�cr����+��9���:)a:����  �Ip$�l6�]�')1t�T�@�UR� �0�ڐ�ZH

�j|�6WĵE�:�@$7E�Б���ltZ'D�n���   �   �$���σ���������jIgM��kN���  9��kn t�I�]��	'ڐ	�u���&�[n-�mn�i�v  �   �n� �`  ��  zA�-��\m�i66ض�h  �    [E��N�N�햀��  �֋��%�бvͻ;kn�CZ� �nm��z�kh k f�E�6�  ��Ͻ~�� ��m$ ٷ` �l5��h�M�m�m� [���b]tfH�J�`$�l�`�7T��m�p   m�V�$�pm� [@ m �m�����v��*& �   � � �  tmٶ� m��)���h ���s m� ,�JڜnZ͹gM��	�n�t��  �nĀ   ׫�R�X���sv��m��\9Ė�-��  I�ζ��m�"Ih�l�WR��U�p�f��Z��ٶ�P�0�++B�ҭ��;qz��\�� �-�9a�	tm�  H ��ִ�WZ�    �  Im   �clI8��|�����P�V��H�T�T�mm�M�u��d����`mݷc��� ���UF��r��m �� 9���(�  �m������� ��� [vqF�   Y\����k$hj��  ��H9�8k�0��u�5��!� n�[@�   ۶m�8�` ��� ��m�6r����m���h$  �� ��u�p2��%P �v�U��gb+�`��D@^j���m-��$�i =c��  -��;]��� ����Kh ��Z�
 Im���[@jh�f�u�k]��nH ��p#�js6N%j��F�uVճ� i�m�۲�[Z�m����`�   ����,��pm��¶�ZIҮ$�\ m&�Z����oi�Á�d��H+�cm�m��lh t��|$��.i%��:���кi1��g� rԒi��  ����$h����Nã�jc�"��M��p�u��6끶�`�IN�'#�/5V8<�ݱ��H��]$�Y��ap��Ò��a��l�v)06���\*�u��k�����z��L�T�;�檻=,#�jwk��u]<�%:�v!�l�,��7���B,kN�pa��.w��l]m�UM����ؼ�w{g�aR�
^�54�m!h��C#a�[�B�0=X.:���nm�v�e@�ַZ2U��=�� R���(m�\��b�H�U�[��h���f်��+���պz�8E�ch����.�ǃq(<��uO*�@n�#;llq	J:P�2;u��[W6^�^��%�@v[k�X�����p-����%�T�l �%t��6��#Uȴ�0#�����J�vÛI�ӥ��U^��]�(�U[Oh�ۍ [C�md΂�0N��-�������3�Z 	��2��m�p m��m�m�2�  6ٶ��[&��M��	;���Z�l^�r��`}�����[��$-��`k����
���p�,覭;S��;iUX�@���v�M�#���\ݥ��9:V�Y� $�N���.6蓦��G� �V�F��kn� ��e�
�Ξ{kmɫ6P��BX����G^iv.�����a�;U�H����}�6͛` 	$�`[@H�N�ɇ[�e�'&�m�6�։�]��  �v�k,�� $u��H��ے�UR��7>� #M�[����eU�j�(9����Ih
Uڪ�ssmJ�[WX�EjU��{Mu   �[v��8���6]nmd�m��-��"ڇ6�-�m[ �Ű媀j�T
Xy�4�դ�j�kh    � o��I$�~����> �J���]��V�U6�U��u��m�Wc�����Q��{x�ŵU���s3T��n���$Ia��vzI��cۻ'6�T�܍�ǂ��M���wH˔^vm�`*���V�F�)햨�Ͷsv��͏nj��	$�gm�ր���P,�ܻ-UUʲ�@T�ヒsvٶ�-��nNڽ���  ���n�[d�j���`   6�&�l!��Y�ӛv�F�L�ڶ8���(������   H�ڶ���.��]ط�d�B�:Z�6��g3�t�h
ͤVDNE��J�9��in*"e���t�Xd���LAm.�N
rM�Is��������_�Z�iV����ks��H8�q`I�*[��<i=�Ö��|v�|-�����8�r���@6��	  vV�����4ݗg����5�,3�f� 2n�m��ll�e�i�` %e����9��8Z�[l0h  -�  p,�����,:L�����6eZUVyG5�W+(��R�5KQ@ ���l�sn���U�j�e;>^I�F4�dgdE�p��G5,S�����+N���i6�m%}�A����<���u �W�k��  x�6��5Uj��3��g�uˠ� ��Z֑���j�mh��H2rAJ  l    8v�E�Xgm&��;d�%-U.v���<����K*@a@m�m-�V�H������l��V1ꪓ;���8��X����Z��Y�Z�"���cn$�i�$)%t�� �5�m���=[�ZX.����J���Uy)癕�٪�v��I�yy�-�v�&�V�|�-��J����������jl�m�!�7,���<��7�շ�u�[C��u[(�pS��gP�Υ��ש is�˹�m�Spm�a��:M��mA��B�{S�x�6����b�|�@U�]7gt� -����T9ع᳌b���e�v�vI ���� �   �t��	��$Kf��&8ɦ��f����8m��[5],�VIU�C���ޫ�ocK�v    k[m�mҮ SeSW2�T��ڠ)	"r�/Ie�a�YBB�5I���Sm��ٴN�gQ��e6~�;m�Ą������ cM��J A� ��8�&s���PUM
U@��4P�?����0
��h(�`�  @�A��b���M�f4T �
|�PQ�<S*
�]*|`4
�:҈dE
�Q�E
�"���B	  ��E�F��ix ��lM
n�"ߒ	�
��(iP��6.Aੴ|�@���M(.�~P���� e��l^�;P�D���t�H����QjlN��O����(ggZ��t�H�8u��b� Z�@4u�[�� �P�6�5 *���ͨv�A����s`�|��t��O�pQ8��O�K��6q�D,�"1+cAh
T�|�
���l6�]"��"<�����!0�'�5Q,��� h���P�A> �iК-UC@8��c�X��A�FC�S��P6�b)�	b�"�"� �  ",����AdA4���
�
U�A0 �苔0
�&D� ?�QUڏP�� �U�1X�A���"�V� 1 AX* H�oh��$V D�U�D�D�����w�n=۽��������U@jU����C����<܀�8�z�j���H��n�N$�]j80%�Pz�;#R�:�m 7������L(K@��TM �NY&eg�N��i]��` m���-:�M,��&�^��IIU]�p�(m��=��J�آ�v
�����m����sr��u����'vs�s�2I�OJޛC���lj�'I�Ր�l�#�Q�p�Ü<ix<�j���ƷZ���+]��1�<��ѭ��u�����4k�uUv���ѝ�<rxR|�\��R��iL�� j��}�)ɱ���86޶��-�.�e��pr!�T����%%�vl���v��9�+]N#7J�A��ĝ�%�����cm�݁�T��¦���uT�@U���J� ���+<��G��`
մ�W ���ك�8�(!����u5R��Ƈ,Ҩ����9U����͍j�EZ4*��:��.��v�<��R��Tڀ�M�V]�Ҳ�"��nCB1f;6��\�#��j8���vPS��tƦ�8���2��Z��mY\��1͌�=N�E���z덭�c�n�]�cRq�r���k��qv^�&�u�ue8���n�α�͐��)�*^�k7e���{&ck[fev�cf�$l8�iZF�F�CS��1���kG��j����/>J�AˬXx�@D�s����dI�Iuq�H*��ܖIQ��;:�[�a8��*�)Y2�0��UA�j�/mX�ݺ���u�$L��=�\�/F�^ԽIÝ�V�
�8%V������d����^�#)XY+�,�챁\���9:m@dkt��[�H��٪�.�sM�%�vW<�vӤ��Qj����Aw5�t�S�ն��n��5��F�p<%�r��&	����͊�۶I���U鲯/��˞ـ�ݶy�L<�gf��8�>��c�j��V:\��h�=�V��7N���Z �.�\$pD7j��d����iڛpg9�Kp)A��Co��ȼ|hU��0mUM�ڜ2���aj(/˕��n2L�c8�,�3������Ɏ.f�۞�[1�-�h�8��Z�w��;ڎ4s�ö������Xz�MHFGv賴�]u�Ki�w1g!�� �� 6W�+<u]FG��	mͻu�����u�π!p���g5���6�r+qm���t=�㈍�á[�����wF�l�]�vחֶct���.��uF�p�����߾��w��_#�]۷)۰*���N3�s�
�m˹�㗌8ݸ<�9"��u�yN�n� ?~�}�����8�a��ذ�D�ay!i,��	�z(0&�遽��hN�U���^]Z/1&�P`M��{�Q����?=g\�VB+\nZ��07��0	�z(0=eK���Y@�AJ�Sz)C ��0?wn���ŀ{�I/x��e�7#��.�x�UVƛm�
��Α{p�Q؍�vW	���Id9@vr�id��۾��P`M��z)Ckp:�	E���d����L��$.8�8����:�UV�[����R�����5�,UZ�; �0��� ��JΉ�wH�}}��ı$	*�)^*`l�P�6tL��~���{�{�k�]����,���ݶgd�zF������3�T��]3�Al:mή=�ٷ\0c�́藈K�������ۧp�v�`\'s�������dR�;�`k����X'`9m�7��,�ۨ��v��ݹ�&��^���e��,mWj�7}|� ��n��ū��$Q�E�* � $�q�sn����>�����RF�T0	�z(0&�遽���^�Մ(2��ˬ��X�ފ	�:`oE(`�&[��JK.��G��[�h-mS˴�p��i��ٮ�n���5˹��-��搲��o���~t�ފP�'tL�����.�����B*�X���g�K��{��﯌n��>�E�]�E��l�3%�&K�7�%U���gf� ?-}�7[n�8Ӥ��{�L�GL	�ж>*�>���ﲽu�U��mˀu��)6��V���`��L	��SVI��p`j[�7k�d7�Wi�7^�ɺ#e㋓UX,L�G��`��r��� E�ۅ�K�n�!�]���T���u�2\$i��"�GD�i\����0�n��0&�l��� �t�]e_n���˃d�3W*�;5Ss�i����cR�:�;�0<���w�,�d�V���-���	r�%�a����2��nt�`zgK`zr�����}��}�U>�f�Yv���-Ә�猚�lp$sW����v����;,/Tl���;q^vS�d���Z�s��nw>��9���d��\)�X�T��"[�&�I�fm�:�$K�e�f���3c��9���.�ϛ�~����]��n��8�㎆q�h����9t���x���j��m9��������̒���3���]<s���i9q�-.pǳ� :��_׻��mqrv��=�T]�{a��x ���nm�<qk��
8�0ƫ�]��gE)+Q��W\v��7Ӿx߶����遻�*���eڻ�J�ˢ��v��$i��*�ɭ02vj�3�p���ͅuE(�ܯ �۸�nt�`:&�����U�-Kcj�VK�Iqs��������\���0'u�a�����/,���`{yA��#��)v��k�G�pV�;T�㊦2A�dnt��\����OI���ή�|�<�N˺ݶ{%�Yy���ދ��ݑ������U|������ ���h:ܕ;-5$���F��!!������fB�f�%�K�0���x�>����.�������3͝~{<�갎[T2�����[ے[��ގ���`T^I]nK��$�N�с�ၻ��Ӕ�`������V^]��X���w���)����ݘ_"*MDF4�ɵ<3f^�晖�c�Ƴ��{��/��6�U�����+,�aW���GLNS-���1����0���#[#�R�ڮՀ}�s����f�X�z0=�0$�UQ�v5j���X���ـ}��L�G8�%�g8�8���L�.v��ҡ@e	e�������GLN[���0���8[	[��c%����Ӕ�`z�L`{yA�����~����X�s&��j����NH�S[�����]���tᅎ�մ��j�SӔ�`z�L`{s��7z:`N���Qy-v9,x����.$�?vo���`~ۭ�k���%wj�X��?[w�����`z�L`{p��w�^U�e�/�7z:`{yK��d�^��UU�U}O��1��iݮ�$�lmWj�>�ۭ��%����&���di��v�;(�t�v㍥��ɬ�ֺ��6Xf���{�l\�,�T��YNխ�T��,�>�~����{��0=���~��*PbWu�f+`n�K`n�t�����M׀w��l%%,d�ȋk�7z:`{z�ܒ���l�}��Z��X�,����A�w$��w^���,{��pV�E䥱�T���-���遻#��A���p\9�p�k;A�d��H�]"k>�q��X]ѭA����b��Og�	tf3H(g�\�*�Y칞:*v3�i�;/5/M��S�=H��.@Lr��+j8�k����ˍkd_#Y1�L\�n��Y�^�:R�z:�����9��Z�S�nw2��69zy���n�;�^+c����Jږ�Hvx��ܑ�c aM��8ţ`���ֶH�O�>�{_g�k\p,Bc��qC�v��6k5�6�7N�[1��u�(v����l�����Zm�?�wذ߷q`�L���&eԣ0X�eYj��쎘�L��3�ݥjI`R�ڮՀ}����&0=������6�R��]��eZ0������1����GLl��w܃+
�	]�������GLl���d�\�f"�%�˺�:	6�!u=y�j����N�ˇؘ���n���R�9d*r�$��Ye0߻��ސi���'~\�9����^�	:n��,��.3�Y�sq�RM�Κ5��*#�G�>K�������e���f��7�]Q�V@���-����v`�P`n�t��t�LI�Fef^+�WE�/0=ܠ������N�?۳ ��\�@���F:��`�v4��쉦���`~̸07�yf�Z�Q�^!�G=u�V���Dd�sΌ�\ex��9bXFܖ�Βh"�٤C[�J��~��7dLw(07dt�����,DN�Mڮ ~��s�l��z037Z`�"����Q�΄Kn����+�Ę"�07dtͥU�}_m_�?R���2�q(3�B\��d�e�9eHQ)�a"�?� B1$#F1$HD�/�l�Cs�E��o(� ʘ�z�7�l\��r:&`@$�R �%���YLU � �r9NO��`_��2\#"���G�^�Ct���&:��M!5����W	b$�HD�\j�ɐb�q��u���@�C��Bo��s?j\ c�Q:� � ^D�pQ�b�w)����c���aH�A@�4�a��~�s��Ԓo�v�����억$�Z�j�?~�ŀ~̌�%�Ը��zM���Mޙ�hAx�,�Y���쉁�ۦ���,��7=Yc�4��km�8�^�&؞5�Vt�rm���.��Lf��E�:R5J�e��m��{�\��� ���/q%��}��7}Z��etZ.�&�(0=�:`n�`�7z\�l����m��,��{�ŀn�`�=�&�GLY[+,���K`咬�{��0�}�}�n�%?k���M{߷�'���.���%V�-b@�=�&W�����;��`~�
 �w�c���q����1b�w�Ų��	���P�xֽ�.��-Gc��Y83��޺#3�Q�RWq����ŀ~��ŀ}����~}������W%mI-���i��di��Q�5�՛�`~�F���9ě<�<�$r��#��U�~����:��Ir��kLɭ0$��j�:��k�[C�\�}�~��&���������ݺ�k�B킰������������W��?0`��Τ��!�D$q���<`��P�E[����W`�s��zn���O+OY�T��Aݶ�����|e׬�M��Le9������v�K>�8:%�v��j9.f͍�5��([���b0����H5Ai�R���\̥ppnۉ��|{vp��IF�b�C�ul������Y��4�M��n��۪��]}�s��ٗ�ss��ٕg��h���9;EҌb��R��!�(��.$��x�6������r�r�C��aq{Sg�;����jő�vћR��}`�����4�Z�������0`�%�?fF��S��աK`咬��p0��ـ{�:`n�t��P��[W��Uh��$�"`{�:`n�t��t`��C,�J(F!+�W��0=�07z:`{�0`�~��u�Z��b�K���0=�0={&0=�0=������n�rs������ ��n��O[/:��<uF����cm�_FgT��"��LwF{�`{�:������Xn�ذ��y�J��J������ĳˉqbl��L	�`~�G��.Hy�W#���+I%�w�ذ�4ͪ��}�w�W����]��NZ�=����� ���C ��ف�'������'<�e�`�Z��#��ԧww��̚�$�0>�_����~�(:8��88�nƳ�x������60[Q�:���bLcg�������q��EZ�+�w��m}��`{�`d��\��?n�!�jzǫ�
)K\U�-�=�=���&�����0�[�8ټ���+J�$�Z��`�{�9�bjb�X�	 N� ��6�AbFD0B@H� ��:A�ZD����8����_�z���,V�z�$q����*�������?~����I�����rJ&�/%��-� d���̛�~n�Lّ�`|���xx����q�Xt����W������c=����_�w�����P�Ug{ۿ&��$�03%˭I%Ϙ�z���88��A�KV$�?���...�����`}_}�X옳�I.s���c^N�v�+��Z�	�{t��$�5.qUzMi����ui�L����t��Z�=�?O{� ��Ϧ���{�R| `j�H-��Ds����g��^�3S��IK\VG��P`I#�����&0?���ƿo�Pe���Y�oB-+s�4U�F���w$��v�g�Urg]��K��M�n+If^#@�?��L	����&0=�u��k�B�AXF��`��m�%�1����:`l��b+���k�5���;ٺ��\\o���`����{�c�a+SN�%�VI��4���r�󊷻���W���v�v;l�7wq`����kٻ�O{�Τ���q�' �E��T�$P@���#	ޘ:��ݹ���oXsm>�*Ū�	H�v�K���tJ.n�X�����ڍ9��mh�B�.��da��BVώ B���u��ב.v1v5����6�Jk����ZI�Mt�z���?���x!�v�$ ��=�[$��ե{n0�F�voi�촼��Ü�htk�Z�7W'�����M�c���9˭��B-���x�U�%���$��B]ݿ�_���n���9��ay�5�1ۖv�Jn�+�G����Q�/.1?�'}þw�+��Z��m�� ��ـwf��I|�}�b�?ui�2BF���vZ�;%?��>\K��סּ�o�0?d�u�I%��1u=^ ��e�U$� =��`d��7��\�����of�9���Z��v[-m���8��8�����,>���`2[�Ir�wv�oM�і�
��4� �v�x�Ǿ�_�=�z���, �:�Hh"�"6b��t�Ƶt�[���y���\7L]�w/P���.fQ�j����R�k�}���D�����(��.tY��t`��R�\c9Ԓw��u�(@O���T�@a�0VDH���%�s�\�������^�0�-���5�d*�$Ptvۀw{����%�� �"`{r���$+Ut$����%�� �"`t���V�"l�WJ�B;%x��� ��`t���V�*m�K�Į���ˮ쀋�);9wlu��[�����V%�˙�jI`�r�n*슲Kp{"`t����+`:&}��(�N��,������,�M�����}����p���AKd�c�4�	7�繺�r��Ƣ �C�
Ą|B�z��=��:�o��I7���s��[���vZ���� �����ŀ}ݻ^ݏ�F�UB��9,��&N��袶\�	{*%�Ǘ�ۏV�.]H6"k<nZ���{K�`�p�����f�O`��EY���nҥ�t���+`uΘ�;�Ln]u8�!Z���j�>��k�:��0�D�����P.[�*ıQ��.違2u�fIl��U6kLf��05��}54*ԮH�rY����;�0=�El:��W�U�}__�M7���רr�V�Zۀw{��$��'߾��_o�`�[fv+We�w�Ap%�@�u�W:��uZ��'�/��֣[��gQ�.9qₑ�V4�;*���ۦT��$����٭0=6�mN�w��]�׀u�vg�\I����o�ذ��c�.qq6o��	�F
�T؇l�{޸w��q.$߻���~�L_�u�c�A�,��.s�s���O��`}>��L	Y��7���{�u�k	��멕ڰ��e0>K�%������|�zF�O�qw�-	����\�:� T#�@#�!!@�k��R�ğ�B7�Ɉ�!ɑ�i���o"b$tch�0����[8�+ خD��,�	?ɔ>!�5 �)Gf¥�89�j�A3��3�cY�0�Wd�&w�4��
a"�i�}����aKe.�R�,��a>��Rs<�L����b'0d�T
�$S��@֬MK��[�����_�UUV�Z��J��А&�gL[[n�z�joO��ۜ�crGg�������Ю�[T��F�K6xH;NDۉ��˟W�����H
ʹ��*&��
1�71�-UR�J����JM؂4E(��u� UT���:	�8��`Dѧ,�4�V-�`U$k�N]��t�]��֖`ݓq��x�{7�:�z6]��h-�k<t��@�nP���ۍ��L;]<瘺�B dw=ū���/m��u�����k,ݝ9���rc�T׶�f�3��J�-�h{E�4�* �|��,V5�]n��X��m�Rt��9����mU+�v��ÙZ��xw9{�c��
�GYe`+�ї#p�w��_+i�æβI�}��}��Ѷ��*�k��(p������c���'E*�[�qJ�*�T��أS�����"��@�,�=i�3�v �r(6f��I4����v%8-�BN���mK��Ă��U�Рp�;��G���˜Z3�Q�-���`m��-V����ˍ.6�jb��ضzgn0D��I��4���jj7`\�ek�퀪�]G��:z��R�'p��(o�u��O�9��X�-�9ו��W<���u�u���9��6̦;�q�n�4���n�j��x�=�{�f�l#�:�$�mm��3'E1Y@�Wv���+�*��]�+��M��N��a�x���b����n��^o:U��kE�p��O���eΚZ�7�5u� m�5cp�m�)h��ʺy�� mp��N�el��7�g���
��QVVQyKm���=U�ͮVnA0VGq��F�=�Λ�๶���^2��U�l�<4�m:�p�ت���*��-���s��9�jȹ��Ш
����l�����u�ԫV���v��71Z%3Þ����z@�$�f�C����/B(��%��	�6�����cm���y��.EyB�mHMUv�e��D�Ym�<n�����֮x���>u=EV�s��9-��@8?�3��ob.N�8C ��Z*� '�:*���  ��6k���;��`���]Ֆ�Ō
���:�MͲ��vu�����F��.�/��DG�L��  ���أ#��ձ#�fv�dɜ�ܛu���[sm���O�}>���4�t������}a��ǅ�:�H�E������r\k1�ڣ����Ƽܙ���:�)D�1����z���0�7m;���s��`]��ۜqpSj(/˽Mˬl��9^x�d���a�h�c��Ak#�ӮCr��j��j��b���V��,���>��	$i�=#Z��A��[LXu�y4*ԮH�rY�n�qg�.s���4����^��RUD�vV����(��j�Հw��X�n�������������_�|�݇���nT6�Rʰ>\U��>��l	�a�⩓&���,t)Gyj��
�����q-����&����J`~��}UtYq�d��nҖHn�vm1p�s�q�ӎ6�Վ�N��2����e�K�2<Í�B�*l,����L	�0&e����K�%������?��{�:V9vʰ��Ō �DF$�$NAT�C�DJDA �����I�$�;�wwqg���&�=�z
�u���`M�`�'�[7�\J�n�Lɸ���Ոb�P�����u�6�wZ`Odi���q.s���x���Q��n[p��X��Ė�����]{%�=��'{ev���rL(㓶L�^�[�]g)��s�^�fף��l�/绽��_6li��W~rkL	2:�K�qs�}�%�s�����X���n;'���w��z��\�ɶ���i�=����...6~��+w��d�� =��ԓ��tjp�dS�C���o{����{w�����C,h�J�m�%�����]�~�Ɂ�~i�3#�����s�I���u���GmQG��YS=���$�fO�~ ݛl	�4�����(Eh�$��'ma+��g�NM�٣a��v9��mM7l�b�V��w{�m���u�㲯��ﱘ��n����s�/�owذ�^�����A�k�ޮ$�Q���d֘쏣Թ�&���y!�dU�m�;�{���5s�*��_F�l��%w�%�d�[j���9�ė�����7}����M��Τ����⁀��Ͽo� 7���8�N)eX��܆�.qW�m�&�L�F��K�GL�˘#"���m���٠�)�Ňn���t]+� g�Ķ�;���WٟM}\��n�~ �Ͷ�F��j\�8�Pg}����C*�)Sae� ��֟���qqs�>��L	��Od��s������D�*��A�,� �wذfGC5.q*�rm�2n����B��I ���vU��ĸ������a�$�ro���)B������ʮ���'�[��ϗ9ɿ}��>��L����U?�u�((/s2�
�1F�Z��ڷk�e{K�H͇��=l�rz�	��r�u���8�G�m�tH��.��`�uVvp�.�qn��l�b"�\��-�F���H�����������z��.�s��|Ym�1&˶��Q�g5��i��;en�����ƶ�랼��<%�]t���S����u;B�8���6���@[bΝ�s�0��ƺ���>���w���=��>��u��4�u֑��$-lj8.ؓ8��)�м��q�q��.,��o�$:슷-�����ŀo�4��dtjI/���`g6Y�۪�vKU��wqg�6w��C =���;��Y�ēa�Oz�F'���3u�`�-�ĕT��07&���ݺF�d�6ժY-���9�߻��o}�|�����q���9�7������ݏ؛�DVR���K���n��>m��s��n����UU�~�����=.ꪫ;�QN�׋g�p�mfV�Q��[�na�|�pل�WG�TB3�;�����Fs��_�6�f�!������>���ݺ_q}#o��|������Nz�@+��[,1��~�w��� >T!q�3��gV�}�{��ͷ�n�3�$����k}�_��� ��@����l���q���������cm�{���o��jBv�vZ\m������/�m���Cm��i�Ϳ���}�\m��{��-�q�m+�}뻽�������ܠ����'��6���q��F�
D W��D�t=���I��3��V� JM�)��N���"��q�[��4E#�X|�o��x���;ۥ��{��/.~�}��Cm�����֣����6���.s�������������������w4��%�����%Q]M;��gv�~��f�e�^�F5i� ��2A6 �����Mn�g;�L�[k���nGY;e�g�~K�N�{�[m������o9�����\c��7�m쇔p�+��Wj��o���}�m�8�#ۯ�UU$���ꪯT�u�UW�J��
��S�m�L�R�^d�]ekC�v���v#VE�LX6��p�mڤ6u�Z�~m��}^6������o���?���6�{}�����my!;d��-�m��w���JH���Sm�����Ͷ�۵����\V���`5�e�:�m_|�z���Lm���~_|�Ē�=�����}�����ܢb,�F��uʦ6��q)>�}��m�s��[m�������(/AU�s�_{���1����x!K!H�j��j���}����w~_|���)�������o�q$���Z�Te�U��kC�՜����[E��;@��뎡b�=�ݾ�AeEu>7m��m�o��_|���)�������\I~�ov��6����=X�d �U�ͷ����9�#{�ٽ�m�s��[m�9ݛ�����s��O���jT�S+�Lm��{���Ͷ���7V�Lcw�ٽ�o/���۾��ak�RKj��ߒ�9&�z�m�쟽^���܎����tp�����@��P��*춼m��w~_|�~I%��|�Ͷ�}�>���{v�m�q$���Qy+��
��|p^�벗S��bH5;�W Zˊݤz묓�sWyG��6��q�+�RM�D�jFp*y�A]�<j���!8ڇh6��NC�`�ѻv1���5bÌ�\;�=2��9ª�fb�2�+��Ƴp�92�	X�ո����tc�}�����g�,��M�V8�����{�Cs�t��ۇRh�wN��n��7%+�@���_)ϟ�V2_������ƈ��YSd���t�u�;���%���*`'�.sJ<%��H�m^�m����Sm�w4���}����%�o��ϛl���8�mmH����}䒒7�}^6����|���Cm��w4!GI\b��d��6���.�������q''f������|����B2�������$��ߗ�6�/}�����]�ݷ�
��s���um��O��$V��YW�6����1��R\���{�UU����UT�~_�UU}���{b�W:�6rmpFz�3vY@�ڳ�]���Kp;��csbm�n�l�|�o��x����v�m�����Is�����b��o���B|յK ���n�o��su���o�A�XE�0E0�,W�)�*��FB$��XE��3+�I��AG	�P�wo{�7�m�}�Sm��i��K�rH�͡`��v�f��n��������~�;���ʇ�V��g��Ͷ����m��opl�%����v��m�ݛ��m���|�o�n׍�.s����~_|�o���]�h�F��m���|�~�\��}O�m�}��6�������:���"�"��X���؎ժ[�8��n���/.�-���.2�^���$�W.¶:���%?~m���SV�{��f�m�s��>�m���_��m�?����8)S�vZcl{�ߗ�6߻��uUU28~�UT{#V��_$���V���������v�*������6���]���{�2�0G�EH`��`�@���ʨZB�D,�H��R�D���H4�s�YI
43w���ޓR��j�P����t�@�d�Mg ���(ʹQ�2&�΅�� �-`S `�(�����C�[L8�&�jH�Z� >M�dD�D�P���[+��i.�@��&�CpqA> C"u@��>4
�W��ؠi �B�`<�]��u����}��6�d�	5�v��ʦ6��'��x���}�e1���w��ͷ��qLm�����Ζ���n�}�m������l���������UUS#���U_�{�������ú"� H4��v�c�w���h�0��c�����$��8�2����vKOͶ������������6���i��?���{��6���`��N�mu��Bھ���>�)���w4�����Lm�������H��;��V㰈��d�cv���������3V�?�y���ݶ�����z�w66�b��[]��}�o��9�o3V�~���{�߯;�����J�����6�黐tU�*�X&�˻��OW�ww���;���8{�ww�m��%��p�D�I�j�!ю�:�:݈�V�Pl��!떤�%n{�n���C��1��v�*�[o_��Lm�����6����y}#o����6�v�8IQ-@ܰe�������|�o�w)����ߗ�6����3�F��'���J��
Q�)�Ͷ���cm��n����)'^���}�現m�˥ePZ��r���Zcoܓ{��z��~u����y�޻��������������c��%_|��w�ۯ���ʪ����UW�I�~�UU�*Vuߟ�ڶ�ݹڧ,<��^�e�.���<�lĻ���\��[��{l{u�r�\DҚ��ug{t�s��::��v��y4�{[�-RЭ��E�^�	���̵������C�}���;�eg�xKu��S�x����(���rN��x�-���k�[���=k0�k�$$�P�vB�Z�d;+���ݸ��O/A`�v�^]�ە�ȗdkhru���ww��?ǻ��O�~�i�E���Xݎ�4���M��0;r����fCnP�q��{�?�����*�m���nx����v�m���ߗ�6����1��ս�X��r�ʬ�S��m���f�)�b߹�l���э[m���}�q%$}��Aҹ��O��k�m�s�ٽ�oםэ[�P?
g9�}��{������m������,�A�m��Uz�k��\�#L7�qW�o����_&���P7,]� ���0q/��?z����0=}��w2fYifSƇh�ٖ���2(Uq�\>����y`�ՌF����T�U�[QEPݔ��ݶ�#Lՙ;�s���$��(J-Ay��qY-� �wqf'ĒX�8�I��Sªgs�=�5$�|`�wq`��ok��W-��V��'X�pf���ʬɭ0=��0>���;j��,����S����̚�3-XN%�_��:�5d�iWY��V�+K�����#��f���� ��z��ʩX6�j��%aAq��k�n��llo]G��lˆ6��_���˙+�V1U
�,������,��v`�ۧ���;��,S���t�0�Rĩ���1���ގ��?�$�?{��IY��6Wl�7�|a'�s�52&BG�t|�y�ǵ�,ϻ�n��q�nҪ�D7e0{#L�#L���W*dz0"����;l�%� �{��../ݾ�������X��\{-nP�Wx�t]g�OK��{8m�8gcW�b��=\������R���I7}��O��}��˃fF�q$��l֘�W���آ�������t�q%�q���b�?{}� ���0]�z1�[K�j��l`Odi��di��..*�����~0߷r;,b�4��`{��$�l�Ɂ�&���˃�,K�\���LOY������Vڰ�w^��&G��&Mi���4����T��ޗ�r��:3Qm۵R2E��R�����˹�m��.Z�o����������% ���d��0?zF��_�=��L��2�KD2!�)�w�wyq.s�C'�4�ϻ�S�˃��K����w�_ES��	��"�J����,훯 ���L������l��UU�m�J�j�\�mͦd��07�\����X�]�������[^��n���$��~ٺ������q!$s�1���6P1Y��2�n��BD�d�&��Yqw.�*��$��|[t�h\�i*�7�ܛ��O���)���4���m�"��ѳ��\f�	�����ڥ8�r.cE�;Y�'��ӌ��:��C��;3[Y�6)l�y�L3�t��<j�65���ܜj�[7d���4����f��[p�����Qx�gnz�ۇs��5�-r�Ka�ؗ���^K�K>}�����>� 2�;a�]0y�[��z6�J�Z��zIkq������_����r���7�0?zF��rS�˃���5A��P��ݫ �{��ˉ&����`L��=���I*�,6����j�Xeڤ��������������q`�l6;iS�#�Y^�\�����5�鑦�q%ϒ]Ϟ�L���<���!��L����>��LL������\뗘�ffV&뭼��ˊyy{mD�e�&�-���!y�F��U���X�Y�>�Dl�[%_�����0?N�L�\?��\_./t7w��g����Fݶ;*�>ٺ��s�\Q.~\K��~��������ڣvU��X�GU��k�7�|`�wˍ������x���[�[k����a�I%���������0?N�L>��M�}�`���5A��P��;V��`}��m���3%���di���O�C�^��l����w5+�<���.�3��)$%tzCLo����cd.iW���?[w��0=�:`{��l�ڛ�+�Y^��n��$ٽ�b�?w�ŀ}���ˉ6{t�0r2��X]�CI���#�}UG�EW�K�d�b2�B!a	)#!(B�;s��]g�׮���/���k*�b��ج��/�.)�８�~���\�`ze�J��Um�e��훯 �\�w<|�����X��u5%�"�
)����;Y��m��V��6Ƭ�u3�5�y�w���̪R���,�|{���������%��kf���e�-�wT*�����#Ox����zd��W��X�v�͛�{ ��QM!ڰٺ�N�}�qUfKс�5�/D7�����[V��Ğ�o���}5$�y��"E�E��P�p���I~�*�9�n��݋V�%uKBU�E}���˃��qs��.%�o�^���� ����>�2�䎕�5Zv�����Q�bP8�ڮ����lF�����c�������i�H������>��ŀ�v��q%�ݞ��;�k*��E]]�]w���F���.s�w��߭���<wqg�I&������Vݷ�]��7&���%3�q.*��Z`fOb�7���H�,�
���n���	�`{24�y�r�sv��� �]ҵwW����l	�07�:`dL&����I�Ƶ$f7���CN�����a��	!�E����+~C&�>!$��C�:$��� 8 �	"ċҔ�Y$�}����� ��5�GL����M�.�hl��L�3�{Α�!�$#ȤB2������	5S����q�c;f�6�m��hh�R��@J��-�[3;X�����Rb��P�8��7 n��򳲵*�n �e��t]m]�2�y.d��eeZT:pI@cb� W����V\B��d�ع�!�n��UR��Be�5�X�a��3dxAU3�[F0�`��W\���Н�/[l����Sv
]b��2�Vcv�ӇQ�Nӫ�i�Z�"��&@�ݙ�-���]�;7��psW6��殳Ľ�\p�<�ۥ��.v���hp 9��*9[L�e��ƥV�m�rm�pT���!O%٩�n�J��W��c����1��n�j�y[��{UJ�����L
�K�*�+����V�v%X
��əz�B3F�� �; ���Q6�T��QUT�ܳ� *�VmV�eQs	֬u���vi!��5lٵm �6m&nm�[�����z��WDF^��',��1 ьZ�īt�p� �A5�!�-gjH[G-��J����Ͱ��&0l�N0�\�Z������̞t鳲�R�����$ ����*�#��W�Cd9��;Qð�l�mAa�^�9��b�u�s�<+����F���FSz2�����vl�i�8�=g��vb$Nͥ�:���,� �q��74���P�{hN�Nk2�����<ݬ���Ͷ�۳��&N��Xk�CnzMg�.)T�u@�W)"��-���Bk�[�ƹ�F�ƣs��.�+�$��9j�Yv�x�2�m�؁PU�Rvz�R��r`�p� ]�P��3T�F�9Қ�^�Ќ��g��sg�lv3���,=i�H�s�tr�ѳ�����F�n�%5ut�p��/\b�%�I	
W�j^
�Б���6ͶCa�ڪy7]l�Z�[ �jPm�TbF�P���WvP���R��1���wlm!킎:d[�Y�7��ل�;d@#m��pK�h���� -GŎ�TV^ݻ1M[E���V[li���1L����� haB����x*J(�C�+�A�;G�	��* ��a�s�;��Irf���EYy	�S�#��9�[1����Z���iW�7<mz�׺뭸
�\89 6\W�:�c=0�.�[YF�n�x,Ҽ�Z��� :u؁��Zۋ��v�9ay3�ۋ��z�c��
rcZz���u!�vV�\y�	wn�id�##&��/H4��S��+7j����e�y�J���[;z؎��$�1T�%��\3���<>U�J*ڀ��)�eڶ��Qs���s]��by�ņ�x��BN�s��q	l#��;W��ذzK`~��Z���Z`E5�����+�.�^%Ll���Ζ������qg�9��;�O��V�UGl,��ow�`L���di�OIl	�E���Tbt�m��=�?w}��?n� o������|��Zʽt䖹����di���&����L	�����먎��Z��EU�uW�M��C8�7[�u�Ӊ�d��m�p�����sb�*۶�ʿ����`vw^�����\������b�=�w�2K��J���f�;�����,I%��7_�`fMi�+�v`�kA���Ɯ���x�������/d��:[vGB1e��
��������/d��:[������C�X�����-X��cݝ-�:GLoGL	+%ʵyZ3�s���c^u�s7nhmH�m֞�^�q��ǲ�O�������Y����o���-�;���GL	{&0'q)��IP1�!�k�7��Y��.&����`}�������u�H'�\�ح����N�%zN��$q�.8�u�WҾ����bv���遳�2��Z�wi,ŋ�L`{s��'tt��������D�//*�Km�ݝ-�7�������WVf]����D*#����HJ2R�Tte&���!�q;\�sv%s�t���y�Gf�>�7�������nt��BJ!2&�v����Y�<�������7�wy6j�ߑ2!�DWT��`mdް?grS>�ܚ��kL݋�-��E\�v�0?�����5��������4��	���I. ��"$R�(D��qq_o�}��n��R
�eUU�Eݥl	�0=�:`Kޘ��Ζ�~������h��r�n��ƑPGcv�jL��cn7Dq���5�U��aW��&�����R�����Θ��07s��&�ŀw��:�Ali�[e��_���U��Lɭ0?fF��W:��݈R�Y%������7�wo���X�w� �����A։Uu����i��#L	^��ʒ�i����W���JÍڰ��ŀsӻ����<wq`����5�Z�)P9c�������:�tu-�9�Y"�l��β0��b["�[P3��lܗ,�(�fW��䝂˻Y�M��.8��^u�i�jõ�[����3�7(I�v�6��͛���n I�w���M;qЗ9F��ΤN�����V����8�]��ͷkg�ya��۠�6+t�;۳u�ϡڗ���{�'�3���.�/e�:8���(�?���&ݢ��S�*�-�c����ج�m��8���ۆ8�"QK�"+��W@����;�n�{�������Ų/FY��r�ۋ�%�$��nI�	rL�����&"'��7H�ܯ ��ذ�{���z�]����?~:&�� 9R����'H��%�7�t���mn,�u�X� ?n��;�n����쎘p�BT��WJ��$;H�c��2Fk�c���f�<����lU�n�mv�=���iʚ���e���M׀w�w�{�����y�w�aF7X�\�RN}��֑v�iS� *��LK�0̖��vJ{�qU�YA}�U]�HZT�����"`v���Ww����I�Wn�mX����gwi���4����ԱVUJ�X$�&nIl��d�X�wn���l�v��ep+�	8�����[�Z;�o<�W6m\���Q�nk!j�CnW�w�w�wq`��$��R�2��,�U�)*�������\\J�3wm�'wi���5�w��4,bn����V }��s�w�Shx�H$��H�HH!�D#�P�H�0
H(1h0�Z����p&�ٮ�ߴjI�s�5$�ӹ��ۖ�,ŉ$���-���t���������f��Q�m�
����-�gGLgD���-�:\���T�5�,���<�ܷ���wm��m�c��XF�3���8�f㲊�::`:&nIl���ڴr9��n�eX���{7^;��`N���[W�r���/$���[uH���� �"`n��fVZ�)۵�T��w~X�F���ÜK�8��$��@���5��I7�9f{�HLc8Wx�*�T����I�0;s��$��,��͒Tꨖʣ�Z"^�f�\2�t�b��#�/./i�iܽ��OgJ��һ-Z̫X�f*`:&�t�J����i����}�
�bX�`n�K`I]0=�:`tL	[��f"�e%V$�,CN#�����ۀw��`���l-,QP�4BU���n���6M�f\jU���w�ÒG�e���� 7�ۀ~�n�	0�0$�� �9s�H^Q.����[�7/2f�:��j���uq��ŊBS�.NN��7��m�]��z#\!��8wglU�|6�k{��
6���2՞��u���4Y���K�����j���R���q���Y�+�\�C��v�����q6z��F��f�:w�C��um.f��#tcDcz�^��;��n�{d=>4�s�[��v�g6��,��DO�
1i��u�e���Iہ��ݻ)�u<�F�<��w6���8'�ڣ�؛�Nɑ�%_�Ĝ������GLwD��T�fV[�)ݔ�7zn,�l���X��\wn��]e�\�UnUj�T��GL�D��(0:WGL��4n�6[vP�� ��n��FN#��:`M;�R��YKX��I&�A�Һ:`I�� ��07@����jؚ��Lm��6P�)û^ϫ��<zv������gOU��3c���%ib8���:`:&w(07����*�Z�!*�>��Y�*�FH��`�  L���US`'�0$��GL����`Yd+uYj��ݸ{ۦ��0&���G\�����/
�I0'r���oGLgD��](�Uj L��S ��,˞���������� �K��_�r�q2�s׷!;]\���ŶKQV�:
��X
!��o��D�j"�UnUj���{��T��	���8��A�����K4�cvƝ��Հk�v`ݺ`�7�wq`�w�m��*��%� �	8��*��}�eYEU����'H�X)�f�gr!#�֖0P4�6��\A��|�}��Y[�0�A�K���i�"��(&`���0�d#JQVc~@D�B���0�J�"��Q^�:��/���`FB0�D�(D�@ �F�q�PNBQJh�F$3�����E��D���d
��0ɅF�хNG��� 8�Rl�t'3�05T�BH��#��^�d؁�J�� o��P� n)b��H$�`,`�)HQ���x�8U�����lv(�Tu�Q�|�p6�!9-�Θ}�[d�B�J�U�K�5%�;����}��0%{'X���ݑݗyk����T����w�7�����f����TGo�O܆͘��ݨ:8H�!�-���i�gD�V���q1��vm�]�w�o���d�0&a���7u����uA�Z[]� �v����M�վŀw��,N��>]]�L�؁2�!�6�:`oH��1���,S��
�%Y���0=s�Ƥ��s٩6 ���FaP�0�I.p\���~X��Gbm�mi�RX���1�������� �������H�� @��!+Mע�&g�C��כ�5dۡ��R+�����k�u��Y�,`zEutt�����c���MNج�u�-��;��ŀw24��RN�?Ip{Ē�3&����}���!IV��b�>{�0�n�z����ڴ��J�Q�� ?I-�&\�F�j\�ٿ�n�^�<�m��J�����`�MŁ;�wF��}�s�'P>"��,h�Z�R�F״��2d0{��~�=�nĬ1�x�\�9^��;$Q+ۡiNp,yz��t�a�Fw[�������;]����E)m�F����-�q/Yݚ��mg���cGV	V���7c;g��'T����zKv�׉Gv�vL��.��d�v�l/�H5�.�C�;�ڬB��8��D��]�Lk/'[�v"P�ڶ\����A!g����%gP��s�����;���?[�?F�67G����u� vBN�<"�`�A�xM&�+Y�r�p�V,G���:`I�� ��z���`���dj��+]V�J���, �2^��ݗ�HkLŖ��j��ZvRYV }�ۀo��0���ذw}� ����m��8U-���w�����06�L`o)��,+E�K�07eGL	�06�v`��L ��Ū�g��9]�i{ �V�4g=t�uڸyg��%����Vln;������ ���X�ـo��=Ϙo|�� ��/ ����s3���}{��Y�#�%(�*��������x�.����:`wE���D��%�	l�7��0��t��s�0=S�`�řt.�_la�J��&�֘�����0�u����k䮫k%X�u������6m��Ʉi�/ =%�S��n��<�5�n�N�Np�	��n����N�b$
|�V�ړ�
�&�]���ٽ`L�L#L	�4��{:P��F�T���0��xw���;��� �����mD�]���ev������/������˜��ْ[l���1�R1e�a���:`l���l�GL���+1�r:r�j�?l��s���?��i�X�w�j�e,��R�cmu�@�<��J���vM�}��ԅm�^'�خ{Cb�*�uZ'-0��x�;���0;yA��!-�Y��ˢ�Ye�l	�GL	::`v�L�lN��B�DWU��X�w�ݺ`gK`M::`wW Ʌfi,�v��0$�J`Oa9�ĵ(􌊄cE'X�B*�!R ��B#*FJ���B�$ -Q$P��Ba�@"F!	 @B1@"�T�1R�!�V0�Y$��	2	D�����q�I8��ok�
�U-�����֘di��˃R�\�Z���Kz�h�<����q�q)�b�&y���N�AL�b6aVKS���(壮�]��=�}� ���w�3��7z��.ՆR1e���::`n��t��7qf󍚻���"7qP?vw^��h���$���䴐*�-Q������%�;I07�t����x˽(�"jK9^��u�d����l��UU�a��G���������~��j�\�'��ėGQm�I!�Mʇ�ѳ$q��YA.��m�.�iE��#M�[=��6�3�ڶ���#s��M=��Ls�6�`�Ƥ؜�(��y�tl���R��Y8z�<�5�ms���!���{uȼs���;//���+h֮#V��IpYmɒ�eu�%�V�=��e���L58G3���R��s�wf��Q�]�Act�9/]��y�Q�K���#���ms�"�Y�ݴ��^�h�pwDq���u��m�Iz�::*�X�T����w:[�$���ޮЛ ;F;-nՀ~�7^ݒ[g�d���왔�*B��/�vIl�GL�:`k��0�-����,�u�+��{��J�a��7u���u���)�=�t�RX���b!*�?n�,����;��i#�n_L�RK,Ϯ���h��l{/d�9�0^��y;�k�:���n(6�:��ԕ�#���,� ��v`�n��GL�0%���Y��2���,`l�}���}U�G.#��0??۳ �n���5RXBJ`��i�$�3j��w�ݽ�b���X��e�<�=��,����7{t�?j���;��\jB�5d��L�d��p`z,�0$��y�.���o����@��Ց�k1��Y��0�ϝY<	��4���Эۤ6����$�i,��E�`l���tt��ٳ ��۪����V�[)�~��ŀI���$����� ��Qj��\�ʰ��,����%���� ��Q@!Z��O�B2@KLav.�_�{�gsRNs��5$��tB�a\���,v���s�O����?~����%�`t�遷�!�,U�ZG{v*��`d˃y�߾<��o�0>��x�of���U;Z�EP+\��8�&@ꃍs�6N���m<�'��sճīK2��ņ�`oH:`I��ݓ_�>a�m�~�w�N��Kai�&F���9Ī�N��v^�dQ��8��ٺ��=�H[Z�V;V׻�`I�|��j֘7Z`eK�l��U���-%�	�A��*:`N��ԙ�!�
�D�
"!i*�X���7]���'N�>n&l+���e��uwq`��X^�f�ۦ��ݎem`�#`��,�v9���cO�k��t��z�tu�#I<rcSIhm�`5H�:Z���,����;�t����Ob�5w��$���V�06�L`t��GL�:��5�}e�;E]	,��}�� ���Xs���X_�� �wJ��e�D�K-+J�+���GL��鸰�:�ҧ#��q[*�`�wq0:�L`{dt���}_a^��ʠ�,�a7����#Yb�RDm��\5I�B�K�I�aN��0!!F�$�i�1KB�����W�"B.`�r��	!x����60@N
J�Mş"0��B�p�!����(٤$�#��2�a
F$jJ"����g�4H�!�K����d�=��$  ���$ a�����E�	�
T�R'QӾ�
`!��z(��Su���E�F�,�I��B�6�xO����]R���a@���^�4 � O�A������=�1��{�m4'��d"�������� �EYb@�H�I&D0Q$J�>���\�e�$BO�8�4ga8 ���9r���m�6�I+nڸr5TWR����n�b��,�t�Y"෵��Z�`W=��U+���[���99��Ĳl�m����Hiwl��jGl�A�0��J���M�[�3��V�2q�q�j ��%��;t\{��ŝ���L�Rn=Y�4�F�u��S���d��ܖr#��g��u�+�"qw�e���<<c9�v�@sV.%G�u������s�=�v]#��k�u��OP�����j�;�61�UV�X�,�v�٦�J�4�x6Q��X�W� ���%���Z��[����UPI���쪫W�8��� 4�Wj��Z��S��>9��Sc��U�X�3l�ji0b� ��7f8����E*����;J�Si"ٹ��]l�+b����`�P�\�,�Cn�5I=Yv�e�z�6ySU֝a&�eW�1�]��2�\�`ۂt9�q+�Y K�����]�3PtX#�I��3�L�]m"�}����,&�@ɑ�W�s�A��'ni��r= ��i$��md�
�n%��	�:-�8��#�.\�hہ�������6Gc����s�����q�v�U3>3r)P6f�z�&}X���,����X��w=�1 NUΝ�_a��KŒ˲d \����w9Az��ݸ��;�\DD�l�/8�v�y2j���IG72C�i��{X�[H=a펬��췞��y���6v�g-T����ƻQv�{6��]�[b��-��iÂG9��f�S3��Kb��Al��s����.�Z�b!�r9^7��O�ۗcS�u��(�U�zl�Z��P���^�e��LA��Q(9����oef&�U��re���:����*�k��>����A��Gt�qm��.qSu�J�2�ݱ/��,u��ӎ�����1:�gr�wq�2�;�<O`�����k{2�#J�/H����s`N�J��ԥhR�]��39�s/�Sj`1�8�z�e(�t'J/T!CJ 4��~�D�h>�Iw���|�7�o)[r��96F}�'��l.�'Z�HwR�UEt�*C�M����+�g�g�:���۫Yq�������������ʠ��]	�w(t��[N1(���ҫ��\!A�o(m�/�Q�x9la]M�.A�E*�3�Zu�]����j�7����{�Wk���SC��/OF�4݀:�mz9����[�fݞv���-&�kK܇������6�vΤ�W)�j�D�]�Zr!���b��r��$�w�;��yruܮ�B�Ukp��t��r�g������3���j���Gm���t��\��;dL���k���J�+���ImX�m���p��M���`����16J�"�u�5wi�g��T���\}Sow�`u{��&ZY#����n��ـ~��0�� ;��p|׫\#r�)8�y��r�#8���n[m�;��eΦ��wl@DkE\�Z��A�r�Yl�>��0�2&�"`m�1��8EܻĂ�1���7��Ns��Юҋ�B�q':4���-��(0=��Ww�����k ���%�="� ��i���B�	m�>ٺ�tP`$��7�&�LȒ���[-����� ���|�����l����j��k(+I�Uh���*�l�3�q�f�Ct�9Q�Mͅ�gM/�{���t��Z�v��|��;��wn�����>a���0w�16J�"�u���&��0=���ؠ�&ɉ��Sb�cu�En[p�;� ��u��\����.�/;�3�$��ۀk�͕T�L�Z'mx�\~ۻLvom�L��}^ۛLBhʾ�ʩ�5� ;��p{�p�w^��� �~'u��u�2�U*x�n
��gvr��[��\�؄ۭ��m�.��ۜU��Ī��VE]v� ?n���L��뾺Mı,K�Ͻt��1ı/��K�_L�g8�����2K\��Y3��I��%�b}���I�~#���b~�~�Mı,K����Γq,Kľ�}�&�X�%��s�c��L�K��9�s���7ı,Os���n%�bX�����&�X�%�~�}�&�X�%��s�]&�X�%���׳��s��-l��e3�㉜L�g�����ı/�����Kı>�}��K��G�)��N�_}4��g8������l��EH�u7,����bX�%���t��bX�'�Ͻt��bX�'{�zi7ı,K���:M�3��L������N[j�*�NZ��=�i�ᐡd�M�����D�V�e�<9��u�ۜ_L�g8�z��8�ı,N����n%�bX����t��bX�%���t��bX�'1���-E��r�;k�/�&q3��[�|�7ı,K���:Mı,K��{:Mı,K�g޺Mı,Kܞ��v!ʡT�5�8�8���&q=�zgI��%�a�8�~Γ�?19�?�]&�X�%��{߱��Kĳ���S��IEdU�is�㉜L�q/y�gI��%�b}���I��%�bsﱤ�K���C1�~�3��Fq3��_�^��֜v��W,�[�_,K������q,K��=�cI��%�b^�ޙ�n%�bX�������g8�����i����Q�ȉcE���t�����C��CF��x�s�k����<y����v�F��m�(��]b�r�1�Q.�X}���mWBzPL�4��Swڀ�`���Sm���'t��hq����q����Z57^�n&K#@���6%��v૫ح��R9�]�W�Ҹ@+��[��962�ҩf�>ϴo9�r`�ˋUvy�8۱D���\ǘ����H���
�X$śF8�4	\K��v;t3ш�ky��2�i�T��l���N&q3��^���L��Kı/{�L�7ı,K�w��n%�bX�{>��n%�bX�;�{8��rGke��ٜ_L�g8��\Ḗ%�b^��Γq,K������q,K��=�cI��%�b{��ݭ��"�u��)s�㉜L�g�o��q,K������q,K��=�cI��%�b^�ޙ�n%�bX���G>q7A\-���8���/޾��n%�bX�ǻ�i7ı,K���t��bX6%���7ı,Nc�ު�Z�q7-�����g8�ų��4��bX�%�{�:Mı,K���t��bX�'�Ͻt��bX�'�$����Q��:��剔�:��&íq�ʨx�6�<�y�h�j����"�`k6�y��qI�gO�X�%�{�~3��Kı;��f�q,K������q,K��9�cI��%�b}�:]>̹�ɜ���2gI��%�b{���&�K	�ڔ
ERN!�P��O�X��}ۤ�Kı;�w��n%�bX����t��bX�'�;�=E	k,�r�ʳ�㉜L�g�_y�n%�bX��{�i7��D�K�~�3��Kı?w��Mı,K�e�z'kb��U��k�/�&q3��^�ﱤ�Kı/��c:Mı,K��i7ı,O��z�7ı,N.�	�
����m���㉜L�g�}�gI��%�`�ｳI��%�b}���I��%�bs����q,K�q����~t;��h:ëɔ�-���ib�t,�qӯKg;V��[��7mtS��	<�L�1�g�n%�bX��}�I��%�b}����n%�bX�w>��n%�bX�����&�X�%������1��[��L�\���n%�bX������P�,K��޺Mı,K����n%�bX��}�I��%�bs���i-L�',,�����g8���o���,KĿ{��t��c �� A(�
����I��%�b^w�Γq,K�秽7��n��1�☸��n%�b�����oI��%�bs���&�X�%�}�{:Mı,K��޺Mı,K����<����Y\�8�8���&qww�,��%�bX������Kı>�}�i7ı,O��czMı,K�$��v����|燒���q�ѝ�(�i����z��$DN�����]��������!�n�}ı,K�����n%�bX�c��4��bX�'y�]�7ı,Nw�ٜ_L�g8�m6xRPN����q��Kı>�}�i7lD���A9��F��I��r����RL����G��I"v�[i-�����+���~��n%�bX��}�I��%�bw����Kı>�;�i7�g8�o�V�S�ڮq|q3�ı9��f�q,KĽ���&�X�%��;�cI��%�����:��{gƓq,K��<zˋ���8�f��3�I��%�b^��Γq,K������Kı;�x٤�Kı;��q|q3��L�ޅ<����Q�^ƶ!��`�pR�iv���݋tq�$j��x� �"�iB���,,�����g8���w�Ɠq,K��}�f�q,K��{��,�&"X�%��߳��K�&qx��>��!T�4Kfq|q1,K���Mı,K��i7ı,K�{��n%�bX�c��4��N&q3�z�(y�KT�8�8�K��{�Mı,K�罍&�X�%��;�cI��%�bs�=�I��q3��^��	�+R�m�Z;*�/��,K�罍&�X�%��;�cI��%�bs�=�I��%�bs���&�&q3��]�zx���l��3��%�b}����n%�bX��Ol�n%�bX��}�I��%�bw�����g8����u�����)r����F�i���mt�]]��t�ɴi�
�C����||̀0��v�t� ��x�f^�ɬ;g5e���*��Hq��z�B�n	���8؃���m!��
�M�Kc�u�����!��Z��r�s8�v��q���wC�h�rv}�����F0zF�=�T.0�.�%ù�9�Sm���v���u�]�O#��mW�w�$Ҷ�Ŋ��Z[
NXǄ���S��G�6��98x�7kR���:=z$�a+U��w�����d�i7ı,Nw�٤�Kı;�{��	�LD�,Nc߿cI��q3��]������UB��qZ���ı,N��٤�Kı;�{��n%�bX�c��4��bX�'=��4���1���m��m�q$��f3�I��%�b{��Mı,K�{�Ɠq,K��{f�q,K���Y����&q3��[�ൕ��+��s�&�X�%��=�cI��%�bs�=�I��%�bw���&�X�%���zg�8���-��>�"�F�v��4��bX�'=��4��bX�'{�l�n%�bX��=�i7ı)��{ޙ����&q3�{�I�jڜN�ď��n��l��s.^�{d��ӝ;�'^����,���3�rs�WQsw�����oq��i7ı,Oc��4��bX�'����&�X�%�����&�X�#8�ո��J��Wl�ۜ_L�g��s�Ɠp�h�!��$ڡD˸��bsױ��Kı=�Ol�n%�bX��ﳤ�Kı9���>�
:���fq|q3��L��=�M&�X�%��v{f�q,KĽ�}�&�X�%��s�Ɠq,K���M^����j�d�8�8���&q{�{f�q,KĽ�}�&�X�%��s�Ɠq,K������Kı>���>PUP�:8Z��㉜L�g����n%�bX��=�i7ı,O��{Mı,K����&�X�%���~�9�L���l���Xz�ͣ���#��d�rG���.��7��V�� �����I��%�b{����Kı>ǽ�i7ı,Os��4��bX�)�w�8�8���&q~�^�εxXIa��s��Kı>�}�i7ı,Ow��i7ı,K����n%�bY���z��8���/i�QW*w8��s�&�X�%��v{f�q,Kļ�}�&�X�;�|B�a>�����#@�AL����,J$�x�	N��>qY
�`p,�1lXH�Q�"�#HF@ �f!�4W �所`45�N�ט�b�%D&&1�`�%�
��!��\�E��.�>�+�W(hL����!���6�t��O���\���Kı9�{��n%�N&qoCY�y���U�U�8�8��ı/9�gI��%�b_s�Γq,K������Kı=ޞ٤�K8���/uj�ŖrU,r����8X�%�=��7ı,O��{Mı,K����&�X�%�y��:Mĳ��L��SG�;\�Q
��֤�:lfW�YgN�
mp�ӝ=�q��-�ҏGHӕ���a�8�8���&q~���q}ı,Ns��4��bX�%���t��D�Kľ����n%�bX�1��G?�E�j�d�8�8���&qw��٤�?)D�K����&�X�%�}�߳��Kı>�=�i7ı)����9�U�Y!j�/�&q3��y��:Mı,K���t��bX�'�罍&�X�%��z{f�q,K8�Ž��m��r�+������&%�{�{:Mı,K�罍&�X�%��t��&�X���!"�~��#܎�c��:Mı,K�_��u���%���g�8���.�{��n%�bX�秶i7ı,K�{��n%�bX��=�i7ı,O���?��5l�ں��Ą�H�u�u�j6M׳��rT�YN��&�[l��q���4��bX�'9��Mı,K��t��bX�'q�{Mı,K�罍&�X�%��I�5�S��n2b�fg&�q,Kļ罝&���"b%��w��i7ı,N㿿cI��%�bs�=�I���1�����5e���lv[�_L�g8�7��bn%�bX��=�i7����LD���i7ı,K����&�X�%8�����������fq|q3��N'1�{Mı,K���Mı,K��{:Mı,K�罍&�X�#8���Q�2�'ke��fq|q3��,N{��i7ı,K�=��7ı,N��4��bX�'1��Mı,K���h}�{�}6ܸ�!�b`�x9nA��J닮��V�΋[g��2���:%]nA�/f걍�:�V��''/CZ��X�Mx��d����lp[z�e	�P��v�h)5)�3�2�cr�V�6(�<;Y�p�=r��u���ƣX��\s��<��ډ�%��1�w�g\u�¨W;��Z��Z<��[���q�n�q�ܑ��h�y�u�M���v}�������Q����q�K�ז ��n3L���ގ��g����UeJ8�b�D���j�-8���'���gI��%�bw����Kı9�w��n%�bX��Ol�n%�b3�{����^� ��s�㉜L�=�{��n%�bX��;�i7ı,N{��i7ı,K�=��7ıL���^	]����[3�㉜L�bsﱤ�Kı=ޞ٤�Kı/�����Kı=�{��n%�g8�����;Pʜ��[3�㉜NH���?|i7ı,K����&�X�%��s�Ɠq,K��9�cI���L�g�5�<��L�U�Z���X�%�~罝&�X�%��s�Ɠq,K��9�cI��%�b{�=�\_L�g8�M�褩�B֢��iԵg��s�6����86.LFr��$��웱ע�/=Zପ[Km�Ks�㉜L�g�}��Kı9�w��n%�bX��Ol�~A�[ș�bX����t��b���-�G����E8�U�7,�/�&p�,Nc��4��� @Z"
���'���4��bX�%���t��bX�'��{Mı,K�=<b�2�'kN�d�8�8���&q{u{剸�%�b^s�Γq,�LD����t��bX�'q�߱��Kı;�y(��6�(�"�g�8���Ē1����&�X�%������7ı,Os���n%�bX��Ol�n%�N&qo|����9`�9nq|q3�ı=�{��n%�bX����Kı=ޞ٤�Kı/��gI��)�L��瞯8F�$!)���Bl&��>w;Z�l<�A���ŀ�I�i�kW2FJ�	l�/�&q3��_���_N%�b{�=�I��%�b^�Γq,K��9�cI��%�bs���̄���9c���/�&q3��_���,��?(�D�K����&�X�%����Mı,K�w^�M������q{Cɼ���2Ȫ�Z�Y����'ľ�gI��%�b{����K�#! �$c#���		I# Fu�`F1 �HA$�
�2f&�w���i7ı,O�z�ٜ_L�g8�����9im���Mı,�D�����&�X�%������Kı>�o�i7ı,K�������&q3��7�|�_#*�Gq�i7ı,O��zi7ı,O���Mı,K��t��bX�'�}�_L�g8�t��Iak�
��nnG)�����8��SoNݺ�m�-T�����Ʒ<Q�`��������ow���Mı,K��t��bX�'��z�7ı,O��zi7ı,W��%$�HԂ�2�����g8���ﳤ�?,q,O����I��%�bsߵ�i7ı,Os��4���s�(����/��_�ZQ�,�[��Kı?c��cI��%�b}�k�I��%�b{�=�I��%�b^s������&q3��]z��2FJ�	s�&�X�~R"s���i7ı,O���I��%�b^w�Γq,Kg� D����( ��Oo^�4�8���&q~�|}AI]pi�YL��Kı=ޚ��n%�bX��ﳤ�Kı=�{��n%�bX�w��Ҿ8���&qo�<6Z�$th�;�8�/��v�����pbkv��>1��8���92Lg#vEc��O��L�g8�����n%�bX��=�i7ı,O��zi7ı,N{��4��bX�'y"���Ph��m��s�㉜L�g����n%�bX�w���n%�bX��Mzi7ı,K����n%�bX��=�$��|����g�8���/����n%�bX��Mzi7��
�1/}���n%�bX��~Ɠq,K8�Ūx��*hv����/�&q8�'9�M&�X�%�y��:Mı,K�罍&�X��T���~����g8����������r�I)�[�bX�%�{��7ı,?#g��cI�Kı9���4��bX�'9�M&�X�%�D_)?4�R*B\I	$�����"bm�*c������C������h���V:#�S&+$h��b؜+ͷ]��g��vj��ۧ���=�<��L6Z��x��g=jv4jѰ]��5�r�݅�N���4g��+v�{w"s�R�,-e��YzK�)wa�h(g��:w�k<�Yn�n��ݢ�H"MȽ�M.��ݺkZ���+�����&qr^��w���=�=��M�M졻J���Y�C���/b�Y�3�՝9J���u[�X�\	-��L�g8�����8�ı,O��zi7ı,Ns�^��,�&"X�%��:Mı,K�:���+j����rٜ_L�g8�o���? ��LD�;��_��q,KĽ��gI��%�bw����K�3��o��)+�;a)�_L�bX�禽4��bX�%�{��7ı,N��4��bX�'���4��bS��_�����b����Jg�8X�%�{��7ı,N��4��bX�'���4��bX�'9�M&�Y��&qoAj�> �%�����ı;�{��n%�bX�w���n%�bX�禽4��bX�%�{��7�L�g[��UY`I�j��,&Q�/-�"s�$+��hݷ��ح�tZ|v�m;-b�&L��Ɠq,K���צ�q,K��=5��Kı/;�gI��%�bs�ﮓq,K��'��/������/�&q3��_��<gЈm�+�13��{��7ı,O��z�7ı,O��zi7�"8�P�g����9-�59-e$d�q|q1,K����7ı,Nw=��n%�bX�w���n%�bX�{�^�Mĳ��L��|���V��U�%�����%��羺Mı,K��^�Mı,K��צ�q,K��LD�}��+㉜L�gb��ܶ����Q���X�%��=�M&�X�%��|k�I��%�bs�����bX�';���7ı,Oȋ�OB���8�5�:���'3V:���^9��o>mmn���ô�9�R�5,�;a)�㉜L�g}����Kı9��zMı,K��}tB�H�s��j	 ���d�z�cV7j����8�~��,8�p�,Nw=��n%�bX�s���n%�bX�wƽ4��bX�'y'd�&� ܰ-�r��8���.��<���g���צ�q,yȋ���+�2n&�k�5��n%�bX��w�Ҿ8���&qn��I��j��e��^&�X�%��=�M&�X�%��|k�I��%�b^s�Γq,K�LD���8�8���&ql?��?�ڢ$�;Ks���Kı>�zi7ı,? �w���'�,K����I��%�b}�k�I��%�b_s���C9x�i$ܻ�Q=�а.a�ncf���-��[j��;=tRn�Ds�g<��w�x�,K��t��bX�';���7ı,Os���n%�bX�wƽ4��L�g8����K[�X�N���,K��s�]&�X�%��w^�Mı,K��צ�q,Kľ�}�'��K��C��]��������Q�7I��%�b~��i7ı,O��^�Mı,K���t��bX�';w�8�8���&q{����[+������&�X�%��|k�I��%�b_s�Γq,K��s�]&�X��Q� �!�D��ߦ�q,K������8p���Jg�8���'�ﳤ�Kı9���I��%�b{�צ�q,K���5��Kı)����[�&{7����yF��v:�kq������us�!ll���2�l�7ı,Nw=��n%�bX��u��Kı>�zh? �>���%�w߳��Kı=����vBff��3��c7I��%�b{�צ�q,K���5��Kı/��gI��%�bs�ﮓq,K��'���.3�&1�\�9�Mı,K�zk�I��%�b_s�Γq,K��s�]&�X�%��w^�Mı,K���g9�f.e䵔�¬���g8������/�&%�b}���I��%�b{�צ�q,K��=�I��%�b}��ؘ�7�c�"����8���/ݾ��/�+ı=���I��%�bs�=�I��%�b_s�Γq,K��w�����w���--�	PȆbFB-�Đݥ�i!��	�`��F @(��0D�i�D�����h�c`�:p�cX2��J8�
֡,%�d-)��Ĩ��CC̆T MVV5�\y�b�p�����E�HZ� �
�R� )�k&[��lP��K�0@S�S/��	ar4�I�F��P��� �Y�)	��&�q���T�[j���qU@Up*ݲ���[�S-ۡ�����ɻ6{:非���c<l���$�X�nP�ړ@F��Q]
�؞��Y�K�5T���K���%r�*����,����R�]mF���v�>�v��D�!�Ya��jnp�}��M��b�b%O����z����G�ZR���M�εn�nǛr���F��p�eq� ���{%��-��0�'5]���;f�ܻ7�[��ΎN�*���g<��^�\	õ*[�`x�L�q`ہ�Ut��gaxu/0�4v�w��S�O;�(/kn��.'�l�UJgc���p-�-�f��ۇ6H�Y�� j���rڝK���F�qZ^H4�qYJ����L�+\G$u��s�Z�6�ԫ[��Iv��m�!�ȵ��dJ֪�y敓�qڃ�n)��e�h�{G�͔���0��H�7dQq7n��^�B�U��U�d4T m#ܚ���dv��a�q])pYVV�uļnp�`�ڐ���7[uB�3L��j[C���e�N��*�YYQ���A��X�c�j�F[ٲ�9���}��J�8�g��}xE�ć.��.BS>����a<�*2V�n�0c��{�]v�`��u��9�;����XX�2�օۅ+s� �vjWrjl��"n���Wv5�u��9�V�wNT^tg��j�rZ^�u(`�]m'�[�t�%r-��<�m�3�=j�U����j� V�*�[�.�-p�9Ԏ�n���iy8��/bvz�ĹЀ��<�*��D�Y�S��L�WN��lb��-s��=���{v���v�O
�H;�dq�Ε�h�]�W���.6��e�)vv��ݐ�f�[/�`���٢��i#nxzɆ�k���vmS���PS�U�l���W�����|e�G��^J��8n"/5n�$�ӷOf;x��pT�Nx(vؽvZ�&�V�3�䮭�5m:������$v�f���HeS�q� ��F�D��P��`�P�p�:�U� o�\��J�%WTg��$�¸Ԫ2�U�z�'6�%C2+̕�[�l;K+�[�ԯ��:{2���y��w9%{�N�I�n�S���콤l�+��n����yG�7��,{k'�cc����@��#&�Q��NJvL����ݟ�+G6�&/2���iT6n����������j6ֆ4۱����Ʉt�#�:��g]��κ��c��w��������X#v��A!�̎�����m��v�֏�5v�.wn+��щ�Y������Kı;���4��bX�'9��4��bX�%�;��7ı,Ns>��n%�bX����1��\�NXZ�3�㉜L�g|��3��%�b_s�Γq,K��s�]&�X�%��w^�M�����b~��A��$|,j�Ee3�㉜L�g������Kı;�k�I��?��������i7ı,N��5�i7ı,Np=��V�	le�;-�/�&q3��]���Kı=���I��%�bsǵ��Kı/��gI��%�bwM�Ϛ
�uYk�S8�8���&p�;�M&�X�%��zk�I��%�b_s�Γq,K��}�M&�X�%�]���F�B�
�jj	���u=p󁜫7<����֎�d'G/�Nv��J�r��4��.s4��bX�'<{^�Mı,K���t��bX�'{�z�7ı,Os���n%�bX����˜�ɗ͙��q���Kı/��gI�aE�"@`�g��PӸ��bc����7ı,O��~�Mı,K�=�M&�~\T�K��?BI�v9b(�Inq|q3��L������n%�bX��u��Kı9����n%�bX��ﳤ�Kı=����T$d-r����g8���ۯM&�X�%���צ�q,KĽ�}�&�X��P���k���K�&q�>���"r�W)�_L�q,Nwƽ4��bX�%�;��7ı,Nw>��n%�bX�{���n%��&qw���W���V �M]N��Ί����N^������UWN��H�q��-nqL����f�q,KĽ�}�&�X�%���^�Mı,K�w^��	>���%��~5�i7ı,N�����)Q�v�e�����&q3�����n��"b%������Kı;�ƿM&�X�%�y��:Mı,S8�u���V�e��L���g8X�w���n%�bX����4��c�Bd� ɘ��{�~Γq,K��ߵ�i7ı,N�z��K���ی��2��i7ı,N{�^�Mı,K��t��bX�';�zi7ı,O��zi7ı,N��ǋ��ɗ͹��q���Kı/;�gI��%�bw�צ�q,K���צ�q,K��k�I��%�b}���ؓ&s�\ a`��{M��V�g6�:w6�j�u�ϣ�㱺�J�DL=�;}��oq��%���^�Mı,K��^�Mı,K�=�M&�X�%�y��:MıL�g���u�	E$�q|q1,K�w�4��bX�'=�M&�X�%�~�}�&�X�%���^�Mħ8�����#�NXH�Y���bX�'=�M&�X�%�~�}�&�X�%���^�Mı,K�w�4��g8���50�J�m;������Kı/�ﳤ�Kı9�k�I��%�b}��f�q,K�.؀�.A�q����I��%�bw��ߕ�����ݷ8�8���&qs����q,K�����&�X�%��zk�I��%�b_��gI��%�b�n�qWic�D�j�QF�N�d��6v�,��:{(>	�Y��o6Z+�j,tݜg78�n�q,K�����&�X�^{�x���\�f��:����[cnV�����u]3��M������}��� �����-W�JR�J`��l���Թ�%U�5�دFBl�Ŏ�+���%�^�f�{���U� ���0kz-�2�ZG�c�#�N��t�\�K�^H�o�o���u�ҵH�����ۨ��Ѹ���_���h�Y)Ŋ)�;���ڗ[�S՟:d�Í��M"k������m](J�Ƕ���li�W���CZ��g	��6bwTS�p�m&�l�v�'��d1��6{5��^������!]��o2�7f0ɶkwAl���'jtK�Ж�rZ��OK@��{l�6�w�lۍ��jcmݏ���=�:>�iz����W����sn8�A�v'8���MH�S�:�Lj�;4턖U�=�����v`{ݘ��ŀ}ө��'Zn�X�T��̝.%ʢV���u�z�%L��k~Tu��a]���_�� ��:`v�A���1��tk0��U��KWic�#�N��t����$�{}0�����r��#�`:�}�s�0=�06���<���@�x0�"m�y�m��ض��ҁϺ���	̳�N����pܨ��U7d�I���:tLwGL�J�&fHW]�"K0�ݹ�(�?.Z=�t��Ԡ���L`K�T�)faBKn�{����釹�q7���`�}p��p�N�H�XTP`z��0�����uXG��c�V2RS ���0%�l��|��b�;�K�׽���Z�U�h���ÐX!M�����s����I�r<���K���e ������^׽ـ}��lW-��Ζ��:V[�"�b��+��������`{���:�L�?'��4)F�[-�`��^�1��O��d��B�HD� J1�D`8�����a"��T`��n��jI�{��o�Ψݮ�^KY]$+�>���{� ���Xw�׀�t�7\vW
8��[�t����ND��:[���լ�7X��u�\jQYkVl�;�St�3n8�����Ŏw6�'M�ڻ^�Α��c����"[ݝ/�}�Uz�_�� �t� �*�D턎Հw{Ilvt�\�wGLq�a]����İV��gK`uΘ��tu�w�ׯ �?CY�l#�ZY+��8�*mͦ�֘�u)��'8.#�D���=�n�I��x��jLd��Ui%w��\��:[ ������7�U%�-�tU� ��ل����9�uh6�n���=��nl�j����G%_�m<��;� 7{� ���X�ۨ�++/%���
���lN�����'"[�UUM�������F��o����'"[�zc\���*�3ēӣ���l��?W�}�&����7�{ �NV;a#�`r%�:��0	:&�GL	ZW��آ�g�B�B��K"d��g*����:6�'�Y�\v�]��j6�̈́��q��I[�H�c�v�և&��ˆC��N��#��p*���!.����nT��m�`c�i���Gy�A(��4�a�����zXȝ]B[��AI:�λf�tpVN�[t��=�n�� �q���sY��:���v6�(�W���xr��A#����*���YZQ����ϵ�X5[S���B�Z�mݹ%�b��۞�ӵ�	�M��o��<m|���,�Z����0	:&�GL	�\xy��l��e�If w{� �z:`v�r�{�[үYe�V�Wx������+���ޘ��&�>��ڭ�v�;I%Xmz��d� ɒ�}^ٿ�۷�*���|��J�^Z�^��Ӣ`ztt����1ym�qy:���m��vr�klˀ��`����\tG#�IȣS�icM�wn-�(�nY���@���,���@���ـ�Zjx/,�GhIm�>��F�*��9E�wZ��ԓ��w�Nov�~&�n��v�Gj�;����zc ��0=::`{��2�W��YbX+`u�L`:&�GL=��ۇ���qzF;m�If l�l������,�`e{'Xŕ�#����;�����g�Bm�9zM#�1�Ia�t�\�,9��b���������L�S+�;��ٶ�����Z��v�J���^���0w�p��� ��w�v��ګ�13u$���Ƥ���s��ɠVM�p�����JB��,�6��)&���4���J&rO��٤֥d5JFVXHHP\-cD�$b�C����8#�5����%�@5CFZ� Y�O�u����B1X�K���O,-�>%�`�`�c�����\�2��!��`�����X! e!B1�!`�����$	�K��i&�}!(J��+� ��R��� ��2�$�0��L0Fs�3 �� �>ᬦ�F��$"3^d @�nMd(��.�re�"�X ���8�>`���4"�)D &B*�%�в8�&�u�C!PJm
3E�|������m�M�dULA�@ Ea�\���	S��!�*!�� @�� ��!5@7~��M�8��1���t��P�(� �@��q>2�z�D@>z��1���H����)���um}Oﾪ��<�'"[ �Iw���;HQ�ܳ 7{� �{����^��Ogw� ��xN���"��ǉ&�GL	9�{��t��x�n:�X���U����N�8�r��k�9�u��5�gr�H�@�8��H5�RfZT���-�׽1�I�~�������b�?{[j�AZ��Ec-�x_��0	:&�GL	9���J�������Y���I�0=::`IȖ�>�v�_�uR"���K-�>�cL	2�L�d�q�q�s�H8�©@P�k����'|c��7��YZv�J���^ }������>�w��q���4z��>�ZĻ�Y��$&���׎ws�����	w/]�ͫyYymU���۾��ݸ����_0�}_� o�x��7S��t�۶&K{ĹĕQ��sn��~��^����Y�VIm�>��&lW-�wtL�D��3�ȨӶ;V�����w}p�ݸۻ� ��^�J��R�-�x��0��GL��l���Q��$�Se���Ȉ�V����P�����Y��L;��?n��5$�Jɭ����c�="[������q������ȂcC^�HI�h���H��)�i,��֤Q�(`�#vU�n����S��:H5�8[����n*�n��Ө�&����w�@un[���p�Vu��y���4�;�wPey�.��òo.N Ș��`T`��~�������̵���rg��Ů�g���NK����ӊ���G^N,���t�,vjc�x�}���$i��,��I~�$�l]��9-�F�N�\� �wq`��^ w�ۀwgu縛?jڼ����%i�I*�7�O< ����;������ �v�V�7ymU�B� �{��&t����r%���Fe�b�Uf�1&���r%��wn��t���Q7�Z����5��=�]������鸯nt�ޚ��(�g\�V%�/1+`{z:`IȖ�=�vw^��nm����H�X�s;t(|@H� >A�t�dƵ��$Ζ����ӂ��+]Zʴ`%����cL�lwGL	9�����YD�������t��#��06�)F^%`����V,V����d��D���3 �8��Q�y[tB�+t�K��&����O����\𻗄�:(mٱ�ۧq��c����;I%_�{���ۀw�u�ww�v��U�9j���������-���d�BL�2������x��ń��=�ચB�?}߽��Ԓs�z�f�lp��]���� �����0`��$��DdVZ*��I� ������>������ ������ɕ��u8�5g
s7b1�n���5�n5�k{s`���U;����
���� ~�v��t�>쎘H���n���K�ĩ`�&�����4��Fْ�/��o�r���S�%��}�X�� ~�v��t�>�u��:Wo��T��F��`ImU}\}_W�I `A�ڀ�Q:�_��RO��H�,������C ;���<��?3u�IqK�3Y��-Uێ ��Y���j��73E��c�����x�δ��uF؎�Pk���s�YZ�m�{��=#L��7����6�F�9\�$v�l��n��;�u�����L�8�Ĺ���ޠ������h��`�_# 7�ۇ�{�_��b�>�*�Z��ԤeF�ʭ�m�7oF�02K�`yx�U��ىR�bL�A�6GL�J��|/����ATY�]�)��~����#Q�T�m�K�H��$�Բ�n^l���xP�z��<����l�춓z�eW�݊��X	Wb��l*��v.��b��M&�ЀOcKɣ/\x�3S�oC)A�ښ�;��n���s�q�m�lX�΅܎�J�#�۴f����ݎ"�Փ�[����#����>��Xؔ��Lk&�׶�Bn��j���6ə&3��l �����3&&n����Qm�7FzXf6m�3�-nnˇؚu�H�L�'k��T���%N�����t����N�"��:�Q���x�nJ���F o{� ��� �۸�ߎ׮��+/"��%F otL�A�6GL�J�܊�0�V��-���P`M���Q���^��m�,M�cr�)�OH�$��3%�2K��%忿���/Q�^:mFm�������<��]����*̭e:��M9ۑ�L���݋���ݽC ��l����H��(0���F�T0�}�УH��Ep��Mk��ԓ��tjI�ۨ�?/�:���+RZ��[�wv���#�H�gD��9JX�fX��Uk�:`t�P�6tXwn�ݝoQ(9ev��ܕ`�J�dt��%�YJO'����q@��Y������s��oG\C�ŧn��G��nL�����;�`wE�06E(`�rUD�J�d����0��� ��u���^��m��D걹m�`M��dR�g���߾H��`vŦ���c���U�~ݺ� ��0;��l���@)����b0���`�&�A�6GL	�u��8��}u9%u�e�j$ק���5�)�yh݇./E-\��q��!�\R��Id���=�o��X��F o{� ��T��G%N�\��6GL�JΉ��$��:ޢҹl���ܕ`ݺ� ��ۀu�����V˥��WK��#*�$��0r�a[u��cH�p�`]�~�4���Eq��S�:9-�:�v`�`d��&d��%;ͭ[A]�ۋ�[����];�4ӷ9�=�9�<\6���@��Du�w=:AuO�m�����.!�L�{���V����֜���J
�V�ۨ�.&�۾��{� �۸�͟����q���`���}&0&�遲)CW��ۊ�$Q�[�w�u��w�v�0{ݸM��)F�$����t����ԒY��Q�	7���r�I�EQU��
����EQU��
��PU_�"����EW�H*���PU�
#��H��H�,�"�",H�,��"�� Ĉ�* Ĉ ��������EQU�"*���UZ����TU������U_�"����EW��*�Њ���������e5����0�%�� �s2}p9|
� ��(���B�P6��* (e%(
(P  P)@ <>�*� � ��*�
 E(*J	��U "�
	HUAE �	JU ��EPD�P��   � $ � �  �h���N�� � S��fJ& r�9}��W�J���R�� gJnϽ�����  �I�ån �ޤ2�����=��i^��} {�_q>�{y5�NMW�ͥU� 8}      
��<�[�#��{��|f��-J�� �uO^N�ӗ.C�����-W@��J����x��� �^�94;� ����A����ɻ����1w1U�1N�[���o ��@�B� !��ҙ}�_Zr���t;��N�*X��i�J����� ���cn��0 2��@� ���;�zL�q��-�4� ҙdS!�d�\���p � J(    �A�ޠɪ13ٮO�W8 	Ҭ�.�]eŇ��ӥ��P=�J��:r�|j�Һ�[�W  �}�G��msۧ��=��Ү�� ����}9t�<�;t��/{j�  �@z 4 
 q�@��˛}���n��,�[�x@�O���S���  h��]�n0Ph�ꇥ�P{AK�    S ��@;���4�  4���:
8�M�t�>���zP� ����@���©P  z�f�J�  �=U*�h   ��U*M�UA���hb'�Jl��@ 4 DHSeJT� Ѡ�3�?���J�՟�F~���j�ffS�oC�o��@\?� ��*��A U�A U�U�(���D�-<z�L7o��z͚��9�~����r��)�sz#��e֍f�͜p�3��p�O�6H�!��ŋ"� D�4]"8Glb^�iW���`"-"��2��9�%�m�#��"
��%(L�:Y$-�%��\�.��}w������&I�H!F���4�B�SXHh��&1�2���7��\&8@!��l1R�������%�0��u�9���B]�r�_���tR		$.J�F0�}�7v�:�E�l �6���P���7���;w�%%�#��q��Ss�J�#f�Q6�@����̙Dp�34��3�IV$���-IV��B0�	��(F�B��IrV�eʅ����	 �X���|�sY�L���� AJ�b�E"h"��ćD��)�NRԪy����/�Za}ըH@EUO2	5����<����~�~A�����q���^��KV�z&_�ݮ���ן�8f�k�0���� ��C?qz�al�)��\]Zɥy�!.BR��!���$�I'��q�?5���)�S5,#�-�"CL1�ta�6�R5�_�p>��Ц,�Y%HՍ�vK����L P��ߍ���ЅhC�W#cX�6C��m�IXS�3f�A˭ܻܐ�"l�����WyyOe�e4��^� ���%a`FX��	��o�d��&����~H3�pۡ�a��\e�o4�$$�I�˃�W�
�悑w�f��{t��"%	%M.^�]���Ѳf��F�6���2�	����z��P�j�
�B�� �c`V� K�������21`id"°���	sS��~:�駬i�B�i��:.UeQ��8r�Ϸ��'�)8	��IU�wV�
����[u�՝|���ݐB2' B5���!��0tm$��1Y 18H0� �e�'�}�C�\�B	%
��R@�BH�B�H�R,�BD�}��A�
H�����1��w/iК	A�lMBB�*�E��!V��`�D�r���?K��� U�SP�JBjp���)��1-/o�ǵg���1���l�Vf\����mIX�ǡ��QR]5j�R^m!6r����6O���d��J���~3�+����CDF߶����^lꊄ(�	��ʠqt�ĩ
%kH� S��3)��a�nHnRe��N8��$�T�a!+V$D���0X$Ѓ�%t¸MH\aX� �aH�Xĉaa�'{�J��n�3����e'��SSW�kS?�����j֥����Є$�ߞ�>e�7f]��k�/5�@�B�����+7�˙y�
u�m.�2	T@���F$0�H�"1bȌH�\��Rc ��\�ʂkv���ҁT{}i�.Q*�4or戌`l 0���8��~���MXp� 5R1�X-��"IґJAH�"B �{��$��ՂUq`4����	$Hm�g �SZԀ�Z���:v��B!��z�Lѐ��(��P�I:tr˨�Iɟ|�B�,����l	J�B"C��z)	{�Z0��ԁ��`?2�H���,.|B捌.�!&�F�3[e�F�7�%�l,f�M������&���SW��K�W���MN�9SI��D���Ҟ��.�+����EBuh�dn,�/#��Ɍ��J���Wj݀]��U�夥+�Z�B{h�5]�{a�V)�6�H�"�kī��B��E9�>��;�����x�k���%�!.�Iy߷)�۸	`B"a���G�?�n����_�4	L$�A�li8��9!h�$JP J�vĤ��Ez��=����k���T����!��$J��2�t�\����H�3��,�Q��nJi!�Ho\��cDa�ٚ�8Ÿ���\��C���Y�O{ZҔ��J%R���Nz�E��Q(R
%����^H��-�i�0HVt��ˮ~�Np�~�j��U7y2�YZւj	)]q*�ݪ�Ǝ�T���}��|f���"hi`W�D�CI��C �ЉA$d���\X�F+�BB_���ؚ������P��81+H�J��K"�b�k�'Ia�����8��0`L#
`���H�@�)�h各L��}/ƶp�u�! K���mb\��"8T����B\����·L���7'B�Elvp�2\#���9�Ne�U�v$	-���^����s_��>4�� \ A��T��3RT�\z�z����d�A�?�(�.��4Ө��D��0ن[>�f��qk��"Q4@�i�\"�A��~&1�ۆHe$5��SA����'�J�/�gQ�2�&>|J�]
�v姩M35�^jm�ˉ2C�S��8V���0!�l-�n��ys�sj���B��B�j�U�5�ez���uD�X]m�X��ؚ^SJ���S�wu|o���B0��$0%1�30�P(���w{� ���5�>W��H�^�t�/Q4_�0��Z�]V�B�^V���bo�B���Q���)!/s8�� d.f~���&~k;��h�WGc��%+�5Zլ�� @���w��)�+*\�da.��"K�.i
p!q��7A��5�Ij�*�J&���A�֥!L%(A
�"��BZF���h!�T�qt��!:!P�7RP���h�+��;�l�%pBR%HDؐ.K�kp�oA�F r!2��s{������i�c!V!�/ܷ�7��\�����k�����~�&�%#��~��h���w̕w��z<�(S�v/�'��?N�"F��#cu����8kG��S10Ig�Y��?|h�D!�Rz����N!{�� B���T^%h	�HR��u�2CwT5.7�ff2������B\XRP�7���M�C���ᄄ1��B�!w�����k��2.�)ɑ��V��x��D���ּ��?i�.�^n�8�7~e�:����럺O�w�#�"�����ˇ#�f���$4C5ąrA �!d
`�

j@�! �
6���[��wJa ��
���!�o���8��, b��� |�BB,F!�H�|�!Ioɣ�F/4#3F�;�I��� \!\hQ���5
���0��x~�T�$"I#$a�\��as{&��SC�Ɩ�m����/u.dX��Ab4�@�����*S,cA榭���ٸT!R]���e�u!�HFJ��Ϗ����vC��a3%�vB��Ƴ99!�p�ja$��A+��o����D���7��9'٬�o���rRQ4h��Is[%\ٲK��7��71˭3z�����%�k=J�/zȁ!	!�Y���Fl�HА!Ђ1�E!, �`!d���%# "	^�$J� @�H0�B$���p � ��@�F�Yc%�3_��_���F6�X�xB<9��:�m7��R�(��4�f����bZ��h���1�J1�*Jabe�H�_ц��+��"��Ij�K�B�Nh�	��J� @���3��&�А@"M@������6'灍	ɟ)EfO�9��!"!	-�{ݎ*"@�X��/�W��\�qٳ}����Ɩ�K��H�mNɋP�a!Mi� ��/$=�B��+��X�RCy�����A���?sl`��ԍp%N���!LD�CI�q���ys�����B�Ƙ�b�p`Q$0���7�����@�
c����0YQ�c5XQ.:�ߥ06(��B�*Ra�|�FҌB�h~ 5�H4D�}���D5ԁÿX�3GO���G0�o���A!��5��h�$(F�]��i���?��)�h"�������Jt�CD�F����)�j�U
c���31�y�p��.�۠��rԸB��4��@���Z�h,&`h�W�DB
@�q4�R��u�D�l461���#\a\&�%0ԡ���ĄnkjB�i���YG�,#!�����SH@��
`�$h�1j1Z�JBE�lX�a��$(��A����,T�E
dR4�sZ�$    H�m�� �@   h6��>�� Z�dt��89�d�WU@R��
���` 6�:�2F�P�n@Vꀪ�ڨ
���� m��a���-��8�n ' m N����@ �` 6�mW@�[B��t�j�M����ͷ%ҪnN�B��H�p�k�-�֒����J�T�MV���6� �RD��w	��d�Z����F�ۤ�5��ֶ� �l   "C��� ��}���Ѳ�-k�  � [v�Z�m, kY  �`K( m��m6�8� m�H�   ky�Cm1�[E� lH �  ��@ 8�I���ثj��*��G]��(*��V�X�T�U-� h �ۀ �� ݶ [I)x�@  IА  -��  	)ٙך-͍���Ƭ��a^���R@�����m�RpJs���[q��� I���U�S����@�z��8h:қ�g���:�.���`Ӛ���u���;��q�����4Lsڷ���g<<� y�7ݡz�6�.Ʉ.�[���mF�Uã����k�Q,;����~��OJ�6N7F,H�Y�`6*�S*��r۷g��K ��&ؼl������׋:٦�9�#�������I��[��3��������RU�� [m6�jI �\��F[e^��d-�d�*���<������vA�[dKh�vؒ�ڕj�
�����U¥��]uf�v�K@ H uK[lձ���J��2���K�j���4�H�p�Ā-����O9omϥ�R��wVm�lm�[@ �/n�Um��v�N�,�$���ۚ�m�GQA�v�	J�UUU�@�8-�*m���lOu�m�tm�l�Z����Y@�[w(�M�)@ �p'@  �d�
ꪎj]�g���IB�]�����cm�ԁ  6M�� ��` kmm�6��Sn�e��X�1��   m[ � ;m��mm�����   �� �� ��ֶ:Nݫm�N�     6�a�M�;��'�o}�����  ����p	 �� m��   6�Zm�$4Pl7I-����` �Q�5�Z 8
P (T�RZ�*��^X ���� l $m� 6��`$�[A��l-��k6m,��]�U�]��Ҫ�U�|  �� �V���t�2�U[G�    �u�n K�Ā  	Ӗ��&�h *ڕj�V��v旅�,��N`� � $� ��a�6��G��7�|���@X.��![;n�;:�R�8�[`�k�Ε��Vs [@Ib�6���$ 	���Ӷ�6ml�Zm���� 	j�NKNۢ�gb�I��I�J���j���O%�������ELz�kb��Z��9�![��*��V��d.vێ�
�s۫��D��֩ݖ�/¡��]��6��6���9)�D�R�j�ZQ�K1����r.V��;fs�fP)v'h$��<m{`z���ڕQ9�IWJ�^�*�mm�]@$u�V�.�&��6�jM���m�ۯbt[Rh�ٷH��,��֦��($�Ē��m�m���zI�� 	�mי�v�m��8d8��[׶�8�I��ڒ�^4�$ļ�4J�vz���k�����Q�n�˰9���֍��k��&鶍�N�2N��,�����3��֦��-� �5܂AͶ
Y�����%$�C�vۃ�튲�R��*���k�	�^@�n������khX֘qU��ԽLUiJM���-ۆ�V�Gl���+Etl������	x4= E ѹ����W-r�v4�UF�7c[	x7\-i��pn�(H ������^⭶��`eۉ]�w��l��82��kV�p Z�Uut�/	�)�j��x�e����N�tt�v����<���R�]Yxj�66)�FK��'u�g �8��l � Ä��$�8�L    ]5���H ��m� i�E� 7El	�0�:�U�Z�y�vVU趜������[@ٶH -��� �ŵ�  �Z�  ڶ YY77n�l�� m� �` �` l  p��i8ֶ��|���UP����U]*�nH�!��lp[R  $ �Ph �i���C�p�Rƽ&n�m ! �bJ�j��d&U�b�GU:�$��6��
W�L�T�]W@UUp��e�+�NIvٶ�� ����T�P�@�zm�	����ӷ@ JT���-sH�]�%]clcA&��3��nr���K�2%���X�4�tһ��u�����zΓur�mQĔ\۫�Uuv�F�)Nt�L�
�Xn��>a�r�j�p+�2����X畣�
	O9z�Ug-T�jy��kb��`y��j����j��VUN �ة�D@�khq���cZ�lPҮ�
�Ŗ�Pl~�;}�@�[S�VV����[v��j[�K�� �J �6ٶ�j�8m����$�m�` 
��ڪ�3�ˈT�rgvm�mt��O���t��	&�,�Ͷ�$����,�hi�� p٪�B���<���6Xp4�Kd� 8 @��۶m&�����.�-��Cm���첄�t�ɶĀm[ H�m� 8�J�W����ejU�%Z�$��V��U@ �` 'Za��섁�h�m"@km�$�NZf�˦�p���� ="E�^�+���@Ul�µJ�UUU�9�ږG�q��m"��$H�kn��r�C��d���U�ڝ���i]#�T�ԠY;Kd��%k����  � 8���-�mt�,�� m���m�[���	��  ��P��̼���`n��J6�M�[�2Ӌ�0Y�9��=U��� �[m��Kp�[Al[庶�j��\�j��2-�Xw �d�ڪ���{
��s;=��sӶ왻vz4s���:v㝺��7�{)4b޴�6P�6�l�f���:�@[g�){(�UJ�d���T9��MR��g.rY�Wj����f�ۜ������M� #j6��b�v`�
��5t���Qo<�r��k� H-�[�cm���.��M�   ���l hںM��v�  �3  	��]��P��,�Ҭ��j�`%Z�*�VVI͐�4��%�`�L��T����U2+P�W�� -� ������g%�d�`m �u H    �6[�H6��  ����UU*�R��<�����ju�:���p5�FΩ��6�� [f�:6�&�Ui�}kX�����:[���tƸ�r�UUJ���X�n8��ݶ����j�B@����5 j��Y-��}�t��f�V��H$$Kv�c�*�V��A ��yV��@8-[���m�N؝���uK�5S�W�*��G"��j9��UUu!-ٰ[�+C��F��g���檞UV�9A6*٫���7"5]e���d��Z(�߯�o����V�UԪ�O%���6��C�vW;��J
8����  �`mP#� ���v�+�HUt��Q�e�ʝ�(��r��Utkiyq��hѺA�).z�@���Ļ9N�l�Ҥ^����� [@�!zKe��Y�� C�ݵ��Ij�Iv��w,�Շ\c�+x�1W)�k�*�����[�� �K��k� �@��F\)om/���'Y�OT�O+O;,�5Tq��·�Ɨ{t�7��UFD!�j���8#i6�9R-6�'@K���d\�m%�fl*��t���    [;��:5l^H|�Tq-U\j��m���ݑ��Hy��^��nnˎa�/`�]R� vRYWuW'fn8㍷B�*�۴m^J퍟�6�(rXɰu��Pi�v
���=oQĢ�6��}U+�+&{6΅#�\4��JF�y��b@I:k@K��j�nQ��j��UF^�q,6��mm�m��I6��l�v[GwY.$H$
Q�7IRl �d�l7e2�6�����* [T��Æ����y���]$ض�X�l �m�  �  ��۴n�j[�| 
����K-2��l�*� �M�I��&l܆ Hp>��r� � ��U�֫g��"jU�ګf�   Hm�  8�H:EY#����� ���  ��h���S��Ы@@$�Jv��� moP�@�n�h2E�Mt�	�e��lm���%���  lp@ [@   f� ���k	͵��ր7m�$��8 '@     �YE�m�     �7����l���x[��m��l�5�����w"��H�������E`��T���@��"��@G�� 0�� '�T?*(�Cc%Atf(�T�`�B�!D�M�)�Pu�_�?
�8��'yb(��E �#�"��/Q��C�T�%8���zCᑑ�$�����m1 ���g�4?(���P_����.��>��@"�GH� 0` E�) �	@�~@�����QE'�����L_� p�i�UM�(�i�~P5񳀀qA�@�.(`� ��W�耏�N??C�6�� �N*���8��H�hC㪅j��T�->A>D0���_� � EQ�0E�)<E�
�G�' 5�#�� ���`��(�
��Q�QW�LSLx�q��\,P�����~ED ������;@��{ (�?
O�?-��@$y{�5D�	������u �A���@���'�� 
�(��Q�EFE���B"c0�������� E��G{��_����u9 j�2>j��wh�t�˃S!#�MK�p��=�x:�#��z�;&6I�ݦ:-��V���h[!�`��H��,M)�*��@, ��'Z��n9V[�P e�UW�vX���q�mm��r��g����ۀ�Hv��Ypm]��5��c�E�훨��cp9�fɓvی�:�J�v��@\����n3�K��]��8�.jӍ�_0�mH=��<S9�]#����*�
U�2��R�����U�\���U��Dn��U*���k�`���GR��n�@�Y\���gEʗ`�^�+��\�R[B%�$f#m����/'B�����:1�6κ�ӵ�Îhnm��ۆ[���v�`r:�h�ʻ���:5���k�Š�ͳ����pҝ4�޺۫!�N�p�n�'#�+���[�/�sg�!� �\l�6G����	�h��V�WY�f�3�6�\��\��r���յ/@��ڧ1�m9U�k�gm�K�u�mm0�MmL����I���c1<�@K��e���މ4��zv^詎�2$zWd�8�u���5��� 9�!�v9�`��b��e��d"k��C�c�=8��<�mcjeэ�֣�j���W,�f�h;3��ۅӹ�g
��*��Ǎ��Z����d��)��{Gev�Y��PI&I���ضK�a��duӢ�[�<���#%u^�$����zl�(�P�6�i���Fm�0��$��Y�5Ö�U�����D���xM�T�{m�ᗮ�Y�nD��G@�]�KNR���G;�;-v���N�[���&��.9�֍�7F�j�� N-�k�Ќ/53���:�`ݱ��9�H63q��h�-TsF�駜��Gn�nN�-	��vqon��[.�n@�p�Q 'JY��.�1ђ�hۮ���7+p�T�� l66R8&���j��x��Ft��j����DLl�!;����0T:Ԫ��MY��3I3�E�&���X�����l@��T�>b�����;  8	�h�=������H6.�bu�p�̕(P�z���M��u�l��m$փN�ӄ�6��"v��A;M��n� ��͆:��mp�:�,�tv6z��;;S�o9,q��g�u2�ݥ�L�rѶژ�(d`���z�۬��[��+�\� �Ojx9e�9�=y����O7mLd�u�ܨ3Z�p�n@�dA�Ck�Ս]C5s-�W06���P�y�C2���\q�
��ϳ��=��Gʎ{n�m�۞�Nɸ�ϔ&LK�����
:�J(A�޸[�H'�f}h�="X�'��m9ı,ON��2x�-�C2\�LMı,K��ٴ�<1ș�����7ı,O�{��r%�bX���eM�R9H�#��{�Sc����RB�_	bX�'{���%�bs�{ͧ"X�%��n�*n%�bX��}�ͧ#���ow���ߗ,�*^2����ı,N~�y��Kı>��eMı,K��ٴ�Kı>��I
HRB���7eQTZ�ww��B��%��n�*n%�bX��}�ͧ"X�%��w;�7ı,N~�y��Kı<(�wrz�f�����fCR
�h��nuӫ�!�Ӆ�ݻEs�R�6M^�]���z�h�MffL�s5*r%�bX�}��m9ı,O����%�bs�{ͧ"X�%�ٝ���Kı9�}/f]�㴤#o�߭�7���{�?'�l�$Rd�BE'@���E�bA�A��џ!�9��~��iȖ%�b}3����bX�'��o�iȖ%�b~���٪d�p�5�5u�Sq,K�����ӑ,K��ϻq7��ș﻿M�"X�%���=jn%�bX��_0�t�kRe�W4m9ı,N��n&�X�%������r%�bX���X���?}�~6��bX�'�B�=�m�I�-�����%�b~���6��bX�'{���%�bs�{�iȖ%�bvg{q7ı,O ({���QFv�.��l�]��7]�Ya��:9;���Y,�^Y�M"��b�o7.m��պ֧�Kı=��eMı,K���ND�,K�>���Kı?~�}�ND�,K�:\;s4d�˦��fk*n%�bX�����r%�bX���n&�X�%������r%�bX�ϳ�Sq<TȖ'��9��əm��5�5�Ѵ�Kı=3����bX�'��o�iȖ*� ,�`" �P�E7�H�Q�K"w>��Mı,K����"X�<ow�~]�����*��h}�oq��K��ٴ�Kı;�gr��X�%�����"X�%�ٟv�n%�g)��ފG)F�FУ��9H�(�'~�v��Kı9����Kı;3��Mı,K��ٴ�K�q����,Sм�T���p- p���նCn�68�e��k�]��n�u�]՚�թ��%�bs�{�iȖ%�bvgݸ��bX�'��o�iȖ%�bw�gmMı,K�k따ΒMjL�j捧"X�%�ٟv�n�DȖ'�w~�ND�,K��z��Kı9����Kı;>l4d�)�L�n�Sq,K�����m9ı,N����>Ea�2'��ND�,KӾى��%�b}��p�A�@D��RB�_�r��G+r=�7ı,N~�xm9ı,Nϻ�q,K��+��"��y�vm9ı,O��;s4d�˦�ˬթ��%�bs�{�iȖ%�bv}ݘ��bX�'��o�iȖ%�bw�gmMı,K�{�*�N�#���P5*6S����/����; Nã�;{OJ-�B�y�\ :�kY���%�bX����Mı,K��ٴ�Kı;�����"dK�����iȖ%�bv{G��3Y$�fd�5�17ı,O߾�fӑ,K����ڛ�bX�'?w�6��bX�Bg[*��$)!y���Su2ֵ��jm9ı,N����%�bs�{�iȖ%�bvgݸ��bX�!n�3!x�$)!IG*e�TZ�.�5&��jn%�g�RD�����r%�bX���\Mı,K��ٴ�Kı;�����X�%�ϵ��C�*@����B������5RB���{�����|�`v�}?�puΧb�k��	��һ5��Q]uΊ�`��<`<�L���un)�0��,�=�p����;g<l�w,��o-�����clI�N��S�Þ�tu�݈�sf�1y��=�ci\�&�����!�����m:�p�2W۳�:`��H_��X_o����������˦�\�t����a�av�y&�.�����8� �^��?v�΄m����k�$�\9�d�����u��4��v� ��d�z�7����~�����|`i��<���7� 7�]���!��Iq��ʪ���}u`{}�;�K�[�Zۈ��6����� |�,����npkj�5���.f��ɚ��� g��~0��0��X�<X}i�Z��Tm��MIVw&�Vf��ͺ�>�۫��W���^r	��q�Q�	��a3H=��:�1�"��9�ظ0a�;�uL�4�"�ir1��Ż�`}��V�yKY3&L�p��Ҁ�k���2�\�E֡�3Y�';�vl�1��.$Z�{B�p-`ItH�7�p��!$��G ��mv�L3&�I�zM��*}���ȭI�;�״���Db@G*����Vw&�Vf��ͺ�>̤rS�!�j�N�`}�J_<��:[��>x�syV�KYZ�q�)����:�5�|�`��`�l�94�ԲJ*��44v^�����u������8�큳ݭ<�wC�t���ԩR1���r��`}��V��Xo[0��X��YWUD�%���`}��Vw&�Vf��ͺ�>�R��JrQN��ԕ`gri�l�:�b)�腋3[�,��X����$Rm �F&�`n=�`}������;zـo9N�ڢ�R&�Wsw8�<X��`�l�Ss�������ub&��_���C�HО+� ��{S���l����7�ػOkD�sm��uk�|�ذ޶`�ـy�ŀf�*��aM�M)%Xܚ_��9ʤ���}���3sn�������i"Sq)!`f����sn��۫;�K��Cc@�S�t���sn�|�`�l���.��1)/K�s�f�ӷbt&�C�U���u`z�$��ǀ;��<���=.N	Z�:d�+��������E-Ȑ���v����юpv{��.��=s]�n�����߆��0>x�m��<�]�ȥ��GM���٥�#��]X�z�������j�n�Jq	��#����ŀso�����`��U ���Q��5�;�K7f�ۛu`f�!���M$�3��sv�Ϟ,�78(J"�Es�r����;��d�(�T�P�v6���蹦{Z�c�d�v����ɬZ��]��K� �=�"���@[r8\�<��I�Hu���*��כ��D�l�V!k�k�_��)ɝ�F���Y1�ܗ7���Ǟ��󋲊�	0;��nʀ�[��4�2vn z�Й]�np�Tݜ;s�؜
n�θ�nq\�Y:���n�v��AR�t�`��a�P�FG�����w����������t���L�ɩ�%�DCj2�yϜ���c� �ꪇ\!)�9(��RC ��<XnmՁ��U��ɥ��[Z)JPM�A�Vۛu`>�s�v�� {M��mVU�Q4��C�qʰ7j�3�4�7�uXnmՁ��NJ#iӔ��Xܚ`i��<���W9�<��S.lV؂GM�������sn���Vw&�[��J�GR�N(�*IR+=�w1xl+��̜v�f8��n�7Q�jl��":�D�Vۛu`n=�`gri���s�ϐ{_����MRz�Q� �7$�����t?D" �@؈Q��z��7M��� ��UQx��4�R+;�Kq��ͺ�7�;�[U�'#IDSq)!�>�� �� }\� ��f�Mhl�)A79nH��6���y���\�@g�1�I�š�l�çu#ȓQ�i��=sٌA����l Py�	ɛU�:҅��(��M�8������;zـ=�� �� {��V��T�9I���ɥ��{���sn�ǚ����o�P�؂GM���?y\����7?9���	��qѬ!	@*\$��M%�Z�����@�_�9���Vl3!�����5����iXB�3!�Ѩ�����\��+8ħ;�L<�wQw8�� �5M�q@�! ��\��!}U��j�;W\�`jh(sW@9� Ca�g�Bzk0��Dd!�p�\�%"2�[�S��>`��qL0�� R��@ˤ`8h�"BB�e�5���ӎ�Sj]��CEl�hp����$�Y��)8��*@ �:(�4��QO�(�-�D��"H��> |
uk�C��D����R�/���=־�؃� � � � ����b �`�`�`���z\�MjjK�.�M[��y��lA�lll}�w�b �`�`�`���ߦ�A��C�R�A����b �`�`�`����\��Y�2I�ѱ�A�A�A�A�u�]�<������~�yg��lA�lllw���A�A��x��_����,F���V�Α�qgb���vQ�m�M�_�}��s�].�%�>�����
�%�wO�@c�2(��$��=��ߕ������r4FSpRB���ȭN�6�������]�k�\�Ҥs�nG����wf�{��K��Ł�?yXw6��N��C���T�ə>�֔�'J23��_'f@�ԙ�d�{��֨��<���%)I!`gri`v�\����w��1� ���*n��E�J�ֵ@v��t^��p]��ܛ���Q�M�C�7�����QB�$q��>u����sn�ݚz��A��Ł��T۸G
�q8��6��I���sg�u��;�i5Hu�F6��U��zx�/�8Q����6(nm*2�t�`0Q������nm��<�|��6����/g�Ł��ȧ�'#De'$({��S7�7��{:P�(Usꪣ�8�R�5�r�%H�t�9�����L�dX��U>^��������E�H'�T�����\����&���ny��֢�n7�-��N^�4�Mq���Y�s)�pѳ
������yՓ�rnd(��-�ʲ�5�u�;Ok�� ��V��;g9���Z��v��|6�;a�6v�#v�zn�5�6�e��Tr��k�wm��'�a5w=���;��|���ʜ�+��u�ʣ��Au���m�1�:�ϗ]���vR���O]v���t79�q�������,�M=ϐyn���zҐ�N��D�8�Xݚ_�76x�<�|��6������!IIJ#m�R�B�����ՙ��%�o��g���z�ʊla#�&�a���`w��{�Kqnm��77ʒw�@S�N;�ͺ��f����s�y�)(��,��Qx�n]��]:6�v�ݺ���6�I���I���
8�C��@M�$���zx�/�8P�y�ə%���(�Ҍ�)7Cdnw&��v����5KȠ=�8P�+�tA�c�QļLÓx��d�9�z(��
9���t�36x�1V�dM��cq8�?.�oŁ���`gri`j��`}��mʌPI�$ԕ`ovi`fd��ՙ���wn���wv�ʓ��i'I�����bt�7�vzv��a�qJ9��v�$ݧ��>~�B���F��#��=�OŁ�3]��fRԒ_8m�Ҡ9�Ξ��S91K�D�'�k�lW2L��n�*ov���K�RF��RN�'Ч�v�{�7$���s�H��	,%#TbB!	@�R0�K@$A]R�'��{���kŁ��>ǔ�!��`9*��?w��6�� s�� �o ���hT����X�4�=�=�?���{�K�W��Y�)H�d��lv��\�j���wu�7mJ��:-WC�++���V�r��6HRpRC�~^��`}���˜5�2��3'J�j�y��!*I�����>��U̗2I%wl�@n��@c��V��ə����DJ�H�R��5%X��fM,�r��������sv����6��'$,=Ż��ܓ���nI���7'V(�_�aTD%1�J�-�����o��9�����*6"(�Cp�5n�>�۫wf�fM,��W*��y}�)�(�i�3�7K�Ƥ�yn�*��rF���8�僎�S����n��I9QH�7B��7�w��Ձ��K3&���v���:�t�wk m�0�`[u�y�� mʌ�*t6(�`fd��ջ��W).�޺�=�OՏQ[*(�jB���ـ9m���,�l��!Ko>,U���h��'*����wn�Lən�i��:P�� ɒ��������A�$�0 ��f��"B'��R�9
�۳���[������z�b۵K�U^�[��G]�h⠳��d��2۝��U����\�^ T��@��kl�C��Yg,H�Ĝ�|�,���,�d�y�5n�i� �6m?����]sb&�t��ӵ��aǡ��X����s�/mF�ay����OFN.�WŸlNr�(�<�x�� �&�ٶXy3�"������G�}���.4�Ѷڸ��nm�Ѻ���Fnr; J�i��)۶-�e"4�s$����sI2��N���>fG�|��ݥ@{==IIIJ#m��ܐ�32iʪ�ȃ������@fd�Z̙ܽ�sI�r�b"�D�����y�n�՞�����O��٪�ۨ��
rD܊fI�&d�}��@wt�@]��A���qy��vu�k�u�t�rU���w[0-��<�ŀl����n��Ƀ�F��
�3�������[>�@�ێ`��zˑ�'c�:��v\M��~�����`m��v��ND�Y73u7s*���0-�ΈP�t�P�8����D� � �?������X�l�;�ـl���L���ի#N9����X�4�32i`j��`}��nF�PR��5%X�4�;�ـ9�� �o �ےn��"�%D��@]��@v�n��{wiPy4�7��jr��&�*R�7*;+�Cm]]g�N�D[�=m������m�4ORn��E�7Vn��ݺ�76i`fd�����-��MЧ$M�`}���Y��A�������y�Z�{#f8�S��MФ������ɥ��U�M�D �"*|/�~��=��Ձ�F�=�T���7g��Ҁ��k�fe*O����EzTJ
5"T�䅁���`z���{��͞,̚XЬ#z�1�$�����G�ek=]Z̊���0n���[Ŧ�>���#u�W)J�KMT���B5N8������M,̚z����+���M)��0�eP�+�D�<Pѿ�����_��������6�9NI
3'J�ǣ�tE�u*sg���k�)F*�9n���X��� ��f+<��fP�����:��g�y��!�
r8�Vۻu@rfeۛ�wg��Ǡ=�a��J������qxrhN5r�������ϐ��z�P�F�U�]R�	MP������ws��E��/�=����c)M�j��l����ɥ���)#�{�`w��Ձ�ɥ���RGu��91F��"fJ_7b��3)Q��3��Δ��*�f��R���F�r;�9��J/���ޞ(��(93rh���3(�G"LQ�*MIV��,�L��n��x}��̥@B�Cc)L�1&)&�2C �����4�䌏�R`�2h�RHA��"I0`�
d���$	,�H�%z)�H@)?s�ؑ��8j�d!������df��- F<��aD#B�1� @�~��$� ��Sw�lN���7	!!#>	���k�eh��~f��E�l٭*Cz���hc"_���D>�p���P���ӡ�{�}R H��X� �FD��Wi��#��"�"� H��B22B0"H�}�޾`���E�����}���R
��u*����ԅ'�6��T�D� A�̒v��Uhls�B��Xz��0M���Bڭ��I�jB`�HO��耀��h�O��+
RY  �j�ð�'dڴn�BқW��]d�g�g����(�aK���n:��\���;gm�5��l��[u�iݝS*�m�n��d,�b��0{��ci� JT$�ٯ���d6N�.�t�<F�{ڨ6䌝��i^�UiN�[���յ[Cb�V�X�&0�!�Uf7��j�^]��^�0n������٪W�Ί:�N赃�U
�SB��c^˸�e�
���*iXp��:�S�;Z4猗i�yA�Ԥm��,N˻pt9႞5m�w*jK����Z:�+YЦ�رȤ��Le�f��,����t:C^��(�8p��c�<ѷ����&x�{:whzh\)��\��ڤ�)\gi�xU��÷Z�PR��vZ�m��lQmX$Ҡ5OlU@浙�U�z���89Lﾷ&� ;����s�M+<�^���]0nŸ{�@cm�Lr*7v�:㛮�d�CO�<E���H@m����4*9���3F�u��\	��<v�,ҹ0S�@tM��Y�'�L�f�l���̸ʒ35�[uas7�I�VL1�W,�C.@4�]Dukd��;i9�mhv�,�q�E�{[��nζv�Y� P���Lh�����G�r�a�V�R��RM�LpK�Öy�할�\5g	�!ȴ�
��Rl�N^�C;,6{m�J�%���>�tZ�d7
ۍ��
�ҫ]	b�<��S��O]��Nm�P����Ll���n����\�i���i��C�%�}�y>�V��`���m��A���k�%m�á�;��nv]�:ún��i��%�+$�]��6:غ�c2eȠ�6�9��ܬ�b�[m�GS���;��uPA�b��Y\c��;�R�̆�{$���[�BV͏AP�R���h�������
�U��a�M��/@��?b�|�pA?*��
"��߯���ڝ=��S�����-��z]QwNQ���nv��p����{vGZa�RX��mv���bga9��ѣ��Y^J�:�K/;ѻ]���uO':��f�プ�n���s�f�N�����Ñ4�q��m��+َ�廀���n9��Ypq����κ�:;��\��SF8]]j��=T� �o����c�p�ˋ޽��� ?��7f�3F���\ՓXɬљFd����6�ɳۭ����M��M�ؼ���ݾ�F��tԦ�������Vn��ݺ�s����<�U�
Q���D��X�y��� ��@vt�@]��Z�w77ɍ�9N!�Jq��`w��Ձ�٥���<P���K�dn�"	R�˻á�U$����3'JבA�����*q��F�� "������̶/v>ۻJ�˹�f���R�9;<�b��]q.n���2'>3�9�r��.ő�J�:��{�/�}X��jH���5�v(�2��s�&d�s&�{��`j�����J@ܤ6�N;���7��� ���#�)XE`ȄR|D��'��TRmfe~.�:P{:P�̊ԙ;����Gt6�!ԕ`{vx�32ig��Iyg���޺�7vjJJi�m���d��fg��Ҁ׽ؠ>��T��rL�;w�(���P�)�wR�#�P�̊Y��ۻ��̝(��(�w���߅�g8Έ.;���(�E���7���V6�aIu�F~~��w.�}��!����;�z���ɥ���O�Lɗ&d̽���@^�t��,L��:eP�8V�d�����Ҁ2�f��{ݛ�(�l��lu2��	0˗5��n�0��Ó[1
>P�$�f;�t�7vx�;׼[!Lj)H9!a�̓73&I�3;�������p����r��o�Uy�2 ���JI`{k�ɨJx��;���w�ߛ~o��psj��]�g��s��#�b\.�.�ͦ�s��=�w|�g�`y!"8|}����2i`����U|���Ł��������)�r����$��6��[����3�J�|���|j%QG ��`��`}�4���U%�zx�;�<X���wD�����f��373$��~‾����p�䔧N�HI}�W)�nI��m}�@~ǿ�
	P��i�RB��vi`~��2�߸����]��`�ə"4�n��;�ju�y7eW�K;�ތ���E7�O=rh������}�}���Ȕ���g� �����Y�&��۳�����1(��H9!`���U\�'=�:Pݝ(��
��̝�u��`� i�dj6�;�<Xn�,�W9Ļ�<X��Xwa�	�۔�D�IA�ɓ�v��=�:P���jfI��~,�^G�D�&�d�Q�XfM(�M�ɣwz|��ٓ�I&�A	"!B���aqVT�-]���]�V�`�D&��],��à�90�s5<�����m�X!s�_�O��q0��#)#a^����Z��x 4��KY��3�&����/$v4sh)g�tg\�Mc;(vzt������g���WF!cOu�����i�Y�Uƃej��Ŵ��u�a����;Aٯk8��gP�θŎ���8�$�;N����/+��{�s�[�Qaߛ�7Bmӊ'Ds�:n�Ln�ո�8vernvN�V�Mc��7���>�+|��D�1�����ٓK�٧�\��wvx�37ɶ�L��%���������������\�H�z�*SM7JHX�O���|���9�� ��� �2f,���!�M8�a�r������3w���2ia�W9�����3��*$Ģr� ��@�ɠ?s$̯w�<�O�sK��j#[	�.8��I��yU��-�=�u�퉢��a��n�oOK����wwGF�2D9L�Fܟ�����6i`}�4�Us� 3w����<�H6�L�"U���2�(^��	!}
����͚�¹&f�Dл��L��%:RB��z~,36Y�K��Ł����k1h���n�b���șm�x����������Ln��d��)T����2i`}��e��d��33e��b�Oh��R��9�$�C��&�z^�r'F��펝��y�"XNw�������r��A��NHt�߭��s� ]�N���ٓ���R;�Z�CüL�@]���&\� 7w�����������+�����H��NqD'/ 9�� ����$!B"-J#�В^��BKu���`��Ӏl��,�V�4�*4��UWsoŁ��[,��KW*���K3��d��mJd�D�`gsm���m��=��ٓK�{ް�cQ(�N�I�@m�h���՝�ѻ<^��,\��'`�V{�b�6]s:��d��">��ŀwse��d��*����E��z/'j�t���N+ �^Mk&N�'J/6��>��z�e�ɢ���J�TBw��"f������a�BJg]?� ;����t��J���8�a�r�����X׾V켚
R�$��e��*��i@f�qȒa�(��nDXc�V�͖ٓK�ʹX��[�Y�)H����3B��KŰ�g3�v��v�Y��23�Ch�Ev��+��uc��B69��8����`{�ـ{��(��zC]?� �_2���Bq��rXw&���r��#���P��z ��MrnL�d�a˪B�"TK�D���9@}�z9rd��l�{��3}?s&��$��9QT�Ɂ�(��o��o��=�l�=ٶ���Z�q�M�Jcp��m�(�[�><��I�{zـ%�\���P%��|�e��� ��b,����/X7��;�N��8-�������y�w���G[�}����=���0���Ľ��J�$Һg4n�����I7I��a�1����9���q��l*�kd۶��c=�,�'I�`ggӹƆ���(r��8�H�J��
=��[r:�ک}��x;^Ip���aٖ��m�v˵ؗ;0DE8�mE ��$%�s�U��W�9�E+��v���)K*�a���Wmn���ۖ�ke\��t����b���k���7�t�>��r���8k&o��٠;��܅
T
lMԎٛh�r���y���p3w���l�@}x�O ���Q4܈�;�5Xfl��W*���x�;����ν��j��7M��5�I�36hfΔ�yNPrL�r\�=���5W�5�J&8�c�rX�l�>�Q����KV ws�]������Uь{�h��]q�/7nWl���1�yN�"��Di��kd,��֦��;\�X�s� ��B���~�,n�TQ"@�Ӑ������~�0B~���.�d�qH5���($ �U !��-q��Q��Q^�M󟵸�<P�|�Z�$�������ba�D����� ]�����G&d��ɒL�E�u9@c��P^>�T���9eM]��l�=���s��!D.%��K���J�Q��������&�J#�������=�ـt�[߃ߎ���i�[+�b�ѹ%���Y���n݇���b�l���wz^7l'�� ��s�-�6(�^M���̹����߭����@�H���7�{y��v���I�l�:��J!~DE6j��h��@�H�1�ܖ{��X������H09a0H�#D�0H�#�LXB0_���N<�BqC�c$�KȤH����)@$7)A�h\)���+�8\ P�o��S�m0�	X*C����������V�+	!c�R�!'���@��©,`�{f�7F͐�!�HɆ4eF��O��8��������B~�SC����@��A�26�)���M�1�(��(!��"��@���,M����l�P ʹ�j�a��\$�A�dQ@�tO؜�YS�~*ߐ >S�~0�U3�G����M�G`��𿾞�>������!��Vܡ�2S*'r�w=�`�� =�� �v��yj�.��(�`����R�o��wޞ,��h�7v2�jr��&�j�����s�lg�l���y�N�:ūv���s1���w}}�>q�m�"�	��s},�f��̧9�K����/y����PK�<�����s�`��L ��x��w�H���	�#u#�������"�fd˒�/7������֝�K���(���a�w��;��`}�l���El��0�j\�YWeR%&��v�se��l�������3]�����im�&T���q$�6�A9j]sX��x�r�ڛ��=oj�����r/zwŏ���ڦ8���g�OŁ�wmVf� �����++nP���J������`=ΰ���s�g�d}�]E$��7Mȋ}��`}�4�>�����$cl!E$��]���;��,��h�:�5�f�.D�2&
PA�%��l����7��x��z �ד@	�p�KR��^w��W�������H=*�նY��qy����%�7���X�[v��M��z�6#C�m�1�B��I.�.��ہ̷U�a��'[���b���1�ەۙ.v7��.[U�&לnw��{rSѻg�S����6��N�p��kD`��[X�V_M�Gz.Gll�'v�rk*<6��]�8��<q��D`�m�T��
�H&�u��������=��r_mNn)�]�u�]�/P�Ņ�.R�l��|s�+*���I��O�Ͼ��Ĝ�K�#����{�h�;�5X�͖ٳK��"�4��(���`wj���,�f��ݴ_�I���R���'�r"b�=y�@}y8Q��2�ey�NX����:j1k%!:�*c��,�f�K�����I,O5;Iz��m�o��$�:��b��NI�ZI/���>�$�\���7���Ifo��$�^�j�H?�������X%+��j�;��,�T6�����z���= y3��z:jڳ�h�����$c�R�I.�6_�%�{t�\�r��л����%�~�$cn���R殷m����u�m⁸�e (� sH �#�U~���k��v�}�{�}�Iu<��$�٫~�Hʉ�P@�O�I.��E�����#U\�SlǾR�I,����:*@����)"-%��*���L�v��HǾR�I/���%�ʮS�^��I%��E]4߸�`�܈��:�T��K��>�$��n����3~E��[XAm�ڑ8�T'DjA-re1v-n����ɜv�u�pv���f�:��ދ�V�T�tJCI���$�f�}�Iw&�-$�����s�i,O|����^F�2$��q1�ܟ|�]ɶ�I%�s~G�$�S�N�I.�6}��\��ݔ��eD�L��E���o�G�$�S�N�9S���6<O s|�o��9m�����Ife�ԃ$
�
�m���$u�i$�{�>�$��m��+���ϾI,��9#tEB�ZI%��ϾI/r���~�$���|ϾI#�5KI������'E��k�Z��׳7�S��M�q�3W\<J�W1��rr}�Iw&�-$�s7�}�Iy�~��L��.����������Ѕ2
`x��DZI.�o���UW8�B��Iw=���%ܛh��_wlMo�鶤���$�sd��K{�>�{��r�y�֋I%��||�K��R�⍎q6���K�	��}�g9m�w^ݛ����w�s��¼��͎�I.��ZȒtGA�N?�I.��E���9\�}��RIc�Gi$��5��ImhCn�J�G��#����{[Pg"�3��pV��]�P[n���{����.����Aӎ#�^�����$��c��K{�?Wz�Y�֋I%�ۯT������eˬ��[m��wY�(�"&�.�ٽ?|��=NS���^G��&M�2J����q���{DF�i� ??�����$��m�K�����I%כ���uo�5���-0�t[�����QMw���f�I{~�>�$�^lv��W9�7�����?_!i7JH�I%�ݯ��K�+�y7���K�7��K�6�i$���Uv�2� �G�D�_�_�gm�Ղ��b:B����YU�P]\�^��$^Ò�Wv�Q�݄�S���s(an�Wl=�E�.��׋lo-�E�ͼ[<�>ո��
�]PCS
�'^o<lf��u5������}�ß}����p 9�����pZ2��u�n:ֻ<$A�[�Ӵ���;��m�{;��i83�(GgN�7jQ�6�z�Xᵤ87=����]s�C!5&fI�)�]�>w���r�kh��g-G��c9�]Yy�'`v;x�����p���n����������n7���sʕR��I-~���ܙ��K�6�i$����$�Ǩz�A��cn7i$�&j��W9�U6�l���I{=��K��~�9�r�ic�A�q"0���_|�Y�֋I%���>�$��kv�Krf��I,�IlENS ��i/s��q�}�~���߳;���m�}�s������"�}���Io���H2T��Q9��I.��ݤ�י��K�6�i$������;~��m��#�<DNܶ'<��7Yԝ��Y�ᕶD��N켜\��G���w���|�F6�(����K�w��K�6�n����93s$���wȍ���;���kRꖘ]2k5����wfn��t �^(��[����s�[�3��n�-�͟}��r�k==|`HEDM�rS��^�{����y��_�ʪ���o��$�-�Ӵ�_em"��QR���ܐ>�%��P�w�fn�m�����[o�����|
7��t>�$�~E?%R����ݥm�}�s�������g-���{�s������$��2�B��N*����uU*��YY�����-&v]''V\�6-}���F%�
S�
�:��ޤ�?z�i$����$�'����י��K2RF�G)
%���[�߃�Uʦ�����I/=�?�B][�N�\�6��J��J���&�$�BZ��;I%����˶Uq��F$(�O℀�$ (R�BAY`���	?  �~�o�ɻm������&�4(�F�$�v��U�o�=���%�޺v�K���>�$����$�{��r
$*t�|�][�N�I{�UY���w�%��_>I#�k��v��p\�5�7f�td�/i6���k�wc��������t=�=���ݏ��&�Ѻp�T�Ԓ[��_W�$�'������u;֒��];I%ܭ�-�Ȁ�m�R��$�E��jL��f��{���ww�����������U6ь�3q���r�Iw�|��$��n������{���I-�Ii$�p�5Q��B#��^�
9�{�3v�{�}�9�m�ﻭn۷�D�q��7�ȝ
��������պ�#m�@G)
%��$gsl,I���3&es���-�(��"���;~H,�Nɡ�r�pN��s�Z7f3�`y��������'L7fqS�n�в]�`��X�[�������f���xОDi(�F$����w2+Y$����ؠ.�U* ��&��&f���yU�r	�*t�vV�^*Ts&w=��@y�v(�2��Cʗ*17RH��6�����`}׺�=����;��Db~e%)��$q��|� ��u�v���5%�0�����N9�"��fb�R�`+�#8�C(�J���i%�ȟ �9a��Gb@�	 �H�#!
\$�����$H�!C@�18���̂*���w��5B5������44��~�3�Q�����Q���ֵ��e���m�ܐ��.����T���eb�qn�ᅛ����E���)���%�Ʋ�g�̫�[uJ��U��uŵm���-��j��
RZ�X�bU��b��v�@t�t�ţ���g����4 l�Ʃ6��-v���m����Nsh$9#n���oc��,��-�h;y�5T� 9�cq��� �CS���N�v|3��y���ڐBS��hT{�/*�ʯj����6��6$��%����<�����"]�c��b6��H�A2��6�v\ihݫ��UU��(6�,=P���:�C(�'V�p�')�̆�z�h����=�V�I�ۃn(�W7X��-;�E��͹jP�am=`��3�s����q�X��u�eN��gVNY�r��kKis����!�eyB� ݎWoNl��g8Ƽ����am]�w<������m���sهcf��.6�'��mvL��g����d�M��m�b0�ɛ�K.ʭfplb��Gp;����e���]��:�U��N����F8�:�:�l�s�i�Z5�n0��$ջ79m�-�����Sa�M4i�^�T���.�խX��Ғ��9�
=�f{jW!�\�8^ӤC��@kmI<��D$3��GN��GS���\hl��d4�[D��ஐt[�C���s�6�0������=�� �m�v���e�-@!4��mڐV#H:��ONU�ATUOY+#UN5��s��GG��:��a\VW��kpyk��*�r��NܛX�l�j��\�8���v�1ۋv+�ʡ��࣭�j��8:�Gd�'c�ˡ�،����z뮹���ضz;D�y�Z���p5�i[#�ՇZ�λ=Iۃc�]n�\�u���M�TPqD�7l�3�5K��C�͢ɉ���Z���n�T��!�����@�6�W�װ%���[�X�Ԍs��UU�n�éW#y
��)U����\�Z�!�`�TQ���B���h�z"g�P���p�|b�N���ܟ�����̫�Y�[4��=����Dv�-nrnN��� �ү\Yye���NѻP�yMvre�l�v5�:�V�����,��K�x⬶��2����E3�WZh�m�;�#���4�-�m#�T�1�6���s���ƞ�M�O0�z�EPݰ�n������]��r��؍k�\�̘�g�q��۶6Z�#'S:��]��9L%���߯w{�}ӿΥ�_Rz��-�l��g�n֎�ݎR�͖8,V%S<�����?Yc&����@��y�-�vf�W��uno��%B'���׀w;���8�7Y�%
d�2?�Dr��QH��C���j�:�u�,�v��-��E#nHI�=��p�n�Os�y�� l���УQI8���v�����������y���Zj� ���V\���02�(��8뭄��ٰv��˞=p������lq!S�9N?���������E��&I/�-�v(n�3Ãʈ���I#�;�W+����W*�X�Vf�幮��w9�C���&7"�7�XY�������`j�h؈7�)5I����v�3]���j����|�p5y�I��P�#q�,�v�}g��w^�XY���J��W*6!�J��@ܤ��&�k�/1����ۥ�6�@=���@�WYb����r�����͆��y������� ���=��~pJR"j����˜+RI;��������1���C֔i(��A�X��v��{�`FX�E�uk������}�`}ܢ&��
�6ND����K���`^l��d^='��ؠ7wi9 <�*�MԒ;���`~���|-����s]�����H��N�P#����Afz��q�\��Hk��p���"x񭊔�R�܌���y�����`j���f�V��G�#N1�Rj8�:�u߸����3}+u� Άkj	:*�n;V����g���1��(���%90K9/13����F���@y�2(��F	�1!�8���!E! ���BF1!����e&�O0v)�LM$	Pr�Cﱒd.MY~ފ�2��Y����1e� �s�g����X�����e*�r��@�p22�)��@m�9�w�;�Əb�z{pa7	���_�~�m�� #kfQq�^����5�͆�V�{�D���SqN;5��T�D�'=���@y�2(̜�A*�m�8���U�����%�}�`g��Xw��A#i@ۑ�X~�-y�;��`w^j�36�Y�q��H�vVn��Y�_��>��[�R^�B�g������Pڶ,���M�\	r�V�`nH��>���ٱ�&zl��.g��F��{b!!��퇝s������88K���×�����z�+)��vt�]s`6b#nx=v`5 c8ݹ���y��6F�.�@����X������tF�-�D��vWCXH�!��i:s�l��x����y��g#f���o^����<�I	)F�E;U\����-��d$��2���[��stX�i���m�SB:x�=/7�������b��N��B�����1�fG.�>�E}	�ށ��� ����l5_�H՞�1o����Wꤏk���Q�
7"���V���IL�X��8����M�M�˹����;�V.�{�{pT����'������s�t�u�l�u����P���'��x���mɛ'r�d1��Ort��bu�p�d����X:r�����zV.��7_�|��w���sx�O���SUuE� �[����KRp����
%BK0�v� s����s�DW8��>zTI�:Pj�R;��`9�u�w;�u���s�$�J��B'��3]��صX�����v��#5�JQ58����݋g s����� �� 6�Juj���y���6��-e9nd;�b����c�p�s��hLЪ�l��E����� �m� ���ܹ�<�m%J���r;�w]��UUT���y��E�`j��`gr�OcN
�7W35u�9m��ܹ�P�" ��#$!$$c��K$��1p�u� 5��=y�;���7rQ�����n�q��˜�n���`}
"~������"	x)(���QX�u�[��[��݋U����pN�t��xa��v.ōh��y@O��kWkn�,�,�G]"�$�(5RI�ջ��պ� ��\�[u�	�Ψ�������[��ԑ��^V���`un�$g�%��a)4��E#�7ދ��r۬e�X��`�Z�VM�&�@��E��w]�ջ��ջ��W�2$#�AH
���۹'zVm�Q�J��Q��ջ��������E�`j��`f���Ri)�[f�gC��ֹ&ۊZ��=iϱW=��.&k(4�G'j�g��������صX�u�[��ܕ�0#" �n�q���V��w]��w]��I�m"������5���y�[��[��݋U��1�I4�
�*I#��8���v���`f�|zI3=�� m���a��I5WXO7X7r� �M��۬�� � H��˗33��ђtzrBM���P	��r�����pi��&\���y��ђ�8%���(��m����8�n^��|�����-�����R{;�6�nѶ۶��l�sP �����A�<OPBU�4쫌1��m�ŉ6����O��7kl��W�����ºlP�b=7c����p.:�^5x�rPp�2 �^d�-��jު'E8�!�7��Mj��4\:�e:����ȶD�ٸ��'��tk������uDq�QJdB'r<3"�`w^�:�u��u��k5�6R�*QH��;�uX[��Y��͆�t���QD�8��X��`<�`��8�np޲iݧQSTH�D���ś����j�;�uX[��̔j`J� �n�q���8�np��`<�`ڞO6�ЭXx�oZ	��y^k��x�a������r��=/��=���#e���y����n�1f�36jV�Ɔ]�T͢U����=-��B��G + #�(t��D�ן|��MJ���`��:m�T�B��Y��݋U��{�����`b�Z����'S��9���j�;�uX[��Y��Ƶ���)F�
(�QX׺���UV?{��5o��݋U����W��pB���q����|�In�8+r�ۣ��vok�nL��d.Y�LIF�Q*�!9$_���1f�3v-^�|�<��`nl��T���I�`b��`f�Z���VV�3%����$vnŪ����qs]v02I$��%���%��@���9�b��WK,�j�BPA^(�
bWxf��h9� cF��X"Brᅗv����&J ��!��F��]��M��d�z�,А�#p@�](@�0,i�k@���[�0��Z���h�Ri-R�BE3V,SI��ң _�P��w3A���D̂� Z+� ��58��2 �`�T�/�G�4
�"1) `Hbh�hnګ�Q�����)>?O����䨇�r��f䝿��`}���5IF	����9UUK==�`b���Y��݋U��1�U Ɣ��j�$VV�n�7b�`w^�>ܤ�Q=���#�S7>g(;	ӟWn{G�`��˭;�r�Jܲ6�ի�6�N��*��`b��`f�Z���VV�jմ�mRl�M(�vsa��U�H�?yX��v,�v�Z�pN��J��D���V�7]��7]��٩X�<�DIE���E`|�u��u�͆���L�0�-iHQS�-�~�+s �ȝj�EQ��1cu�o;���6y��ԋ�M>�����;+�e�g�ۗYC�=�q��ں<?��S�\�*�S��b%8�Ө���>�]78�n��n�r�L�
t�܌����`un�1f�36��9UI[�yT�R���RH�^����7]����`w^j��N�D�IS��D�1wu��Vu�,~������z���M������٩X�M���{�����rO�?$��$ a��8
DT���C (	��V�2 F��e$ԝ�CW-�&��L�ڔTjhˮ$�Nq�(nέ��bN��'��)B�a0˂8e䈙N&،�m�f�.� !�L�I�sp��Y�dc�#t�h� ���'���n1xy�ܩ2u
n�u9�<wk�h;\4����@$]u�G*J���W/=�Z��6�nv멎����Ns/���ӹ\n�U�	J*ƺܻ������wu����$�F�����i��.ű�͛��(��K�٭���(���1F�(�r%��uX-�v.�|�w�<X��dID�!9VVn�w_���{�`g��Xw*'�'D*�*�'������Qx�jL�N����>��~�Q�%8�Ө�vm<�`w^�1nk�1f�>�e	T
�5Bq�qX��:u��:y��5��8S�G��cZ����׊V����1�:��6<)��6���R��^"���%8�>�ّ@[�dP�������z �7���$9�5#�1f�UT*t�c�I�u���n�f��`b��1V��5T�'J+��5��8�np�n��n��F��LQ�
B���ܮU,�����=�`b��`wi�tx��%"�NI�����ś�����Vu��:�U9"u)R#)��N�*���b׳F�8ɹ{Q�#(�=6}:N��N�FT���Y���<�`w^�1wu��T���*@�m���`wUs�]78N�XO7X�r&U�qSrR��SW8�np�n�Ē���x��3��U��1�NB)IJm)$V.�n��O5X׺�pŴ6�$�
�R;n�ԙ5�����z�/"��on;�/��+�p�^��c�ѯ/1���ˀ�L��<=��9��ں˞�rJp��B)�m�=O|���V-�v,�v�pNP�IDQT�Vu��n�6�j�7G�[QPB(��`/�`<�`�s�]78>uV�q8��Ӝdq��uX��U����n���G�
��,�B7Æ"��l��(���H�D��B��$��(X�Ea2H"��b!��/{�`mn�)yS%HI:Q�`f�s�]78K�XO7XВJ!����5�{kǵ�=ir��5�q��v9�g�@����M�����֎��<�~��?yX�5��u��SKVc�:�R���RH���v,�vf�����s��Ғ`�$��ڰ:y��7yZ�=��8���Ҝ�cQ�Cd�iE#�36��u��w]��7]����jJ1(��7N�]78�n��n�歘(��BI�A	޺��*.D\�3��rKM�:Y[<�P�$cV��M���T��d(G&���zi��Z��wm1.���^{c�s��!Zۉ�6���@U;lQ�0ո��nT�kH�m�CrN�7[��7n8�h�R˦��U����z¹�vôը9�y񳧎���j��#�;��p\`]7۲<���
��U��[f[8J��n�;�d2���M�9��:�=��3��@m�9,��6^�>źlpp���׺���#��Q	�"��5��u��SK��U���ui� �:��G��7]��ճ �M��۬��jF]̧(���vf�����`un�1w5�v��P�P�I�rJp��*��[�p��������[0N�jE)JRR�JG�ջ��;��`fmM,����V�V�ߒd$#)<���E͕�Lv�4�v;vG�q��=[�K�M���BJ(����g�,m[0�np�� �Ny�SsR��������9�lʕ	
bWB���MX����7��`��;����P��t�`w�uXn��q#3ޖ��<Xa�F�*�r8�7v����ڶ`��p|��Ysde
UE$���,ݩ��޼�`����UU/o��T����]�0N��rE�\=1�<&����x|p��s��H�s����L�눒5NTBL�9:�~���;ך�7vX�ݖ�[�(m dC�ܔ�`w�5_� �{��;���3v�����P�ӕ)Ԥґ�`���>�칀'�j���A��1�'Ș�ER�bx���k�nI�g�������)@�qG���W9�q,�zX���`w�uXn�1V�Zۍ�M���)�f�l�=_�o���~��X]�vܭZ�F�:(hDl�sΰu�'�]w��!��3���
�;D�(�P���RX��V��,��s��}���;���JJ�DC��3�y�5ɒL�ܷ�ؠ�[4z�U������RW�Hl�ʨ����� ^bɣ����7^���ؠ/�T�6F��%$�#��;�[,��$�~�sr`.����#B������� %,G��y��{ٹ'�x���%:N��%�޽�`uf�:��������֐[�u�N�K��J]��h���r�NpOV�x�x�u��jT�:R�:��R8���vWw]�w6�{����+V#xy�P��uu�l�u��;�7i��6y��1V�Zۍ�M���)�w6�X��V~�K���3=�`ndأp%"�]��v��g��g[� �ke��=b[)�er8���v�78�Ӽv���J�Q(���3���!��G1�
�������t�i)�
��tP?�����&j(<?K�T�"y��d�A�vf}
���e�7B�J�� lHA��(�h�"Da"ǽN������9H6_���K���P�H|�)d#!
�,c �����ִ\LTnh�0���[L H�Uc���r�Y���0M�,�p�jr�?K7�%>����y��ځ����Т&�K�:�Vf��m-3C�\��v���H�ư��K(o��[%����a�I��Nh�8#�����G�	�s.U6�@p"�R@:~᠌���7Y�[�GIC��wZֵ�W,�5�kX�E�R-;�\����¶m9(e����\\)X��N��պy'��RZ�Z�8Be[�Yږ��*U���iVUU�� �x�-]�
RZ�H㱅V�T��H&�I�s�#�̭�賎��r[��"�V��9T�[��U�wX���Pl]�A��;�݋��i��m�{��ϖ��v��mӶe�% 5<;vh��8�A��C`$�H6��()8���䗈�[J���2�宦Ӳ�+T�����j����୫���y��(���Aݚ�@k]R� h��kծ�Gn�m�.������:��r�crORj<��c��n��ct�,�I�t���*˪��qݧ;Y�95�혭�c4��s��I�����7E�=<�J���v�;�C��7��N�t׮�J蓢qI�lI���nŌ�{oO
90�tYH����7�iz�]�����K-��YN�j�b�T�[&<m��[t�a�"�R�J+̵PUI�4�F��
�z0P�\k�<��Ѱ'�$�gj���ٚ�c�U�n�q�Y:-	Ï��VKms�яU��+�v��ϫj��7n�˵�Y�H�N��E�8��t(b��
�U�m�a����R"��ڐ����H�SJO8��+r�5�d.��[���h�G����(�t�6H��xA�Mg��� ��Re�sN�}�F�6�f���Q��\�q�m�k����eU�
���Q)[��R���J�d�������UM�܎�i�<�	��h��-юj�ۅs���eyyA�c�vu�n:�%��\p�3۲r�f�K�;jmu�٪9�Kc�����g!�ɛN$�Gti�ۦ��ʽW�`�EW9絡�Ƽ�f{9j��Q��ä���]�ϳ��E��нv����nH���571\�we�a�c�Pm'�24-��i嗜�c)��XW�����g�U�n�@͠�vxݠ]�"�@H�*�AtS�T�pʪu�f�8��E٠:�"f�����Eш.� ��.56҂��_������EX
��������QөgV��]*���G����Q�,��sTxy�e�d\m��Gf]l/�E%�h�ɩ����]��{���󚍢���I��m�B F��Í�EW`�c�;�=���β�g�h�eڎ%x-ORN��K���қ�u�y�:�s�r���㆝�]K�b������S<�ö)t@���E���8��u�t��Fc�����������o���vygs��I6.�NbۍH�<�T�5�>��k�m�����LC]ټ�`y�s��;�7k���B�K���74�KʤJ��RLN8�����ݦ� ��� ݦ� ��RIe5@��IӒ��;׺���v{�f?yXo����wM���>F�$qXz�������K �ml�;ך�]Fp�$���8����Գ}^��������`z�����$T�EJ�9v�o=�3��k�nՍ�؝,�r�s6-��S�5q�I�q��|����;׺���~���K۱�����)��Uڻ�7i��P�$�$��`��� ;we�w6�X��-��:(�pr,g�� �n�y�x�78�R��H�6P�$I�`������{�����`fg%#b��*!&G����`{���_�}�`��>���ߙ�ƅ��V%7	�^W��(�d�2'[��O�}/��ru����q�j��93�:��3����v�wg�s�o�������*	�D�+�7]�{[� �i��\� ��:D��̓Sjɺ��kw��;�a,(Dx�
��D9����ܓ�����SV�m��&�Ld��ܮW��zX�|���v�we�����DT��*�ݫ�v����� {[� ���`}��5��$��N�D�؊�;s��ҁ���n�/b�g��6�Z��Y�
�v�N�E`uf���,�����^j�7�Im�B���NH���>�l֤�;�歚��@y�2(��S��9Q	1�#������`uf�>]�vݬ��5�*1�ӎ��=��py��=;ΰ5Bq��yʑ���n��H!(ڢG��M���u��;�=��po2O��p^���4��vS��;z���O���<�]��-�7���'������==ΰy�x����M�Ҝ�Zq�M��ʍ�`ͭ���U��{���fk�7�n8����%I`}�5XǺ��9Iw6x��W�����M0(������=�`}�8P�M�33'fl�x�#b^J��9 �VfM,R��z|�{���=�`}��#[��q�@jP�����b	U�A��dK��:�2�4k�A��Q�.nd����QC=�6̫�8Xi^{/]��7�[�C�0�U�sܽ[s��A#t̸z:�Ң�FU��n�oVEŷ>��\࿭�\���]��Q�9�����;]�.�N{%�Kx�&�E�6#X�m87�=�y<���/�'��6�ȸrM�t�DݸݰV`��9�hv]���������~�v�ӣWu�qQ��<��bݮ޺�㓷MƎI��;}]����z�%F$�9�w}^������U��d��������)M�u%�}�� ަ� �u� 7�w��29�}jȓQ!)M�����~�>̚Xske�}�������e	A�D�6�=�l���������)�Zیbn!���v���`fl�7���=;ΰ����hL_Qs6T�s\���\�0n#[/���2uM��<8:+��n���H�nD0�JT�'����:�u�.�|���zX��i2��Y3Zַ$�~�sy�$F A�����5}�ܒs�����,�Tml!Q���'���u��;�w;�6y��;xWE9VFJ�I�I�w6�Xٛ,��VٓK��pJ�|R�8�K ��� ��0w[0�N�S�D�jDV��Vں6a��l��g�ǉ�g�m��N�.�1�d)�ց5�9&��>v���� |Ӽ �s��x�	JhH�अ��d��76�Xٛ,͚X�V�m�4�%A��� >i� v�1ZJ#RH!BDD,H"8J���D���F$�-۷l�7�ـo;�N�l��T�6)*K�U,ɾV��Ł����76�XєnƓ@�D�E`nSs�z_:��;�;k���객Y��pZ���
���������=�8%��Fɵ�?��ݾ��5���{�������;�7k������%8�22Tbn��; ���}�UUr�1o����`|��y]�QVq2�M�u%���`n=�`|���ske���6T�h�B�ȣ�������������Y4��$�\NS���e$�
�%8'"�>]�v��� ݮs�>�� �Iss+�R����	qnk[���ѯ/1j�&xŨ�N�<��s��V'���R�Z��cI�r5Q8��߫��=�z.3��|�]��y���$��JTi�%I`w�4�7��vX����I���zD� �"$�ξ�p�n��N��l���OaF�)ȣqX[��ske��٥���U�������2Tcn�� |Ӽ��0�������\w~q�6\��S\��S.����Au�l��Y��v뇰���X�ظ�*8�8.M�;��n2�kv(�+D���T枨���/���r����\�\?�~1�f��n�s<�Ҙ��gM�&^���7�x����f(��F��k���9��v��78�ɲ/'$㴓0��e��<��O\uòOZ4'S�� ֓�rx��8R8�t1:m&ܛ���M^�{�����z�MpN���n��k�Âׇ�4�
�9�<��ձ�ۧ��7m�����ɞg�|��\f=���̒��?r�?-�:�I��M������U������u�=v��J!(�>�k�U��I%8'"�=�|����g�S���X���X�V�m�4�R�ģ���w�=v��78��8�1{R*�JTRT��f�����7 ��x`�2�UR���ʬE�q`�@a����[o퓅�[����8D��׺�����$:(��HX�uX�4�ͭ���{�����F�R������[3��I P���z!%)T$���N�u78�np��Իa*1�Q��`�[,��V��,Y��Ҍ95�)A��8�KK����������Ƞ�Y4>h��Q6
1�G���K �ݖ�����{���Y�)ߒcdr�"5Hj�[�.�I� ����9�Nǒ�Lx���R�(�R����)N
Ht��~� ��x�np�ـ9N\���TTҕ
��%�nml�7�76i`���I�¦��ES�J�jJ���?}8�aj�(X�Bh��*ID���#�L�FV9��n�����	����)�S�2�ҹi
�M��JB��� GT��l�A�	&�>6|֒SFk���F�dP��UF9�d�E!��c��!� ���m:m>Q��S�����DqE�?/	�:�?~P?pߦ� ���`fAVȑ(�r"Gw8�`{�`�N����r7�
%Q�T�$����U�w6�`i��7�� s6�W��F,ƞ[ٌF�LQ��"��S�}��w�҅������(Qȓ%F4��p�7��`o[s�o;g舄�!������$����RX׺��H���`{^�Xske���'�(���0��`w� ���Ӽ�78N�I�B�D8����q{f�Xo������f��M�@h�B$`��W+�{�,*ի͹M�5*�0y�x�l�=�l�sŀv�1ߏ�'M�	Y�&��ڃ`}qהc8����������P��G^�%u� ��0o[0��`����x$l���@�C�B���4�W)#ۻJ�=x�h�N������Q2<���*S�'��{�`ͭ�z��Ľ��,��+39)j�&J�m�D���N��l�7���5�9�7�t�M� �4:qԖwf��6{��;�N o4� �蘅11�z���ɮ�8��i��B�&[��ⶁkOQ���N2�ó��@{uk�N;ID��a9��{M �7=�!�;��g:�\ ��:��.�)AX@���߾����-�m��{*=�޷"g��起`t�9t�```�Q�r^@ ���g�74��*�J���E��ܝ�#�#N�.Q����^� �؍]��ڧt^id��J�fcQ�(m�����w��c�$��>Q�+�R]���ZŇt��N�P�ە�&^�F�GX�4`��V��y����Ƞ�k'W�{:P���)C�%�)!`���>�V�z�U��ri`j�Z��)�l�
��%�}ܭ���=Ļ�<X�},�ć�%N%*	�*K�*�K�=�`w6x���`w+e��3u7��P9�Xw&��[���sk���^��Cc�i��Q�H�'IZG�E�[zl8�v�SDi�6Z�n����3(D�6�N',;�,��l�>ך�s����f�yX��[*D�*1�R���nI?}Ӻ�Q4C� 𠘨U7d��,����f���F$T�$
C�I`f�����g�q-^�; ��zX�֔�m	Jb�B��ęrL�:������.�d���zWsJU(qШD��+s&��Ӽ�78�l�<���]�r�6Un�8j�nr��4	�	��m�1�^h*��<�6���ԩ��Wը��)�l�$�> ��}x�x�kx��`=�%;.*��r��r��7�u_�s�ʪH�{�T�N��ZɭI�rQ���L��eȘ�z��\�G+d�)!`�BH��t����`o�j�7snI!"U�Jqʫ0>Q;��� o�����8�l�3�ͶT�BTbn��E`�[,�ɾ_���`w6X]�*J�"'"�m�&���m���|�x���gk9�w�;W��n�:��DQ��RD�PH�O��=�5�f {y� w4� <��9SsT�K���zٓ�~2fK� /7��7yt��^=s2I���4u(��:�����,3ke�K1���`j�X��)�l�D��������Y'{����~�uٹ6,`���G�TEB��IB���w��9�)�w*�T�PR9RX��Vu����`�[,��-���@��P��Q0u�Mi	8�y��y���7g�r�-9�/YF4�(������V�s]�fml�>ǚ����(�F�R�q8��c� �i��� ��� ��r��Y*1&F9�w�[,�f�~�+�Ļ��,7},�F�Dؐ
C�]��l�=�ـ���J�s_^ w�z��FڈUDR�ݺ�<�]M�^ �k��=�ـ5�BV�p_A���K�5�4[�����d��˔Z�j��C��Ƅ�q�8z�k	����Ʊ�d�Bcoh�X�\<gP�:N����n�xri��].�gI��K�u�q�p��[ݵV��ۉ�9�Mn�ӻn�۲�k�v:�8d[�ѻ�Z�.�a��� R�U�S]���]�����V��.�$q=��<e��0u�Ԙ�()li���d�8�������{��`'�5��xRc"V��L󲜶�m�{u����=�\<���Bۭeݨ*T�9I�X�g�`�V�;�O�ʯ�g�<XU����m	�S F�ͭ��W7=<X�O��V-ԍ�H�Siʂ�ʒ���������X�Ӽ�]-\ܖ���HXݚX[��3ke��ݺ�7slnH���*���`w^j��N���`ݳ ��4�ei�����s�=�Zvx=bt�8�ۧ���r����z���c�:���J?[m����K:�U��{����o���F�D�$,�5%+�Wxo[1���Q
.��l�1nk�ͭ����W�/R+�&�>N(9�����nk��+e��ͺ�5fi��1�NB��nk�z�M~��A��O��Ҁ�Z���hi�H���;ܭ�w6����4�>[��r����W�D��\�!;(%�	��ke���^5h�����:�4�j�q8��iʂ�ʓ�77�V�v���֯H�Հ�U�U�Z�!)"��������{������_�q#��Xܒ:Q�UI�*���y�I?~�� �"�&ȠR��ġ*W��x���`��w1WE��j��n� 7y;�7[ŀ{[Ł���&���z�����!<)�S4�yJ���37�w����z ��d���8��dD�9�jT��%8���l�c]k\�:��X�FC��0���Eq�!m���ɫX��X��� ��� ���Ջ4�6
�M�X��W����35l�{��fN�ə��Z��ۈi��"n; ��zX�۫��K�s]��uR����1H�L�rI��~T�n��Ǡ�d�2�u|#�f�{[�{�;�d�I�Kn�]UZ�=�ـk�s������`o�~g�6�ư�qL<�9�vy�x�^ݑ���9�;�[�  �M�5�Qn$��ݬι� n�w�v������3~��?{ߓ�#�)��Ԋ�=�Y5��^�*׻J��E��y�w%�&&һ�w�v�� ���ȉ��fmzXږ��n�:�J	��5�f��� w4� �o �⢵�S`�Gru� ���`v�� �M� BX�!-H��)R�����,�_����b��#���q�jq1yG2"8)��	���l"$�,bRlXb�� �U����
�����z����&�(�u�@0���JU��D��H��	w�tdJZR(d���bCn`cf"9rAAJ)�P�x�9��9�Ca"f�F��HP������ڰՕ	D(8� ��#�1V��#@�C@�.}� C�m�T1Ьb%�"e�Gh/ �/?s�kZ�%1 j�Z�ʣ��h��!�jA�S����x8�ktrpl��1��k��ķMR�X�s*8�ʦ.���Z��r��K�($
��%�Sv1Y��!�,P$2�T���n�2c�
�V7�Ԟ�s7g.z);u��
3Yô�h�Y2��]x4�V^ꖋ\�ʅ�Մi�<���G3zK��D����/$�5HO-"��m�`�k��n>��d6���+�P(@b�m�W��5� �R��m1����UZ������W�m��bK՜J\��UK{�m�˵V,C�t,�����4�WV� �J'��d���+�z趵1���.t�4�[I����n��[;E�Ю�;v��{-P��S�����uU�p8�v6�ہ�ܧi\��O-�	Z�N�!N�w`��L��8��.:�*�pO`�aHУ
Vm�Px�2���:�j��|�l[Pk������-�����3�%�'F�{okK�4v��i`�G_?}U��N@^,���"̰�v��S�.��vr��5���4�^�9�դ�X[��Ms��e��,��^��e���v�p�;:J�;J���@�͵��Mb�!]�^��B�r�*� +�l�4���T�N����� �҃#�ݕ&F�Y:�uפ8K��Ic9x]����3�I�n����AW\����)۝�qS�wQ�[qlp,�V�nq�N���<s�f�P%Z�[��zN��ݪ�B]m 7R�sp"�J��l�E��y�>�<���]C=� �n�'Lչ���y>����X8T�,�vkm������*���՛w`�u�Z�:T����\=�[D�g�\yb����6�*�nl��E.�i3�u��25U�"����%���c[�la�=[κ�ף \�ݲMd4�.Y孥y�4�Q�XJ8)V�E
F!'9e�SڅIbZ�c`��YM�.4��4�Y�A���FjZ��[mPK0T=��ffjM\�Z��Z�b"��"��^*$�<� ���G���C��C8(p~_� �?��K�����n�H�+Y�h�뮳Y��9�Dy���VRBrC�'#�ga{ca-5�[/=8�un��Dk���jN��Pک�YѧC]�\��J�
���pR���
]֓`�[V���\uۡ�W�[��	��a�&�������vl��s4��8뛑�W���Sv �v�>ι�ű�.��ys���}�$@<��>�
WD�6|��2=�~�w{�o����ߥNy�j�+Y�ݐ.�yy���N֭ŌF'9����a�\��w|o�F2*\n�Y�m���_^��,]78��X:b�v�U�)�G*K;�u`}�۫�o"�=�Y5�ə�� ��(�	R��reLDJ�3�x�=�(�M�fR�7rm7$P��J�)��`}ݚXsN��x�nـ=�59w%]�QUv]]Y��;�7y��5�f�sK5�V�"DQȒ�)2S)�$ɮr\8��g��v�E�Ea��)�B�z{/F���c�JiM]ڻ�7y��5�f�v� ���`}�g�&�S�N	ʰ;�4��H Ŋ�����̙�o�N}:P���@{ה��2w<�j�<���R�&�,秋V�;�7y��5�f ���jl����˚���N��x�nف�Q3�������T�5D2R���`w���nـ�� �w�k)�bS��W����ƀ�Y$�3���v���Oj�9�	����
幝��$st��`�������DB^�|�ŀ}힦�J��q�Xw6_�\��$���h��T�'
��m�T�����9
NI`��K;�ug��p�5S$�2I��*t�/oiP��F)&&¤��Wxkx�nـk� 36�Xk�b��t����`w]� ��/ w4� �o�m�G,]�sT�Z��F�a�W�%��<��c���8մ�r�ĩ�&��k� ;�w�v�� �v��97E)A��)'*�;�[,��Ձ�{�����X�ۅI#D%6�9$�� �o�M� ��, �i��OtnQ*RQ�9Q�*��=�`nf�nI?}Ӻܛ@��
T��K�����`ork�D�Q��&��"�5�ŀ�;�;[ŀoW9����.�9-�Mr؍��b�xͲ�̄�|`wSù�iu���We�dj�Wa�4ʠ�M$�,�ߕ2�d�'8�����9ı,O��p�r%�bX��vY�&���噭a�m9ı,N��p�rȌr&D�;�{��9ı,N�{��ӑ,KĿ����r%�bX���9l�fjL.�Թ�iȖ%�b}�w�iȖ%�b}���iȖ?���/��?���Kı;���M���G)�r��m*<�plJ�q(��Kı>�}�iȖ%�b_���m9ı,N���m9ı,O����9ı,Od���.��-��f�sFӑ,KĿ����r%�bX�����r%�bX�w]��r%�bX�}�p�r%�bX��Aw�I�mն��2�ɮ`fҒ�ɮn��D�n���Ch$:��c��/��� W5��G���8͙�&Z���pw<��=�i���ͳ+��5�[��������a�l�Ҟځ!�N�͉�q�-���7�m��reʻ.�Z���s銶��L��.�췜:8�:�.��������=U۶�]���s2���_[�-ù�e�e�(��T*�nr��L�.�8�'����Fp��\��9���ȇFɝ�\#�����Н�����?/��Ou�bX����M�"X�%��u�]�"X�%�����"X�%�wǵ��i�r���O �)F�9Q��|%�bX�w]��r���,N����ӑ,KĿ{���ӑ,K���V���2IC�������I���Lú���sY��Kı;���ND�,K��kiȖ%�b}����Kı>��ٴ�Kı=�}y�����.5�u�h�r%�bX��|{[ND�,KｿM�"X�%��w�ͧ"X��̉��~6��bX�%�I=,�@HJ "f�2�d�'8��w^�}ı,K�{�m9ı,O���m9ı,K��=��"X�%���e?�_D��ٵ��.dظ::�
vGY쩷��GRnW���V|ױs��^��;si��ߨ�%�b_��kiȖ%�b}���iȖ%�b_���m9ı,O�׽v��r��G+�u��'4R�FܗÑ,K���{�Ӑ����Ȝ�b_k��m9ı,N�^��r%�bX�����r%�bX���w��L�nf�4K�6��bX�%���ӑ,K���{�iȖ?�2&D������Kı;���ND�,K�w��2H�PR��J��_�r��G+2{�ӑ,KĿw��ӑ,K�����iȖ%�b_���m9ı,O{^��'IF��G$W���#��R9K7}��"X�%���~����i�%�bX����r%�bX�}���9ı,����o��N�����Y�7W�W�������A�9�-����ъ��Xl�;���jk5�m9ı,O�{�6��bX�%���ӑ,K���w�a���2%�b^����r%�bX������ֵ��\35���h�r%�bX��|{[ND�,K�u�]�"X�%�~�}��"X�%�߻�ND�,K��vٞ!5f��f�����Kı?{]��r%�bX�����r%��F	�@FKJ��+S�1!�F	���0��j|�PZ���O�w��6��bX�%��=��"X�%���鐦{0х�!���]�"X�%�~�}��"X�%�����"X�%�wǵ��Kı>�^��W�)�r����i���)G#nkiȖ%�b}���iȖ%�b_���m9ı,O�׽v��bX�%������bX�'�I�7�ښ�!u�%����5��=��A1�|]m�kv4��5�v%n��·gVf����s4٩.h�r%�bX��|{[ND�,K��]�"X�%�~�}����"X�'�����Kħ+����D��6�7	%I|��R9H�b}����Kı/�ﵴ�Kı?}�p�r%�bX��|{[ND�,K�׫o���2�)�33Z�ND�,K���[ND�,K����"X�%�wǵ��Kı>�]��r%�NR9[�|H��HҨ����+㔎S�̒��o}�2�d�'8��yt�.D�,K���6��bXG��'��`�&	�+��=Qv'��1�+㔎R9H�fW�*���r�ېY����Kı/������bX�'���m9ı,O���m9ı,Mͭ)��'8��Y�)�1.KĊ�v���+��/�q��iuY�x������}�֎ɢ�g��5�٧��������{�������ND�,K��}�ND�,K�{~�ND�,K��kiȖ%�b}�x�S=�h���K�M�"X�%��w�ͧ"X�%��}�M�"X�%�}��r%�bX�w���r'�(e�;�ow������
C�0����oqı;�����Kı/��[ND�,K���6��bX�'���ͧ"X�%�}=g|fh̗2i�Ff�6��bX�%��|kiȖ%�b}�o�iȖ%�b~ϻ��r%�`,ȝ�����'8��[���	yDDJ��_Z5��Kı>���Kı?g��m9ı,O���m9ı,K���"X�%�P�A|x�L�kZ�F���mA�5�vq[AI��t����2�u���s�PvM��nQ����O�ےt�l���e�re�k�}��^�au���g�	�y�Y��;���xc�ln�v���=�͚^5�D�!zX24���{q=��aW��q�^� muO�-n����'c]u�+�m�+t9�q�x����Xw��K�� JM�VG1�	��W+��9�w���PB`�i�qb�Mv�u�+C�9e;/>4z��
�vy�'.��l�% 4�(1�R9�x�#��R9Z���iȖ%�b}�{�ND�,K��ӑ,K�����ӑ,K������TFT�����G)�r�}�m9ı,O��ND�,K��޻ND�,K�}�fӑ,K����W���&܃NK�|r��G)����iȖ%�b}�{�iȖ%�b~Ͻ��r%�bX�w��ӑ,K���v̅�x�Vh�5sND�,K��޻ND�,K�}�fӑ,K����6��bX�'�w��"X�%��x�r��FT�5n�6��bX�'���ͧ"X�%��}�m9ı,O��ND�,K��~�ND�,K=��w�����~��:ȝ`I�F�n�\k�)�Q�E��ݽh�9�Kt�'j!5��u���a�!;��K�LǓ L��ot��2��x�lI�}��7�%�b~��ٴ�Kı/����fL̺lљ��r%�bX�w�8m9 "`EA�?�Ǒ?D�;��iȖ%�b}�wٴ�Kı>��ٴ�K�G+w|����6�7$R�_+㔎R���ߦӑ,K�����iȖ%�b}���iȖ%�b}���r%�bX����_h�0�W&f�k5���Kı>��ٴ�Kı>��ٴ�Kı>��m9İ?��;��M�"#��R9^���B8S�TFT�����ı,O���m9ı,?�=�����ı,N���iȖ%�b}���|��R9H�#��Z��
G�&'J-�n��(T�I�p'ܶ1���չ���:��K.Hܡ6��r�r��G)������Kı>���Kı/����� ��dK��{��6��bX�'�׮R��Y�,�SZ�ND�,K��~�ND�,K��{[ND�,K������bX�'��M�"X�%��y���f0��3R�SiȖ%�b_��kiȖ%�b^���ӑ,hpT����{T��8(��N>�%%� ���������0[�B<8��2H�}�؉��	A5W�~��:h9�L0�w���P�~�S�~8Hj1ՠ���"kHL0 �k!V�`@�؇���,@��ƒ0�%49k�VQWC0W�,+��2%Q�At�(��6X3��w���ٶ�~�xm9F�ߠD�BI@$dc�!6��I"H�����V��K+�󺚰�f�	"F	"�"��` U�T�̱�-tH�]H�?~�1�6~F?{�)����F踒!��b�� D�
�J;��Ԣ�U1D�#�M
!�U?"o�=��g �PDqC�l:�� �h�Y,�@��Y��~a�(�@�+���蟢w��r%�bX�{���r%�bX�Η����e�[n�Y��kiȖ%�b^���ӑ,K���7��Kı>����K���;���m9ı,K�?���n1��e"H�����#��R9Y����r%�bX�{^��r%�bX�g}��r%�bX������Kı>�����6,�����v.��n�7\�/,a��hY�lhNb��+p0�I�+h�+r�u���Kı>����Kı/�����Kı/{�ka����L�bX�����Kı>��)�j�K��3F��j�9ı,K�}�m9ı,K����r%�bX�w���r%�bX�{^��r%�bX��w��֋���JMd2�Z�r%�bX���ٴ�Kı>���Kı>����Kı>��ٴ�Kı=��^MkZ5u�.\֤��ͧ"X�%��}�M�"X�%����]�"X�%��w�ͧ"X�8HAH����
�� ]r'�{����Kı=���)!��j��e֦ӑ,K�����ӑ,K��;�fӑ,K��w�ͧ"X�%��}�M�"X�%�����������F,�1k��q˒�Xsn�\�	h�8�OV��pA������/\����j�?D�,K�����r%�bX���ٴ�Kı>����&D�e�;�L�8��N2���G0�
^�f�f��ND�,K����NC�D�L�bw����ND�,K�����r%�bX�g}��r'�eL�b_���r��!ȉqA1/3�ᓌ�d�,����r%�bX�{]��r%�bX�g}��r%�bX�Ͻ��r%�bX���9��ە$�H_+㔎R9H�g��]�"X�%��w�ͧ"X�%����ͧ"X�%��}�M�"X�%���;I���0��Z���r%�bX�g}��r%�bX�Ͻ��r%�bX�w���r%�bX�{]��r%�bX�C �)�}�i���sY��Re�I�rn�\& �[�@T��d���c���G�".�A���N{+�i�(�Ն�v*���Mx���v�z�]ym�{mu�?����6bQt��Ġg @��;��X��ӷ^t��;DuƊ)�/F,q�b�ci8��㭧��nݫ���+����(����<n8�۞�]`�֝nm�;/��܌d���!(��.{���w{��}���XNתZ�vn���\�gd��ѱ���-ۋ� yO\'A=4Ĕ�*6��R>��#��R9^~��iȖ%�b}�o�iȖ%�b}�w�a��"X�'s��ٴ�Kı?�{�g�*jJN���W�)�r�����6��bX�'�׽v��bX�'��{6��bX�'s��m9�ʙ����e$0�&��l�]jm9ı,N�k���9ı,K�}�m9ı,N�}��r%�bX�w���r%�bX�����Ra.R��5v��bX�%������bX�'s��m9ı,O���m9ı,O��z�9ı,Of�i�NF���n6����#��R9[���iȖ%�b}�o�iȖ%�b}�{�iȖ%�b_��kiȖ%�b}�ݿ;��.��醂�G.�Z�\ڧ�u��s��H��/g]n]��FnYɖ7;Y��fӑ,K���ߦӑ,K�����ӑ,KĿw��ӑ,K��w�ͧ"X�%�{��f�f\334kZֵ�M�"X�%����]�!�?Qz����ko蟢X����[ND�,K���6��bX�'���6��bX�'���'�j�Mfa��Z�j�9ı,K�}�m9ı,N�}��r%�bX�w���r%�bX�{]��r%��R9^�ߡ$�!Q��jI|��R9V%����ͧ"X�%��}�M�"X�%����]�"X�%�~ｭ�"X��#���'�ӌ��' �|��R8X�'���6��bX�'��}v��bX�'��{6��bX�'s�{6��c�������������i4MՇ.n��H�����y��v��Ϝ\��s����ISo=h�K��jq?D�,K�����r%�bX�g}��r%�bX�Ͻ��r%�bX�w���r%�bX�����Rd�0�3YsWiȖ%�b}���iȖ%�bw;�fӑ,K���ߦӑ,K��;�fӑ,K��v^��sZ�pչ����fӑ,KĿ��kiȖ%�b}�o�iȖ1W���"'��~@
���M��{��m9ı,O���fӑ,Kľ�Y��Ɇ\�CYu�ֵ��Kı;�o�iȖ%�b}��iȖ%�b}�{�iȖ%�b_�����Kı/{�a�֬˅��.��kZ�ND�,K��}�ND�,K�U�}����ı,K������Kı>���Kı>��Y1�\�-ۜ�\f������vip{���^��9�ɂ��E���Ҽ�B�6��bX�'�׽v��bX�%��{[ND�,K��~�ND�,K���_+㔎R9H�{�~���e(�Ɩ�v��bX�%��{[ND�,K��~�ND�,K��}��"X�%��u�]�"X�%��{�9u�ɬ�.��j�3Z�r%�bX�w���r%�bX�}�p�r%�bX�w^��r%�bX����2�d�'8��9!�@&A��D�m9ı,O��m9ı,O��z�9ı,K��{[ND�,"�� ,����$ �X&��D�o��ӑ,K���K�ڔ�.a2f���iȖ%�b}�{�j�d�'8�h��eᓌ�d�,ޮ6��bX�'��m9ı,O�;���?X��k�m;�8f�pIX�6�^'��C;��G��	�*qT�&.��=��5���ı,K������Kı>����Kı>�}�a��?DȔd�-��ze���N2q��<�>kP�]k5�m9ı,O���m9ı,O��p�r%�bX�w^��r%�bX��}�m9�  ʙ��}�s$m$�4�29$��9H�#��V�߾��"X�%��u�]�"X���/����ӑ,K�￷�6��bX�'���'�j�MffLѭ]h�r%�g�$��o���9ı,K������Kı>���Kı>�}�iȖ%��r��~���e(�Q45"�W�)�Ŀ��kiȖ%�b}�o�iȖ%�b}�}�iȖ%�b}�{�iȖ%�b|���F��@/��l�֭5��6�mLf�$D�\�ˮ,Չ���c��e�lIdV��80ٻF4�� �J�\L�m�p�vA�ɹ�I�ܛ�{Zp��-B���Y�Ͷ���wgt�������vY��''2��Ƞv�ɸ�Ō��[9Q�q�h�Ɵs��Obt�ݔ��2
����ܚK����J<��_^گNR8v-����B�
Xs���LL&K��Ma��?�/��ߤ�ѣ9��k���Pn���T�u�e��H>ȝD<�����aљ�\F���������%�bX����6��bX�'�w�6��bX�'�׽v��bX�%�����"X�%����e���֤�53Z�ND�,K��ND�,K��޻ND�,K����ӑ,K���ߦӑ,K����g�n[na2f��Ѵ�Kı>���Kı/��m9ı,O���m9ı,O��m9�R9H�/y-�ʐu��9�9J%�b_�{��r%�bX�w���r%�bX�}�p�r%�bX�w���r%9H�#��b���ci78�"�_+㔢X�'���6��bX�'��m9ı,O���m9ı,O��{6��w���{�����po��i8� �U	���Of��v��nxݜ
��/&y�ub�ܺ�*�m���5�ֵ���ı,N���6��bX�'��ND�,K�w�ͧ"X�%�����iȖ%�b~��{F���fd��֍�"X�%�����Ӑ�@��D��@�m�Mı7��3iȖ%�b}���iȖ%�bsyd/��$)!w[���WB��Qtk3Y�iȖ%�b~��ٴ�Kı?}��m9ı,O��m9ı,O�w�6��bX�'��\浬&�h�]kVL�fӑ,K���w��Kı>����Kı?}�p�r%�bX��{�L�8��N2ݜ� Q�������M�"X�%�����"X�%�����ӑ,K���{ٴ�Kı?}��m9ı,N�{-��٬�j� �Z˅q&����<\�`��;�ޤN_W+���O��.�pe���߭�7���x��}�iȖ%�b~Ͻ��r%�bX����6��bX�'�w�6��bX�5�C_���Q(�brU�9H�#����{ٴ�Kı?}��m9ı,O��m9ı,O�w�6��bX�r��^��m&��R;�|r��G)	����iȖ%�b}�}�iȖ?�Q5�߸m9ı,O����ND�,K�w�sZ�m�˚$�ִm9ı,O��m9ı,O}�p�r%�bX���{6��bX�'��m9ı,O���Oh�0��̙�SZѴ�Kı=�}�iȖ%�b~Ͻ��r%�bX�����Kı>����d�'8˙3&���DLH�D8��:.�+g�d��'E�6nt�s5��7%,p۬��tƬ<U��$6�,�����oq��O���ٴ�Kı=�}�iȖ%�b}�}�iȖ%�b{���ӑ,K����m���p�5�&f�iȖ%�b{���ӑ,K�����ӑ,K���w��Kı?g��m9ı,O��rC=!5�2ɫ�6��bX�'�w�6��bX�'﻿M�"X�%��>��iȖ%�b~����Kı=�%ٞ�%�0�f�ZѴ�K����>��6��bX�'�����r%�bX���m9İ(��'k~#h�-�!A��҂j%޽��r%�bX��}�f�d�E�35.����Kı?}���9ı,O�w��r%�bX���p�r%�bX���)��'8��\��q�~�%Оnp1���ñ��q�y���v���i�|�Ī��r-��D,��e&?^��{��2X�w���r%�bX���p�r%�bX����6��bX�'~�}v��bX�9]��?�m��9AI%�9H�#�b~�}�i� r&D�>��6��bX�'��]�"X�%�����ND�,K���atkFY��4k5�6��bX�'�w~�ND�,K�k��ND�,K���6��bX�'�w�6��NR9H�w�R�l������|r�K?�D�w���Kı>���6��bX�'���m9ı,O���6��bX�'�����S&��ѭY��]�"X�%���{�ND�,K�%{{�)2�foK* L��1�2ĉ� �*�� ��� �*��A Uj��  
�� �*����*��"���@�TP"� � HE `,E �A U� �����V��*�@@_�A U�U�tW�@_�A U���U���d�Me=�d(�Wf�A@��̟\��|�  UDA$E�R�� ��T  
 ��l
P�� |EQHH
R�   P*�          

�@�$�@�RHJ�"�IT*�  dJBT( P � >����wϷ����r{� �J�Y�(���L�ҩW;� �B��(U�� R��      `  @    � `  ���\m(*��MR���(U���1 ���4� 8�PH�%$P� f�Х14,��0h)�
�����1FmBc^� 7B���������J1��=hd�:s2���QX�u_x �q�R��ϙ�&�mr��>x (TB�� ( 2 �A�@b�w3���� �K3�N�u�Ӟ������� �s�{���s� �x�w����� �y+��s�����<s�%w �u��Wst��<w.�wy�]x � %B��   ̀ 篶{����9��&�nl��x��,[�S�>Mŕ,�:\ ;���ޞ��|��iw���[\ 4��)���&���{���_< q�3N�1Ӯv髽ޞW�| ��� )T <�&}���<��qezr��� �[qs��'_-9y/g;zf��r��o{Kŗ�  /s�N�w�/+�B�t��݃���o.��q�w ��X��95�\���w�����IJ� ��jf�JT @�=UH���&  �"{J��H@A�����j��! A
B��" <S�N����?���i�y��{�C!)�Og�=���cw��
�L�9�"�*�TQEO�T�"�*�����*�(������F���l?���x^sM���߼�A�M�8��N61��3_���X,��M}x��uc��#�˩yx���Tj�Q��h�K��6���/���� �|$a���y�E�|�6F�Y��'	�^^Y�4����GG���z��Z7��><ꯛ<����D�0���u����y�$;T1��A�@S=���5�н��Ff�7�9��|3��B�s�d�Ќ��#�dDa��K"IY�e��6Y�sI�c��C�8��LT�3���Ip����y����m_h�F��O7�Z8h��8�S��v��lf�0�gֶ�}��r��`�@�]��1I��BXJ
	��m3�y�#ϑ��EB�&� R8�:� �J� ��f�zNki#�����k�k|9�t��~>OO�lw�g$��FfKDbL��x�h��A�ꐠ��s0>��v2a�f�X�`���MN{&{"��T��+�ii�M�9j�ͅ}β��L$�G��DJ�r�盥)	�}�	�5kE�l�y�a�y�=��#	)!xp���u_	bi�"Rq1J�s�L��$D�*��!51
́9��ӥ�U�Z�!�0�*_M[ij�ߣF��T6J��t�[ˤz���xZߞ�蚨��X��M.����Qg�a��F�( ��<�f�>�.!��1�E�[�A8f�1)�uFV�G.��4��m�Aa�K���A�ݧ��c�����4a'�N2�$᥂ ��19���{�ﺍ��H�}_W�T�E�p�gyn{�~��MF�z}6�8�6l�����=�3~�2�}�|z���aVDƂpKTp}ٟ:mu���{�㴘7�;�{�y�@�A)�#�*@��|^:�;�8�7��K޾ͣc�u����Bj���3��h��_Ȥ
�|τ���k�}�~�.�R��c�H�bB=I��c�'�ϓ�Ư�i��6�k�о���^	��T�}�R/sR}�R����FU��Nr�%�O�T!�u$�k�S��#�z�vs�[p���l4l���BNY��ݹ;��`�^�O~N0f������<}=~ߞy��9A��V]���}�z�%��_�nR��I�X��5E��Hr�d\o���xǇ�8l���M�p=%� �$�Ya#�1a�'	)"L�3��������?f�ğ)M����O���ۆ��K&&k=�o}Y�A����G�B��j�� M�T	!5%Da:����j6�[tc�޼���$�Hd~IY�j�8��H@��!�^�*��z�J~kϜ��*i��kQ^�h�h��p�p���4r��D`�����f}���{͜�'�� ��,��}����a�E��:�xS��Y��|N`Z��l4F�>l�&����~���e�ޢ�.+����I)8$�`Y2�X1�	MF��w�����3>˒W<����샳׾ǎcX|FjfI �2=����qբOnp��4ll4C@N��[K7��4m�ۘF,�ha�"CD�Xt��a&s����<����Ք�$ā�I`!��p �R$Ĝ�
1�
�HĐ�vRZu�u8Χr1�	t6f����0�٦�l#5��5��5P[�4�A�da8���[�i(7D3L�r�i��[������
�σ�&���7�E��9�ʅ%�H�$ML��3թ$,_MN'ן%����Z�.�E'�|��,����1'>�8kk�L�!��D��鰆,�ǥ���p�#�~�c�k	�3��2�d`�@D��m���]�3-��oZq&�I3A���Ĭc59���g,����y���^k]7�գ��H��8�c.�=�y/��Zg�.Z��ך��U�j~�|�^!�.)��@����Y���,K��~�Xy��כ6x@H�Z�f��##4�fϣ��jt���6+�$yi	���S!�#{�xTP����Ӣ޹�fj���<ۂ�W�r_��+!4��o4czAX5Z>�7���0�Fl���}�<#����3l&�4I����ba���f��9$Y�XPU#[�C��[���b���L#��p�j!�O��0���������b��	8�H��J`��Y���fE<	�14l8����di �i	u4��#<d�j���HD Jq �u(D$��J˲��&l��OsC4Nh��L�aMI�A�T�1�$`�i#dÇ��}�O��[瞚�/�4!$�/�L�ɈQ$�g���>ϵ��`r3N���a�a��f�f����4x��Bt$RV�����ӷ�{�	�[��֤�Y��꽏x���}~v��PF�C&%�af��"%���N��MN���o����.���/%�+�³�yg���b| �E�l��i4�o��m3C��v�5���h)A� ��������|��#9R}#!��B	*Rd�52o�#�^�5�g7ɬ�9�}��Jj.���:�TV���s�+��áj�c�0@L1�'����h��~��sο|��IS4;H1�F5MNk���3T������0�9��f��'���V�?/];��w.3|��Y����X�=4����Čb�0Ó�3�MN?!�$��ID��H@a��8y��i�,��y��Gf<y�I�4�t46h��R���!�=)�v���ux{ÔU���Ri��~�l�})'����!�i&	pCE	�FM����`���x�S��Z��5�̈́����-��G��y���zzf�v%	PI���C1�B�o��fk��<������DxFPI�3~oN�h,��ɮz�� �Y�U�y��_q��0 �;xN�6��Rd�� ��`�� �F�`10�J�f�;��(��vDF�7}}�]>ݑֳ0��C�Ǐ�#���c$����4l,5��N��Aa���Ώ����FRA����!U�� Bū�|}Mn{Զ���YHG�:��߇��<��	I��d��Ͻ;� �)L߾��.6w͢��׬�--���{��%k�V6!�S]y|�� �!�+!O���G�燉f��7���g<�'\�f��l���R\�U���k����*D��[uͺ��F��Γ��e\	�t��$��i<N:�ѝ8F�1!���.2�6xTF����$ƈ��$c��Y�.�5�:YhvTf�F�(d����U:1�4m�X���kS~y�Y�y��[�p��#3�\f�z�b� �YUOa�H�2~w蚭>M�ȅiМ�j�2�f}R�����VVE%�H
@�I)�!���!a8l�+��j�m8�"���kcR`�JPD�C�*��Y��L��L���l��@`�Hd�ȇ�wW	�Z��j=,�~�S��G��f��t�j�=����߁�9{A������t�es��SHdCR�!'PԂO�����*a�S$H���$��lá��1�n0l���o�3.6N;76Z%Ą��lf�+����	&���� �c&�S�̍���솦���e(��!"��(,��B �U �C`�Z�t���͞��ּ�;�:��|30%�+LBJ'�{�:w�ߞ�����|8   	 `��_ �  h  ���  �$�  `|�<��r�ր6�[F�����Q�ہ������   -�          m����0m�`k�  ���ρ��l     m��i6 � -�K$m�6���n�� t���n�H�"�%�dP�ki�lL�T	J�t������|�*�v�ԫkL� $p�8	� 6ݍ�r��$-���` l� �u*孕�MƮ[���vqRr�h	@ڳl�������-UWmU��	-��e�h��$�I��-[����     q����P��U���>�����mf�,�8�m�ڤ�Aΐݶ6�@N��1U�6^ʖWln*��e��l�s�S�,�l��L躹��
Z5�,Rz�Y{8[iV��v��m�M�0�7l��#6��.����7ZӀ�4 �Ce��#[j�2�(]k�gP/*�Ãd
���"j��u9��U..�6�8�AW/sfj���S�=.�э�0�V����ԫ�;m�ۗ-OF�����[%eH�sm"u��{]�]�ܗ\�ҿ?z�_��|�}󛭷L�YN�y�T�n�HJ�z�3��pc�*�m���شa��)u+������_R �4�S6$kՍ�e�����f��� +es�������]X�v�3��h
�`�RZXF�j�n��U	��\�I�M���@$s�"N�k�-86�Nl�d�(�9���mm���A�Í�9mI�� �	���r�Z�������N� �6�{ p6%gm���'Kh  h��ŷi6$+[]�^���� l�mnգI-0  ��@v��lX����l�r�jz�B@���0-���u�[f�p  Fٶ �  �ְ   H�R(���n�U�@ ����޷e�� 8n��6BC���[&�l[��h�  �֙z��N$�����`���Fݲ�  d&F�l[@���`	m[� �      [E�d0�ml �    'iX ��6�           �r@�uö�;U���m�H9�q5T��K�[��
U�)���l�]�� �o��     8���m�ǉv��% FצΛ[Q`  �	  l�tͧNݛlĚ�|;�I U*�[UZ����~��:h-��;]7KZ�Ԁ�JMj�y�h
�B��i6m�r�W%^�*���-�ʲ�J�j٬SI#n�[O����[B@  �a&��`t����lI]���v6�1�$	6[� m��N,0+U�ޙ�  ��!�[[lɱ6��հ��hhn��� [@  [{j�         ����  � �l   m�m� -�Io0 �   h$    0�v[\ m�R�8[MȖP �    l � C���@�� m�v�[�^N t��l�MV��`l           � �� ��       ����    m�m �`  -��okp �v�`   �l�-1m \��m 6�  nձ�K,�� ��^�P�� m�tͶ�m���Y��  ��ρN��h�ܙ�C���*����  ]@+�U  $ ���h 6� m���D��imI��e��	��0A&m��.��	� ���[@ �  H  $kL���H�M�6�  t6C�� հ	��qͤ��Z��n�l���h�N5�)d -���a����0&۰4P�۶�7`����  � �     p  [M�gm�@���   m     � m   i� m�`-��    ��    ��H �  m�  l6����H    )��c\G|�>_�O�-[nJ  �  ��&�kd����  -�n�` mÀ	 �` ��f�.��H�   k��M��m[[l      m     k�� �o�  pɴ�m���  '[vؓm�L���   ����t��!���<�m[�`h�	�۶�i0�i� h�p  �   	 �ֶͧLֵ�l [I$8�]��&���f��`  8 @ձ�սD�  �f�m��tS` �;m���a ��� d 	�4�  &�)@$ 	$[M�V� �Iz�v��[@*Z m�@6�m��n�m�	$��m� �����rBX�sl m�t�L��d�  �nC�d�ųN� 5��      *�VP�jmS�ҭ�P�     h ]6;���rޫoh��K(u�b� [E��lE�Η֒� 6Y+���iy@��m�;��Uc��[9����[2�7 c,n$������$�݋�6m��':��d�٥t�vɬ܏H���5� G-si$�^�SF��n �\u��
�i22�T�T���g���ge`m�WtV�,[�Ͷ kF��جÙWl�Sǎ@�qV�����[��VW��һ2�u�u��j70�/�RJp[`I�5δ�-��Y�crm{*B��M��+�Kʞ6�{{*�[�Z*��UmJ��	��g�?�����׆s*�O-j�z��m�].��n�P
��@U�mn�S�U�le��r��8�:�U�)�,�ĸp[��¬��V2-W���3�����C���Uۭ�I�H��l��S����a�������	�X�Dv�wm4�����+[Ƭ�E��_Z�v�鷱�R�����(M���z8Cd*ڶ��I;A;=����\�<�(m���]"�NYx�q3��f5R�����.k�YX
�	UW�j��Oe;M�ܯ�7QbZ��JÑ�ŶN�m��e�	��[z@v�vƷ^�u*���T9Cd���ڪ�Ulj٥Z�yXpѵ�� �����ls��4U����G����iv9� �B�W,���Wj��WҵF8�� ��m ɑ��^��b:k���R��� 8�UT78kfC�x�Fa�_�����7 $�nخl�5�ۑ��km��3]��,��s��5�GgtJ�UTF�:��p��!�gѸ�%��SJ��R�M����V��r��u��L���cm�Ȫ�VNk�a�T�N0���u����۰ Kw\�K��+��W*ݴ��!��Q	p�MJ��6���q�(n�l�ƥW���R�uK��mU�d��68
4y��x6݀�l ��m�Cl��Ul�l;&ۊ��c��  l�f���������Y�=t�*�O;����@@ t�m�-`��l�`��S[�i.�    � ���I�CFK��ɲf�ʶL�lm��@  X6�d� �ln��-&�:nix[x��
Y�� 2�VʵU�pg�����E�HXrK]���[�$�Z/M��jn�%zk�NQ����Hlu�\�R�5�c����D6�;y���E�&ڠ  *��)x����U��s���d�-�C��$H	��DHk�lsV�ڕ@�+F��%�p [AŻ�g|�O�v՚�ji@�T��d�6��R��w.��p.��I�ۆ�nBjؽh/Y��6 �jL����>U*�a�������Q��YT�8�i�*�WX*��u��T��nj�ST	۱m��m�۱�bYp���Zl,��c���u6�8�-�m����xР=��;se%j��8+jpԄ�ht�	R�p,0[bZ[R 6�Ÿ[@���͑{l-��[�Ue�j%*ѥUK�ҭ�iVr�P���r�Qm,\N�V��\��:�� [ �S[mmԅ/clk�nK�T��.ٶ;v�YE�`څ6�.�� K}V�X��,���[s����q�M*��#nө$��\-��b� ��[��p�^$0!gO3F�{�;-ʁ]�ݞi%5A=�k�r>��BH.�O@���� [wh�ඎ$�T���J�Eq5=��U{m�P����m����b�gH�e� �#��K�9[x H�K��;n��` ���X��jZo`	�z��݉6]��$:�^��6��iWV�-�4;XU���1[.M���  k���8����<W�����ڲ�-�{��{����?̀'�> ���7�^ ��� '�**�FF����`_AA�*��<}`@= 8 z�)�<_N>>'WH��a�Uv�aY����HFX��^����;�@vG�)@�Ni��8��q�
��6������`4�d(HH�m��<:�*�4� >��&�=}_6���l�Gj?
,��*� �T 8������1N�����K�@<T���� ���"}��H��) L�*PE`�x�>��NǪ` {�U���iP�D�QS:�*:�4 z|����/��κH�]�x��@L1 C	2����'����*���!�
0�k�QQ�v�"��!�2���I�qAW����
�	(�0�0��"0����! �@��P"�"�*�߻�ox�Z����ܙ�� �`  �i��l D��i���Svt�kL��S���:R8�`�ә1��e�����U�f��;��3<�:⣣=)�GI��Y�h�g(����/�oC>�4�<mۣ]8�` wE��on��`��S�crsf��uF.�۴m̙��E9�]N1x����f�w[��:6�:�9���g�\�M�Ԛ�]�醴�$C�8ؔ���t3��EiN��a�΅i`j�a,����m�  �g�q��1�Sb�v튪W���5��-�m�M)����EkcbQ��.��l!�
ڕX	P��,��lu�P�j��ɛ���Z���6Ѻ�Ͷ��!�K��I �/Z� �[p�e���m$��Y�кک�f����n���V�X9Ю����R��,��a�,;��1H	%�.p ��e*�j��-4��8l۱��M� m,�d�fnI��$� T� +k8�U��� �`<I���,�5��Fwg�q@�� ^ej�U�r9�Y]��9��n��OԼ�n���L�u�x+OI��y%����[�'69D������`� �����7! ��F�u�:�r��]��ۈ[��r�n��`yt�Rx�=�^��Ό�`�9��u��v���;�Z�	�ȱ���=���cgz�ˈ�p�e���R��i�;!�h���U��)�@;f㝀��ܻ`wF����^�T���N�4�Z�k��w��*b��<�a8�{p.^��z:K�(6u��dHR[q���h���E��N�ฮi�.%x/8�y䷁7%��	5���v�`�.�7j;=E$ l�#B�ؕ�Vx6���U��i��ئ{0�	��Ln��z�\\,�N��������J޲��Z㱻D�.6����iιg>VŨ����#�!٫c�%RqI,& �llk���<@fQ��!��A�~w���޽���w�����l���U_�w~o{�d�^���,��V5ƌ�r�ڻ\�����T��97�=h�g9�>*�ݭ����H<zۍ��͝���۔nP�p�@F�n[b��3�lg{`eU�h�k�8&m0�أz:���j���1�긢�v�-f�Y6��4�mz�Ϯ�9뮶�jd�I�çV��4s6��3!m��,Fnz5͐�ӭ���&�D�q
.Ԧ�a,R刖�'q��yݑ�EL�Ó�ʛ�p���.�l���c��=�h�����/j�h}Z��)�s椙�|۽W���� ��ՠ�4�+��0YH�I)&�[l����m�{��;)�k$cƚ��@:�@-�h�@-�h����/䠱�I�4N���})�I��S�K�;���v�<ѹ��n��@�C�n.L�u��7E�4�������Q�@�BT�.�� ܞ�;��z� ���oY�\Y�U%?L���8��z��?`~JȆ(q�HIR^_0���{v�k��ₘ4�S D�$�o+4޳@�^�@-�4
���"Rdň�	�@-�7�������*����Vh��"ȳ���un6)'�t��`uN��&ʘ�:t���|����������vl������/��f��u�I���d�g��u��Fz:�)���_��y�+4޳@���;/,��#jH	ɠ{�� �ͫ�͵`��}���G2z���n]U�woU��fڳ��B�P
#�T@H@�:�u��*��\�<]�ǉ�ck�҃rh�]L	/�0ޗ�N����%\�t̙1ē��Z�� ��\�z���h�c�����"ō�"Œu����3Ӎnܐc���v����-WT�n���Վt�1��"p�- ��\��f��e4���<��jț�A�BGXnm_$ٻ�Ł�;��>��Հ{xiY=�n�����~���i�D$�=��VٽV�5m���j�b�2�����t��l���/�$��Q3���-ƵXUI27.��N= �s@-�4�ՠUz�޹V6�8L��	�X��P�5<�����n��[�,���wk�6˺y��)�`I�4޳@��ZW��:�4urLpM�s#Jɠuv�����k�oY�\_��LɐsrH�
�W�Z���H����>]�6��[t�2K�ANB���P߻�U�gwU��۳`f�i`|�t��)$I�BF���f��Ͼ���0����~�����~��R��w^T���29�S��ؤ)�X]sul�/y�������a!�G����Zs��$nѺM�#�ђ��-�,Μ� R�V�<:-:�����)YX�HN�J���+\��jU�.��]�mѰJa=�u��!ƫ���ˮ�=yL�����9o=�������YvZ� ��\�m���3n�������h:����Ө������ß׻�yξ�͝ՓX�8�s�vF��&>���s�B]v�6�]�݋+�nl�I��T��Mzn�jf�U(��!~���8�)I�{���JR�gw�)JQ�ͥD �^�m2�5*������)JO��#�Y���s���)C�����R���s�R�������.]UT��E�"�cڸ�~��JR�w]�qJR���]��B�x��L��7RJ���\B�A�!�����R����~�)JRw���R�����|R���߻�Z2]:TU*�麪QdB���q"'}�%)KϾ��)J��v<�A�$�b۞rۙ&J�S-�j���N�49e�c]��t��k�L����ۯ�u�vl������)JO�~��y)J^w��|R����wi�QU�JS��s��n��r�,�ANJuBy)J^w��|��':8�o��ѵ�����m)C�߼��R�����┥'��{��JS�����i�����jj�D Q�ͥD"S��{�)JR}{��y)J^w��|R���ӥ�w��o��ս�c� ,'��k�R�����C�JR�w[┥~��JR���q�Z��l�[�{���)I���C�JR�w[┥~��JR�~�w�)J��r���Q� cL�51�H�.�'fnF�-��
�7��FxJ����V�e�z��Zއ����~��)J{�v<��;�w�┥'׽��{�!�Z���d)755q"(��ҋ!)K�w�┥'׽���~��D ��Ქ�IER�n�UJ,R����s�R��^��$0�
R���w�)J���y)Jt�3i���T:SNj��B��^�Qd%)y�s�┥'�{�%)N���B�
33F��cr���#����JR�gw�)JO.��JR��{�qJR�ﳽ��)߾��7oZ5oY��0h�[`��ݙ.���sy퇱ӯm��xRu�&�j-�9˹!����=�����C�JS��{�)JR}�u�y(�q�\B�
3 �m~��s*�-o{��)J~Ͽ~� �Ug%);���%)K����┥'�{�%)O/lmĹ�R���UM� �A3gE��/;�w|R����{��)����B��[�6�7(�*��j�.R������JR�۽��}�{�R��^ȁ�N�}��R���cdα�A2��Uq"B�l�<��?+>����┥'�����P"�cڸ�!g�d�T��ML�SSV9�5l��Of\X��{b��	��������SgkΖ�p��+/{���O{�/߿u�)JO���y)J^}�w|R��a���ȄSXf�aJ��U$�UU�)JR}���R�������)I�s���)�w���(}>�u��e�ޢ�j����JR�ﳻ┥'�ϻ��JS��{�)JR}���<�A���%��j��n������A�>�}�JR��{�qJR������)y�����)C��w���k-�5���k{��)J}��~��)=�}�JR������)>��t<��3�!	YQ�w��ٽֵ��{�l�YT��и�y�q:#�
�.�=�%�yNC��=\=Vή[�־�3��by�734���ڥ8��W� ���֩�4Tj����H5�c�yj�*��N4v��"�h��n�Y�W%���α]���c>�q�n���:$]\��ٹ5ι���Ƕye��,�[϶�NMZ�C��jRI'GV���v�7/\̦ۓY^�{�㝷g����$v��������F�uӮW'�s���Bt��'�9����bjS��]T�B���ߥE�"�û┥'�~���{��JR�|�j����L�UC��D �F{�R��]��JR�}�w�)J���ʋ"D#`<Z�ꁩT�&��)JO���%)K���┥'��]�����~��)JRv��WJ�����3V���y)J]����)>���<��.����JR��wC�!B��&�*\�ҩ&����!B�����R������JR�ۿwCdB�g�j�D ���Ӗ�d��5{���E���$�
�l�ׇa�u;sWl�rs꧍h�s35*`�ʑ�u5dB�}�{\R����{��)}�{���˄B[��dB���[���*���Y����)I���CȀ�/�@x�J[��o�R�����y)Q����!B�a��v�Uˠ�5��|��.�����)I���ג�����R����t<��==��\u�o�yo{��)>����R������JR�۽���{��Ja/��Z�[���LӪ����"D#}����)I�s���)w��|R�,�ڈ�!B����:��X�C
GA��0��ㇱn�`��c�=;����p^8g)�2�)R�uRƥR�_D �A9�1�)w��|R�����k�JR�ڸ�!i�[aT���T܎���R���{�)JR}�{��)w߮�R���;�JR�0��WM��������o{┥'��v���.����JN���#�ںSH�.���B��<Xu	1����I�X�0C��ε��sb���d t0Z�D����'�h5��8��%�����4�9�M�#&i1W�ǉ���l��M4V�)�ZM`���������x�v�3�-:�1pӉ�D$��l/|O��
���6�����Ŏ&�����
O���y)J]�{W�!���fhnIrU�!UB�!)K��w|R����wc�JR����	�U�N��C�JS������&�StJ��D ���J,�D������)I�~�a�)y�s�┇�hJ3�(J�����۟����q&�z����<���"�@zx�-�[�׶�g�k{0u�Kwܔ%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg~��~x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	Bw���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&{����<��(�B!"��(JY�P�%	BD%	BP�&f	BP�%	����8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP�?����kY�њ�������%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	��w���(J��(J��"��(J3�(J��J��(L��s���J��(H��(J���(J��"��(J3�(J��߿p��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg�~ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�P�B/.�K��r��uT�o	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&{����<��(J!(J��30J��(H��(J���(J��;���8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP�߿~ߞ	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP�~�a�(J��<���(J!(J��30J��(H��(J�ý�;Z�n֍٪�f����(J��J��(L���(J!(J��30J��(N���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&~������%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	��w���(J��(J��"��(J3�(JL�!�]:��(J��3_�~ߞ	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	�;�?do{�e���f�5�	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	Bg~��~x%	BP�%	BP�%	��P�%	BP�%	BP��%!*�������hn�~?��A�A��{݈<�����wA��I�Bn����1L�n��/:gSt�n����ݍ^3���h
y�����|�[�kzٽZ�����	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	�~��pJ��(O3�(J��(J��30J��(J��(J>�����J��(J��(J3�(J��(J��30J��(N���8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�������%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP��n����5l�o5Z��P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP���P�%	BP��	BP��%	BP�%	BP�%	��P�%	Bw�߹�(J��<���(J��(J���(J��(J��(L�߿o��(J��(J��30J��(J��(J3�(J�����8%	BP�'��P�%	A�ː�%	BP����(J��
(@�g~�H�n���R�(�����J��(J��(J3�(J��(J��30J��(O�����(J��0J��(J��(J3�(J��(J��3�~��<��(J��(J���(J��(J��(L���(J������%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�&{����<��(J��(J���(J��(J��(L���(J��������ћ��%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	�������%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP�~��\��(J��(J��(J��(L���(J��(J���v��<��(J��(J���(J��(J��(L���(J�~��	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B|~;�/f�[�fj�[���P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B}�_�g�(J��0J��(J��(J3�(J��)��J���_���(J��(J��(L���(J��(J���(J��?~����(J��0J��(J��(J3�(J��(J��3�߿o��(J��(J��30J��(J��(J3�(J��ߌ�j�9�9�I�v$I���H���Jo9����Yx6x���#�</�pmv[R���E��\�d؊8VV�`��/���T�ł<t�7;���l��V�.��4)Nۡv��W
DԺ�`÷m*�v�2�Ц��/cUs�9����c�x��^�m����	q���e;N�37Y��� j��.�q�+����(�`�M#�Y�ɴ�������|0.۞./Y�ڥ�2F:����g�w3
��;b�h����� ^��{��v��(O3�(J��J��(L���(J!(J��3�������%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	���ÂP�%	By�%	BP�$BP�%	Bf`�%	BP�	BP�%	����~x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B}�_�a�(J��<���(J!(J��30J��(H��(J�÷p韲5��ou��o7�P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'{��	BP�%	�`��	BP�	BP�%	��P�%	BD%	BR�~�����(J��"��(J3�(J��J��(L���(J����	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�&~���~x%	BP�$BP�%	H�`�%	BP�	BP�%	��P�%
5������U*��ҵ PP�'��P�%	BD%	BP�&f	BP�%	�%	BP����o��(J��J��(L���(J!(J��30J��(O�~����%	BP�f	BP�%	�%	BP��%	BP�$BP�%	Bg߻�ߞ	BP�%	�%	BP��%	BP�$BP�FI�����"���8��RQL������ ���a�)w߻�┥'�w�JR�~�w�)J��n��F���U��<��.��s|R�����c�JR�����)I���a�)�^�'����Y��^:Q�R�`5E:ۋ����LA4�n�D�Y��X��)JR{�{��)�����)=���� ����߳���)C޿���mR��iE�"?nͤ�8�iJO���%)K�{���"�v�Y�!y{�Ĳf�RrRuU<R�����py)J^{����80'�w�JR�g�)I�ؾֶ�NQ3N���5D �G�׵q"
O~�v<��>�{�qJR�߳���)_a�Y�F��U�5����)I���ǒ����{�)JR{�w�<�A���j�D ��ݡ��䩕\K��E���r��tȅcB��Xs��l;�<:;:�WH;��o{�����~��)JR{��py)J^{�������u(�!B��x\����5@���{׊R��~�߰y�2){����)JRw��ly)J}���⟃1@Q���E4�EJ����5D �G��k|R�����c���`L���@�@��4�H�c$��@C�<-	) I"B�ED
Dm9��O����┥'~����)�j�n�*���\�ꦮ!G!&B�����)����┥'������"!����!B�r��sM�R�z��R��}��R���;�JR������)>����R��t��i^�u��v�^�ڮ[��K�#�ݍ�g ��v۳���_���g�-qS���)I�s���)y߻��JR��ݏ%)N��)I�ؾ���k[�oy�އ������? NJRw��ly)Jw;����)I���C�?  Ò�һ�/ڲ�ƵZ,��|R���~��R��}��S������JR������JR���N��ݻ{7��Vkc�JS�����)=���y)Jy�ϻ�)B|�UC�M*.�L����)�;�l����z��y�)JO{��%)K��w|R�����c�JS���)J[��{����?��d"��bT��`��vQF1���]��n�g/=lP�e�t�vN��޹�����U�o�JR��o�┥'�w�JR��]�qJR���{��Ja}��[���eI$�RU\B��;ݏ%)N�)I�s���0��W�!�̓QU"sM�SD���)�����)=�w�<�� FJ_���|R���~��R����-�*\�*N�����D ��{�E�)w߮�R��}��y)A� ���鸄!yp�B_%2��sT9�<��/=�w|R����?�l}��?g���)JO{��%)O�|d:t�9�]��[��Z�l�ѡ��ܳ�O[-ō��+n��l����[��-���9k׫!�gK��Suw9aca6qǚ ���N�T�g�	J搈�mv͕@W��B���F�Ø/Z�uL�YMF�s��C=�;�]�k�t�1��<n�S��2g��\C�6�������}m�H����a�Ǝ;��[
%bۖ�gے�hy�ݶ����y~��#g�S]tv;k���n!�R�l���>�]n˻2.��9wO��Ռ;��ѭj��R����ly)J}���┥'��'������?o�R���˦jb��*��ҋ"D,{���rR��ߵ�JR�~�~��)>����O�Jt���_�U2��MUT�B���xQdB�g���)O�R$�~��R��~��qJR�ǽ4fkVh麵j�[����#���&�~?��)JO߿��<��>���qJ� �'߳��JR��˥�$��$���UW�!,��O%(�=�����)>�~���D#7�� �A76��4H�ҩ�2���.1��]T�ݴ�e�l�i�gJm��H�bn�1�N�3CR��sJ>"D-}�6�)I��{��)}����.J,��QdB��֙2�˩T�S���)JOo��#��:@�# ��(`�A ��!*
~6�JZ�����)I�~��T�wf�$��Aˎ���Je5����o������o�R�����y!�����;����┥'g��%*!@cX�F:�J��Uq":��w��%)O����┥'�g{��J�.w��┥'�����o�7�z��f�<��=���┥�����������o�R�����y)J~w￟�H�;nñ�BZ(�d87��A�&e��nz�sk��6��qѺ/��N��{���)JO{�vJR��w���)I���ǒ�����\R������,:n�Z����)}�zo�R��}��y)J{��u�)JO{�vJR�{Ӻ��k�f�Z��of��)I�{ݏ%)Os�;At �lU����_��)y�ߍ�JR��w,�f�kZ݆�n���%)Os�)I�{���JR�����)>�{��)�������of����oz┥'��%)K߻�|R�����ǒ����{�)JRw����s��'�U��UQ�;��3��)�M�I�=`zvy6 �>p�-ܽ�üJR��w���)I��wc�JS�����)<�w�<��=r�ώ��7�i���|R���ﻱ�)�}��R��w;�JR�~�M�JT�Z�=t��UJe��UR�"D#~�w�)JO;�vH~c%/�����);����R����wq�{��ٛ����R��w��<��.�ޛ┥'�}ݏ%(>��U[��w�)J^�Tfh�麵j�[����߻�|R����=�l|��/���|R������R��{�f��1tt�D��[�ĥ��\uGu�m��+{a���\m��9���}�v���ﻱ�)w����)I���d�o%)K�~7�)J߿fg�[���Ն�nֵ��)w��|�NJR{���%)K��ߍ�JR�߾�Ǆ.���(dB��H:���E"i���┥'�����R�������@d�w��<��.���|R�����73�L�f��K�Y��$�	��┥'���%)K����'���"D,�n��5-ȦQ15;7�)JO~��JP��c�����┥'߿��%)K�w���)I!��'�X$+J!�tE7Ȣ$Zd��1ȩ�f؅vnn�f��C���4l�D�c�	�:UӾ�^p�u�Sy�zFY��u��$��v6���6�QJ|!��kÒb�ӨRK�@��H�Bai``d��b"+J&��1� �x�#@C2El���R~{�_���\��RIeub�ڒ�m� 9�j�,�	$q�j�m�Mҵ�M`ڷc��csѰ$aR8"�f%IC�6�a
U�&f�(�v�-��e��p$sq.�6%��|j�]
�����8��s�ȁ�ήM��X�:����	��&낧O^��әӦΝM�ab��#�Kl�+/g�mcMra�3��=Xn�q��u
Y�b` (��P �Yl��ʸ�kf�[�v�fd�	5����( m$�6�H�%�3lZ]���&.����ڳd5k��%YUm�H�u9qMQՒ2�HL���7e�y��X�e�����V��\���j��j�ۥt�2�UUa��Q=����m�m�m�I��mz;i��З&ĲC`�MgJ��5�pm����gT3E]UT���w1��ք�I���&��`%g��N6�m\K3l�6�v��jU���5T��=�ke��5Ht��G l �X��rX�����mn�U�*&F讥^{;/UO͝a�R�;U�Y�۝����e]���u�z�8��t�Y)b['Z�	�dcj�;k��p��s�eUrv�m���ȓa
�8�$r�j�q��[�3�^;g�/����l�ۨ{/�cq��3�QŒ�Zl��]<�H��[�ضӻ]���ެ\�2f#�O����}�v87ɯX�֝�,]�;���[*h��^��_o����,�vذ���;�cu8qdv8���K��M� ��F���	;�������غWQ�ORu���:��Y �Ɍ�ؠ��Jq,5��T��!����Jn[�c��V^�i�YΏ!n��K��v��1B ��㱲�R�4{Zm��u�Bl6dwE�u�vݶ]j�,aQ+�{O7Z�Y��DB�d^9�捓�F�	�B�^̫uQ�u>:)�K���l�mgF�~����[�v�*�9�=�SBK+��	��`筞e����e�f򵭠�~:��M� ;�t~>U@qP�@߽�{���w����! -�M+N�+e��m��]f맬�v�NY�ݛ��I��뚛����R����}�Jʘ�7���P ���c6�K�����.ea&�xT8�E�)���T��R�y��l[t�vfy��8�k�l���Fs��jN!,l��naw��{ �H��IZ7V���0�k��fS�g4�3̛�;v��s�ֱj��!�m��n�&�K]u������w�߯�?�V����`���M��%��IM����1�&q����	�k}�\ݏ�v�{5���,��|��>�����)<���<��.�ޛ�~	rR���`��!bxp�Ku"�T�:����'�w]���/�����~���)JO߳��%)N���s����VkE��#V��nJR�����)JR}�}�H~D������\R����O
,�A��=L,uT���4U�R�P �;���JR����k�R��w;�JP~ %����|R����?�:�SJ�ԩ����"=���(�UY���~��JR�����)JO�����;Q�Ѯn�sx1p���9(b��AJ��)�a��؃i�.n��{���ݟ��{=�?�{�����ߵ�JR�~����)C��wi�"���R�����\R�������O�DJ&i�T��E�"��U��"D��$��EG�	�%);~�懒������qJR�ϻ���?��Apu)�/��?�e�F�Zu����);�?`�R��}��S���=��~�������o�R���Z��rP���uLuME�:"B�����┥'�����R���ݷ�(O��@Lԝ����y)Jt���k�޳7��͙����qJR�ϻ���J��~�[┥'�����)�����A�ےӑ�*B�LM�jiC�tGR�ʍ���8��:m�{��7PkjX�������dh�V�	�74(��A��� �)=�>�%)O���\�U�T�ԥ'�����������ڵV�Z�٭:ݙ��┥'�g���~Ad2S��ߵ�)JO߳��JR�������ET3�����۹���f5�[��|��?g���qJR�����zi�
?�(�ᒗ��<�����sQdB����ZKR������)K�"(��jO������)~�o�R���w�<����
!C�����'H��3Nhni��{���z���������?~��qH�Au�D �_{wNd�۪mU(�7cna����#B^�=���ƻ��s��Y؋�����kv�3U�[ٽ��)I��~���JS���┥'n��O¡y)J_�����)I�~�Y�[�F��5���Y���R��~�8�P����~��C�JR�����JR�����\�I
��V�|���JT����R����~���JR������w���<��;����)J�]���Z3��պַ��J��EpM~����)JR~����y)J{߻�)B>+c�?�2O����%)N�~����:)L���J��A�c�i��@g?~���JR��ߵ�JR�};��JR���-Tk���Y��N������\��.�ۣ.y��ϣ����IJ^�|tDB�7Ҿ�\ͩm�Jh��j<D ���~���)<�u�y)J]��w��PB\����hy)J~�sx��5oV�5�oz┥'�w]���������o�R���~���R��}�7�B��BX��s<ۇ(��UOZ�<��/�~��┥�}ݏ$?"�d�������)I�k�<��:e�{�-e�4om��7�)(�d?}��JR�����┥'�~��%	���� �A��ԩ�7�Y������%)N�]�qJR��?�1������R������┥'����,�A�%��W+f��PU*&G-�#jq�KEH��{����n��t��t����\�#��N���71ql��+���-i��e*�Tp`r�S�YUv�U	�t:/K�vr�P�ą��N�;Q�*�1ٴ/:��mrqn9z� �ز:�snKu����״��_��~�!�;�Skkl�����s�.��6�Y���5%��q�s\�K7ww�`!ͷc��l�!�TQV0ڛ����籜˩�d����@E��{�r�Һ�m�5�7���R������<��.�����)I���q? ^JR��k��┥�#���a�~4F��ַ��)}߻o�R��{�w�����{�R�������O�C����~ժ�3v�i��7�|R����߶���>���Г|��l{x� ����E�ږ�T�����~��W�����`��Xr���_�:�nhEܹ�v��f��K����W�����7gu�lg�:Ћ�{U�n3��G#��<� m��C�N̼#ۋ����{����<=�*�?���y�6�����wM��e�P9�I��Uꊰ�ڶ�HQ�K;���}�6��U��
���~��_�S�RM���-�mz}�}~&�k�-�T�P���ĥS�������<͛O����[�/�$�|Ɇ28�ޤ�=]���V���^�{��6�0K�[֕e�q��@��IKe��2�{uhɈϿ-�BkZOF?����ߞ�k�h.���I����[��7A553S�����M���l�x��3f�l��GX�4"hi���`y�t��iVLRV�JTD%�"�=ߞ��ߞ�{*X�&/Ƀq�)��$�v�V��;^�͇��NW�ߦ�����!�t�
UQN��3kK�D>���}�6��U���h��2^5zL�Y�����9in\s���z�z�z^<6�d�q�0Nd�"S�ܚ��`y���ni\�_03{����'�@�	���4WZ��ؐ_������ڿ�	/�D�w�7-~����\��~��X�6�����<��l�5�6��&&��aВM��U���������X�ItDDK߯��o�?���[%���*���^�u�M��^�������-�f .{lbv�pS��b��{p��n�����Nݝt�/��wr|o}��W�c�)��c����niV<͞�����l���7U@�Bf������ү�P�1�����l������!$��ˎ��*hj�)U)��V>��`c�ٳ��
)��~� ���Ձ�5�Ω���R�T���IB����`c�����٠{��,ieQ9�#���vlP�=��_ wwU��;����wu��g��X�4]��rL��v��Å�ҍ�ݺpu(Zt�A������ۉl�s튭�m�Sӌ��#��y�#&��`�=�r m�J�[4R��Mg��؊ ����ճ Q��'T�Hؙ�r�2�I�p��3O; J�g:]�3�����Lq�:��Y�3r��M��7nH��T ��Ƈu�ٵ��j��S%�tA��͵.�'�n~���=����H)a7��K��+����.2��v�uq�n�*n�yn�������}[��0'u۝D����w�V��Vl�P�a�{�{�������8�4�lߒ�ٽ=��|ß~�6����75����\�M�UNj�z{���7f��l��u`��`{���ꠚrMS��P���M�no:�n�XBQ�#1����Z�ϒ���x�rF��@;ٮ�Q�;��3���{�6a�~?e�ѣu��b�(��P�)۩S[#���_1�v4l��9wO Z�*]=]UX�;d�˒�S������	��c��˪��St���*j�l�p(�����0p'6$�&�hGH� �!	�8�Ʉ��'
"?(������M�vw�V�ݫ��5<��d��jT����zl=����!%�BJ&N�ߪ�������Zm�L2Dۏ@;ުh�,l��
NwM���D�EIN�d��US�������uw?�ǝ�@;ުhz�Q�	����7�����j����������� �y��V&����M�f��Ȉ6����������`fl�������Z�7y3��MC��/2�[%�oK��F�]%�ߒ�?~_���i4D���u56�������w�-�)��	��y��ӄAJL$�B�V1���O���r�1Omq ޼�z��&�al��P�b�	A�k�l5�8�Rp4��g���[��t�Ź�>4	�J]��8�<P6���}͞�P�ݏ��F4_k*
i<&>HBbJ��t:�/�x�����t��� � �:�(!�W����'��3��\���w%�4�����1�������U~��+�����Vv\�F̑LhRd�f�˭z��z綹�w�w4�r�DM�&�lY"Ib��� �-K�a{6�Epk�]�c$Ľ��tN���|���kd�c�9�z��= ��s@�n�С|Þ�M�fkgT��SERS�����M��hu�@�mz���ڍ�?��M�k�*�^��o�wM�vo:��z��n���2��O ;ﾚ]k����g���u�@����(�� �'#�*�^�}�Z�*�^�WZ�nPL߇U�D.mr\ U���5,h��n�h�f�uʃc�����NݍqB?m��+Z]k�/;V�U��T��cqD�#�ȴ
��@��ZVנy�-��q��H�4)1'��T����)���*�V"��~�8�����@���h]�@��z��bQ�D�H�q�^�- �٠Uֽ�k�4�_~����Cl[Ck�sC@N�t���!u2�a��j�:Q�떌�/NU4Y{3��2��q��y��ލ��v�洬N�Yv��j��_V���]\~R� Y��,��9"[4hk5mU+���<#���/8yx�r(n.{.���ܾ2O1�ۨ�]�N���y2�ˑ�5�-$	;&�4ˍ�0OF����A�����d7Nh)K�QR��r�q
*�c�k���g��n����̥��R�s����V�H�enu����Y�A�Zh���}4
�נUz���Š�Y��1MȈBI< ����*�^���b�/Y�^�"������&��ٳ`}�[N��&�v�X��l�8��0DD��z��Ǡ^�@�[^��ޯ@/V�I�$�@�^�@�[^��ޯ@�wY4=��$�Ȣ����fk9�y�N�����n�r	�I��^\��R㬼s�$���)"r=�mz/z� ����<A������ϾM����<p�G�r���8���JrI�?�<A�}��˯��=Vנz��"�Fi��y�\�<W���ٟ�._}��*���<�pij��J!�p�G4>\�)��wM���t�ә�VmGГ������<��|���u�4���:�1W�`�����m��9�`���!]	p+8P8L���N'u:�3�%mMۧ,LsB*G.j��c�����uM�ff�|�wM�ڸ9���F4�n=�[�@=�@=���m{�$|�O쑵$����۽V�ݫ)@�!(��TG\���lW��ge��@$SI̍ɠ�ڰ>~͛n����=�6���.A�A4��L�U��ٳ`rI-��S�7��� �&0=}�t�*��v!e�j2�ބ�ݤ����Q;I�͝�ϛ��Բ&7�#��@6�q��nM�͵`�������ޛݼ�n�T��9b�	�U`o�m_(��l3����u��u�4ڋ	?���#8��_��`k�l��!(I�3yU�ݽj��,�L�D�
��sNÔ$�}=�6��U`n�ڰQ�?f́ݜ]rL�Q&���=�@��~P���_��`k�ٰ7�k�s"���"�֣��P�xy�.�h[��:�<>���v8.6cT������|*NJ��Xn[o�����������ݾ����XUR���UU`}��w��~�IL��~�6���lsv��$�~ID���?&K���R�:�v����=��N�7wj���j��V�H�q �iǡ�b��[��guXzw]���
Ww�?�����b����2'1h�j�?�/ew?���`{Ӛ���!��
<�߿ -!��dK���kYາi��q؊R�A�*���sEn4à�&U�'������qZP�"ʯZv-H5j����t/3�8O�����l�-T:/R+\ru���U�ѓ;�݃��N�(�k�)1�v%���u�9�E݅�趄8�sq`��m�ݠu�Ãct�ؗ][Qg��@E#�Ɖ��ie��%���n]j�����w��&�}��}oprպ��;��)&��+�m��Ƶk����������{�?|o�_�����R�����r�@����ym��n�mӖ�J��sN���ٿ�ٙ;���z��;��!$�=�Nm=M!dD��H�]~Ǡ޳@��j�9{k��{�	6�&HE ��aДCy��`y�t�~ݛ����e�����~Y��kq(��<S��6�K`uoElvL`{�*�[�Z�R6����p�s��Kjɝ���nz��&���f*����}����ӵ�T�<��T���_�/�/Hg���@?��/�d� M��^�Ǯ!A�J"?nՁ��`y�vo�l������$D��#���女�}U��ǝ�`nN�v��S������SU35_��z�>ޛ}9��~J_���h�?��	�BA!�h��lСvV� ooU�����7��v{x��Kr����g�7Gm�q�/x��q�]�^|Y����x{�a~�8��	�@~럕0�1�7����^޸�����s�[�oىs�-�wM�����l狓�����ji�UVgu��f�K�@!�`&�B�	 LJ��B���#5�vJW�k���[��;��$P���J�����|������f�}�M ����UBh�s5S`k�l��w��;,��*�נ_t���X`�D�N��%�g�:���!Sp�	�,Id�ۮ��7}����b#����a~ }o�@����W�� ���o#��ۛ#1c��5_ٵ��DB�2s�ߦ����M�^�4�.-�Fb�Ȣhn^��~͛:(l�ޫ�k��X�0��Щ�S-�T�tB��NoM�v�U��~�nWP2�9�p�XP����5�� �ֻ$hm<x� �zV���6��K�(���~�m��߿O�6��J�����Q��x�x	LBh1
+gIӞ�)i��a�j���976�v�;���y��@q�7'�$��*Z�J�k�Ē�U��P�_L����_|�z�z���I�M��9ԒU�_�}��~�����Z�O����ͷ�U���	DD̶��\�Ss���܏�K�'�jI+���x��1����$�����Ē��q�G����2'Ԓ^޾g�$��*Z�K���<ItOV�K��o�S'���f&����$�����$/��<I*�Q�^�������W��i,I�w�	]������4�h����*P��E�!8}�f�jк��h�!$r"v_��!�с�H^��i��$��2P�`��XFCN:h�%���%&h�	!�^w_o3-k[�m�� KCQ	k`�` -�l koB�ӛ�y� �qc>K�ge8�AT���V0��D�z��`2�4�'��[t�4l�0.�Z%�'��l���g�װcv�/c3c7^�ٱ;p����ݫ�����ۅ��n��w�v�6���ێ��	�ضG-m�ӮWt������Vۜ�dw�<��=���i��0�[�ֆ7Z�G PV�U�d2TpO$�쭙wXK���-�J��SZ6ٺL� 6�m�����UAg�"�rnE��u�[+8A�p%�����8�����f S!\�vj�����Z�֛l�ԛm�#��6�ڪ�Z�}+J���$��m��I��-�6ͭ� 6�6��vݻoN�ȶ�p[�mC��ݭ�c�J^U&�R��s�ܮP A�j�/*Y���uqXm5�vWZ˱�(J�R�T	J�� m�i	l[@֪�U6+�j�kv�x�:-[���6!Q� [@��ֺ6�m��u�K�yە�DWUOm�-�v�-+��/���n��6�H�oG.��� ��6�e4l�;l��Tr�N2l�`H�]ҳ-���);,!l3���ݍm�ts�m�W\���Q�n4�U#T���N2=��=�E�c�,��8^bۄ�tu:pl,K��Ekt��m<���1ۇ�p�V���Y��\�m�g��Qp��'��.��:*C��fm��5�Gٜ�쫌�i������ٞ5�mл<(tEM���.�:qJZ�����ȉM^��ն;m9�H d�cq����]�ƚ��G�f��n�*v�@<����Օ�ٺ�⍜S&ͷkv-����N�" i�ݴGl:�W���\pf�[Ds��R��S��<�,8t[��S9B��u1���؀�и�vm.�e(����]����'VMS�u�,ݰSk÷6�ٕ^S#�!��-�d	�L�m��ڞ
n��wK�ݽ�H�����O�4,��x'���/��R	T4/�w������M��.�Dh�V��k4l�&�lNǳ����r�8�<����mA:'VҾ�rݥ�<�/1��(�A������l����G]��q�Ͷ������v�̽��6nT�Jp��r�U:#��%�8�y�p��xT�lɹ�7a"����S��=h7X��Zgc�&܄�{qr�6�f`�O���tƚq���ҧk���n}�}��/�JokFR��60��Z;W����'a�WF�p'nκf�y�֓Y���#	�&/I|����IWҵ�$�����%y�-I%r�IT~Y#q�#�Ē��kRI{�_3�orvӶ�O�g￡B�T�w:_����Ǎ�	Ƶ$�����<�$�;��$�}���I+�ũ$�����r�8�H�y�K�Y���$��ߟ�$�}+Z�J�o��%�k��bȆ�P�jI*���ĒW��RI_m�<�$��(� ?;������-n�7f���0	L�V�i�6f�N밻��-��cl�;/ju�LM���$�}+Z�J�o��%�9E�B_L��wz~������UJ���M"8֤����y癏����(�$����<I/_J֤�V�6�?\B	0ng���W>�����<I/_J֤����y�I^�5A���$H�$�}���Iz�V�$���3�K�r�RIy��*���"$n6�~x�Kޖ-J�o��$��������<I/x)-q�:;]e6sL(5׆5m[mW]��	sλ<�u�s�r��R�r��'������x�^�Z�J����Iz�V�$�yy,Y9p$ss<�$��(��?fcl_?��|I.v|=I
�o��$�1��BU��m�1IԒK��y�Iz�V�g �P���M�ow�xy�fg�o�| ����ȷ�ҍ_����ZԒ]z��x�^�Z��w���Ē�}�34$�x��dR#RIu��y����ԒK�Y�KޗQ�$��
5�T_���3񱛁�T�Ԉ�v��ڵ�vU�l��(��j�L���W�cj�n�J�'�Z�Iu�<�$��u�J޾g�$��] ��H<�D�$����Ē���jI.�|�<I/zJ����/!e~&�dD��9'�$����RIu���Ē���jI%���$���q���T�U%���!%3����ͷ�5ö�o��������7�_�4IGtmD�E���C ۲�� �Z��us1%��R�C$	Ĥ�<I/y�-I$��<�$�}u��K��g�$���5y9�@wH�\���X���dJ^�;[Fc�����ڐ7�\<`�jʅ�X�I%���%��ԒV��<�$��(�$%�C)�Ǆr9�$�����Jf[���}��DL�mW7m��=�?|�z�J�ǁJbFL�Lz�K����%�IRԒ^;k�Ē�u�z�I{ݍ����Ȓ	��}I.�|���^[g�$�����#����QbX � �y2�I1����F���L��{����o���D2ڳX��5Bi�=�Ɩ�j�/k�ؘM�*u1U�-��g\B۞�r�5�N�X�E�g���Aܯ��DA�J�p�4U^z��n�N�NW�Ex�2;��p,��ۮ�H��<wg�O��ݦ2��i`F���N��5�_��鳋j��%�иo\�	I��v|����9�ج�M��B�gn�ݧ-�Gm�/绯��H�0M�f��<�C�ƊX̜���CN\���*6z��y}F9a8�Ա~�����0;�i���6I�P�U.�&'�A�h��hz�� ��4=빠z��*�H9�I���J`�c'�UoLX�0=F�G&�Cm!����M�zS@�n�篪��.8B2!LxHԒhwH0$����S �&0:C
�]����m������B]��6�������krm�ηf�x,n&FLBF<q�@����}V�[l�<������_d�ⲷ�k5�ʽ��9 �i�5]�����V���	&�}�zH�mf�/)�~��coF��i�6�;�ٷ-5I�9�UUXtC���X���o�0�1��\�"�1Z������L�`M���7���w4oQh�S$kӘ�Q�Mf�勭m�%�1��u�ϒ�����T��(�k˪X�#����^�M �l�/��hm��=G����d�m��'!�m��Bl�޵`owZ�72��I&�w��D%�	rM�������<~��CC@B�3 �!�%C II	 �C`��~���r���~ށyܮ6aQ���L�/�w4̭,}�V�;�V��N�_��[�@�M����}�4�����01W�İQ>�q$h<�K!T-�+�s��	8ms�ڳ������b�,��Va��?coF�ti�{�4?wa���Y1H�C�h�wH�wd�c��\We�̂Ɏ8����������n���l6I4H�%&h�[�_w��*��V�Q��(q!2"S;�j��<��'��eL�t�s�L`M��΍0'vA��Ï�M�xҶ�g�3��6{Q-=q皻�a�=^rs��6�.�盨�]��&�`M��΍0'vA�{�����ڌČh�f��u��/t��{���`$X~����W�wx���`�1�7�L�0:�bҘ�I��U:����3���X��Z`n�i�7�O�_�
̰�XU�Vf0&�i��wO�^�L�0l���Y�z{�=:{����v�h�ͼ-7��&��f�7\u�`2����틎u��m�5M���#�&�b����4aHp>�kUJ�j�Yٶ�]�o�[�T�ف]�v�P�F���)�I�^"};<��n̦+Ͷ7& u���<<�%��5��<䳷�ݘ�d]�Et���8�ݔ8���۱q���N���qڬnl�h-i��/H	�R�S ��P4QUI�!(K�{���g����b����\��u�V,�Z�qܫq[u˞�7	w/�ι����]u�+���Lލ0&�A�{d�ޠ�������܍�M��8F�hz�������V�zՁ�fڿɳ��� gF�&�Q9"�{女��h��s@�{���z�4�b�M�wmX�m��ٳaВo3��t�MU��30�t,��vF�[��������# �\J�U���'�V��N�dtg�3�qcsq\\N�)F�|}���?��y5�bq&�z���{l�<��4}빠r��b��#S{�Uy�{�
�R!QP��I~J.���,ou���`}�/K��x��aWFfc{��g�o�=��3;�����4�BtTe��ݑ����&0��U�?���������#�nf��;V��ē�������mX�f.l.WU���ut���q� ��Ku;K��ǫۭ"n[�a*�;��Żq�ԠCQ��$����d�4��\��4$����DLC"�I�{�)�fbGw�nh���@=�٠y_&�1@P&4d����j��'uّ
�@bhc�[P]f�A��g��x�c�'�@6���]DȀI���	P��P	�D`I�C\��y�$0I0�!0A0��2������3JL�$7���8�o��؛��
�<p�ݏ��W����
J�"$Eщ�.���|��K���lrC�F�pB�I�h��7�H�#6"4*��Bp�@�&R �e�d��QqQ>D�P�P@����|�I}����{��ݙ�'���%]�19��i|�	�W���3;����S@��w4
�;,F6Ȇc��fS ݓݐ`n���rSK�~b�����M�ڮn�� kc�-Bn9eOO`�9}{B�Ǜ�.o�7�nݘSU}�{��`{�J`�c܉�6UP�
iMPꝁ�nھI(l��s���=�����^pӓ�jiT��љx�/��`�1��})��Ѧ�ظTF�m%�-�����]����~�W��H,�,/���o//�@��~�Ҳb�h0n=޾������rSղ[b���}�r�=xR��1����'틢�(�����i,�{]����>�O�űmrn���?4��\���l��޾��6I��uv�j�:*f��y�t���<�6w����m_�B��z�R�n��������f�X��v~M�7�X}�6��VƱd�6�RM��Z��i��[ �����Y�V+�y�fS�Ѧ�Il��ݐaxx��p�	�R�
A��w�{�{��ߏ�'f������E�(��V2���!���#����%�3�2��\:uN���܎^f�L�%u�]SYT�Rգ[��p�p+�\����j��gG���.R)��ڴ�\�Bn�ᣆ�.��xu^q�:����ƞ���)�h�z�h�ɸ�ٵ�u��y݅۴�u�vC۶�r����1�I��1��{��<��x�*��A���{��;w���=��8��m�8�d-�ZZݲ�M�ў�V����$Y��K�H��;Y���'򻥰l�����i��9R�
�5i()"�=�4Ϫ�=���}v���eM+&)�& '&�;�ލ0%l��7d��ʑ]�嬥t,Yw�vF��K`���Jh�o�������F�x��߭�nɌ	ݐ`n��˦M�l.秶�S.�uv�g���j;px�;q��:�^��m�[�#S���nՁ�����n������`{�/e��N�SS2ʪ�s+K�q"PB;\0�P�۽���ʯ��wʭޘ����n��2�W��
̦�0I1�nɌ��L�Du�1�q�G3C��|��女�>�@��w4ظ��Q6%�= �ޘ�޾�������[�r���RW�nɫV1�c6\D�(�-�W��.U:�ܶ.8��q�v�S��v��m��_J`n����[ ݓ�WC

̰�v,YW��ݑ��왠{Ϫ�z���l�COpD��� l����2���+���Lލ0'Y�H�d�#�I�{�h��;��y���pj��b���T���v脷7�_��`|�6lhtO
I���!""�����A�p����q�j����lb���:mкۛG9���@�z�h.��+����
�d�&8�s4Z�������]��jEbQ�#�<Vנw>�O����+oۚ����=���e���``�z��ܫ߾�U}�{�W��`T�	�;ؙH�`K�C��2LRSJ1J*��a�@�QC�����B�Su	�̀��H�C3Lp��$FaP�|�Vt�8���Hi�U4X��V茝ޟ�=��`}�ZX�B����X�z���A��w���n���۴�ю���f��Nyb�L$ �$�?�fj3S�1AG3������`�1���F��p+��d�1�br- �z�β�����>�}��#ۃ��$� m�<�(��v,ս��7d��T��ej��y�^N�06���=�1��e4
�\E�H���9������0;�A�����K��H�B"D$�y�H���MU����4����:���\�]��Y�ێǰ7nx��nmû=�����^:q�����7���F�g���^�Z 6�%W6mL��aUmO;dn­F��[4l�u<����˱��.��T��d���N�@�X8n9'�m�鳺���{t�f��׷�2J�[.���9I��x6;	�vBmͱv�Z�M[�(v�N��{.d��ɰ��qm���
��� �sl7G�U����+ێnqp���3j˂YW��oL`wL�w�L���֨YO��rh���=�����^�^�4�R����.�`M���IlwL`oL� �۪J:�S�C(u4�興M���V�O�����`NWԋ%#,Ibdi�4��hzS@��s@:��{��:�DH��9Y&1@��;uR�f�9��<،�z�¢�=B�<���%�O���rhzS@�n�u�4��@����b�A�!�)�����%��t�wL`t����@��&�"qG3@:���h_U�u�s@���La&Lo��&�t�/�0:H��ʺ�K`t�B�)&28�)$�=�)�{��h{�6�ͫ�"�K�2Kt��;�4��c8���]r�g8|^�e{\7g�3��ηX�p��Q0D"������{��nh���7�c�d�u�&�3*��73�9}��@=�f��e4����>YS�C`�ۏ@=�����r�j@Ci*��Ё�"K���V��4�ڝ-��D��s/-
�R�5V�I�u�`f�Z�1����l�/a��M���rH�{��h|����}~���h[E��\������6d"�����&�M{�����v��8�qu����&�&����K`:c��0;di��"�.�R�L�ꉚ� ����BI$ٽ�Ł��j�37j��l햵��UEJu5Tw���߳��푦�L`�c���X�#�?�4�{�׽�*����*1a(z��2��BQ	��ŀfw9���WeL�j�*����~i�nɌ�`n������"�$bX���Dh1�dZ� B�-�U��ϳ��k�I�:q�m�i�˵��RR�3��f֖��k���=�z�>"x�Qa�����?�~ߏ �޵`y���{v��l����j��ԕTX�֬<ݛ?$ٙ�V_�Ɓ˂�*M�b"n73C����?~�;��`oL�gF���E?!�ĦF���f��YM�Nܫ����*�G�e��b�|�n�n�0�,<L`�|~��Lq �Ă,�#���)������H"��2ċ0��Fh�S��``n�L1=<w�Iݰ|��3�8����xl�<8S��D�Gg���V��h�##>��ۨ����r�0Df0^��zux?|����9�~0�Kp���O��Y�bOE�D����f�ic,5̍�����Q�Ƶ��`�c!5� �6��W[X�# ���$�=|C�sD;8D�LJ>�x��ߧ���*�]�VL��km�  -�6m�h0�yq�2�+;u�n�or�f�e'��P5
2�I���)P�&�`ذm���W`�t�\m�u��̈́H�QƮe8�N�ʔ[���;u�t �Ǳ�8��9RՎưq�WV�v��[&����V:�5�O[i�\z�w, Wm��m��h�]o=�Q�k���d�􂨩�l�Ʃ��mۖ�ւ�ce��i����e�-UP�\�++J��( ��]l���^ս\��Pk��wT���n�W�����D�r��djYN���p�g==UK�J�"KP�UT��ٵ��x2 �����Z�j��e�]��m�l����V5��`�Vݖ��W4�mN��E��v��/R[���j�jPYV�#a�궥خ ,j��Ƹi̬��*�UUU*쀲ʪ��R�<Ԫ�R�UP�+U+&iv�� [rj��7j68ʛ.٪ v�� m�<sm�5��.� ���j�,�ٻdq��y#Q����C���2+��m:6��k�mc�f�t�it�uQlY�µA�l� ���`'$.˵P���u��-��.�t�zن��D��N�c�.�M���{e��ܜ#؈\t7mp��C:�l/uau1�w3=���uaL��m�.�O� t�������H[m�k�zU���7g!Ϋa��$.g8�e��"0˹����R�]ut�s��,(�;q��C�M��u�b)�I7d�v-��!�[�K��i5���vh[m��l�V@ͬ��V���]�H T�-�y��B�Y	vz�]�����lnQ�Ks��x,���1�s�.��mN�#<[���ea;t���,A��g�:\�r�Uۋ+jB��N�tL�ے���,qXE��^w�ny��-�ʃƣ����rX�����Z��v�wfmʵ���J`=��;����Nc���{Sf[�� ������AO�=����҇«�@<D��x=��~���ӻ���ߛ�̑��Z��T���g:��ڳ�Ԥ����b�Pm�BVE���U�Y��6�\�lY6��K�m,�l��qL��F]�B�eSsm�-e�m�D]BS�P
���E�i���M�t�[RIˎ봋<���q�j���{yoS��x��rm��HU�%׋n'P�[a�.�6����͒cl�<e1�[C�X���]�}�{�G��P�$ѡF{8�*����k���jstz����λZ$���"^{:�nJ��hzS@�u������>�K�#�?�#p�:�����[ �� �=�U���&ٗ�$H���r�|��Y�{�S@�l���YL٦!�)U2�sSa�y�����?�`mt�����%e(�(�B�h�S@�m��=Vנ޳@��*q&� �&��ҏq"�l���t�7J�b�Wk��q͓l�*ļg�`蔉��ȴ�w4U��^���k��1��.�55D��s53J��$���i$}����`z����Ѧ���`����ĦF��9^�@�mz^��+k�=�"�'!�dr4D�z+k�:���9[^���z��ieȒ1���"n=ηs@�[ ���%�6D`+�+���b�{$�n��f�4:��v'� mfs\]r�iQ��`����weMSl�S4�_wM�{3j�͝��G�=�֬5l��P���&<iǠ�Y�r���n����8:Q21&6�$�9[^�}�xr�I�Gm�������y�h[f�n#%�h�4�c�h}����X��l�ݫy���kxϚ�d���z�נ�l�=Vנ{��T��+�)"������ԍI��b&��+v\ �۷u'廤�f��Y ����ĦF��}�h��Z�۹�z����!S!��D�%*�zw]�BM��֬y�6�ݫm��J,�T^|_خ�)���L���l��ݹ)�{�Q��l�y�ц]��]����1��2>I/}�I	$�}�ױ�&:E��j��Qw��;d���0'ti���-���U#` �~��L���"��:�'��@6#��{������i�ѓa
�ِ`l��kz[ � �d��Fۄnf�{���ޯ@/�����,�ehX�dk"��jIl�L`wH�gF�Eα&cr<��@-�4�w,��V�I��t��I�TP�IDIǠw[��^빠z��@��>�O������犤���C7Z�T���\�ʲ��g���H�n�)��r�ꐧex&^H�N�l�hUMV��i�[U�;4�Om�I�5��<�e��N��3u<e4+ʰZ6�8�4!���:�̀v��=�P,�3��:�����j�Fy8���7��)���c��Q'��5�u��#���GDIj���'Q�In`YP7<kTo׽�r�v~�r�q^N	6K�be�J�b��Т<�vTm�����S׌��Q�L�U^&���L�%�%N����͚�$���� ���=����w4z�o�$�)$`�I�cƤz����;��h���<Vנy�thuE�B��C@�s@���궽ޔ�-��7C��m�f`���L���vA����w��~�O��w$�#���!�J���Ѭ��V��ʇ\dú]˭ɳ�I�ee�b�]?[N�0=� ���LG�wǎF&%29�o]�<�`�`&�\N[����W��h�z���
2%$bhPSvdti���[N�06_&VE�E�17޻��ޯ@��Ll�0l�/�ŋu������:�~��`{fA�'F����y�ڍ�pv�m#��6x�#q�g�i��n����)a�:n�&�k���̶��`zvA�'F�[%�=�thuE�B�N`�4oJh���9{k�-�M��$����mEQ`n�ڰ1�vlk�
RB����ZIB�
I$WwU�wV���Tɑ�h�5&h���z�h^��-빠z�h�6$�X�Jdy���F���`I#L��l}��'�W�'7
�f;6h��I]vF�g����:��.x)�m��y:! i�Mx���`I#L��l	; ���*$Ĉ�Lm�@��������)�yψ�w%�Ɇ'�$�w��uw�����l�0$�� ��䟓q`�Lxԏ@�U�y�`{�4��}�ʒ[w����j�^PXVeU�VfS�2wF�[�����=�~lQ̍D�o$LPV4�ܺH�`c�܉GZ�㒍�Jl����hCv����������kz[v�W�K����V��pL�Q$��T�?Il��L�`{di�(�L(�WyJ�
�Yw��ݾ������#LW�^���q4	�1�q�N�0=�4��ޖ��ޖ���T]J3*�
�,��������z[kz=��s@�܂��9#���6cG�p�$�h1Q���� ��fpWH�
�c���9Zgv:�Y�Ł�P+�O�~����A�L�N�!��v��U���X�L�e�hU���4uϞ�h^���� ���c�g^����=��n]�.+.��=��F���q��x�S���PGk6��lE�w�=����y�{Y��:�RۏK��h�a�b��$���������K͝'������u�"�Ɠf!4p'���=�9�]�sP�?}�[�t:�Z翿����l�nm��K���V��*��&��R��M�癶�����#L��o��|��6)�C�LYRD�܏@�����[��r���=]���E54�mB73@푦V����lN�06�] �L�"�$���^���z���׮��{kZ�O�G$���c�T\U،䮭����v#3��x�6��]�m~��8�(%27���z���׮��ޯ@�貸������&��^w����@Ij�h�ެ���ʹ{���W�Tw%L)�jD��ѦV��T�l�`muv�����ݶ�&�|<��3f�ݑ��F���Ҽ�e"�Ef&�t��0=�4�ݑ���#�7�\,N���㞩�{Z���ם�1����T�y��o9�Jk=<k�-��ݑ��F��4�����9A�����������H�vF�]���4���T�UQx+V����`{۶�<͛%zi�!T(�%I8��5��V5d�N���@�-�;�4�XX`&���Ԑ��Lq ��b O�f�f� �+{v!�)�Ѡ��pdO]�
w\�> 8�mP;� |+�W�O�#��WY��o�*����*�/z\�N<�	LI��=]���e4ލ07di��|U�Yˣ*��*��`ñw�Lލ0=[%�7�Xq��E��ؔzCR;��n{C�.x����vzM�>Vu�SEi�볂����07z4��t����z�{�~��D�񛐚��<����y]%�=�4���� ���і,�U�h����t��ݑ��F��5�^�؈<CD��r=�ߗ���f����Õ{���ʃ��B���(N1"�ٰ7P-f��72�7����Ѧ�F����:4����o�hxʹ6cl�ll���7�����;�Ǯp��ۖq��u�N:��]ny��3�F���l��`{�4�����i'E�������;�,n��=�j�Jf��r�'U6S�2	����zl�6՜�I��}��ߦ�Q�2���P�&���4�푦��S��:�f�u2~���ª��nwZ��ڰ6�K`zti��B�������++32�q��T��}�9^����u��d���u�֖����Ӷ��=Zv���FMR�Q���ٹ�(�� 쬪�.���s`��
]S�g8%54��I�{��pN��n�X��&޵6]ٶC�.8��q�1�Er{I��Û)k�ຸ�]z��H�n�.�F�0n������ˍ�sZٌ�Z�ZWM��%n�
��wm�����wO�m�W��N�~��-tZ����ڂ�ɧv�˼�y պ�����$��pxG3�z�4U��/]��x���nhߏ���L�8ܒh��L	�`v�� �&0$Ar�bJc��E�^빠w��h�٠{_U�r�(cɌ`�,RL��$�{��+ ��ە����j��{�ƜyF6�h�٠w�~<�~��;޻��H&V�S<��Cf�+�YS�;m�浺!�U����%���$q����`�rh^��/u��3ٶ�B��}�6>�9̓RMH"�sE��ݵz���Q
<���E�}�� �~���4�˂��z�Ȫ���noZ��6��oݵŁ��j�=��6��BsD��+P�K�����������F��`z.��,)�fU嗙�N�0;di��Ѧ��4���l�I$.�C]��{4�n.P�����ɶ�䉸�����D��$��$��_�ۚ{n�u�4oJh�JF�cK�drf��ݵ���6k��3���7wm_D$����uIr�@�f��ϻ����o�/�̒�MJCA|	���S	Q0D�7 H�I���j��oZ�32���%�)��SSSa�?v�ou�=�j���^�W��0��Bh�8h�w�4���-����w�����yʭ�(�`v3I��r\��ʕA��PM�5�T�獀.��)�?�B�������0�1����`�.�u4�c�)�Xf�_舅��,��V{6��DBl�[��Y(�UN�������Ld��ݑ��&0-�u*�&ƚMȴ>�ľ�礪���Õ]�{�W��%c䱂�E�$�T�M���@��U2�3�4�$��%0	$����;|�]�E���J'fv��
-�V�:$�۵��㌷t��JjՅQ���+���$��%0	$��0:��"dȌ��M�]�@-��4�$��L��]��Tә���ڰ3۶�脡&��t��-��r�O�dkY��&���}j�כ�`{g5�~I$��� ��m�&5�!0�f�^�hw��� ��=�j���$F�4���	#����ݴ���CZ���6.��/G<L�n�#G��wkr5n�=�-힤y�nې�g��֠�<�:z��T	X�>X
C�n��B��b�Y-�VGl�3H1\+\����\��֞Ÿ�6�ٗ�{�9�����;p��0��N -yع�CnY�������lvam�n�Q�ny˩���[n��_��}�~���ݼk��f�li��f���w����w�";n:ۭ�L��S�u:�3�a̚��Ypn��h���m��=��\��lvn��i������X��_�Q�}�6r9�>��#rʧN����_DBM����}�6�s]���`�I�R�*")&�޻V�U����h�f�Q�i����#�hu�@���@=�@�]�@�zĒh��-Ve�06_J`�1��rS �I������O�9�h79j��XYֺMM���66�r�n�Nót�y�U.!3�8ȱ��{�f�޻V�y����h�+��O�n�ޢ	�'�w����<��}�mOK`zvA�ot����%�Pog�`���0r-�~���ՠ�Y�{]�@�,C�"s��3+K �fՁ����	?N�N���|�'�HM	�h��hl�盳`fei`tD%�k]/�4V�Y�3�q�WZ�d�0�ge���fԝ��ݔ�ɇt���N��FF�[o��O��ֽ��=���9��<RC�y��h.� ��g{��<�S@�z7����8��;� �7�c5%����ɞ[%�"��cj&���Y��{�f�岚��zw]���r�Cin��f���Ł�B�ӽ���\X�]�Ӯ��~$�D�b�DlɆ���y"l�t�h�ݴ����M����fH��uYx��0=[%�6vA��Ѧ{e4�cQ��L�9���oJX�m�=�������(�l�G5I��m!4H�p�;���;�)�x���ޔ�;�\��ɈX�4�4ِ`�1���?}��/�|��/',��@>��1<$��ȌnC@<����})���m�L	�+�e]ոa4�L��������y5$���:���3�]ۯ	�� �4�����=���=�,��K����}���n3E���}�M�v� ��f��}V��ҹ9���r#� �߿[ղ[e���d�J�-VU��y���l���#L��hu�@��0�ؐ�H���zN�07{ �$�V�l.��U�6��a}��c�	��0���0DWGffabAa��f!!�Rx���h4c���5����) x�h��0�"��H+oJ�xC l]�AQ%vv�A>�y0L�a�bl�Bl4�����f�'�ؐx� �	\H�
jH�i�� +�}�k��h��$�� Ѱ6�р  rm�m�
Bm�. r�>�fM����f⛮��(Pb��Q��]i�T�Ek�2*��(��(0�w7�����7\a�n�b� ��^�K6y����Wm��{I�Aɠ�[��^u�ˇ�ۘ���ܫ½;p\v,��%���.��N�����u�|v�ŋm�����x{%��v�v<�a"k}��~ڪ����V��D���;��0�R5�W�b�m��ڦ��M�m T�7g�� ��	vvUj�^G-���[�>�衷:\aӌ�ڦeQ�:��x��[g/[EȲJi�i��N.eZ��X�p�bG�m�m6݃Id�� I��[�J�h�tm� �� ְ[�.�\��d�K�R샢����줶�d��e��yeP<j��$mC����d��@܍2�UUT��J�UWJ�-uR��AKTe)Z�U��]Y4�\�@: �����U^�&� �`k5����X�j�l�T��z�j�����m�YoY�@��{Er��7;oK��M��M�tK�0�u� 	gVj�ޞ����Y66��[m�����Y�I:������9�n���Ε��u��T��3�<*��Z�d�a^���#����@p��9z��5e-��pݧ�C�旉�!���c%���Y7:�v�^^50 ��n�md���iA͍�i�s��L*Om��d��;�.m6��V�bB�������؁]2�h��&x�[+��+�4M�	��ZV8�:ȫT�i&icM�du�ñ���=�Cx�%z�qV��H��u�m��\bsJ,;'�;k����[$�g5�z���*J�p않L6�I)#��#�f�3W�򽬫��I���	�g'&�qwkmO+��
g�P�^���8yR��_mlgvV�ڼ��)�=��#���S��WzɊ����뻢�.�+�Ș��x�iz�mG�!�C`s�NmNy��?��0���l�I�Y9�@�D��c����׮�Weѹ�Y���!��I��j��j�r�J�8�ڰ�Wvj�h�q)p�����rc�P*�����q�ʽ��Si�:3��[I��!�B=�[�G 9z;6�u��׍"�Ss�Y�.�6�B�1�Fc��s/��/I�+>;m�بn�uې�ѫfl;���[�ۡc�+l7ow�=�{Y�<�Ae6�p���	�V���ۊL��k�����
�Λv\�!�M8P/�}����^��zS@���fLBɒI&h�1�+����`oti�$��_��c�Hb��I4U��[Қ�F��1��`�Ad��R�2̼���`n�i�I��L`u_ݖ'4�1�R9�z�h^�@<�٠u�M�zU��d���`���a�����������m���m�r���6֧��n�QL���S��^ ������^�ץ4}빠���8aS&���ʼ�]�s�4����x����ꯋw:Հ{sj�!��K��1�i�̫�w�l	���07z4�6t��mz�eYTA	�A���w4ۛVޝ�aТ"�w;g��1&F���޳@��j�;�j�=����mkT��xG$ps&�C�V�zѶ6�m������1�	���ŷ�+���D$�@��j�;�j�=���I(����`f�#PI�H&���������6foZ���>��Z��ul�r�'!�{�]� �ͫ;��(U^��v����̖�U8�	��dFk�g����<��hzS@��h��l#��E##�@�wK`w���~���6O�0�1�96�s�V8XQ�r�e+�ۛ�#Z�L��"Չ9�B�Y��Ÿ2ms���7.e�:vA���� ����l	*�k� ��4;����_��@����:�����QX����d�&Ӧ0=]��vA�����u�Ǆp�5	$�<��h����w�+�/<T_��w^w|��a�R&�Bd�-�Jh���+��z�Z�H�M�~��7m��H"WaP�6\j;���^wk���{>|��v��cq�)�nC&D�9 �޳@�z���@�Қ#���9�7f�5�rO ����������@�Y�^�@=�9�E0$��R=�}V�ە���!6{w�����`b�X�{�2dN&�z^��}�h�f���נ[��E�6�!4�m�N����-�ӲI|�������$gm;.ą�c,նܼ�
+�6�u�mrW=<s��hղ^v6� #;��ۃ��6�Uv���	B����Z�A�V��m�`�5���p,@�����#]�2��۪����$�]љ]�W����mh�v�=vٟn��6�u�R�r���&u�^^E�r����ەx�6@gY�v8�Ǵـ��WJl+͝��>�?�{�ww=[��g�©�m�ml��By{;O�Xn�7>����;��Y�Ȟ!�123��Ɯ��}��h��4��}�4��."I��EUU���ٿ�
!���� �� ��7��ؑՆ\C>�@ǉ�D��>���`�c ��[%����VPƜ�<RC@=�٠����â(O�������2�MYR]4)����?ckd�ے�����km�;��:�%&�C�k�}���Ie�H:���p�<�&��Pq���u�Q���������})�wt�7�0'���e`<&L���z��Z�g�H;�� ��h+k�/a�;bOCl����`�ڰ�mY�""���=__����yV6���,y0NM �z���[�:[ �t��޿���ʩ�EUU���ٰ9B��=�? {w��f��%[kXƿ(H$5��q�ʾƂ;n�ۚ����7kZ�xϳu�fy���m�Df,��1��ⶽ ������>�~�����H�&c��5�ld���0=�Ҙ����:�m�sE3b��x����}V؀|�P0��!i��FH �P$e��1C�����}�4Ֆ�L�?D<#��v�J`�1�M�?�U�?y0?q1_���L�#�h���}�4=빠__U�{��N$��A�0q�	n11�N��u����ܷq"��ܖ+�v�4�ɋ�$�I4��h�w4��I%��z�kgH�ujU&���nھI��w���w��73j���Ie�8`��Cs4�h^�@/u��w4h�m��cN��sSa�	B}=�6��V�m�.�|D�W�^~���k�^v��hO1��"�����-빠r�נUz���p�_#�hG�4��C�5�<Tv� j�Lv�[j���*�����'-L��h�tЦ���~�߭X��6׬�oY���\�����!�q0:�K`t���6t�l�?�J��}��hx��P�E�w}>4��h^����Zv:��lҕT杀o�j��͵`o�5�rJ!C���1�-�H�j$jU&���͵`M���&ɌoL`r>"�2��W*�m0�#a.6��jڠ:k�. D��㵐�X�W��b2%#�&�r�ӳ�n�����`�;���)A�4�j��z�:��c,M��k���`�"�7�ʎa���2�;@S��8(��w/VZz^�A�O.6!�-;����ڷn����}=��[�[Up����ێ[nnř�гpl��8�ٮ٦�4UK�'СE�E�.UU!a�v裍Ӵ�Q$�>,k��мfݭ��*<�5(�&,`L�E��m!����;���1�M��`t-u�]J3*�*�0��`�c ���`M��@:�\�9�m�&�_z��Ѧ�����	,�]*��l-�B����?4�����=�1�v��j�H�!?�2'3@�@=�c ��ލ0)l�ԫ˫�h:�N�0jX6+�����y���f�����8�ݶK��6�$�n�s�����O߿p}���ŀ:��`{�_Q,�˫�j��5V�ͫQ
=��	L���V��^�y�@�~�֘ħ�,y1'������$��&0�����Q#k������ڴ�l��@����:�"Ɣ��LP�32�l��;�cgF��%0=����C�gTn��a����Gk�'cm��nq9z����ڴ�vΠֺ���v^f0���Ѧ��L�L`\��q5>[����I�����v� ��hwY�Ֆ�X�H�8��L	; �:t�h��*�86z1�pc�v ��������3 (J)���}�v"8��z�,�Αӣ1`�22̐1����6��ɈNH|�a$��&B�&&9���)LWhvh֍�� �"
4��k,�H),
30pS13���	����%���������M�u�E�R��IN!�f�Ch����;�k�@XF)�$l}ُ�L~������I���ҚH}�_#�`�0���vb'��{��ۀ@���]�C�klL�l�D<^{q��x{$�,Ć&��$�}��� ��<X Be`	b!oz/��M���!�O\(�a�J D� 	�ka�3�+ʃ@�@>	�IBL��) �h�"��=DUC��lA���p:j@4 >�ZV�}Ez�h�@�����/^�`n�i�4�ڢ��ڬX��2���o�z��z���V�!�m�`}��|�Q��I��oY�[�s@��4޳@�r��jp�����9͕��^S[�	��8�4/kD���O�&�A a�?'������LIɠ_m��-���������z�3��9�N[��'3@��4^�zo+4/]��#�yZ_F��?L�"���
����T��F�nJ`"ʻ���9�@/�Y�ym��<�ե
�ҡ��*�Qr����U��Wu�"O麦	�b���=����y]�@��ٰ�V�Ifw|T��pUEL�v�mγ�F�6�d�O7����n;n+��b���b�,X�ŊE�GȜ� ����@�ޯ@3�mr��f��0��`�\�J�9�j���ٳ}�!Ca���`{;�XWj�=�I\4)#mŠwT���L	�%0=]��_r�KUK>���UWY�wF�nJ`z���/+4����D4���'3@��)����=:�0;z4�/���#������-��'SH�i�.1qn:�8������q�@C�����9��RĵQ.77g�X5��Z̐)R$�T�%�C,+M��.�*9\��٣�U;l㍉cN���¼n�����pm�r�3u��綴��ûu��t㈎뗍�3�$��ey����=�?W�wlb�b�5��;��ȍǷH�0&+j
�F�c���������}�Y2!�ڻ��ѶeާZǬ��c���1������I-�uס%�W�My\����=:�07z4��rS �qCJc�jG�^Vh��Sm�LV�l[g\U���˴U�YyY����m�L�&0N���r�,JG�����/�ՠt��=:^0����VAuj�fF��Z�[4��� �����m���o�=�3G�9��f�1�5F��Zm�;[i��ָyzn�0(�:pN��&RA�&�yz���Y�^v� ��1k6Sj�F�Rnjj�=��y%�|�U�YEKn��L`�/G����dB��nM�h���/+4��4�=�i51$��- �����f�w�f�}v��[~��D0i��� {�_M �z���Z��4�}n��B7�����N>�!a�m(;���s�����ۮ��'ZG�1�������=n)8�����/�ՠ޳@<����<�,JG������*�נ޳@<����Y�#���\�)�#b�= ��wʯ;�w|�=Dz'M*���7�>��>W�Z�"��M
H4��N��ލ0%l���l�����{*S�5*�r�{6Ձ�DB����W��^Vh:ֵI�#�)03�h3�d��Xq����ƶ��h6NxͷV-�$�(�(D�K�h�j�<W��N��ލ0"�G
�ŗt�c�r=�z� ��@�z�h{k��~o"4��Z��f���L	[%�;{ ��*��-��
�!]�fx�?4���[��S}�ƉZT"�(B`ء����sT|�����`�x��xG1�+d��d�T��0?�_.��{�m�C�c��\]n�s2Tr�F�n�ˮ^3۳D�<n�4�C��y�3�ll��uL����3:���Ձ�n����>��}�|�#�6���I!�^VX��_�f���k�JJl#c�����T��U`nwZ�7'5��ՠyY�UJ*�(D�Kt�9���3g��n=�ۻj�Գޯ����I�8��j�y\`l����l���E/�(R�X��m]ev��������;HU���/�=�q��v�켙�Omɸe���r��m9"���������ӕ*GK��]T�ݙ��1^��iX\��]��3AKe�T*�� �m��+.�9{�=��H�{@�ks��z�zᗳ��n�qt��}�}�|���<pN5��6��8'p����x�ٍGݼ�m����tR9��K�IdDD/�Q�3��~s%qBs�Җ�(-&F��q�m��{�_>V�Z$�.�u�GN�GS����O�`oH�e����L�u�Y�vݶ���O ��ۚ��Z����[�� ���)'��C�9�������6T��F��(�*��Yw��ї�v�S �*c�#L{�4�VDX6���G"�$&0=�4����ݾ���?~_������/�9vvôF�ŋvS��y���d/iݸg)N�ς��ѱ�\�����߿4����ݾ��=!1�+� ��I��S-�敁癳x�B�QJDBJaѻ=n�3��73mX��c��I1L��z��4�K4�]���^�^���8�1I ��ލ06���&�A��λ��ku�H��!'�}�����^�}�M �����m��#��@�nr����}	F�A�x�ڌ�s�!rX�֎ݒG�!�?�8��xm�hޔ�:�h{n��Sr4���Q���`n�A�{�1�푦�����wCM
H�q��K4�mY�p�%�'F��X��6 �<�&�&4&d�^����h�W�u,�<T��4���1������S �l���4��_/���I|���,ơ1�� � r6�j7[E�v���A�9�ڋ���7[Fg�n,�.
ݝ\���/���^Vh�� ��h��M㌁R8��+4�٠����Z��r�'�n�HЄ�I��}4Ϫ�=�ՠx�����Ɲ�����m)&�˺�^�́�Kݛ�Q�Ѕ�):���~7 <py�Qɠr���Kݛ �ͫ ��j���[�˜�s &������Է��юҲ��:���X;;�8�s���j�:��<���g�����~ ���L`uN��<.��D���	����f���u�h���@�{J�Z�@��Lm(ӓ@;ޘ���[հ��'I�T�K+H`�1��@�����@:�4��4��S�x� D�R=��6l�	Owuxw��Ǚ�`(P�*��"�*��
���
�"�*�Ҋ���"*���B*��� ��!�� Ģ�4� Ѐ"���3"�3
(*"���EPU��EPU��AW�����*�������*����
��"�*�Ȋ���B*����
���
������)����" �"/�8,�������_���02?  5*4�gR/��'��   ҃  w�z� [�>����ު�{���Q�U8֎A�Kܻ�ڭ�� Ͼ���m*��>��޲�-W��{ikoz�ʥ<s����ﾪ�{t��Z�[��-����k>v]�}s�y۴Ym�O}�� 3o�/m�-�����Ͷ��s׶{�қ��-)Y�ꪣ�O �ީU�U۞�S�#{�:RwwU�/��$    @��M �JR�z�'��i��ё�a��T�I       Ob�UOPi�hi�#C&A����EQ&��4h�     �H dM2	�<M'�����&�ژ��D����Q��  @��(t�=x˧z��8~�D�AU y��O�aAP�#��\���! ��@L�E�I�e���*���i1(�C����p?���?g��~�e�����I$�I$�'I$�I$�I$��5UI$�I$�I$�I$�I$�I$�(��KN�Ix` � �0��0g�{��$�I$�I$�I$�I$�I$�	$�I$�I$�I$�IwwWiBI%i$�I$�I$�I$�I$�-P�%	$���$�%i-��I$���J�P�I$�E$�KPI$�I�J�JRI*I)I:I$�$�Kt�I%���Y��<UL�R�J�I$���I$�I)I%I$�I$�$�V�I$�I%	$���I$�I)I%H$�I$�I%�:I)I%H$���J���hH#����N����P�UM�O����&)~�K>�g�Vr���N�8�8o�v��c�z٧���w.�Mw�M۸Wi
��4:��m�em����+,�`Y�5ӣ{��c&�C�/��n�����;w]�ީ�ٽޖn���e�FKeQ�s�3um���{e����ڸHI��D�f�o[��Ĉt6;�zMX�1:u2�j�R�m�i��a���ĭ6x]yؑXc ����9�RHfB�ʤ���V�nfx^�L,,!!
@H��21$H4#0,&F�+)5(�M�R�y}�6�V#�Yc~∉$7�AE�<aMƋcRBƂ���Q�f�[��FF!p����Ba
�A
�
єl�F��;É�5B���@"���3p�Ҙ��ù�F��%�8JaDJnH�(Ä֙5 �!\���6s�]q4�W��R�e�ԭ��*�9��doa�Č����a<x�{�x|#/K(��'2�K���s`@��Ϡ������|��-��$�ۻw&�8DξB�x�
�UpF/�*I�g�� ʺ$=s*nb0XΞVu�f�2'3��MiJ�'��zB�6��w&3b����Z�RļCUaD*ǁ�&��� �u@[�.IjZ�0�zԸb��%Κ�s"y3�6�.	�XMX1O��f$1s�XƎ+.F��X<!��b\�#ki4�9�o�y�Wl[[r>a�i����[is2�=9���k1-9���V��YFuS��ZmG�&��o�(ݜ�y�
�z��MU��sx�˙@��i|5��2�*ۄ/E�s����z�i�skq��H�rY�.]ی��.� �jI#M�i��cM�l�k{�DJl��8W�[�h\�ù�[����4�gB#Zb��ޫ(Ȫ��ǉ0�4��ʂM<.8ܙܜuu+ś6��*���%��Yy�0�s�&9�duUxg�ҧ*�$�d�
'���i�� ��Nq!�L5ƀЌ����F�lAp�z���g�����M�Gn�c���2�䍥�vʼc)�ٛ6i	3�{=��y��z�v]L�	t����7%X���s�z[�U�rK`���tz�5�ʻ=�E4L𻵰��:���:�O5�:�i��-��s�''a�h�G
�2�[��k����	�j榙�CY�b&�ч\��a
ݙ�VL���]�M�=����vUW�T�+�4)����IA�yvF�����U�cZ�g         W-ڗ��*�����5��ĥ��2m�.��jہ�9v��k/-��UJ�����$e-��S���;�h&�K����Z�;#���������,���\�׵��!qp�H��9��c!�Yw9`^�R=l�nƺ��m�`�,��[k�y�c��jjW�qӮ�m�1l]!/Wm��r�M�d��-v�<� qw���oN���C1ͮ�/d�Nm�{���fyV���\��rY�aB)���.��S�벫���Ʌ��g7';ٶ�v*�;m��Ee8w�ǀ��=�vtl�UUUUU�UUJ���EUU:%��r��kM��ݑ6n���q�π��u�m����F���eݓ9���W��j��{6�6h�P���JEj��������U].&ej�^���U t������h6 ���6��\C��]����
��Z�c�Y�xpn�+�ד���2�,�j̱�����	^v���٬b��,pKV��>=�V�y��,Ҩ ��z@�]iCS��J��UR�/Xí���ڪ���:	�`lJ��r�W5�C�x���gf�]K9S�Wj��9lQ�`8�-ƅa�u���q���]V������Ϥ��J�ײ��g�ZKP��.���Y�2���؝��̚ĎC�UU�U�U@U[UUU*�UmUT誥ZU��������V���
��٪������
����UP              @$�     *���j�������*��
�5UUW!f����U��Vꮦ�UR�X�bnk�k`)�u ��SR�Z\���^��S����lr��s) ʵUUUUmmUUUU�U*���J�UUUT5UUV�*����ڪ��j��j�������j���j(��h���c���9�C�N�b��z�OSۘ�����Fj�D�c=�n�Q-�vW/.��X9C�Y����p@ O�?�DQ�۠�:Ni���aÙ�=둦�RTcQE0E5APMQTDDEDQ5ME$QE4DEA�`�"*�`��������"��f(��cD1��	���0UDErc8�QPP�!�:R�! ��E�d&�f�Q��dRaY�}�ڨ�U��X�U���"�*"�*"��"�*"�*"�*"�**"����*"�*"�*"�*"�**���������������            
�����*���������������"��Q��X�U� �d�w 	��0 �djY��	��T�@�{^�4+G���i��.�B� ��#� xpׁ�V���K^,�h�3��jip�Д� qG&ӎ�A�	ށã����B� �)��>#������-�2 �<7
�<�����Z;�M���)��I��,bJO<ک��<�Qٷ^;q�(5|v���CA���f�j�)���Sg{�"-�&SZ8dO<_4GWȝ4:�bQ�A�M�U���i@!����@����<D.���W��-Ar�a��P�;E�UQUUT������1UUUUUUU*��������UUUU@��UUUUUUUUUUEUQUUUUX������������                        
������UUUUUU���0	?�C�,>��ww�~��wt�#wwv�%	��P����'����A*
�D;�HC.�Wz�`Ձ-��,!�lI������t��' ��S��FU��8�3�gW@�n��;ahQ�e5�de wu��6՗���Ɍ���Z,$!���q ��iq¸�rRH�q�l����uJ:��� :���V9���v]�$K(�;7.՜N��]��λCn�sW�h�Ma.�i�kIi��T)�������v��eP� ���Ѻ��pv��l�q��mLu�C��w����t*)
��$���3�Tx;��c��tS�� ����"k<����!N�y���f;d�k�-��6zڎ�\Ԩ��8"�3=q�w����M,!%��UYlr;d�K���o>��(���}�!�fN���T��i��\��*m����	�YV�E7�59�����d@f��������G��Q|��̤}�گU+]�T��7�)�[�=�\,�ݢ�1���5�0��zs�5�:�8�f�u�<��J�݁e���%������=�\�y�E��2h��bޭ��0p��t�p��4��EA��u*+���m�)��Y�z�Ѧ@�ziU(�E��O4!	��(K4.��6rmU�/ �N|�8@�j�f�Bg.���� ��ز�RA�K	4�/{kz���t�vkT~�{�����๜�o����:n��L��@��9�P������
'��F�7�FY���V_"�Ƴ �uN�ZYKV�^������#�DDrв�>i�&a�F���uQ5s2z�>;3w���)h�B�^�Y��4�DO4�.�Em��u`=;YV0yt��u��]�;X�Em$��r�[�v���Ғ��Rt�Fs�Q���Y5��Ia{��ì�����vx�n7S� ��ӣR�w3���q�fc$�y��	Sr��B�|�ns��Jت� fʹ�o�X;P4"�`^�6.�/^d�("Ь��N�c�fyN�Xxf�كD�*�A�����<������N�:G� ЊE(.���.��-�s�g?��fr��www(���ww}ݜ�tDwu�Y���Ҁ`���;� ڟ� W��FO����U}����U���en���z��6xp)8�UOB/�����/���-��@�����q=���W�p����KǬT>�5�ko�@��os��=��1��6�=3�Er*YS���H�� ���gx������Ǻ��e�7�j��_	�v4[q�e��x#����z���7��~&�bO��l�[y�_� ^��=�����:�)�R:t�Ɩ8�ޮ��k?��~�Px��}�!ɲm�ok��ǅv<�{�뮸ǰȅ� y�NN3�`��䌆�~��ܽW�t�
�ygf�Y�����M�B-3��턍��j�U<UXܾ�}���W{�.��3,��]�8���t���~��v'�5�P@�ƶb�X��"&⊽�OzV��S�)QW�?@��E]o{�����b���;�"*;����>�J㲃�K�ax.>��.0�ĜŒČ� �)�@�J�3��Y�Z��ߏӠ�d�j�J���Mj�K��E�m��cV�:cX�Vh�eN��3w��ľ��h�����"�bD�`#��Kq�+���\Tiz��x�S��Ic����1��}Ц"�e�	g��O}�X>���o@�,Fs|�w>�=�ͣ�[�m�&��oYi�)�H�W�����y���~<m(�x�����ڕ�i�i�c�K>'�����;�>K m�	��K��Sv?�W����h�1975�FCG�?�������۴^(|:����;��ns�"''��>̓��m�����5���e���I�f�Yu�]��c�#&�&E����_�.{8���	Bf�M�3 0�a^���\�a��x�����ͱ[J���D���fj�[�g��y��FCc�7����H�������Oߍ!��ʩ�u���ь�ֿ݆��ɖ�C31C2�İ�H��J�o��O�W5t�����X�W�X 6�q&��5|�{��s���2��KE4�1˭�U��3.s5��>���[��_8��{�,HL�∠����G?x`�[�D�����(VPn�JT���9�Q�-,%�k>��5��PL+x�Ʒ����%�;��Ooə���ﻻ�DGw]������WDG{�����~��{�S��� z;��O熷>h��e����á�E bk���O!��Sʲ�5��
U���HJ<+Q��v�5U�C�F�̃h!��SvӺt�ss3�V�,�3�3�u��{N4��Ly{u����XB�홵F��nt�Fs��v��9n�-�f.�e��=ȇj
��m��A�ʀ��5������p�g����r��b���m����6M�+U@UP@�R���!;]��b��l7Q2,
�.�l�[PQ?�c�'4�/.B�eܫ�?9?�L�����0@�b�_R�bD�'[��М��C���Tn�h�Wq�6��&8�o�ىLQ��v�ls]�ݾ���F���쵕A�lT�����X��g�e�h\�Ľ
�C�����~X����r�f	�5Y�7Aΐ�x"t�݀.�78>uZ��R�P;�󫇗}5����e#�(�`Z!�3�f����y�3��'+���56�g����p�C�y��e#Ò�e^��k*�Y����!����;��������S�o[�#!��q���!vP���<���j0/�?[�⥤!$,W/1�7o{K��"h�=�X3�0uU, c3�>����$|���`5���C�^	�/�WFL��L�����M�U$$��d絶��;�{έo}���&߬q�h+ A��Kx�1��'��\�1�QmEH�
팆�q!�s��L6P����%9vm�'c�����v�WR�N�b3��������;���5�"v>��R��7  �P�"��& �'"�xE,�K��m�rQ�T[k��	bD�[�� >ޫ�t������g�=W��0���	�+���������� �A��y�Ś �v=�r ��|U�#�S	b�%����|��[XJ:���"D��X�'�5r+�P5ț�y9���	"���$mG��"9H?��)_b�@�* v � ����{PDD;t����֙]َ.�kGhwGqS�dr �=���E�N@I�A�����@rDND�}�_^ �&�&�nB�?�$l��l�ڬ����u".��<%�����Y2�Ye�����)ؔ��L�>OvQ� � �y�7H>�~�4��A�A�Dמ�u`���Jq�6�>$���|��~b���R�B��M"ɺ��+M�Dv�o4�*Ҷ*p���}��c
�e鸭L<ˑ=	�D�i�e �C0n�X3b7�\r�_5���8 _�И �O>�7 i��aa��g�Y��B�o�ӎ 8p����hx���k���;�1������.V���L����u�9B�
��U�5��Z��]}����[_�8�]�����b������#�������jz5T���4�Z�RU5UDI�dX@��-n�\���I$(�KI�j�N���S~����Q����!e�,O$��C��8�p�<>Q�B��`O��G��C?�>Q����<g�?�>�2�eW���{^^d;Ġ�Ъ��s��>"�߯}�cl�,/vgG��\\��`/��|8.9�>�y �Ii�Z����n�O/Dg'rg���XTGP��r��	b�3_��I�F��6��T�f�Qa@�:��蝣�rձR,< �%ԱR�\úi�n�:L�K�^��#6��[���ϼ�޼���/���F��c4Z����H��5粎w�	~CO���33�uO��+�?*OC&��%�U�e|��X�ϟ,��QZ��)���|=����,+Y��q� ���0�����S�����i{��/dc��$r�`�r�e,Un���}�o��i��}r�٭�r�<�fl�s􄎞$10��^s�I,�����3�QR 0ɜ�l�i�/�����/v�VtQ�-�Ejּ�=��9���4
�H	"�{{���[��t+l��r�E=�2�o�]T&ښ�-�i�v��"�h��)G/1�S-~�r��9�;;��>J��{�̭Շ~S�7w���a�A��f�d�f�^������F�ʽ��^�/f�i�+5F��ׁ���m-(�Y�lΏN���o;������/�� [3<�X���v=�F�W�]1��2{�X�A֝�ݷw$�>�bs�s����@C�3fe�3y�`%���y3
�;	�_�e�&L���p�^}Vu�%�h��O7;i���Jݸ��w��o�/���限�O{�.��v.�ﻹ$z;���]�t]	d�ʣ�MQ(eJHCޘQ��@�YE~�B4y��UMn%���&�ߡ�f�iH����.2!���mՓh�+IJ+˖�<pI`���HJ��o��k�-11�f�
�%`H�ۗ:sq8ڬ��<B�G���Vm������͇�ޅ����ʣ��|��H�u�\�׊m��m��	�ݵ���y�kn�m�;�5���yιSӦ"#V�f;p�'")i��*�Meۭ��j��eZ�8��@` ����]��t�(������sV�k�md�9�R�G
��������}� �BEQ_W�,���(�j*(�D Q � ֐e:�
�4I$�EEL�V�"�a<t�x�^{��:��Ս1Ӧ�cM��?�0i�m�����s'AУ�y!��;:�Y�����Q��夀H#=��W
2��+*��t�*��0X��[5ZQ�JF�U���eɛQ+�bZK���t��P����5�_��tw`��ɏz=$X��;�Ebkm:"�E���!-\�o�	/\��k_��K	~� ^GE��n��Ɛ�{�>��k�o_���NK) (����p����z⼖����X����4@�c�ݱ#ڶ���~y����;օ׼�K"% �fd��5����]\E_�.��l�{�v���#��́��_ s��3��~�	S�TR�0�Vw�v�X<te��a�n�U�H�r�.|z��[l�|�y�uCs?�S�ɠR�aY�w�!
�����AWbM5�bh0��3e�jVZ��#��N�'��Jgq�	Z����Qiy�K3O�i�ߧ9n��$�Ç��yZ���`#�al:l��8D�4E��F��O�$r� -}XY	��9���zx�u����sEC�]v?_ޘ�(��[རF�#s��N>����n��|g�mK
;`�&V��{#& � 5u!-��`l�DKJ�'�#�����ډ��~-��uFS��Oi�D���Ql�mZ�z3��Y��y��:�%@��oj�i4<o��@�zaZ� ������Á��,���,v��d����(����<�l"�?~��hD�t�IJ��nqƹ�DvT�b7:�q��5	��"\v���IC�-�^�lٲ�E�OX(am�՝�g&������'U�]I36W\h�^9��b��z��ʷ��s� �\-l�c���E谼�1�$��)�J��,ts0�`�(�|l��@5����E��-0����C��D����V4�4�#\�q�o'&��^��G�w�UfYu���3�y����ó������9��8� ��4%j��?C���!�C%�3��D�����Ki&�i�ykJ0���8��3�p�&\���l�v�,��n'"���Dc����]�E7�� ���Gߏ�~�39�w��%�";�����wv�z;�������n 
>������%��[�{��*1�p(ԑ�F��!����%Y��d�0t7L�S P�%҄:w����!��wA��*�d
��@����@��$B�H[k�ȩU����4�+�]����Ló8a��fwpa<��$����q�aO�Wa�P�F�m��H����=�Y��3v��dt�Yc���D>���_�d�-*2n�VW^4���-:������|#H�v��<�#M��KY~p�p�w����qU?/<�s+?GOڟ<oq�km|����D�)\��|�Vd�����!2�Ok���9�#Q�#`�,�h����q���
��<F������� �����Q˴�:�qu��u��P�]���=p���5qb�X
H2<$,c��r���Z 7`��dx���\�°Ka�gH$m�_WD�-$Yi#)�ds3"�i��`������\��Qq�m,,���&`�,̩Y�;��&����Y�Gg��AhUB-u���F�1�8��v<�-Dai!�u�k�nݮ0���w�%u���-	r̮�c;��}|�ϢN�l{4F���h����4��~wiz6	���Z��ވ��℄Y(�h��[m�T]��K�O�>�88�v��/#N0v8��n�v�p��P"�O&��{Ұ��o�;���|��~D��1yp�ܯ(�~�ʩ���Yx�����)IJR�VR��<i�-wQ@u92Ak"Ye��Ԅ��-�Os�-�n�l8L�"���ij#��Q�~
3�߇5U^��Ym\̐�В{7b��f,��c����ԥ�iVUV����V�O�R��B3�Ev�j,��j5�OyS�P�r/���uR��|��,��21��ݖ�qS30;�ޭ�i��񧷗�c�s�'Զ�[c<H��YZJ=�xp[��0�)��3�z��oM�v�m	m8H�l�͙�{�-DY��N�Ļ�ɗ����Kq��������,��-�x�����.)���x/P�$���{��
��9�P�{[#�n;�L�/=��8K
XUW�D���ش���~�-�E�Q�#��4���8��.Wһʚ��~o��_�£{�����Li�1�5��v'; v�c.G����W�'!S�^��S�;A�=��0�DA�V�<�����	�=�e����5�?�H2�Ȑ	��y��|�;�&f~�w��%�";����ﻺ�=��www�����?C�9�D�x��$X��B*��LV�,4�� �v#9�ZI�Bi��؄����J���x���h�M�V�y��o�$X��S�-��O]��
�/hƆ�BVGԫ���`�f��o����T3�Y��*nYz��6�]q=yXl;��:��Y��y�dyR��k=מ������Om:��4�������-Y�D{� �\!����C�qq�#�-/kvS9�q �j焜Y���KC�\f�]=�u��NC�^\�ǈ��@5mmm�*����J��
 
Wd	$2C\<�]�PT[N�N�[Z�U�ܰfꋋ��F�c�ĸ�p�O��ּ�ᾃ�}h�:;���qz�-+���ǝz����g��-��6�,*X��k�l�U ƻ5���`�@���6��-���c�%�,ecB���,���6����3���aeǉ��$�6E� �lZH�$�t���D�-�����"��J��e��`�o�8,$k�Ϣ�|��a{���y?��i0����x���HE�$��~�#�;v8�FA�䁌cS>0�Yii��Gm�B�7
93�Vk3��;>a����w��7�,�
�4t���Xa�<Y����7���7��L9Cq�0ɗs�*<I0� �14)��-�1�<;_�hqj�N�d3�!�����l�w��)���~m8p5�����vn\k�^��ֿm���xp\�ek�y�=�j��l[O�o����M���<�-F���s�l"��p�&3��V[Q�2j�е�9�8W컪�P�®��e�fI��V� ���I�+��Um]K�NW^U?ce�6�";S�Pi���^"i�hC��h�X��0��'ɇv�Y����56Bt����I�y4�4�x����}�y��H��pw���9>zKu�]��g���?r��ɣ�]a��l���z���.:�Ǽew+o��rF�_�x$�%�'q(���a��n	q���%�OdN���T�����:��Cp�?~����;�",����:�q2rl����HJ��Ah��W+��<F����<^��,�Ǟ��D9�4��$ l���f���k�s�F�A���? ~���T������&2ֳ1|��-G�&`��2ù�$�oTH�܇!^�jf�u�,n;���_FOC��Z�K5�t.��!H���v���v7	�޵W*�9✺.��6㹂aN��
ļ��-$$�@��ZȂ�D���ik?�\���8�#��;�5�K}Ⱥ�=3��Y[F*��֞�:ċ+�~n�@In"L\@D���n��5�TÑ���^�G{�#�ѧ�sϚ��mAam#�����kǪ��.l���P�|H�Z�g(,��D-N��ܒ���{������㻺���㺞3Ѓ���,�ԁ�)�m���7��dLk4U4J9EJaQ01��#Yn%����?�N����h>RP�>ќ<a�)�+��C��-\���4��7�|�`�a����g�K�[��@-�n-<s�Yk�z�p��H����X�Qi-�jݨ|��]��Ǵ�T��OJ*Lk�5{(�!Y �\�<e�<&�	6~����w"=��xQ��qe���Ɯ�%�%�z�뵑����*��x�����P�ayfT��̹���z�m=�=n���h+-�d��B#�L����RgV;G+(��i��<!���{�+n��h�-fF����];��P^
�Xz�0�XIoq���L<Ț�̓0��4r�� ;�n:�p���4�ɑ�(�����B�G!P?Y��"�p��ڇ��$Qm#9�ӈ*�LK��Q]������}����eo��V�E��`��c�#�n h鴶���Xah��*����q��:\Y�]��'K)`7�kϒc:��-'�}��0��$�E����0�� 'a��P4I�H����`3`�-~�\�,���+__�SL�IE.�1�Ȳ��֋a[ä�
t�ȵ�\D0�>=o�q�=�ñ�s������c�z�&C���Q?D'��_���e&yu!'n��e�\rv�ݎ�Hr��kd��n
m�A$԰v���N�U������G�0E��N��&�,v����2�'��/���f���,nPd�����۹��������Oc{�g�=dھ�v��v.�+�ZV�~~�},b`(ݶC�Hy��ic���>VH�]���2 5�/a���ڽ�پ_��3ʷ�AۊQ�R`��/,�DxwP��H+.���}S~o���>I�dI~mA>_}�*�#�DɈ|9�j��yt:VK��Fs5�e��4c���DB���{�.w�绻����\�ǻ���麟 �S�v X��������<�zUL뫬�'B0��ߎ���0;�BHHC,6xAف!(�rT��e0�A�B��,Ƽ�8�dB�:�bs�[�>�x���W�Cn)&�!��+�w=<[���r��7˾_%��VZ͖9.�ݝq�h�4r[�����#]�Qِ(�,$8�^I^f�{^����۰�1�*r�;LTCƮ�ծtY㶨�2����Jճ�qz7i�y;n�����UJ��R�����UY]� -��rQ�qvv·P
P@Elu�L��[�n�:!y5ۈ=�<@4'��xAAJ�v�/G�t�����\$�>��mo�ı�q���L�K����O��ێxԖ��5Y	�"�{~׏�ώRn�1�������?0^��X��+�?7*c���-mvv���Ю"9��y����i��!��2f���b��m#���}���֝ic�r���P̮_3=�{�(U��C�2c����� >`�nQF=�Gټ^�T�U8����E,�,�Q�����6�g<���r�;Տf����5��(o���\-�z&���h��,����'��k��+6{iP�{��Ղ&�>j0`�Y�_���~���!l�GB���*NcnӓE�d{%�j�l=� X�%�"���t�
M>�����zc f;pT�̉��p��� R�7��W��QIp8�e�D:tp~�a#r�k����j1J����V�~ﶍ��_�,%��{Q�WS�(؇����&k��?�ǿ#�d~73~0��,�A�?�rv�6��6�B�y/�0&`8��{���uӔ�m ��v!�+Ϟs߿=��u��+U���ڬ��e���߶Ѿ������r��'����^� v=\�ڢ�>i�� 0?l|H8f�j:��/	m���٠r�=�㞷2Nҹ�\Z���d;�N��� SL�B�U:}3��'����U�@�y�.k9��\����>,�����Ѡ*+Xp�.�k�qØ	K�h4�.r�x��s-�Wj�Z�3�Ϯ�� GI+��^�������i�����DbN���K��������wt�w��븻���ae�, �	����v�@��,aX$(&)���X��(��d���[mt����h���s�eN����a�fӦ�qI�2�	�Mj,Wh���n>�C�5Ά�m��y��h
[��k9!�n/���ؿ�ip����&\�x��K�����?��|G!�ރVmQuPb~d�<��c��fI?}&!Ƭ�	���������YШ����y���a���>�#�O͠ ��aǸϱ!-�٭&�Bس.��e:ϤN̏[UU���F:�B'�%�{����c\}�,ThԂa�v~-��ւ�wW{�Wu+�竾wOR��c���L����7Q�>˧K��5�35����0���xV׿g2�K�i�=�����;�9<�S���.U���*��ݮ՟~��Y��I&����Yfޞ�W���Ay��/�aX,�n�>��on���أΧם�;�ؼ��,�}��Ǣ��!=~�t��l�D�3�ýV=pc ���C�^7��&��%�����`��0r� ^�!�R�l��f�F``K@ ̔m����b0�V��g�˨ ��>pO	5	�D`�qYH�"f�_D}iE
p�b���P�T5��ݧ�(T�g_?���{��1- n��,<Qe��~���Q��M�/O���m���(;o����]>f�����������]�`��'���_���_�ikYwc�:���F�ҙ��9U�.����!E�����i��x|Pfk`Y���چ}�p����?���"B��0.w�?{W�/^�W'�h�����{��=�ӗ,jr������ʉ�몪��E�h��>�2!�;L�A�����٢����¤4v�T�*:�T@�2
���
���RJ`�8�¢�JH��P�_�R���G �B@RR 0@����V ����$gR	�C&B�E�$h0H8Ua��p�@�JᔑB�@ ,D����B�VU�(m+�ŠZY����H�*w �Ӯ1����O����z9r~ N�2�ϐ�DrQO��0�g��U6��wn�����D�؂>�����٩ϱ���#����C�>���p�@G-w��y�:�O��=!���gxy$@|Åc���G����fg��0��9��t���fvr�x'�>ň�!*%)	F��E��C��	��!�EƠ�S�{�W6�(|Rj��c�_`�a��l�k*��.��R9��*����y6漳��� �0L(L�@�JPLD0�ID�@A31(Դ�PO�a&a�Y`��������
B!b��
�Xe@!DX!@`�
�(�h���R��
�JB�(ZB����$���Æ`�h�(��)A�) �	b	h�d�Uf��X@i@F���"��"*	��"�)Ji))���(���	�`��bZ�� )BiU(�F(h�i��`�� �I�`�&�"&
��D�E1#AIDK���*ly�4�pZ�X�A���?&f������<�ET9L�d�e�i���u���zO:��N��7��0d��g�O���?�G��Bi�g%�@y����g�ͽ�a�˄0� p�������=�k�J���y_������ÕQP�N�7��4~�g���7�5-��{�@��UT�<b"�����Վ6�����^{�P����$Np��y� ��J�:MDx�����~�  ��6���0k\��P�����" !�� �t�I�d�'@�G�v5A<�ͪ8pA����/8s� �3�=ۃ��|���H"y���ӛ��wG��=&�����&h"��|��S�$@z����?^���\����� x��@��Г5a�8�L�9\��w�wg�xo׽��?���s��"����.7������|WV�w>�ۡvDv�Al`3��M���̝D$�(�����9u�D�T?-4�ɰ��<^��1�w�C3�50�6�ӉLz2Wȑ(oːpx��)����