BZh91AY&SY0��9��߀pp��b� ����ay  �� 
R�!@H�U(	@BP
  Pz �AU@(�@�	EPRT�  zEEI"((
�P� �!
�($P �J��*T �Q(D�B�(UUPJ��
 <     �      =���>����}����������fo�u<F�s� 3 �=/���}>7��E
B�J  ��aTu�j � ��R��L�P���8��>�:��)̀�v�aC���:��;�$�   V�� ���ҨYoB�W�T,���熕���ޔw���i{:��ލs�� �sw�mJ�[^(@7/U��`{�0���f�yC ��� _^�S,��3��9vs��z}@      c�G��-�{yPͩ}�^g�� �gp�����.f��>���У��'��{��*@Dr�rq9Np �����x<��t�0;��x/p �xzw;�d��ǛW&��9�#��     v����]�����Ͻ��h��} :\������c�c�I3��(^ǽ#��'��q�: A�g��z�p ��cvp�����:�p ��&Q�%;��,��>�U@^>     � s��t}�;��f���*e��rt,��y�,�]+��ӖK��ʻ� �&*e���*s�E���>� �9W;>{t9]őw � �ްr;�����^(      ����J�J0�����&!�&���J�4�d    '�UR�#��	�L�hd��'�T�L�*0 	�  ����M�T�( d    
B�L� Jm�y��4�44�O�?�����_��}O����}{���������������QT��PUW� �����Uo�e� �������U��}�@UV���9o�v��U���X�.�BAr(^(H5������xM=���"FLB�#��-F	$�\�Ρ�PZ�u�an��K|?n�BOݩ�M�r�CɅAB�\R�*qY4�X����7��7�a����^�gä�N�]]�<�("���BͲ������rSVT��X���D?]�6A$���KLDWE%[^�E$U*񘖯�|������i���qCYpCX�	���|߾��gI������u<繌�j81s�!f-Xە��n���.�MH]o�E�������x�蟇W{�#餶�x\��V?q`�ߛ�w�v	�MV�;�4a�a�2��FZ�%O�P��o����&u�LC��!S�D7�f�#��W�ƚy
'�,,(���N��(Oe:��$�鏇��p�fj��憉����8�n�a3>>G�L�ɘ�E�l�I�ܪu8��rlg��Y��]��p�z'gc� G!;���!̲�.�V��,<c�+��x�8\��2�,&���\��<�$���	o��n����%5�������8[��\woK��xT
cS"gJbs;��,C��j���*��L �,�+J�]O�H��3�'O�o���B���NذT�B�����N�!ݧ�6����;�p�7~�Z&�^N��:tg~�1��Rֱ(���p]FYh��>���|Z���K|�cF4`�ox"�Ν4�*�"���Ӭ���p�����C��|&R�D*J��ő�Q�r|}*�˕�r�x�/Ї�c���Z��"0�2��mON�0��C�	��:�6p�Xw�X���!®��yl�׿t�{ϙw�0��p9�g��'�uߝy�����뗩RK;���������g<,�L�c �ɉ��#�ג�!A�$$�a�9S�PkL�sGW��޵�d15�Gl@�7Mޔ�J��Nr�j�VI�������;��V����Z�<��0�a�# Y�>u2��Q�b�lKD�J:�k�v�͆��NCӣ�q�3��%�@ļ�&&TQD"Bj��g��>�w�y��9���l���0�0q֧5	�˔F��'��8��5Ù��5c�Yy׉m7���{��;)��!�[���R�W��sy��I7ɬ�w{��"�Q$�!d�;�Mt[q�'f�^obꚚ�bB^.N]f���8:�����h�����n�nj1}�H����{7�Y�cp�ھ�VLLǋ���V�L��;�"�E�1��/!���\�ma2���y���q�0Ov{�7w�T:��Y�H��3�p��lA�\��VP�O�fnF��]�{�ϻΧ�ǱD��G �>�5%g5���#(&#'$�FW2�jlNH��_%�p���&����$,�T�"������y^��8�kπ���}�F$�M���qr��,��F�5Շ
Ώ:��>P�c<��ʥ�<)yӧ��E�hb�L��KL�����]���'�F�5 �B�r�b����u�o1D��c�����N1ac:��7���]Mi�k��mJ��_r���$���'��^5��7�w/��{v��K��CP2����ue)Ξ�3ז�'�Ɗ��בD@D�)j¡���s�nV�$k�k_9��q$;��p��j"2Lc#r�&�˶���¼ꚜ]�Z1̣��Lkz����`��S98,Bx��ĽÑ��X��q������}�3]kZ���JM��ɬ��*V�¢�`r2�*+!1���֖7���oݘ!Dß�a�ա��11���6k�=�	I&X3����r�1u0A���"	a��o�`p��dA��Aj�2��
�3gS�KS��ua�a�'i��$Mc�$L���ict�$h�J(�tp-h������ �p��^SX<bН&$��4$���Q�.\�Z�h�q! ݑAd�E�Tl���/9�u���k<o�3AYL����*0H��9(�=k�u�P"h�SOC�8�oW��34I�|����j��O��x!�08��դ�
UVA^f�q[��I�������4Ij���<�k��D����ub��`���莼ۻ����Oa��d�N�B�tkQ칧7Z	�d���H�����J2���2\,�%�0�8LQ��1�*"$,k wD9Zf����R��bf�'==Թ��c�$��[�&8���(JI�Q��~yκ��{���%7T8$$�niO\f�B�|U�߫��5|q4`���d�x}������3R{����LZ�u�h��:�b��_n&DWN���$%���8����c�m$�PU(�`�^��>�9�Iq
��%���5�Ey$ܔ��ƥ�r���i�ݓ}�|����9S����oΜ��ݷY��О`��r:���O��GZ��8���B��l��/o1�L��Ww��q��uԦ��Y��S"s_o�8�&������/>sXE��ĒR�"2�<Fɕ��ײtq�)��<k����.��돸*���}� ���>�F	u��v�0Z�Y+zj�Fq6�]�vӏH���BU`�1}��Y�^�%���TD�E�!!�I1(����l���1X��1���ڊ��k�Qs��C�,�髝��Y��IŚH�Dke�l�L�8cGx.=5vs�A�`����:+�?�'�\�CPn�{�c���H1#Q�%����F	f��NN��ז��f!�^��L�I��P�5�~�I���s��Vg�8��e�.��y��H{wCz{�j�3v惘�5	Z	2�Q��,jQ��Nۂ�r�S" kWd��^�*�1w��5���n�����<��\���|?snX0��U(����%	LM�C����,�n���y�5jſ)�Z�I�ƻ��d{��&��|s�1���/��9YV�`�
�F�i�j1�E	P�����&BG��P[�}{� ��d�&%�>n�W�k8��<�g �Ux��3k]p�|4b�:4.���K�}W�J�^�`��}F)���<�}�{6�ʁ4	VR>CU�������$�i�XI��%�΋'�5�*�LL�dj7d�k�ړ@�2�9V<ư�X�]CGVI9&�7W������CM�jX0U$�o�����~<!pƞC"1�B�8�-���ӝDˈ��9�V�����[���PD���[ʱ��Y��b^����Mō]���sc�<8��؜֙�c�}����t dh��Y ��+	p�i"�\mt��&�(L����N�)��8آB��8���u�*t��
�eeP<�q�h���k�k�����b=�]OR�_��q�.>}�A���_k\{�SY��B��%�*d˝�Vv�P���R����ѹs [��I����,���@��Й5�q��`��p�n� �-��R��`�L�N$drZFG�դ����^�w�ò8پ�SO��,��Q�����nC@�bWqa��O1&�c���£�vw��f�4�U�Nr勐X3���?]�	��>��q�7��q8���k}Nrp�lGx<��$x]WD���	s,�6�0�[�C�3�50Ղ;;���&�y��u�GGw�7�]�|{���#2��Ds�"1����>(��jU�@�'���ћ�5���s�1���H�'���e��b�(��
�WVz�K��G0��|�iB��D���
�wǓ�|����E蹠���ܺ"D]*߻�����vw��w�~��]����u?�u�᫞V�ۇ8�RcM�&���̉��7w��]k�^�{�Zy���F�b��P��6���&�n#j�=^@Y��݋N.fE�p��`�qug��X<�m��c��״�����q�������'$-�m���w����uq��ﰞ��}��i�O�	uW�了��Mٻ��$ˁ�<�\��:F@*x���Zj���C�ey
��=@���G��Fz038�c�<�f���Z��|}�xFN_{c����
#6�����75	Έ����1D(�$#P�YӼ��,C��
�o)'�`�Wuc%�c�Ɩ�1��!��:�Dnq,q��4�V#K�4��>�]O{��������'=�Գ5f�%�3���1�D$����7�dXǈO#�?l��c��{/,���__��ΔA�ӻR�9��R`]������m�����
͍s�$��N=�ѫ����6w8��"g���Ϝ���I	nx�j=�NS�7�X�<p����C���ŧ�iӝ�|׶iw���&�>���Hc��R�|j��Pp�T_g�FBu	�M˼��1g��D�0\�D�c��#dX��L��$�N�����_K���q|��d'���=�>���1�E�t�u�z9�]^PVR�ڲr�C��21��	ı�G-f�z�֎���$�'�n�܊%;S|z�=8"�lV�uPP��lX�Wo7�}�Ԯ�*��q��7q�%Ҁ���A�d��H���'*hB�,Y��F�N�P`�84���i2C78:1l)`!��JI5 �f&#�5�g��Ϳ�1���72��qL��(  ���C$;�Ph�4�:=^��J�a�2P���TdF+;É�Vi�NlѬ#��i�5��}�ĉ����Ld=�BR�Nd\��
�� ���� �7[�ZtiƦg2\r����7�4Д%	PN����FMDBFb��HH4�C%�Z��w�Z��,��H�,X��ۘ�mw��{��3��$������);3f�r&t[ ��ANN$�,k-R4	�D��ݫ����S*��s��ٺ<H��.�kQOSSIY�Eqw��a2�,s�%\��[����3/	q�06����O:�c*z'�BkH�u4��h��֓Z�b�PC݉��d��"b�o�i���S����m�H#�\:�<HW��𛀠'��F�}%Ndch5;���3N�5!a��N�b��
�ѐ&�,I�4cFbj �q��D�F�Sjs���c[�8f� �fcϡ�wt�)�N�NpF�ֳ͘ňY�$Mz��@\�ūJ��<i���R+�p]�T	M=I��ż�o���Df����`�O���r1� 8������2 s�Z���O��IW�1�t��ʅ�j��z�!�f�e �]X$F��Ѩ�H�b.5��C���cXňl	݀v�����7��韊>���ob��fU�   �kik@    �      ��[@   �  h� 0`)A�  	�  ��      i��      $    H�  �k�)g@      �lm�$cm�8 m[����      ���l�;�|Ht�R�����$%�]�Ep[m�E���N� C�k��)@Z��I�P��n�RM��@$X�N�[5�o\2mR�$��q�5�q��L�/OJ�Pci �Z�s$�U+i	]�vj��&����lm�$����n�,��EP��=t��V�m
�m�a�ԧ�c�jA˦��4�NI$�^�����[N�U.��j�-uՔj��6@�� :����l8�m%�Ò�̙� �;T�mUU��ԢvN$�Z�&�+��8�ni3m�#�5Y��l#Z�.���[���Ƥ��J�ӽ��C��kr���;�mv�$�):H�K���[ckn�u��.ْpl�`i�ڝ!+R����UU�1�-��m[Yqz�ۥ iL��_�m���4�T�lsm��u
V�F�:.^�!&�ځ�N��l��US��s�/����#v����e��]�pg�a�Q#k�3���о�Tf�ҩm�{0qT��v�6Yi	���K)A�nθgD�v�E�Ґp�6��c2�tv$j�m�yM<p;g���h		�r�gX�k�Z Ш���*�U&��Nd����\:�#�3ع�Ij�*�n[B�mu��Z�V8�{D��r��I�"�6ݸU�*,�[V�����D�$ppH����K'^�8ᵺ�&Zd�Z���^�9�]�T�v��۞��*���|l[�E�U�!�ኪ��MbpA��
�Z�n6�3�L�գ�V��] =n����Y-�i6�t�GgL��箞@Z2e��
)��:�h�eb��!V����l��gcB�T���
"��,�@��'k�tY�.լ��b���e]����Z�f�mB�M�rF�Us5ɦ�`ԉ	�]ָL��x&����Fi��Z�G�����������c�[i�������������;k}�a����I[ɺ���Y-��Q�Cz�X�#&G�˫z��;լF�=���Oo�6݃�-Zs̨۵�1\����(@j2�h��X�;8X�p����rs�T�ׇ��ݬ� ��\^��M�N�6tU��[ԲA���.&iy��[g�p��Gn*v��d	�9+UK���������ӭ�n�"��k��,`آXM��y^�m[J���J�W�}��+�!rSN�Z6�$k�U@rY�U� �UOG��ޮ,sJ���k���L����[VԀ8 p�ٶ K���[rM�%p �h���M�Ғŷ�:-�����*��_E��]mVy�j��	Tdy��`�s���0uV�t�R�lq���8<�d�'g��݋�A{M� �aӶ�ʮ�$�`��VQ�;Pă�od�M�f�vs����ГKLH8u�:U�W,Y:L�;]��k� �9]mK�e�b�a��N���;9.x$�F�v�TJ1��*�hEڃ�8p`al$:+:�j������V�sJ�epM��7�N��d��n9��gA�9Z��fx9��Qܷ�P(9�Y����[���p��)/A⍄kӷU���W�����6��f����ѭc�����U�­W����=��b�;דvƚ�jG�N6�������Od�Ap-ꓖ�f��G,ǴJ��;uU�6���ҨmN��e��&Ʃ����M�-Un܂��Y��UU>�2 ��n5��p�U�(�$h7�C��J�V�e�X���yx�m��,��K&꫘I��6�m�x䛒�se�]t�`�m�M��M����X��ЍZN'�T�m�5�lu��<�L��3����d8*�_U�)W�Z���.�Hm;�$�rE��U���5\�U]*�P�Ԁf��%	����յ�F�����:���Sӕ����d�n����2;$�2m�&�r�:vĽ��b���ViV����V�@�c}�rdWc捆��>We�cnZ�����$�d�k�| 7[���I`آ��3��P3�M�%�����XaTL,������M��+�r����;r�V�uU �e�����J��]��Yy���v��4�ڽ���ld;f��0n�C��mSPu,���/a�^�3�7b�jc
���vB�����]���h]�"lP���}.�lq�np�k�v�v��x�!NL��On70<e�7:*�#�dH�gL�k@�P��뢅T����-u�1:�u��iW���+:AS���.��"pI{k�64@Y��q�R��j{�y�c������:9� ��UҜ[ru�rI]�[��e@�*��Y|��������8��\@+q;r�����U�	l��|����t�jj��V
ʵ42X�L�.�뙶��L[-mJ�T%�<�����ݶ�
_We��U������ڕ��m����2����qNyYi{&)�]s7��?>��y�k���{^|7����T�# �}���0������ �nY�UU+��\�ʶ9bV�55�\���$�6�h-���/@ʲ�*��ӡ�y'm0��\[wm��� ���� ��X  5L��孮�dtE��;v��m�8'I�OFٖ�a�-�%��SsuPHm�҃�x,N	�lkGk��+�num�7[��]Ûv��Si�2vŭب\�>�lan�7V�%q��l@��kZk�ݼ��N�� ��)γ��p
��U�#�GJ���nҰq��pjlWo���m�Fܳ���\|����n�{b�r5Iٳ�u��Mk�;A� ��0�Z��U2V��;4�lv�Sښ��g�GmT++��Hm۰ r�H[M�m�w�e�$	ӎ$�Y3�K �p���c6�A��8�Av�qt͑�Zwq4ŬT�vXF�f�u[J���*کt�ۀ��VPn� 3���c�Н 6�B�-�A�;4p "�vК�D���mm��m�H�]���R��*���j@k�6�K��[M�m�1]J�]A���U+�R�8�k]��{d&�[MU��%���g�kqiU+��a�E�TP����,9n�A:6i&�Hdp���K�#l�m�J)M��l <��6�$��gFN� ɀ2��m�t;C&���F�\��v�+j��]R�Jp-V\2v�^���iӀI��-��^��6�M�H�.��hΔ�	kF�jմ�\ �̎ٵ��pk��l   �ձz�n��Yt�$����hN%.ݨu�>�:�����yn�,H�nmԞ��oa�E�֖�Y�l8At��j�mm��6�m�u6    ���B��U-�����a�l<��J�ۜ �I	$ *RZ���G�-����j����v-�� �oQ�תL��ֳ�� ���K�J�Cn����8� ۴��h  H�]�ggC S��hv�b��'n�n�5��h   k�-��9�`	-s��[\����B�`<$�8�q')��UHuB��\���]^�� ��]��rK�i�Z2�*K�����U [[i�1 ��[\mv�����?�*��5Hܠ���`Zm����v�5�m"��FlKm|��>[d�`  W:�iPAUn(x�4�X��j���-��Fձce�p r��2ڷ[��-�m��m�����h�P)�۴��kp�[B@8�$N 6�ݶ඀ 8�׫@�>��ϟ  ��X]7d�A��`l���	lb�{;hw9�z��{r���F��@�\��)�PC5$����#��U�)-T��b����"��pu- �敨��Wm��A�]��� ��lC#*��uA��KT�[lN45*�<4�K�c�trt�S2���^�f����/Z�h6]'�j^���d�vQc�����P8��W��kj�e�zʺ��$m�z�C4� ��1�U�`7ݹ�磛���.��sˡ^gD��NܽGb�r6�R3���wDCk�+���۰n��^Ʒ%W��Kg9pm�U�C\�G��N��!���NHU�"^9o����*GbYXI��f�4��{+Uu��T���y[n�,�ӭB�8�^��<��M���F��԰u!�M�������#ײMc�E�:x��1�vݶ�6������#��vHu�h�>J��9I�(�l��.�oa���Z��x�m*�TTʁ!��� {hi�91���8�]'��vXr�WWmJ�U��;�� �ĭm�Γ3v����j������K�h��U������r�Weq���u\�ml*һ5]lSg�mf�`�������  [��sm#l ���O]$ÛWl$�۶�ږ[jA�� $竫�*ԫuJ�u��=l�@�M��� m�H�m� p�l ���6ݛl�n���m�I��l 8l 8[@ �8H�  ڵ�-��  烇� p  �h�6ۀ q'6�8�`m� �` �#�i6��   $ -�� m�l�R��m��gm����3��Zɛ����Lۅ@R���v�5WP<
������ʼ�;H�Uu:��޵��U�_㈂*�����������o�x������D(�LU%t#��(�z�(��$J�	C���( "_�%ء�Fa]�p�CX��B���螄LA�h�Nls�T;C�Q6�`�r6 ����D�=S�� ts:\ ;*��*iC��'�t'�����3@�`����/���/����&"����fhA"��]�:;@x
mOa�W�x��}P:��6��*�0�"�DH�R�� ��7�.A<*/�W������]b
���=@<�����T�������N(�z0x"�0�+)��]����&�=SH`/m/��EN�;�D�6�����B�о&t��W�������D��9�9 B����{4N$�@�!"J��Å"���Ȱ8b�����b� ��v �想C�i]��*v�z+І��;���&.HcN%N&˔�a�b�f���6HC��FE`��a0d��6VaR��Q8��9�K05�˘�I���a`8�)�Pa�zQSA�3X��B����A�*���!�d�!PЪ��@pS�D������E@UW����ݟ�����z��Q��@�(�H�JHU��T@$�#,��3V@k%@��!� � ĊÐ�"L�df&d��(ѣ$�)�Z���F�h��=ޒN��������h�� ���!oϟ��gm� ������-6 ��]�	8nMjz[l��Im�t�b��͛�VNA�[gj�Ghk;zЬ�eN��P�z�W#W<O-�.�k��q��t��V�rkq�']�i�[5n�N��y��4��r�sͶf8ѹ7i����7h^���ch�Y/2*� ��I��N$ۋ� v�����t��E�}�(���c`,Ib�`�H��㋷��l��9gs�OoM�D2�ud@��lՍ`�vs���{n74���9���=]g��Ii�ۭ���uخt��݃J�k=�˶�������t�7e��GvGi�4o<���+��Oa;��6�W����:|��:��ݹf�ݻa;���iwd����l���Ji��we卌=�v�V3�8����A������5�l������)k\)���<tY؇�]Ű��v��%8��ܷ6"m������m�m��*v��w�,�u��Zf��]����N�^(��[v�1�wYt�V0�B�kg5c�� �'�F�G�j��j�pt��ݭ���l�Ugt(ڋ�s���cje e/<��<���V8���7QK\��̮^�Oy���<v���<;Y"K�yً��N���8Dڲ�@��f�q��cl�8{��.���B�v�`����f���!n�E�ր����V�G�v��m��ѭ�K"��ؖ�I
��v �itTp(媦j��m�	n��2�)���I��2�!��ɮ�q����ͱ�H�ۛ���:�H�k,�#R�5�۩@ƕm�O��m��]��G**B؁ۓA"O`E�JK�&��_\�rm�^5�n�%.�Xn�r�t��ۏ��]˔����� x\������we�݁ۍ�p��u��v��/E����k�W:-���u��f��ʒ�$9�(s-�C��)*y�2P�wV���#5�J怞Y2N�/���2�T�MR�VS��4.���Ŋ6�����=�`j�`ڠl҇Ȧ�5�� ��N/k�x�t��;P>;�asa�|���-�V8ڮ �*�u�[˖��@�>���ne%��n1a�[�g�6�=�c�[�H���S�l3S����l���&�=�/�Θ2�KOI�,n�{F�=����N�1��gu�q\N��rbcf��D[��I�2�HAˢPn�k��yr.�۶631�М<���t͎��H���4�k��k����LB��l�?��ww��Nf������RLLi9I�6���ϔ��9��q�6;sJ�`�XU���Q�������=�����x���}�K)��զQcbi������w<����������i�M;i��ό �{� {�� �y�wy�	U�M]�jƙ�u��`��xw��]׀u���0v��hV�i5�ws�;����;�`lo�lgwwx���ET��&�ڌf����L2�U�;�Z�"}q;?
Ք4��wcCbo@��V�.��:�ܰ��x％��dd�v6�ԗ�>���KL¨��X�� ;��w{��}�
����iP�;�:�ܰ��xw�+ ��u��W_�lh�Bo =�ڰ3}���;�`�ݢ7ڪ��jK)��%m�,N���7���>�|`��< ���*��ʥZ]&ڿ�-�l�S��v�<���;FvTV#�׉!unś3�wn�t��[��m�i��p�}�x�w<{ό�G��7V��wv�j�0�{� }�� ��� ���~���_]t�����h-��� zI�U׾o۔�ؙE����5����� ���:���m]��o ��� ��������x��\�m�ht�Wv�3 ��������z��޿-Iu�הq�;�1��|[�6L����ZV&Z@.���t��hA�9�6Z�춓t�L�}�x�w<{ό����u+wM�*�E���ݫN���|�"��T� ���`}�u��e��������|`�V�'wv�7uU�y%V��F�[UD4M]��ݴ���� {���灿�t��8T\u���]w���V�f�[��m�Ӭ ��� ;�s�7��w}�������ߛ��m��lmZ���k��n���VѨw�Yr��h�*ݰ����ՃNՠ��&�{��7��w��+�~����=�u.[��e;v;m�{�{��{� w�� w_P���Wt�6���0�>0��<%]��x�8`��%\�vݖ�t�3T�	ݞ#wUXԪ������oe`�Q�R����������s�7��w�����<��U˻�M�Onlk�����*��l2��6�::�-��&-�+����Rۛz�q��qκd̗�A�;\�Ezӵ;�ݺ���h�Xt�Oh�l�p��܍��v:Z�]$��7f�H�Z{����#m�rF�:W\�-��^�+�%�=m�6�ԉ������]2�7]$RLh�``c1�ӫ�cw�u\��Ѻs���G:�QSI�4�M���l�˽�w���㟭����8�n��nd	���e��qQ�X�Y<u]����*�h'	\a�+o@���ݕ����w>0�{�+);w@�ջv�0wvV {�s�=���7��Ϯ��G!1![��m�m� {�s�=���7���=��X_���`ēJ�&��x߿UU������+ =���|����$��N��-� ��� �we`��<���jK�>�m5��i*Ңq&8E����1ȓ�8�iz��s�,�rp<��zĞ��Ξ���uv�M�b����X�� �s�W���l>�2��B���m�,v�d�Ԓ�}�ӿ���!�� ��$���%���D�N%3 L��̮�.j�`|�[Xn�x�R"�4=LO@��L�X��`o{����+ =���}�x���+�	������3�;��V5�䕵�{�k�=�|`��/�)�J�U�v�X�ό ���{���7��X^����6�8k5�ٷs�;�릌�&�fF�W7.�Z�s�:�#8���i[}����{���7��X�ό�Ew
��&��Mݦ�{����ό ���}��uv��N��-����i`{v��᝙١���ڰ=�����.�ۢպI�]�`�|`��<�ό{ό ߸���m�tۦ�u����w>0�vV��MIw��!��n�J���X'J���`�����[�E���.���ZƸ��q���2�$�����������}�x�q��ի�خƓL�7���=��X�� �s�%]�����N�,Ujݻi��2��{��ό{ό �]���]���ӻm� yߞ�{���]w�9[CG	V���+ ���v���J�v��;��J�U����$�+ >���}�Z�?�d�]�D���m �P�dof8��;8�-�uݮ��t݇[�����~���;����� ��� w������I��H-��;����� ����we`��J���7@�i����w��w���ό��QV;��X!&��>0�ό�ό �� �޾�n�a`��ƓL�;�>0	S�C@'�<�ό�Ԡ
!�!(J��e�9���l���ְ���a+� uS��5��q[���-���:�l�Gn�������6���X�OW#n��ukź����[
J��t"�Q�L6"��l؎��m>ݍ�'ssب��y����L�K�tػ7��:x:�D�^�p�ە�������,S��t�Ż<ڔ����~�vôX�.۱�/c��T�`=�,�K����V4��P���;Sw�|p ��B��:;p%3�ך�l�]\����#�	GX���;+��(�cv
�mѩR�Uė�{�� w��w��w�|`�w�r��һv6� ;�s�;���;�>0�vV�+��X:V�+i�o �s� ���;��X�{��׫�:�S:T�ـw�|`�� �� �s� ;�W���e&ݤ�����ό �� �s� ���=�:���M�=�3��.6յj�ډ�;�^�[j�qH�U/�X�Gf�Mħ^-d� Ϸj��N�X}�ӝ�� �E������hi����ж��3<��K82b�iS�������Oۿwe}�_[n�a`����������}>Y���i���<�N�S�*A�R%V��ܸ��{ݕ��������~��:�t�i]��g����]�\~�{�+�ˏ���T�����˧;�pl��
����y8����w«q���+=��]��'k�K#�-��}>Y���i����;�}����(�Z����EP����o�t����}��ga����F4ʴ��$	���C��{ݟ��~��'� �+�ֻk��ѝ�5Dw�l{��8��fw��
�j�K-���!�AsnN.Z��Z�}�#�>!>S8���؞Σ�`p�B� ��X�#Xo�10;����/��᧦Z繩�<+�N�z����I���Pu����'�y��.���B3m��(I�d��i�Se!P�66d84)$�AA!��"DS$� �B��1�ˬ���$%�&⭥�ci��Ilfg��D�d&`� R�d�ᒹ�f3fFae�c$wz�Q%��,Q�U ���!N4���(�B,X�"�,�Zjm�qsD�I����ЕdĐ�mԱ8�\u��0B1�f4���mvj�՘� öq'-Q�v7���>)%h4OZōu��A<�VCF"�7�A�='
��{ɏE���1��z���6��&Ad&<0^XH�`���LVYn�1�@�|�@#�2�k���3-��Ap֝y�$�l,#0�������F`���%V�Z��@�2Dcc�%������
�sz��5i�Ezh��4E�4�W4$�P���c8���	VkH�� �
�0LL0�����'l-%&%�3�Y��7z4[MC�jH!�LDй.@P�%�[v0��6X6�M�u��lu�剮�42de�g>���?
v�]�P9��*z;܋DʠD�,��(�"��tj����C�A��>�Ғ)��J}�[�┥'_}���)K�>�Z5�٣[2��5��R����}��ԥ)��o�R��y��pz��� �����qJR���Z!4��T�4AuUWl�;�;��_\R��:�߾��)J}���┥~{���)OO}��E���Xn, ��<����[hJU�$8L�y9(8����s��TTiB��%�n`�`��߿h�)J}���┥~{��O¤w)J~���\R����߫_�ٳVn�n��[��)J}����4�~}���)O��\R���~��ԍ)w�g�~+�H�v�e[�%�$g}���g%)��o�P'�����)O��-����g߈ۣ�:������9)B����)JRwߞ���R�����(I�&������#�4�P= �
�>�ζ|���eĵ4K�T�ADN��)I�~{��JC�8(���������ϻ��0�}��Q}��܎��P-ͩ�\�C��#���^��ss�ܚv5�`�D��]��JՒV��?�`�a��}ÊR�=w��pz��;���)J���ߴ�,�,�~��H��:��IvqJR�����R��~��8�)I�~{��JS�}����������f��1�9o{��JSϿ~��)<��~��)Jy��┥]����)O�}�9�v���v�՚���)I�~{��JS�}���(z��~��)Jw��s�R��xy�h��l՛�[�{��=JR�{����)G�I;��߸=�R�}��8�)I�~{��JS��,�ʑ~����HݒR[Ь�P��	^z��jݤsնF��uv��`I'V��q�	|��;9�	/kS�=+�Wc��d�N�;P-�k��mt��Ӷ�+�Awg�CYc�����j�Y�����aS5��0qd�eM��m.{t�.��.6�YA�Qv�/V;;��C�y���!�m۝�@�x���7�z��b	n���pp5{i~�MtY����k��n+H7Us)G5����)�l3����E�k`�;]kP��=�mt�#N��mr��	f	��~��8��;��qJR�����ԥ)���%�%��|ϿY�;��ݻ�qf
S�~��JR�����R������)JP�ߟ}��R���ߍl��[5���qJR�����R������)O�!L��=���ԥ)�߿p�Y�X}��߫�W,V�[�L��)@_=�\R���>��ԥ)߿}ÊR Rwߞ���R����֋_�Q��%[�%�$g;�ߴ�,� ?�<���)JRy�~��)Jy�p�Y�X~��?ߊ�ⅱT�n�PpwM�q��9�5� �8J��m��������=w��65mli4�l��qf	f���70IJN��߸=JR�{��8-)C�~}����?}��+��ʢdRJn`�%'}��������7)�����(}��~��)Jw�p⟄IL�����گս�Fn�o3{��=JR�}��\R����>���!J]���┥'}����)K�s>���k-귛�����)��<��R��߾��)JRw߾���R�{���qJR��}G߲:ԒW�v�Ř%�.��빅)@���pz��;���qJR�����R���<�~�G�v��f��o���������6z���W0�u����Ijݢ�ojl\���֭%*�RT�����)<�߿pz��<���qJR��<��"'R��߿}�)JR~=���������[޵����R���p�
R�=y��pz��.����JR�����PY���Ȑ_���Ұ��i��Y�Fu�}��R�����)ӻ� ��C�5��	�
 �8���(I*d�$���CI� ���߿s�R��~{�)JP�xy�>�[��,˖s|��)J]���┥'}����)O=��R�(z�Ͼ��)J~���+vJ��n�����ý���=JP��{�)JP��}��R�>Z������-R��%5UQELko1D[ɮh�[��^UȻ���c�5p�vI,h��[n�ZC�E[�]3�0K0����8�)Cמ}��JR�Ͼ�)@v���l�;�;������b�Hj��{��)J���=G��rR��߷�)JO<����)O<�\
R��|��du�$+�.�ۺg`�`��߯�)>�Ͼ�� Ҟy����)C����������M4SQAM41U�)B�}����R���w��)J���=JPx�,�@��L�`I�b.`$) <��Hh�SX�4��T>�����]��ß�Ϣ��T�+V�f���z��<���qJR���>��ԥ)w��o�R��y�pz��;�3��?������\6�4,ۖ7U.�lY��&��u�+9��B�`����ܽ��/@޵�kw�(~�Ͼ��)J]���┥'�y���)O|�\R�����������z�]�8����~��	2R������ԥ)��o��)D���~��qf	f���7lu��ۣ�{���)I��{��JS�=����!	����pz��/?}�|R������Z��(�Ӷ�Y�Fg�}�MR�����~��)J]����'�$2O|���R����_���ֳz5������R�����~��)@~D�3��~��)=��߸=JR����8�Y�X�?�������c�![,U8�QɔZM��0�c5�磑��ͳ[cM����g�V:���vs�n�b�r�Oj�pf�<��]�ȹN�;�z�n��9*��]�8'p�U�u=/`ۧ5�8�v&�C�yd�K.�3�[�RΐzI�۞V�͹]�;V8*�,��H���.��ݞfqF\ѧy�H���;�_Eؑ�q�������i�<:գ�����F�(3͸.��Y6�n�g7m��b�:�m�5��v�uH*�N�+X��5�q�,nIbJ��v��%�/����]��)=��~��)J}�p�JRy}�S8���7�~%%L��[e��)JO{�߸=G�B�J~���8�)I�j�g�݁݅�ٙ��݁�۰�g�Q�2��n�t�,�,���~�s�'��{�ǨiK�>�|R�������qf	f�~���\��eR�M�_��*)�{~����)K���o�R����pz��C�=���+˧��?ыmBi6潻L����=�|R��U}��~��)J}��┥'W�{�ǩJS�5�5���Xo�cA��jCK�<��3��zZ����I����c<�rn`�k]�ֆ(�RSs)I�~{��JS�=���(~�߾�+ԥ)����R��zyl����f��Y�o�ԥ)����t�,��
Lx��Mc��DT�XD@PQ88	�@�$�@�,�L��	�z��C�J�κ��)Jw��┥'�{���`bY���~_���;�cVU��X�?y��pz��>���qJ@)>�߾��)J}��┥'���}�[�f���2�s|�6=JP�����R��y��pz��>���qJ)>���=J%�|ן��*+l��H�[�%�%���[>����H�vvd{R�|�>���qJR���s,�ߌ7�l�9^3մŞ�sv���y�+O2��4�B�]�&('w3 �jSmjY��"�ۦqf
S�=���)>���=JR�y���"R��y��pz��/|����oZ޴[���5���)JR}�{���������)JR~��߸=JR�y����N	a����6/��qm������w��)JO}��=H`�@���`3/��!����D�ڢ ��ZV�	� %31g�pVT�u+r��������K>���ځMUf�3y�l�k{��"�����pz��>���qJR������)@�{��f	f	a�Ǿ���mJ(�+NK�qf��{�)JP�����hz��>���qJR��=��R��w���n����Ÿ�Ȍ���[��ZV�k8p�"���]�꼩�Л�����5�;D��v���qJR���߾��)J}��┥'�{��@�JS�=���)=��Q���D���n݆qf	f�����(Hd�'�~���ԥ)�߿p┥'�g�}��UF��/3�}�e�[��ku�f�qJR��=��R���{��)O�Q%rO��߿hz��n�\[���d�ЕU�Q55�R������ÊR��^{���)O��\R�)!�G�lJ�#0L��BtYjq@@w���kf���� y���|���R����Q~��WRv���	f	a��߾��)@~%����qJR��w[>�콪�������2�jX��U�.B�k9��đYv]����D#��ө��Q�š����(ص=�Bb�9���)O��\R����~��ԥ)���È*R�>���pz��<��?��X�l�G�n`�`�����=J ���{�)JP��}��R���w��
R��|�F_ovn��k2ެַ��R���~��)J���=B���{��)JR}�}��R���/��7oV��V�����R��!�y~���R���~��R�����pz��� �����R����o�͒�����nݦqf	f����0�(�(	��~���R���߸qJR��~��R��y���-�G|������(5���@�VK�ٝ:L2��i	I���IbJ�!2�7lS�
��]iC��(@��%NE�+s����\�!�ptb>u�^�К
fF:@�'�
h�{ΈM�FXl�;�	
V`n5�̍� ]�]X����\�gf_����Ҷ�ht�����m���-��l��	�`$�-�: 3��zIl�GdЭ��ois���KJvy�y�Z�/�w[||u)Wc��xm͖l豸݄�tq�흺��܍e�i:kW��x�6�H�q���n�GF���hnɻ��y�dr��Pu>W�v�3::�M���s6ձԀF-v9�v��q���0Aչ���nnФ͑�Li;{n�W�qu�Fk�� ��{u�pm��}�x�=/Ip�}�@��]m���=x�l�I`�'�oY\=��ټ�A`GJ��dQ�s<�ۙ��{�u�+֠�#U��7�:�.e�/1�r�U^+μ�-��nC��&�.�<2%x��n�][(�]D�6,�nW#U�<Pct�kvl��%�⇅���llt�t�2O\�&N�(&*�ۡ�sKg�Lx;<���<2�r���	ے�rF4�����n��ҕ��F(:
�[X܀���6�3�n��/Ml��D�8��Sq�a�����q��h;.�G�����w]<��[b�!���ˮ�v�b���/\�1�.�e@L܁�GP[r�JN��|�wk�v[�X�-T=)z�����\�5��!.�$��J�T��G���qLq�璕5�p�Y>>po�<o}�ܓ�.�g�z�˃��l��]��2�H[�O'D;ܱڮܘ�D��r+"YK[�7j�F�yŜ�Y�'��v��cp=�L�b�j���R��m��2k��)��M��xv��1����-�9�˱��@9�P��Y�GU\ѱ��8��;�gy�B�&;m�Z������H+Z���� Wl-���w�6�`d�s�:e��v1t���5�J��F;cZ6CjP�K��l宱��n.7v,r��K��p��ݦ�H�[[��P���x�[I�On�;�v����[��"���@^)o]�������"}�/��7j tⴚy��ԫ��ؼ.ݫ���igeZ�ج��5�Gn���]�vix�u��54P.�&��b�t��i�mi�93730����`�w�!����(~D=���"����_@��EOa^u��KӹW�65���އl�c�3;&}�����k.����[�s�����j�f�����c3l�u�-�-�����C���kc����u�]I���������Ҽ��e�>�+jķ<��n�ui�qv�<�Dv�[Q�p�벎��)��,)��4Q����k��Ý�Mm�W>"Й�_�w�"}��mi���B{v���k�1�S��'k�30� oߌ>ƻ'�v��7O��..��a���i���#V۠�Fܷ��}���c�~g]�y��F����)JR~��pz��>�߸qJR��~���R���{��)Y�X~;�/���b��J��3�0K0��w��?����}��ԥ)�߷�┥'�}��� )K߽���Y+Q����n`�`����ߴ�,�%>���qJAZN���=JR�y����%�%�WOѶ~��)�����3�JP�����);�߾��)J{��┊�~����)O=�e��m֢��f��ow�);�߾��)@����┥~����)N��\����ߏ�4+lE�i'*������Pl�����q�6=�V�+v;IN���o���?-(�C�F�nK�qf	f{��n`�({�߾��)Jw�����D���ﻳ =�q�R�%CTT�SE�}���g��fe*(��Se!�V*fAJ��%����Y!R` �+I%2��L�D����L�-�X�V`�[��z�,l�h��x�4	�p�>�t��'�� >�4��Q4�t��M��f*�s�Գ ^�E�}����=�T��(�Ю��ݷ��4X?۩^��E���Y�c7���oà"�O�7]\��Y�r�f�a9�{�*z��֞���gJ��ݧ�}s-�����,�j�崋�Ա�� �m# ����"��c�T]�[y�����8n���i��W��3�i�US��h�Co ��M�;���~�V;�C�;�K��4����U`n�fUDP4H�UDL�`s4;;3�Wŀy.�����L;���y%v �	��KTEHUKASE�{۵`3���ڰ>ޓt�8`�K_�&U�]ZV�1]˺5L�<�
y8���"q�ey��$]�#>��ߏ{��+yV7CBUn�����hӣ�>�I�{�2���t��u��D۱�e�۫i����n�T�p���f�}:<�TT��j5t&��v���}�� �ڕ���UX{R� KdT�J[F�V�eZ��f`�}���x���߷ʻ�߾�����	b*q6����U�xg���Z��n�"�*��媬wffxfojZ�� �ڕ�۵�*��b�b �5\���Xض-`�(��F���M��7<nv{'��
xZb�B��n����>�I�{�0�t�U��������4[v�m���U��>��=#�=�I�~��IR�5N�Ҧ�[�� ��U��U`��{�K0�H�3}	7Nեc���i�hUG�G�{�t�p����:f��뾉�n�-�*����=�K0aٟ��,˗^ OH���S���w��N��	��w��J�w���θ|�ʰW]�v{)��w\���q�&ywG6Ka1�0�hy��4Ms�=`��Ju�"��ع�	8�W�C�i����3��m��2nՖ��/��]�p�`ʘ�Y]��ݭ����f�$�Ì�[<u���Żf�Grr�.4�'k���2��'����{v۱�f2��l���H��t�	-�$䷍"Iҏ�>�a�\��n��Ub���Bx+������\�%��Z�����Kt3\\=�]�cO� c�h��
�-��]�ė����Z��W��U�����Y��ji��Bn��m�I��N���<��3 [��ww`>��0���5T0Awwx�J�o����7v�`j�zw8Zb�B��t���x��W��� ��E�}�U����|��~�%�ECM3UY�n�"��fyݥٝ��˗_�=��`{|�`��,�^�\0	�5�ۭ�Mc�k�ɝ��zk%��:�S�t),����a�eb[MyaStVB*&� �V���U`{|�3���>����%�7Nեn��=��f�}>�|�؈u ��>V N*�6�`ʑ`%�󙙡��ݙ�ۗs�6��e�۲۶�'n�;�,ݝ݌��U��U���hUS-UQU1SQU�����_��� ���~��_�{�7@'��N�ui�mݴ��m�$z=#�=�t�w8`���S*me+j˻t't��6܉�ɹ�]���޻3�(��$q�UhP�ZfUE�ԛ .�bx�zG�NN����P��=���L�t��4�V��U���fs�;�4�q`to.� �(�~����(ݥE�um��;�˕^���s��t@ҁm0Bg��0F���fI�#]��,*�Ͼ�*��~�����})~wN��ҫv��_�PozL�	��{��US�K�'�|K��i%n��=��f�OH�Uu_��tπ�Z��3|����s�ES/A2��hŬ#�8�=)S��Ѷ�C�y�G�b�M���i��BcLi]�m�ӧ���K���g��Z=#�$=gU��ն��D�V`gT[�8�� >IU����������i~���qV��AKesQ`w���X;��/%����M�Q(�����������ϒU`}�K0����3K�;A� ����t+�Z�x�w.�`�J��X��j��)�i��ݬ��S����n�7E��8įpe�bL�m��n��s3v̚�U�����۽I~R�,7�^ |��wg`>�j� L(���AREL�T�E�f�+�ݝ��%V��Y�nΨ�wgfq�٠;���"f&��������wuXo�f��˥�}�3@���D�h�;�UUX3�9����7gTX�o�J�y'�Hz��J"�1ڻb��@��^ ;;6�� ����Y�[��G�����V8�a�E����[.��c���������w9g��� ����'Z�q�&�GZ��N8���^��o��Nd�t]<�C��0L�gs�M�Sp���2>8�ec���Vۊ�:��`"�\�PY,��3�6s<����\��rM)��������ÎN��P0 ����|�U��}�8�V��{nM�bɍ�4��:�U�g_���#��n�9A]���#��V�Z�\=ndӸ�y����xg�_�w�ظ.��)�UQ`�{� >IU����fv�7g��r��R�-6�Wwwy��3@>�U��o�f�:��3|���4A�&[�� $���**j�-��vuE��P}ޓ4�#�;�r��1�K���ݷgTX��� �%V�;3��]��t.iz����������/%x�3$���-Y�l{T�%�md7Iӝ5��h�l�쳓�;�7@��ӷ66:$�ʥ��7h��dA�~%����j�|�f��Sl��^J����m �Н�o �N���_�( �e�lll�,�)
,�"�"i�H��A�� �Y��\(��������(4�.$`,ceHDET4l�@�Rb�"	%�����-,b̑�J@��lD�18��=�����E���;���[3~C�}E��M�i]����}�`�%xs�0�����;yv`�R�4�;I�cM`�I����Ӧ�UU]}�`�]z��[m�]��]����J��������67T��I�ܹZ*Ԡ�wL��V�X'�R�ֿ����<pscE�ca"��J"���Bbrs3�v�X:`���$i�����t��o��vwl䕵��{e�0��ot��wt��&V>��9� ��K�_ߣ�\EU��*l�]x�+k!��a�."Z fǃ�$�9x�!�9ǉJŒ�	9e3TF8d���p����W��%v���#�0����5!�xsh�V]�TkƂ�E	� �Y�n �&g��`h�mL�r�۱��т��	gz�˨Cl�e\�;�7N��f&���U �(�����n��Mkm!����"��9����Xf�,қ6�im�U��UaYu��X%bf4�ŉ$�1�b�l��=J�xs��^%4�����gx�2PS��t���)���s옱	����hfg7D�C���9��Łgq�0L�3�hL.���X:\0"��c��bK1U��@�T	�uۚ�Cu݇y��VQ@X1�������r��rj�1�/:3|8Z�lT��*`z�pTODN�T��6#��
�(�P�]"���3��L�E��0������T���ݧ�c��?~�I��w�M�:���	�����M6�!����0	�՘��� [�W�|�"�_z ���&��.8�iK]pt%��`m<�Ղ�,��/l2u��͝ɱ~9�}���֢v����9J]8�.���������	�E�S�i���t��X;�f���I�_tX�W���m�����������%�p�(K� ?��٠{ʎ��X ��h�l�a|��cuM�-�W������3! ���
�LLw����$�(v��V����@�� *�;�hH�wӦ�_��*��v��m����v	q��'�S���Hݎ�]�R9�Ʒ*[�,�ʖ�+pd�&~�o/j����f����ߔ2OLЮՎ�OZǙ�}#��N��u�E���Pz��mX5Bv1*f��7@�� :{�htp�%BY��
bv������	s�����ޫ��%M:VէM���%�tz}9� ��n��� ���������K�:�*j�vȝ/�����'������b�]���GU���M�pm�Jq��nM��-���mpۤ�q�3=���m�wggN�^-��eJ1˵ը�Ӹ���c�1cy�ӼHL�S�}��l;;4,h���٪;�MT@8`�qn�X�fs�����cM���+�.�k����C���s,ۍuG�p=P�g9�S����b��z�6�$�9���.�8fJ�$*I��U�J�׎�s�Ah	�]��k�h�i�qn�5�w��� v���*�]��o��?���	=&��"�%�����]%wL,I��'�MҀ��<_wG�}˥����:�]�݅���tx�����<�tX��� �-!@TU]+v�m�_wG�}K�'�M��G�w�Ԕƕ�j�V&kǏ@�.��O���� ����і�]��N�wQ��t�t<\�a��w�Cdɝ҄k=����y�ՀY��<���m��I����	}���]/ �K8���\q�ܷ�I/��봡�$,@���$44�L�L�H  �ҋ!��3�{���K�'Ӧ�=G)ISM��ui7�K�tzyIx��N����?��_��;m�Pm�v��_33�(�՘���;���ｵ�	C(�;+`+J�n�	���������R^+��e�˧h_��7C���֧^.����u��,�,�d��x:8�%�{&�w�
�~�C*��7ai�ztx��G�w����I���:*�%V�M���=�R^>�n�{�<�q\����[�L׏��)/ �}��upԁ&��N�K���������˒�WCUv®�Ӽ}$� �tx��@����uJ���g��-'����	}���)/ �I7@�IE��;�v��-Zmؘ�e3�{)t��]�vM��e޳�W���ۙv�Cu�i���c�I�_wG�}�K�'�M�wG�K��D�m�`��ym��>�%��&����%�tz�u#�P�Ղ�6� �I7@=�/���>�%�ޮ��N�Wv&��0۪��V��Q`;�fgN��.����*���o �����Ix�t� �tx}:�Z�*�;v9뺰�Ԑ�Fڼ��t6��ˌ�]���[��Wm��e�p�%*�۷�.�)E���f {uW3;��@tv�V ���U0-1@�5T�X	n��fw���`tv�V��(�vx�777�P�7B�M�wO�K���yIx��t�R�*i���c����~�������F�M����wv�Ժ���X�"�j@���*��R��߹.����`(^J��ٚ��wx��RI�	P��_[��0�j�fQX���r�vL��Z�6�\�c��v�Rrq��y���32��(�A�}��O������H��rr����y)�c�\ˉ�ٮ-��������/@����p�k��3�S��\����&�rLkg�3]���h"��N�:�F賺e݅��쬛6ݡ�n��i��u�d�ms�۔���	Y���:�U��%��D�U䖦�3f,����s3�d�;@Z�8\t��ŉڬ��Xѭ㗇r3�n|gg�(u\=�c�����K� =�U`(^J���M�����PwN�"�7E���tx�����E�I�7@<8��T�j���o �=#�>��`wM�wG�mz�Nڢ�4f��z��,N���V�������X�鞊i�
�-�
�M`wM�wG��I���,gT*];�ۻN��]7Nݴ����AN��f��a�;�e㛃�95����q�]T�[tX�ot���}�f�����;��.� �h]DKM9EQ-5V�jW���3<;��{���jɰ3�՚���	~����m���Vf[�� �R�/j�9���� Ժ��W^ z_F��Z�J�Sv��'Ӧ�wG���4�#�;��k�l�iP��t�=�� '{�h�G�I��I���2��V�)�G+U9������<��p՘MWn1v���ǜ�;kn��zWj���o $�L��� ��7@;��B]�i�-STU���34?��~�]6v�� �j� K�^��L����M]&��$��U[��
Q)E�G��?{��:������wgTm���;�����s�U�wou�B�6[�0y�UDL�w`��Zo $���}s��$� ��;%1�B�ݟ��Ʈ��<k���8^�\U��=ETPz��ܙ�����u`*�2���>��`Ӧ��E��&h�IEe$;�"ݶ�	��t	s��	ޓ4	~�`�wZ���hE�n�����w��9��:7�l�]��(TKT�*wm5��&h�"�'�M���A�B��m�k���Uߞ^��TT��,4Md]U� ��M�����˾���lo���7b/EPC���.�v��n1ڕ�V��8T��{l�tn���Ȣ�J�WE:�M*M5�ON��K� N���K�Жtn��&�wM����`�I���`Ӗg3��@v��������
���j,��^��M��� �T�F�&0�ӫ(T��f��,Ӻn��0��f�{ܒ��J� �V��݁庳 �T� ߒW�IU���w2���|B�$�u}N���a�Dŉb�����CD�(zI�!	<�A����b	�J�.fR%�v�ބ6i^Gh����3��[��Pp�rZ0� 0Z�t����8 M�H2�>��Vꪀ���Z�੶oU��� pn�)�����0I�v%��\e�s�X0�@�Ү�g`O=Nܐ[gJ2m��[��@���3�ɫN�&�f���@gv�8�:���Z��Aېv��C	�F��-r�jS��նNa��m�����-����[�ٰ�Y�L�jvnۃ����a�r��`v�F��R�7l�bUH�z�G���������K�t��tl#A�Z��7d��m�8�c=����a��aۓ�[X�j����Dv<0:�l����(��˧�s�ۺ�Nt�=�������܇L���':�b�N�ۆٷM�����XrO*qؠ�M�.{�eʑi�ض) P�cE�F���9��%�2����R�h;Wb �Y�n����{�c��ڬ��t�dX&#��:��]��My�v�y����L�ޣN����z;xzD�pG��ݞ��AY��+s�溉yYb�/hn�H6�B�}>pN�C��6��r���g��Z�>�m�x���L����ΰ�'���if� /3yVK��QwVMַ���sv�N|�Xx݊H�]'g��9ص�X{��h�+n�)}�۸v3�^��'C���v�����NjOg,��%�.6& ��s�dB3�J˽�͹�m��F6�3Κ���іZ���	����Nz�ۨ&6��c8���%�Ѵn4Kn�j�#�<䍠8�eU�F�Ar�fݻs�^�i��;�(�y6;tD��F��d��T�-gl��m�Tb�C�W�#E�A��U,�6�^u��l =�c�	��+[��$� ��M�'X8ݻ8�����N��G�uҮ�����m-���v�p�,5��{��Иh7�$O���� (^���<]��3�ֻ[F6�؍��yZq���^RV��-ISyÚu�%e[��θ�W5N�p�D��J[;B����j��"�tF�-;Zߨ�m]�b�)�S�zC@��>
�M��C�*v �j���:S� �M�� �SޞV*�Z��� ��JZ�`�-JGgTug*O`��{Z-���Q����r�Dz�K��c�b�q��v$C�^c�n��+��k��%�����kU�;���a����k;����5ME�sf�0�(�]��#)���V�;v�����g9�)�]�:;j`��Ύ���+��=�q�X��G���nf��6Ҽ�6x���i	�m"�ZR�(�R�>�`��}îæ�p��-�ո^gm�h�5%� E�v玹s�jy���[hs�UQ5K ^T� ߒW�IW;3>@o%ـ�@��KT�KUUUE�o�+�$����Y�n�E�3�D�qU-RMd]U� owU�庳 �0��f���I\J�V� Hi���n��8`zt� �#�:΃m�t��.����p����G�zzM�>����Q��C����ks�m4GP��5�rA�=�s�������qn������:Ɲ�xޝ3@5%V���gf�t�E��4k��j�AkuۻĒ����i���j��7@�)/ ;Ӧh{�QU�V�۫v�x��n��Ix�N��$x}]֪�:Le�m���:����t� �H�Ot� �ʒ튚�T6ݴ� wӦh\�`��_tX�,%5wb�
J�7tݴ3�:v�ٝ�r[֒:H��g;E1�v��=�1B�T���7��}rE�z{��}�3;;>@ܺ���陖�&�BZjjl/j��fvvh�B]6 �˯ �$� ���i]14˰��@���7���wg����IM�庳 '��mՎ�cBM`}:f�����n�����u/�&�X]]��Y���$X�I�wL� �I3@�J�]5L���ݲ�+M�h���:���Pp�yՅ�%u(��4g�n̤�)0T�SU8���wU��o�+�>�"�;��ʉN��0n�bOt�V���� �w^ {����jY�a@Ж˧J�&�v�`zI��$X�I�wL���Wq���Mi��wx���ywf����3���?��M6N��h�IT�	��à}���%���dj��q(F��=:M�;�e`zI��$X�{�i��%E��DF��-jIm�Ùx��Ջ�`'�,��[�OlYܛ��:�FRi�`���$��Xޒf�����n�OW"7i��Cn����vh�ЗM���� �gTXkK�t������b���>��I&�r�x�$� ��(��� 
i������)]�����S`o����J�*R�kr�.�>��%��K���=	t�I,�!���
�����XMg"�xh �D<�1�4��>��5�]���:��eƶ������֝��nZ���0����\ZQ]U�Ų���Lv�rW'kթ�4����N2�����3�#�Sq���{stn��P�p&9��X�l����L=�x�&��Okhb8˗�F�p�6�.N'^�s���3Tݘ��Hpv,��k�Iij�|fa@pո�l�x�Ovf6֗��k���Jn�!v�<�-�c��
O�&wd�jx����-��~��3@����=$��@��K�>������%�B&�*�� �7T�3;�˻0)]�I^sD�S��5U5D�����v`l�>w�>�U`}	)�=]�ZV��֕���^����f����wM�	+�F�2�j���;���4�H�wt��t�w������'XN�z	H���ܮ��nK��`��yE
��n+ͤ�5Kh�cn�ͻ��IM��� ݝQ�� -�׀ޞ��&f)�i�!�*����Y�=;�43c3�8�A�8��3���%7�����/2��UE1QU5�R���:f���,~Q,�0��Q54�Qa��������=�6�w.��}'
�&�-SAv���]�BJl�g��%ـ%+��3�U�%����S���G�X�EZ��F�N:X��ӷc&̷@��}�iNy��v�V��<ں,mh�۠w.�����$XB_A����;m�ܺE�;���׀z;�l}�Y�	6���1��hb�� 7��4�H�_`H�F ��P6�����`Һ,�֗�e5R���Mw7wx�$X��M�;�K��t� �\J�@Rh�[o ���t����/�g�˯ =��`&�cT�MT�AS35�%����{��.�rp���	�dV;q���ɒ�j��m:(lm[{�w.���I��$X�wM���qQ��tZT�Q`����� �wt��0��x�p��m"�4i�����,ﻦ�˥���f�$j;V+��tYv��ﻦ�����t�/���Q�@�W_{�}����}�l��:N������x�W��ܺ�l�E��jY�yk(h�*
�`jɘ����mn˷&]uRd{-W��s��^6�ȼ�R�)-�U`�%���z�]����ܤ�~�7@�.��}rR�Dګ��u��34�Ix��n��]/ >��f�}���DP�.����I��t� ���ܤ���9T�`�`�է��t� ���ܒ�vwh�˻� o1�2:�����j��� }�t��^��7@��E�z"�JC �1A���2��I^����B�HwGVs��c�jyg���o,&�!��vK�om��Gk����,��]ڶۧohq���`ɨo%�[��8�gW͜vLm�g�;q�5»�7F�|s��*���B�;]D�u�h��>�y%�Z�gh����Rú�v 1K�K��-q.���#h�s��6�Q%�������Zn�g�;dMIk�Z��^ha�b'��?[p�n��F��䬔k���x�1�\ ����2��ö�@�&$-��^,��=K�7�M�:�"���f�=��Z�m]��{���� }��4	�����D�V���t�	���tX�zL�'�K�>�I�Һ�n�6�I&�����f��:��o�[ݘF���O�.���M]]]]㷙���x��7@�� >�I����H�;tP���C�v5�rBs�6�f��i��N^���k���sD��6
�x�t��K� >���yIxz��R���o�M�է���k���L���*`�3�: >H �B��=�u��L�%���&�}GY�j���7M6��zL�%���>���_tX}8Wq;b�J�X��ffh�"�>���\�`��L�'u�ҫ@5USA5S`gږ`���<�p۫� P�M�����̆��*(�����B+�;��%uU�7CɊHZ%\���j�B�D��n���Ӥ�m?�������K��t��+��5N��V�Zk >��f����7�t	~�`\�)~�ЛWWWWx��_tX��}�V����$!ᙛ	����A	%&�ݫ3#v�CF�mYo&5d�a�1`Qb�.A�ƃ�Bd�WG��2g�^��$���3)0�c*J��DK�t��Ł�2&	�1�aF`�M@w����ֆ����`N�N�Ԏ)H���	� Ma2�1�ht��4
�b"ǉ�����2k1ބs[�-�[��!
.�0�Ma�oF�X�68`�fcZ��1 a��0���	&t2$ֳq,�8]�!�x�l�֎��p4�PR���B�T�u��t`c�Ȫ��23 ��S��r+�U���2�r29p2�JX$E�X#�`��bOAI����6��܇�x%^.�D$H��L�j��L�o��� `[�h�1�-c�"u�`D˨�V��&�f�;T�����bIiR@a`�"(lN()�;���ؠ��� ��t�� ��#;��̮��yj� �F̴�"�
;-�k�t��K�E�{�3@�� 﫺�F;��
�=�%����Z���WM��� �l2h���j�e�B�wY��B8�����ݙ��g��1�cH��u�'��Χ�59��~�}��4	~��t	~�}8D)*bbd)��Ȼ��G�M�<A����?������3@�-�j�T5M���I��o�&���`��L�%���:�N��CE�����Ot	~��y��꯳�~�+�>���J��@��A�s z�t��~c��J�ݦ�t�զ����K�E�o�&���`ꄛuk����.S��r��@OXCד��	�9��eW��A��{<^���b��8>��h˥��I��tX���4�wʕ"0n�Z�i�x��n�/��}�j�zuE�;�@��S�D�UM UY�tj���W�(���3}&�|F�ӱ1't�k >�t�G��7�f3�J]6��1%T�L1LYuw�(�S`w�{����\���=��U����%�tR:ē����k�_k�޵��j�\؜n:��5n�Ӎ՜Y��vm��F<fx͔�jN6w55����՜�F��C����� �z�y��ok`$;��f0MiCX�'0c�&y�9�D� \u=Y]��ٝ��FK�z팴��i�ѻo)�m�=�.�4��p8�|㵁�OnÙ��(�n6����m��N�;@i�&��-s�e�9���W�+��S�,v���?a�f���L��%�u;J�6�܆�8�fvKn�nTN�n6�`_\{k�%"���)TҺ,��\�t�^� �}��������s��v��m������L�%�E�o�&�t�Jm!S�V�4� }�j�y+k9��#˗fЗM�FηHq-�5R���qUw��v�cX]ݺ���$� �]�J����U2LM5��If�)t���y+mIw����B��akM	ʱ7D�u���T&vn�4C/q���m��/0@S�W]=L�TTUU���6�I^ ���;�]ݘ �ꖉ�ij��j���}��s����l%T���J"� A!���#Q)!��@:փL\YMX��K:d��@#0P�ia�x8��\$0L3j��4�8��}�s�X���_tX{�Q[�����ř���Xt�t	}�`�J��P�Xxj���b��kgfwwxK���:�$���[X���6� ���7i�/�, ��3@��+ �I7@��uj��j�I]
�0��Ч�qjM��'��핍�vݗv�U�����hLmRL-[j�6� zt��N�+ �I7@��,��_QR��l���o3@�&Vޒn�/�X��f�z]�J��;������XzI����\���G�����~��U��+ 﫺�MSi�Nݺv��� =:L�$�+ �I7@+�2d�������� �ԯ �f~��lowf �ڦ�^݀TĄL0AAG"���=�y���cb`�֬��C;z�x�hLC�v�J�v	����z8`�M�%�E߶����t�-�?*j����-3 �n�9t� ��3@��J%�`�[TЛ��@�� zt��OG�n�w�
�wI:��v��M`mW�wM�z8`t�t=U_|A�L$��VX���6o�rjK���_�?�`�7�����H�#�I}�
=�l۩^��߿��+߮����vs�hܷ &:����\71�k��e�V�)�ovm<�p��]�ݢ{��������y)�n��@rUŀ�R_�MSi�N���_�X�$�wL���w�Uv���H�Z�I[ �$��Θ������{���j�+e��{x�3@��I&��"��L�$�b�����\4X�Y�/JQ`�W�-�G;e&��0�)$?}��������+����\�v�ݎ�)0=�����:v�M��PVHtg5�g��5l��vjM��jLtu5���㥰����Zz��h��0/lhn�޵὘�/g�+�y7%rd�g���[TX&�i/4q�F���l����S��)rz�'v`��p�c���km�!�(���Y.]p�h��`ʽю�H�68D��[of�8J�%��;S�`ݑ�)U�.5k%>�f�z�c��m�4�z��X�W ���;k:�"bzsi���m�������L�'s��I�_qV��v[e]�m� t�f�;�0�&�˥�����*�m6�.��-��{�0��t	~�Ӥ� �]Ĩ���P�2LL�����]��ѫ�`�I��8`z��ӫCi�-�-=�%���t�4	:e`�&�%�~���/�T�*�bu�Q�ڼ�c��]���Iݣr�ѷK؝f�=2��n̆�i&������ ��׀%������ �t�{�T�[UhL��=�Y��I�p�j�
�����못�_}x�f�$jQH����u�{RY�(Z��g�5wu�˭�A�l����"(�&j&�����M�j���$镀{����r�Q��[N��6��t�4	�2�t�t	}�`���{��� �𓮵\��%JIj�qX�^Q�>5�p��4����<�����}���[EMECwW��m`{RY�-����&h��%B�c�I
էX�I�����$�zL���)Ӥ�Lۦ�Ot	˥��I���y���xAly�	��9
�� ����_s�A��Y�����((����� ��f�=&V�I����{�T�]KD�T�5�Swx�V�;�.���)�x�I���T���ںN��g��ڻl��jv�b�ׁ"�9ii�n���v��M�P�����]�� �$�r�x�I���X@�Juv����*k0��/��� wu����I&��U]���X���M;n���k Q��X�V���`
5)�6>hmeq��m]]][�O�:L���t�(�٭���gq٘��� ^���Q_��B�� �$�E%�I&hI��J��O�m2�j���$]� eĦ��r��I�;Wc�7.�6�z�l�L�j�&ڷn�N���)/ :I3@�L���t����#i[�wI�w�$��I&V�I������յV�5e�{mff�'L���t�v��Uŀ�����U�!RT�4�SMa��_`��`l$�`s�����Dw54D�4�$QSY�j�E���U�j�m`j�Y�Mlڡ�>c{3x��8[��ȣ�ef�y���"#�l�f�ݏR��K䞝łx_y{� ��4�dI��s\i`c�g=OB"!����a�kG���E��3f�k�pN=���2nhb0�6�5�%L����+���U��=��PY��WjƁf���ǻ��Iôz|�3|ݜ�<�F;te҆D��|va��0m��B;��|4A�O�IT� �|����W%:��Ù�1�N�` 3�DaD1	jȈV`��A@%1�\�a����.��p�V&�{��[K$��ڐ�[FٻslH� �8v��[ז�M� �N��M��l���f�|dQ<kV��isv�R��24���Jiz*Z�h��e �9�{lI��Z��*Mζ��C	��۫�X�GC2����b��;���`s��ǎL��B�8`t5�%�;9-�r�6��!f�u�sӅ"4/U�ћ�,6D%{=	4��ې�֧�81	�
�e�q���K�%c��Y�R�:�=sp��:Z�[Mi9�c�u��=���������ɯJ��t�[AqyډjҝZ�V�lk۶��X
�I�g�;�����P[u�x;�ru[�[��/E��`���Ӳ�:���khS�ݹ�u:{{1٫pƶt�ĝ۞�7k�P�N�e��1!�&����۲M��:��1������.!Kri9�ƣ�㍘=$��1;oNSap�i��˓��i
򍹈�V�Ԗ�v筳��m�G;]�۳�J���]f�� Nzq�d	�v�:s��l��7D�Rqu�e���;E�wk�v��=�D/[���t�o66m\6�oC�n,9��OmC舝�	��jj�U���'	��[�C�n��ا��+΍�1u��$qF"���ۤ�9�C��*q�V�Ͳݡ�]g�;����YX�Om�in�'C�w>�#�1��Yk�Q"L��;���Z0�rɧ�����,K��ũ�ɯ�E�#���a5�F��U:ɻmk��>�l���6�uLn��.�C�&'m; �ʗ<�mP ,�:gl�\S���#+���v�nt�{t����qs�������"VHi$�n %�ĉ:��Iݮod��sm�@�]Ė袠��)qQ2���^����y{]����u���˸���uY�u�G6�W��
M]G3�MF��Ѯ��n���B ]�lh3�g!�C�3p�88�s\NG�N]0[�ױ4��n��t��/�XDI�^��U�V�Ol����e3K�H���.���k��@�������it�g���Ѧ����{���{�@�A ����~�*v/���/e�`���z�����p�d�3g�r�Z��鹱��e�ݡ9���1��u�R���t�K��ivVl�t\�;�f���W��-�H�nhG!*6��5�'#v��{rZ:P�5Q�#��4 m�]���u��$�!;MnA�[��]����mۺ|r���Gil�v����P��n}�ø�P��q�E:�4���|�\\�nh�ZH����z�షs��*i�H�9��k��]Ī���p�Y����u1��Z�pGH�f�����nN�a�C��ui���ݷNҴ� ��H��2���Np�:�W�$`��Ε�����2���Np�:�= ���ڈb�v+�XOj�R�Y���
;WV �����7�T��m�v�	�M��8`Ot���XOt� ����������&� ��W�s;��.���j��5%mi/�0=������B�T����{�N�IƜ�nբ�θCj�萺䧺�$yn�TD�T�5�T���.��5{V`	*G3�d �˯ 䢺��Z��������ڳ<��;=㳴;�P+J������E�z��)�ڰ�cE���wL��{��%�E�t�M�:]Z��i�mҶـu�tz�H����p�:�W�$t�jdM�`
<���w��WE�����K���/�l��)-�"�\��Q�ŭ����`K����X7m�k�p��vyh�ʃz��`����v��l�����fg�:t�[{�)����**&����'G�{��%� �N���}tF�Ӻ��6`��k@�$Xx�T%0b!�Ͼ����_}���K���:XՂ�4�Q�É`a��wt�yv`	*E���h��J�%�S�uvZM��:n�:8`�r^�/�Xz��t���Jն6��qX�kn2�B]����n^p��m^�˭q�vv�	ӫ����է���zy�z��`��t��W�v�uv�:,/RQ����B�o.�)J,_U�	n�*E�e�� ��M�$R^�����BB��SX����N��H������6�� ��~��jK����)m�ښ��ot	��{��^�.H���t����I�ܖ�+E�4�i:�y뮔��ʝ�y�5�&�"�6��/Ϯ;|Go��;17Cn���\�`Ӧ�)/ ��-TWv+�s/@褼}:n��Ix����	��v*5N���Zn���E%���K�:)/ �N*�E�V�i�դ�@�^>����tX��n�I|Y�I46��	6`�}/@�����������@�s��WK�r���IS��Ҡ��);m��1rJ3�Q�:#�:�J��ml��K�;�q��n�q؎ш�s��}��`>��=G���s���p�q�9Ŷ�\��6M�b��T큸�[)+�v���Z.��e��v[�v�i�ΰF�x��U�ga�;x	m�l���^7m�p�尻c"���|����
��[��]\��V�^�C�V��f�<�ʆ��G33�fa�պ�����EK.�6������ծs�nU��q1G��B�1�8(75:#v�[J�Hq���������������s�z�������N���k �zM�>���}ϥ���~��30���>�������ڲ�����`}�֨�6=�l��� o1,��C
i�-3 ��r^�]��,�����>���<j�+��Wl�����ޓt��x�y�����g�~��H���PQW!iU��W��nz�<���c�r{l��ƻ�S�V��vj����M5�}:n��]/ �������@(��`kr;�� i����"�k����}�s2�=(��Be��$)!�C �e��ai2I%@��%
!����"C�LSvo�y��K� �����(����V�	LT�Xo�р(�Sg;D|��0��苀tt;n�����4	}�`ޓt	�%�w�!�]\�I
3�ӻ�4��7�&��K�>�>��K�MIw��C�a[qXAV��T��u;7l�T�	p�ٔ�o#��<7�F�� )�릕N�ݵi��>�K�>�>��u� �����@��'V��ۼ���z_H��I��%�8:�@MQ�34�q�(Ԧ���Y�5�ߛ`0�U_ eU�ݘ��{����Z� �ڕPK,Һ,m`Q��7@�0�ϥ��E�z�rS��I�wm'���}�>���x��n�zu���U5�90#���P��V(z8���:Cc�f2Xˎ�z,gn8����F��E�ne
��s��t� �ޓt	�K�>��Ll�bj��$���F���ݚ�I��8`}������G7��]�m`��t	�p�>��C@��S`o�ڤ�
������"j� wwgu�X}�р(���N�vgwf�vww�n�W�J��ګ������}�L���� �ޓt�8`�J��T'l]�ytGs�zx��o�a6]lʻEА��	^(�\3��+5	��ԒBYt��6��Y�|�����]��{��lt t�~�I��������wM���U~�rX�X��M��i=�>��}�t��:�"�7ޓt,��BN�N�BM�ߪ�ޓ���ot��%�:ݤX)!�,�M�����	~�`�I��p�>��mh��s����!�5v�@j��rD�<�5�66� .N�V&�Ӷ��Ÿ�7!!�e"S�a�{X�=ON��F�I��9禹�����9q��&0�#\k��׆8�;������zz��!4%e]$n�t"+����}�n�r�8����.���˹݀�,;�hȨ���\3��pk\�;p��=�F<���'d.Si'i�鎽zI��$��*�7����fb3ɮ�!��:���;g�q�m�7������k��R�M�P:�v���y��F�AwTx�2�����_�����`[�����?C3���6��t�L6؁�6$���� ���_�M���9�� [�����$�i��&h�<��F /j�:#�ـv���ڜWZ�
�۲�WM�e��G�ozM�'�K�>�vC@���C��m��4���7@���K�>�vC@'t���߾s��AF���X���u��7t�x���:��N���tz{B�Ѯy�&�ݴ���K�>�vC@'tx���\	m�ݺI�i;�>�vC� ��,�HL�$R�R4��`�
��M�� ��M�'���}u+�T��aE���4wG�ozM�'���}�Ս�l6�UND�UUXs3����-���{���|�6 -�V�=.$��mX?��i��'���}�I��l$����K0wxn�G9MU%A�g��A'�Åmv�]S��c�jv���;.Q�Ak��FS[smuEa,�;^���߿�hrE�o�&���uN,����t�	]�m�hrE�o�&���}�t�ҿ~�����@��B�jն����T�[�C;7�o�a��$`cXW5�d�&İ�����2�:��p���8Y�cVYc0�9�flR�ɂ���ͲgV�����N6���p�\��+��a��ۤ��7-�ce�X��kz�n�Bi�$��a&���ֆ����	A�u�ݍ$�{у�a���J{�=�1���fa-�5f�<[`gV� aH��(�ZtDU%4g%9v�������qd&Hd$������3[=�W�!��by��;�&ӊ�=��m^
�C�^��BLAW�^�� ;@U�:@}P:A>��{��^�����R��J��&�ݴ����}�t��	�U�I����SE�mګM�i��zM� ���w��yIx��J�uunݎդU*lN����\�B3� �<roNp�9�x���۰��t5�[o�aB�y��N����n�<���>�I��u�Y.���P�m���zM�'���}ޓk@'tx�=.$��mX?��i��'���o�&֟����{�7@=R�D�jة6캨�3�K ��{V`ck�����`$(�߷MI~=���#-��$4��{��>��n�=�+ ��鵠t�t��N�]4���i�Z�#��U����&زg@�۱A�\j�H��Ԏ�l t�U�4�����Os���2=����(6
�j�n��Ot�_3�;�D�W� v��=�8�����JO���mpr��R^��|`���3�K0��СĲ��M+��k0�	�����N]/ ��솁�^��+)J�QE��o �y,�9���R��=� ��C�L`4f��m���-�U8Ղ+�J@6�mu�.��n��F7��E�g���q��e���t�۲9���� ����m�uųb�s�{FW"�+8CB�F�	Ӵgs�a�n�S�x5K��n4j�l����oe�.�n���(�Iną&sL��Y�ટ#���Xk/a�f�'7P��S�(������ˢ�m��kh��5@l�@�v&����TRԦfa�0�a��ո����G;�[�h�l�[�����:�*g��탠����uq�l�NqJ\U<F₯���~���x��!��>��j�M����n�n�	�vC@��>O.��z�_K��]]��7�h��`����X��!�z��6�5EI-�SSa������K��;{������n���h����j����*k�����_n�0�l����̊�t���j���������Ӯ�qm���ܝr�9<:���ױ�/f�c��h����,��T`�U`g۫9��ݛ�t�E���,(��"jjf ��"�� 7uU�٩����ڙ��m��<�+�7���.��t����E��o ߻���K�7�}/@;�x��q�m�)�i�m�褼{ݐ��>���WJ�j&��]$����솀wtx��n�<�����ߖ�M�N��X㝱�ݚ�}p���v�6ư���Q%`�J�4q	�22ȜI6� ���=&��K�;�솁�]pn�ʝ&�Ui7�l���߿]����W� -�W��{�4�M�DQU1SU�l�E��Z���;��������3���Vv�f �,�T�TCL�4�5U5���yẁ�������N���UR�M��WWCO+@'H�OI��%����A�~*�H[�u$�c�I�pF��d
�$U��=�;����ɸ��#�ڙ�\�*�i��OI��%��� �#�6$N�+m��J����')/?�� [���]�`yy,�v�2�fzjf�f�"�,��� Z�Y��ݘ)������i��h������٢9wU���ـ-���;��gvfd(%Y���>)}��Z�u��?*t�IU�6���7@��������=���Sihf)*�i�K�/Ei�pQ��cl�pFl��;�WI�v��vڻ����0�r^�N�����E�*�Ui:��n� ����	}�`=&���\_u*��E��B����2��6�%�s�4F��krW���u�4S`�����k ��7@����F34)��=�]4�5U#E[E������_H�����Iw>�X ~�0sm��G+pD��&&K�q��ctW=��s0m�@lth�ֶ��'
m���3�^�%ݔ��Au�hmɵ�z�t����O+.���������m��í�q�	�cs���V�'ډ𸤱�[�J���j��@o��8���s��L<�On�l#p��-v6�������Vx��[G �v����B=�ў�'=�d�,Ub�v{L���V!ڛ�י�ن톒&[kdN�:�x�u�X:��!����^7L=�@u�78pK��A؇Z$�Y*+#�'k�K���o��
S`j�Y���@wOtX	6��OC1CD��EEV6 �%7��or��;����Ӧց�]pn�ʝ&�Uj�m`���)/ �6�	rE�l;�W-��ͦ��&��#��:mh~�`���*��U�T�uui�vـ{�M�_�X�t�w8`�Ć�̠�I�M"Ք�V�h�kp-�����v#��=:K{/@��cJ"`���}�j\�ՃO+@'�x�t�w8`��k@루�h��E���o �N��ivhww�ٙ��H�5{V6 /j��vh��ot�EQEIOPEV`���=ӦրOtx�t� ��~I\b���
�,jՍ�ڪ���Y���گ�%�=-Q-QS1U��ڪ��Z� ^�E�"5F�l��&���k��ЇD�n�x�����-sق�g��6FkB������(�Oo=s"�\UX�]���,jՍ�� Z���:�WJ�ͫh�M��;ˆ�]��{�����='M�%®�.�n�um����ڵc`Z�����38��;34C���?����՟f`	N��{eԲa&ڤ��`���	:<�:n�"�ѫ�|��DT5KQ5V�j���ۺ�F��c`IU��|��F9ZN+�N��Tv
)�3�K���,p*��Dv�Xnʳ�WZ�H��lVF�հM�"��t鵠tx�t� �x��e���M��x�vC �V�j�)����$�b'�"e��%��f*�����%�0%����k@��pj�ɂe�Wh�݀��f�:����`s3�0���,�N-�t�詉x*�*H����=#�'�C@;�<N�_B+8|��<����2v�'d�ѥ�7f8���Wmb�d)v�ʷ��J��9mb��F'�����V[�9����r�,��_������!�ኛ� 7ڪ� ��ـ{�q`%�X��<�iURČC�v�x��Ӝ0	=�k@;�<}��lwJ��:M��>�� ��Z���=�t���!FX�v��f��mhwG�w�M�>��r�q�9`w����Bt���dɭfHsA!8�������������v"���ۉ�1`1�
�n���gaDPQB�`.�4 \ӝ��*�'��	U���\�!�[����{���f��ݢ3G����/ �/	��W�"flD���T��ذ�O1��������{����Cݷ��4��.�{�	�:�#�V,�X3�,��uaHQg3�$���^s<��*Lt�9q7K0�t������5-��pF�1����zObz�g��xLGR����шF��f X��q\�s�����Ab� ��[��PpkՃ[��1�����AA$B��bYa3��d�S�t�8!f$W��"p�ώu�����o\s~�Y�ZaÅ�.�I��P������>(0������L �k�]m
WW��;�tZ5D��f0�=���d9����Da�����h)j� �X��{M�1H1v�́C�p�)��?~Gn�Vݮ�j@5��n���v�Ӳ n��6����"� �Q$����K�b�%-�+�3�k��JV�
;t��U�n �4��)jB��=�cJ7l�d��p2��]kV*�gm�omJl�g^�퇛���6ƈ�6�c��ۈ�.��;��� `����.xݴ����Z1����ٷ�9�:$
�^""��r<ٹ������-�7k���7kp��si{$&wJ,�/W�K���<�3�/Zہ�e�c<��L�յ^(��%ֽ�'�M��Yh33���>�E��>Hٸ]��ځ���dL^�m�m&�؍�Nt ��'$W`�y�֊���574L ����q�a�ڼ��v�\r9���g��&uU���<��X���g����k�|6^�:U���D�8܎�VY����Y�<�h��lγ;��ۘ�S1��۷m�y�a:��,sN6
;��;n�0h��J�L����8�QٻaN;lk	�.ދn<a
ܽtxc�7 v�j�ʛn��lm���Yr*��w
BRnA1���u�mrŹ�6�N�ۭ�k]��=&�� %�o|�_k�EVUT��F���-��ܒ۞Ұ���������Gk5m�cXVۥ�.��9"�3'!٣�&��@�kn*]ۭ��;myKӣ���f#�$�kɂ��ԕ1�D��=�9���a��OOI�s\��g��lOoV�U��rJ���%޽5n:��(<�va��������][nQ�L�RmS�H��Ʀ������ր�sb�U�$�X�cv�cv�)�Cm��!4��#m�`����g�M�ӫ���h��(��X���<t��8�1�닃;�-��I�B�m�>]�y�w	�`n���q�c�7ۯA�ۗl��L�ok]���R鹁Cñ��b�۳��x��3����nƸK�\�k�m�҆X;9b���#A��fU%$	6#̹_\�
u�'3�=AKR-6Y	��#u�".Sn�u����N��
��'mDq��$����g�����(���D<E�
�GB�z�\Lڽ�Qz�b���ޞ:X	^�e8ۅ�XA��n�{z��j�5�֑�����׌Ӹܑ�vN�<�M뮘ئ�vW'����nh�ODn{m�تa4�I8�����Ǎ��kM�y�\�Mqq�@�Vێ;tMts5�$,��L���)�x�ӡ�y�pa��.�c'8�梞�`ع���gm�y;k��m�g;������OK�+5В;�QhՎ�%
ڈIM��� �f�k���y6N�7&��{[������ӱ�AW[MV�m۷7n�D�;��an�y��[`K���-Y�y*E��䱰�;�TSZe�Wh��ޝ7@�����������~Ct�ГotH�zzM� ����t	��˦�i�M66ـzzM� ����tH�m�/�T�6�h���O+@:H��t��p�==�kR^����[N�8�b���@���g}� �&s]�y������;�{v�jz{<5L�5X�.��R,/j����{�t�:i�Bt�OtI2��� ���NިbV�o��uU����`o�Vg;�;�4@&Ӟ`��������j����] �*�7�0n�,	<U�
�+t1RlV�և�ߤ�xӗf��"Ý��V�t`�Q'KM-i��]��x�:n��s�������=�ֿ]�t*)��~V�v4�}
�:�vt�,�ٺ��NN�X����>n�v8��Z�)1[��ot��0w�C@>����yv`r��&�*�j��bh�<�����K��[˳ �gT_33�B��8�&�F��xb���%�`}�Va�%�٦��#T�E���|`���Rڦ�TS�N�}Ӧ�r�,�h�[�� j]V���h�
��覝��ܺ^���h���t�_uq?;E;��U���7c�����P�n�2rG[�ø���r�ov7Z�y�j�I�Jۼ��%�_H��t������]��#��SLML�e\`ڣ�>��tr��w���}#�-Re:��ҫ�Zo �N��{����%��G�Ow�R�-U���am���+k��J0�*��voS�����߇F����~�޺��>g�[��4ؚu�{�� ���t�t�X�.��'e��h�~B��i~ƥ�Q�XTB��7Hj��+���aǬ
W��[�ɴS�������<�7@�+ �y�z��T�;Ct�t��M�jՙ��K��[]р$��^�IշN�N�E�;Ot�X��K��� ��M�W��H�M�T�t�u�{�� �H���n�ܤ���#��V�Wi�Ik��I����n�Q`|�IF�q�w�ggn�M�W!*c��bh�z!�m֟<L� �s[�ڷ���^�b踾s���%�t��`0����cY��<�C�����k���{;)gc�5���C�q��Enzv�:�J�50��]�ެ�Oh:��ɇ���GV�l�¥r۝�.n5��f�n�`�v]֔��i�g�im��}��w�N�"P�uQ	��kc�r�H��d�dU[-���E���0���a˳��HUH�rEr�S��˰7-f��Ѷ��G��Ý�nU�$��{j�0�x[�j�BM����M�;�����h�� ���D�j�5V�i��;�E�;�A�|`�uXo���w�:��QL��5D��X[�� y%V��7@�+ ۗP�%	��Ww��ww�Xo��wU��;;�G��t`�%��J��^�*���|�`�X��%��#�=_x�~��7Y{�������s�^�v.��q����s��;�n2
�iZi:-�-�N�4�{�{�� ��� �tx��7@��Oή5l�f�,����w*��7��ԦĐ���G�{�M�;�K�>�*�?J�l�5Q39W媬��f���g�,N�נ}ъZ�o�LiX�o ��&��%�w����=߹Gj	h�%��"f�3 �JQ`s;�$���;�<��7@�W2*j��v�M���M:t��Y:t1�m�M��βg5b��a�v2B�+������b��N���C@>�����w�K�6���U(i�n˻�� �tx��n��]/ �zd4	~�
��;L���v�x��n������$)fa���%h�$]iP��7�>���H��蓠�趐%n�Ot�8X�+F |�U�3�G�{��<��M�wlݶ�L�;ޙ �tx��n���}"�t�(�6��n줪��l�oa�Y�X4F5*aQ�f�6���Ӎ�E2��bn�Kp��� ��&���9��� <��� ��OD�E<�$�̓5V��9ݢ�tX[]рI=�R�݉
ڤ�X���Ix�����<�t��N_��-\U�UDMTXs�;;�n�� ���>��?b$h'�_]��`dt7tK&������p*�� <�xޒn�ܤ���%�EW%1���u��b���7l�k� GO �F�����o5㣑��;<�d�t=��5���zI�r��{����<��$���V�i�ܺ^�s���ʬ����w�<��MSS0QUS5M`n�� ��V�If��m`|�)�e�n�-yz���I�t��kwgwh]\�p���y��V�$Zo �:n��镀tS����ʾ%Ȕ��DP!JbX,@!a��~���HV�MF�r<4q�v�+�(l���n��l���6�1��Å��N<jL�۬�;I��kҌ�u��0��3҂m�y��ݕ�ح8�#��q��9��&��f�iW��,l��@M�h��������<���6�f�u�qG%l���XUҦՙ�m�����]��V�ܸ� ��>��y�9�i΢�m�Lhz9n��]�=�������{���]���i%˴f���9z�n��]0�*�v�DyX��qV{"m���R�E&��O�����n�_��ܻ0�麊�&�j���")�"�@;�<N��L��뮻$�Wm���P�3�w�x���8`/tZ��V�;�h��;��'�n���N}/@>� ��D��n�uj���i��s�"�@>� ��n���ܪRT��6���掮{[���&z���W�w뚻j�ټ�rAUn��V���e�m4�_tX��x}ݘ��e`����wc����ʫ� �R��ww�vyvwgf�M%��U�����h��atL�S��,L���U�ݽـ|��`%;�p|�`�8��4	][C��=�=9� JwT��*��v���� ].���&����i���- �H�	=&���K�x�e�#�閩*E�t��ވ�R\�0Z���m筜�m=��1�3���&r�4�ҿ�b�� �t�Ӛ; ;��NѰ������"`�(���Z�%ݢ-�X	JJp|�X���?��������Ӝ0	��.��dQx@�t}�-������<�]��C\��]bS�1>�`n9�=9�P����/L(��c��[,�'R�tv=�s���6թ�a^��A�.;�	1�1ٍ\xƖ#Q�
�"���h��ց��fMe��̲ɬ���{�� A)�� ��n� �µ�L��2����0c`�C<��%S�����Hi=��.�2CN��Ch0=��t�CFȐ<|Έ��,LҎJ�G4kZ���!����&fB�C���)	�څ��SW�=�%��4�
D����XD0>�y�O*�ʇ�Ţ
1���&��Nj5�Q2#wPh��!��Ksƀ�� �	�*�xh�����f2d1f�����%˙1r�����8�T�֑
.`=s�MPLn�&��.C���	�՗�������8J�E�At��z ����������z*h<Pڇ�����y�U���X'"�TISUT��a��IE�o��wyf3<o.ư<�CsOCTU�ww�ހ}�<�����+ �N��{��Wwn���S�7���e��a]]R�IΨx�ú\k��v�#'@�y"ڡ&�6��twL�E:����|�>Ԫ��']MM2$�ALQY�{�e`)׀��wt��H�uF6�ݷI�X�u�����&��X_�V)V�N����/@>Ԫ���Y�{v�a�����3��3J:��H	~%BB@��L3�3^�~z���s�+��dR�UU���Y�{v�`j��`�ڰ;;����I�b�I5X�#�J��c���%R�v�^Y�ٺn!K^̪��Wb�i�&����R�,^�X{v��ٟ 5r���9n5EU44UT��`j�i|���jU`j�ـ{v�|�������ꆊ*(�&��f2� ���:n��镀t�� �#�v����mQ3SUV�˾�5.��<�ZX{y����`�"���I����0/V��ݫ�j�;�����J��izC���c�q�)�ll0�>�cdM�j{t�ZM�jR��ju*]vKm��q����nlaau!�٨���r����B0X���{/V�.\ �B���F�ՑţwH��>"��aɶ�s�'�����}���3�qآZ��;V�N����1A���N� ƫ��]��|��ͻa�OVێ.p;\n�Cϔ��Q��[Wn�Yh�Fy5�٭�w����w�F����J���M')Zq ��p<]T�������
^��K��Ly�Th�6���>|�^ o�������X����\�6:b��x���G�{RY�y*E��wb���
#Z%CTLC��UT�X�v`�H�5Jذ{����џ�am
��ē��R,R�,�nՁ�Գ O��
�j��۴��tS� >�s�=�&����5%��>���&���W���IeUbtqR!BƱR��)a	��1�m�ۭ�3��Ph�B��In;�t� �I7@�I��t^��>�{�T�J�[�&�m���� �!04T̲1I
��/=���Ͻ߷*��ݫ��S��	�����jk������� }��zN��tUķm��i:i�f��� }��zN��{��/�U�Bt�2�*�4�XKV`�H�<�ZX����R��6�z㎷k%jļ��}�����D�b�9-��ٹ|vk��a3ᎄ1����~/���=��`|�ZX�ݫ��lg�N�wB.����8`E:���� ��M�%x������7�m�Lʼ�_{�����u��5��z�� /�M�=#��Ю����t��;�̽��X��n����xy_��I����v�k ��M�=�� �S� ��ܰ}�Z�v����T�k���Xq�ƥ5ӚЗe���8�;��:���H��l
@��(m����x���{�&�pF66]�馨I���x���{�&����\$J:o�ʇ�/@�� ��&���z/K�:��/ֺ�ڻ���k �zM�>��t^������	�`��7�{�z�]w�(��V�X�i=�>������z0F�6�ܳ �wvhm�]U'k@�F����.��AQ�Bqo,1vp��	�c���u�+y�7���������|��ٰ=�����@j������45V��*iݭ�@��E�{�&�tp�:y�?����vNW��I��Ӵ�NҪ�V�f�T�T������|6����������vwh��ŀ�yE��{vln��T����*����ڢ�0�u�_����7@�G.U���$�0����Q��n��8��Μ�J���ܘ�$v���8��\+u�U�.�k�g�w�o���u���sf��cڻfr8-���ڸ�.�v��p��Q��M��Ux��y;r���&��y黷�	\͇��l�������s�y�nL�k.���@�[V��F�^wd�y��q���4v:˶�s�;*en�C�͎�v��+�hҍ�V0:MV=���u�����S��gs0&f�kp�V����R1�1n�>��2x��28{q��ɭ�9�K�sc�����T��S��wt�x��\��X����0�u�|z��]t�]�WVƓX��n����x��r�=��F7l�����ē����x��r�=�t�q))�(m�Zv�0E:����{�&�tp�>�BcUj��tӻ����G�{�&�Np�=��?�T�֩
?ä%���']���g�0��˃G<c#h��7�J�p�F��%e�k��������>�� �S� =�s�==|F�������b�� �*E�@[7����㳡0J����-!��D?�
3��`�uX��,����5QT�t�;j��`�u�����I�H�8�R�j�:t˥CǗ�$x��n��8`�u��qԿZwM+���&��t��zG�>0��x�Wq?���n��ݢ��������뇱��q�(��C�p�/3�g���d1-�YJ�+��O�����`���s�=�t��b�we;MU�v�0H��{���tH�};����MҺm�� ���&�W���ڒ";���o�w����^����S��
�V�xwI��p�$�� �w<���n�����lwm��R,�i`�ڰ7ږ`������߭�ߏ���JZ��i	zx-�p0l��m���	\���m�3�9�����jZbh�9O(�n�X���H��8T�$4˶��f�G�w�M�:Gt|`�Wr
I�4����w�M�:Gt|`����ܔ�'JէWE�m'�H�`-U��{wj���;�ʡ�pe�- ���BGP$0�>SZ��*F8&AIB@P)��pҁ�.��۠uIr�YN�vӧI�i��:�ۻV�H�9����/Q������(p���"���3�����ہ�.�2J��7JE`�imk���!r�=��`��`j��`lz�Põm�B�մ���7@��E:���x��Tn��v	�`��:s��N� �{���7@'��J��i�)�jb"bh��wgh]\��5j����t��!¨ċn�ڵE]\`�U`_3��]�����;��_���y��` ��iPU����?��D���9���DQQ���G�A���w~�@UV���g�6��_����/�?�߫�_���U�s�_������y�>xo�ݙ��W�����������?�?�U������(�J����I����C��o��g�{���������?�����y�O�^/��������^�������k�D�TH%D�(Q"H�IQ%HQ �PaD� P�Q"THVI!D�E%D�Q�eD�D��Q"TIIQ%��@�VTI�RUQ$P�IQ%!Q%�VH`��@�@	Q!eD�Q%�Q% "%D�Q %D�$D� �IQ$BTIeD�RIAHQ$UIYQ$D!FI@�%D�%D�!D�%D��VIVTIXQ `�%D�Q$BI�IEeD�P�FI@Q Q	Q E� Y T$�D� ��Q�A�QTH IQ T`�HaD�THT`�P�BTIHQ!YQ$d%  $!��FI$$HH ��BB	EI	%�I	Y	d $$����BBP��  	BVVBA��	F@�HHT��U��d$BU`%EDT��U��@�$!BE�� $H	YB��` YV��IU$!B  BBQ$$ �	��!!`BBBA��Q��$%I�%V		Qd$�%BYd "B�bB�&P)@�H!%$Y
T��ErQ�Q)VP�P�aQdQ�e$ ZPd�e	F�`XFE�e�iF%@R!D�Q(Q �Q���E	Q3�͟����#�U@UV>?������_��>�</�}?���� �����g���<�����O�����ƹ�� ��y������}�Z����� ����U_�0�l�
��/�3����lDU���;����t�_ď���K욾���ӽ:fb���o��_�U������������
��Q�� AU_�_�������"��������?�����;��?�0���*���������f��v��=�������U���������@ ��_������������o��(+$�k!�n" ��{0
 ?��d��0'���Il}f��:�`h 5��Gm@ C� ;�n{lZh]h{��裡�@{�  � �  e�@�  \̪��a�nځ#@j� �@AУ� )�� � ( ��    C��@��� �{�Xz��3o}��ty��Пc_x�����`T���E<o���*��   Myh9]���ʛ���_Y��Q��Qj����DyuHy�T���G�|N w6�}��=Z�������� ��.W0t�x��t|�������}=O6z ��= ;�Dzntҁ�{����uϠ w���� v�2�N�=� 
 � � )�`t��� 1��Wn� � ��������P��J59�Jz[� 
M�G@��)�{� 4�+� =:(�]��:�R���Aӥ��}�!�gv}���n�@��C i���=���o��w�< } }�&��זͶ����ϣ����`ro`;�{�ڊo������A�}��)��>�[TU7�8�����P/a���o��xI\'��:����=��,����x4�sM�=筴'���=�A�X���z�v8����v�p�=�k� p�l�}t� h��{zY��� ��C i�`;��Gm��n�݇��`t�`�����k z 9;}��A�
U�$��y�� ܠ�}>�k��A�{��   ��SmJR�  D�*�J3ڤ�!� 6J�G�@  S�j��%T� �Ѫ��*R�  "B�&�@�)�'����?����MI��g��}���򠀪�w�

��TT��
��P@U���T��~�X~��?�%��lÄ0�Y�0����RV��HR�6oK��\�����k�f������3�HP!YL!p�.k�������6�<4���X��H4��({&�^pwg)53z�*@&d��ʒ�c�{�����! �VR�@&�ɘke�m�˺I�t|�W��������]���Z��\HA��Z�6l!La���2%��2��*D�kF�0$0M�g�{�o���,�He*b���FWC����Io��J�
J�BK�/&�k3bH��ȅxD��vh��	L�n\u7�a0�z]y��ys����#X[��3L	cK�n�_�*�3��֯�*���WU�uuOM��+.��M0��3	�6H�Ƥ�{�$�Mc�4c�V݄���ϹC����|XXB%I.h�3Dѭc��i��T�Q,B��װѶ� X�Bod��y|�M�!�C��_��	���fK���<K�%����>��${��$cRJ#(K�'%��g��x���[�\�����x7��!��	![����K�Y�Eʮ}��Q���pt�!�T�L�=vFx*Ŭ��c�5���h�9�n�Sh}��!am,)��xl�\iB�,�md�fc1����d�4-'��FD�7s.o7��5/8{�2�\��5`�I��_n�9UB/7j�W����Q�Wzt�2�����{I}IS���k֕����s��c`��k�+1����O�,͌ѐ	fѤ�?4�XK�%��Y�!)�8�B{�d�d�^KYe��u��P�+䆂5�R1X��\X�# `@�Ȱ�!��\�C�C{׆��l�_�1����	tx�f�f�2o>�;����>qs�]�K��7���{�K�6y���BFH!Ld�L�&�L$��n��\+"�Ȕ�- ��#���p,\�%�d-�2!@�50
�$	B�%Hd�`F$c[�!񫐚)�8W�\7�����̟��^�a�o8�g7�l��Ǉǁ.�2�4��dߜ��m��-�҅��Kڻ�e*K4ɜôU�.���=�p2_N}�Ӆ)&M�m��C��L)F�y-<�C#i���d#D����w�/7�p�Ã�sz�ƷP��A�,��!cKna���.�x�9�>�y�rB�S�$0�1<�D�	�y9B�����'w����rᄔ(�Ӑ��1+(KH@�Il$���&K��!}GJ� Ѕ#XP&:���Il����$��k\hF��5�$5�H�3'%��[N�uwS�6�\�o��Li�'{�E���9E|�S|8�Q�[��>O~=p����dtlx��LR�`�9�5/��&��˚��.��|$��=bVZ;}�U�}����#��Mq��/��by�w��O$��r{6jY��5緜�>��R1| ��[����<����f������Ĳs�n��s�D��eP�ɷ˧o=�s����$BX@cϵI��E�$�>��fD6ʑ�)�i
aJƄ*D�k))�5�W�R���Ƈ�!�w��N���.r.�H�1�p�,�
��rf����d���7�����m��j2k8\����#��!	�E"0�)e2H�$���%�zN[-��B}J��ԂD��'�x�0�&s�S!q;I���za�>C�^3�$�h�.oe�%�L�)�f�R�$�g8l=PŲ��	��a�1�P�Ir�]]�����9�od���,�I	p�l���f2��d%$IY���� 1���P�A��C4Ħ&�y䞰�]�crkɁ4Op ��3�$ad�%-=��l�_zƇ�6D�:5��oZ��/ Lפ��@٧xfY���BF�m��u�s��w����u��:vϹ�s4�f�h��>M�xV�5��'�%)�J���HIB�C�g��22� A�����d�����(�ך @�E���Nh)k0k
L�s5��=��8I2��C&�X�F��͛ߑ��r���v�]�Y��k)<�ϵU�w�}�+�l����h�6h��,�z{�kd&�N4�14���)I`��o!��	N�&��V2�RP����f2Mm)��l�D���G��
����[˯����?�NÚ#+N�/a��K&��|�9�	s[&����p��OFz��o����,��.��1�]T�F���.����7�r^Y)�%�k�3���[�Hw�>���qPq��U|����*�Ъ�ڄR$��n��K�,���G�G�b��-�_J����*�v�՞�p�.y�s����g��6Y��L3�Zh�sR�7)�X�C���� BBM�y�Ϥ5u)��1c)FsZ����]��[���G�'>&�LI
�B�
l��<�$3Va�.�h�֏8\9��,��㲿�c��wd�bP���"B���F6��X�nɑ�!}���9���9%'	X�9w���� H��f������FF��$RA�1$�-&%�.�y��;��y�<Ϡp��U#0%bFR"H��Ƃ{��
5���a�ٽy��/0�>>ci"р�		윅~*F� �RRn0 R,�"�Xf�T�=`�=�`�`5�d�iaa�sI,��(0��aC[�.��{ϽӼ���oY����9��"��^�9���8�Yf�n�
e!,��5BGd0bX�*���X��!1�LbJK��4�6��J!�ͦ�[���!�&rƄg�E�a�Y�50��˰�z� �i�K-#˔���zI�{�޻�/򌄀��4��<����&��OhJ�
y�d��{��ח�!�Q=4l�20�I%��r\HF�I$H@�c���K JD#
�*���0�F��"K+���\7�9�.MM�8E)*±� � o�j��,׻asAL�^{���0��y�5�@�u��nȵ���as~rxj���`B�"cO�ă	B`B��+%�L��.Ʉ�Wq�����5N�QHYT�Z����/h���(fu�wwNMֽ�%�4���F�H���z�,�c*����˺�>Y*>���iI����t�E�OE���+��B_,eQ��4�}ߝV�y�<�2k=�����L/��Bo9��#	������Ւx�53wSe�y�Azf�B?�K��<%<��t˿�����[��XuUo�W_c�G�yB����C31�����8�J�p�[A��)<������y�=�#��%��ަm�n��{^���8��m���RC�8��(밆SG!ɩ4�1��)�kӞ�T�)gN�,Y�`,�����*��p���&�,��W��п}m��n�g����Mf�|�|�"H��Le��Bf}�>�s�,�ĳ��$��B�ٽs�˞���S-�n�&3G</	r�����S�5�y�/	����j��ĉ(��`����XB���3�\�>X�������|��
DO7���$HB�֎1i�4@�b��՛��f��/���&�f]�S�&[@�,H��`�lvR<8V���1td	,l�K	$���"�ϞE���v��t��48�XKwB�����C��/��>9v��c%��-Ё7�\�ZR���x�t�:��JXK�!'����]��Zl�3`l�-�%�cK@	�l2�����	�sa�|�sR����\l�d���Md�	�ȕ%%�2�(O8{^��y�p0�ф��$n:.n�9��3�4��
F�*�e��>��A"H�� 	�4 %|��4l��B1 X$�p�2$���	�i�a4e�Gn���]{��;;����
y����ܖIo!{����h�VǤ��n�@��̃�)�@R>��a�!����<d���BT8��t6Iq*jk��!A��a�D# |;H�!!�4�7���C�p��!.�Cw.2��L$Ӿޡ������{Ҕq��;{最�f�/�L���y�I�d$�F�}�i.kp�c$�|��6{���0k�}[ 9��^�;����}�p��5q�a!XR���ia#m�������q�pԦM��'ϔ<�"��Ѫ@�B�ȐL.��ly��В������ؼ�Xk^�r��!iB�L2%`����G��V��"B0��\�m�y4�V�B��j$!d�n\�	g��/�Y�Y
���X�6}���m6�M�E��F9	����X�"B��KIg�ss���j�aF\���k�=eKp�-��>�I���i)�{�=	�{�am���6�MƩ{�e,.�osm�I�mSP"���^$!�R�#e!������!/��Bo�5�=޷�bB��R�s��f:�S5�6F��o!I�l`I��i93��f� ��,-���"�Sx����4�N^��f\��ֶ%<��h&�Rg��HP���tI������Je�ӣY.;��{	�2�kj�		L�#	�jx�o�讍�
�����Vz�ȫx��%��t�C���F�_sܺ�.��h��K�|�}��O1!�K�d��$��\�͜Wg��0��iu���C[ݡ���#$�#%ނa�0�%���w)�$ s���	��\2jfk�XY#���y�F��'��)����561+��I3DKa,
,�l��b��QM��9�CŅ��i�W�R�^��$!�C��	%��b�q�̾yw�y���k�^_)�4�F���r�$�b����\�=�i�K�/2C�7  ವ�*OB����)r��V�US��ګj����W���1�����*����V*����������UUUUR�UW���������V�ꪪڪ���Z��������������kj��������������3��謵R���_UUUUUX�UT;l�-\cm*Օ�U�8��� ����d���ySM@�Cjt+YV��UU�ٶ�`*���*�
�V�����0n�S�^j�R[n������٪�ڪ�����������V��U�Uꪪ�Z�4Ĕ�{[=����~��@UUUUUUU<��/.ҭR��mJ����R�5U*�tl+K�UUm�O��j�^Z����V��nD8�9��v1a��vN��_n�|��>`	���R���[��$X� �,R��UP|݊"���W*ҡ1mO1�.ʺP.'�ȼqaE�9�F�
��¯Rr��粸<�kԭUU ��T�,p.8g�W�]�U���)c[L�E����R��l.��j�U��\� �kj��͐��S l���Ī�R�`���SHk\֘��)R�����֩����n���;T�l
�yypõBm���E);u����Rp�,f�Rc,�[�-f�.���ez�x�l�UJ�uQ��Dz����Cb^em�A�cbR(-���	�V����A�fU*��ڎ%UU[k��ڀꪮݕf�3���U-�k�X�,���&UU�V6Z���P*���2&��ڀ�ڪ�66�n��Ԥ��O5T����UUTn�Q�l*�V�V2-UJ�UN��UWU*ҭUUUWU,UP
��]�k�h��j���������YZ��h��T�( �V1aҪ�*�V�r�62��3�UUUUuT�[��m�VQ�VͩY3/5�J�qU]UN��Ȫ�UU;�UUUUT�QF�� Gjj붹�ZE�������f,�\����py�>^|Зl�����i�j��
�)�-��ܙ�g��a�R�
[5	�*�T(B�ͪ�#a�;V�5��}Jp�����A�Q�sr��s�o6�u{��v�U��]QQT�,��jV:˲���RU���K]@�Խ�๊��֮U�[q,������:�m�����5�E������]Q�Q�g
����ps�NIͭ�-�vZ��B�^��e��y�������`�evj���UԨ�UQ�u5U!¶�]U@kQT[R��mp9b�Uj��#��Yv�x��evc���	G�n�j����FJ��������j�J����ڪy�U���$��`6ڪ��*ڪ�������5Oe�ڐ������j��[bŤ�6�X�5q�#kTM�n�ò��ʪ�)VV�j���L�U�R�͊��Vڪ��"�V�m2�V㎩U�y�U`'�.�[QY��ԫ�UUX��� �-QƝ V���U���e����T��[��kv.�V�EUP6��JGLV���3�:lT�ڪ��;.�uPxUzZ����ʈmm[GƧ����U�UUT�UI�Y��}O�R�@U�UUU//UJ�ڙYZ������tP��U�te���d�; �+�[V� ����H�0
�J�UK�*�Q�{��%k��ʶتAU���jZܖ��7+�<hb��X�
���.������b�MR�+��psz���K]UV��P-�%�PA�V��6�޽��� !�ʵ����V��WEù��ʴ�Z���qb�X� �yЄ�J�H1�yn{ax��8�.ʱmcN�������Ó:Z�r���t�ήѮvʱ��!24�����f�����V0j���a��Y��,n*}��Od���� ��Nɞ�Ұ��Fj��RU��qS]��G.�"�h�-7Kh�*ஔe�)h��`Q��ʫOgOKz�=)�������V�]�&�Sp�h�4��1�aA!���L���2�
�)^��ڱ���*���.*�mnqK1�����*j�4�u�z��!�x��UQ\�k�Ұ)�eƚؖU-��>G=���'�΃h�hl&ܬݠ0bк�,��m�s-���ڰ�6V�P9\��\T�ٴ��VRU��&mH��
����"hFi`B��؛$i��*��E�����g�	ԫr���D.w-��6����Mp�
�ܭU*gU۰c��ب�b�i`��������<�cr�AԅD��X���Ռ�Q�t��j
�7V˦��Ul��bl�W����N1��W���PGmiʠT�f��`㮮۔�y=�|l/]R�]
mu)� :َ.g�YE�eh�a�Ό����(إ��5��R������ڮ�И�
��ea0N��GXn����s�P����&�5�8�k��c�p
�]F�q,%5�����\i��tU��82<R��6X��À�i��@]�oZ�ݙZB��X�%Ś55��/h�>��8���ʘj��m�q��!�U��mV��5���p1�4����6��+��Q�gn�1f� vfy_[Y������M�����4Vʶ�c�@�`ڙDcpV��"
vl��8'��|�,�]h��PA���mX̍V���v`*��5u�UU@T�n�UQڴ�1^׭�U����%�ŗRda`�ʪ�iU]T�[UWL���[U@O>2pr���]PU@P]l��+�|W}�j��e�V�j���]n��9fɫ�һ]�����Z��m���I@�H���Wʭ\�Ml�	�-T �Gc�����!m�Ut�,]/-V
楌�6��)�5U%�AZ�U��*궩^S�՛Iq�Oo%1�����D��u�6 +�m�l��O6���1�{,�D��PU���-��F�m�{(K��v|�����TcϷ3���L�S���xw��Y�S3CUJLm��]m۶�yYIua�,��ƛ�Y�N�m��\a��c���͔����R�myn���]pWx}��ꪼ����)9�M��R���r���iNڸ��/�rM4� ]��*�Q(����T;�W[*�TF2嚱��] a�����:�6ˆjU��;j��.��A7UJ��m�+�Ǯz�� u�;a��z�]��gG[%v���X*�j�nz��p�E6�.�8�[�V��ڒʒ�UQ\�P{l�3T��3<웎j���4�l��cu�cb��N���Sl��O-�l�[]�����Q��Z7J�v3��NV�t@J�l�VQ�wd5A��� UPs�5LۤA�D��cF=������b�ѭٵ�x���F��R�6�sb���;��Q�&�����8����g��5n#u lMK0��fK���-�q���7iP�&�ݲ���Q�v�xU����F��H�U!2d�V���W4p@<�ܼk�Smv
�"tUJ�UKUUUU@V*� ���UUT�9Zծ�ҼQu] �ӵUP,V��^�A� UV��=�y�23�TD�rDZ�5��blu�0��&4�`�mEV'	qUm�j��)r�R���s����`'��Lk��We�m�tjUkmڸ6B�u&pfʪs *b���v�5[J֨��xU���Y˱�F�)��ϥu����5��U���U�+aN�䞒�]__}��Y�ƃa�V����Y�������S�U�3+/-UvW�f���ܣ+/l�/uJ�:A�Xݫh �
�����V���v�U+�rT5H�ځU�^gEQ\�u�WUTk�ժC��Mj��v�R堩�m�*ҨUU]UUζx9^:X6*�[
�/�wb�K���-v_�UUUUb���ԁUUUUUUUU[UUUR�@J��UT�ml�b�� 7���t��檨�HL��ィ�.�KV�����r���Uv�'*�U|��UVP��X�Y�UV*���GEh�ify���Z�+geV����e������
<�UUUU�l�U*�ԫR�A&*ꪵSEUUUJ�U*�R��\y�5T�UUUT�UF�UP媨��q�V[��e���n��V�U����W��^uD���TA�$�]WW*eU��V�ٴ��l��aC��mm�*��[�骪펢���@�U�ꪪ�j ���(6wg��X�gfک�x�ʵ]��C�UjU���UU��n�۸�vk`*�*j�
������YG�evj��Ov�S���՛l+V�	P��z�>��d����1K[<�r��v݁�%����5�x �(Hn�M�R�`�@��!T�r��m��PE�[9Cv+j�s���v�f)a�ݐ���Y^:��%���-�7\^���S1;��V�/[��#���V�[UUR���ـh�j T�i|�����'XѱU1��a�,3sU(�k64ݓSt��5pV��m�Q�+j�iє��j�ۙ
WI�۲�jZ�a�
�������.b�UU++r�UUT�PUT:
���jT����U�MU]UUUUJ���F*���UUUUUUUUUUU Z�V����������*�������U����V����]��Tv� ����
�����n9�-�@� *��UUv�*��U�UUZ�a�������zꪬ�=[��gun��{Y��6U�B�����W�*�������`X*�� �UT�UuUK�`*�������������U�`*����kj�nZꪪ��j������V��������h
�������UF�@�ꪩR�UP[_W��ԫUUUT誂���j��ڪ�RZꪪ� ���Z�
��@UUUPUrm��UPU���U�����*�����5 ���?UԫY� *�R��fUV)1Vmt�=�]�}��j��	���������s3Z��
�*�*
� ��;�ES����
B��F D�" A��HĐ�b��B����XQ�d��wE �D�: �/ 	@�P ����\P}DZ��	O@<^ �:PLU�Ch� r��)�|��P0a��� ���p�� ��� ��
��6��]>DN)ĉ$�#"��"�;@��x�G�OE}�����@BFR1 � 0��=��	�(�SB' ة��C�����
����h/�!`D� �HR���G�E]"�Ջ(�~ү��b�@�f0E@�j�(>�	dQ� MQ�Am�8��S�=~"(���EH��@'*�a�0 14m 4LW��Z	�.���U�ED|��PH�
�S�؟%b��5 ��+�{�.�-T⵴V�B@��|J�F �(��BFP���R*-*�j�V�bm�W�=Q}9CH�� �@>}@4
���@�,�RU$�--�-���������#J6I��$+!B�`X��hYIX�K)D#HU��JQ��RY`�2�T�!E�
Ə��xz
�n��J9*? HA���4�� 4*)��Đ�G� �$F!�(%M
�"E���&��EW���G�C�T(X\R������
�ZE*j�V�E�U�R�@Gb�yug��� +j���VqVZ����r>j�j }��֛<O]��q�����8UPV�ڲEZ�gNCP�X$���cc�q�6lg\�r�e,�݋l��	�N���il\f�a!�y��Vm[ˁ�0�0��G5��tp()@�Fi#�X��2��ҵ�&��+S�m�+[V�F�$�{0�M͹؞.&ݻqpK���U��!	��.�����S���z;���\��¦9u�=����	��#a4������"4�Y�� �66&�g�9��nT��,�Rkr��m:��3��"S�S[�4��8�%�b��ܚ�7�nMR�֕݃u�g���f�Hݸ�n8S!y�y������Nw)Ύ|qN61e�* �>��WpOMl���f8.&��3*f6�7��Ĝ�=��W���CŸXdLv�/d�-L6k"�ccg\(m���զ�	�-k�01��\��)]�k���uF��"k[=�����b5��x���˝Ƙpb(������6}���g^�gIƦTɂ���ͭ^�gVUpLs��-�[/c��p��e��)�&;*lv��m��X���eN�u�&|�ɥ��������K ��m����&�b#�BL�M�'\����L�\i3q�V>�.���qFn�ƜT��#
�n6�Z�n
�k
Qu��v��hZ�`���\����\<4��ڙض̬�]�����2[kT����a�)F���LA㋬�vr.��Sn���4v�3\(&l���KUj^�UH]j�\a��rks�v%"S�^��AM����劫��3�f5�#S�8D���*N�m�\�<��us�v�V@�f�|��:�ʹ�� ���E�(k`M�u�ֻr�	Í���ۤCj�9\������Wt B�t��(,��WP�i�.n�p,/6Ҵ�E��I�s���q���j�BJ�����[,V堥�ؔ�8.d�y��6m]�c�5��ܻ0���̂�U��
��ނl@�����] 'S��X�(x��C�c���#�FY0��WY�(-�%(],Ƌ
��ؚ���z��9�d��7U�5�\�XZF���1��WFl]ere�l+�SLuYT���*!Όː���6�$R�����7lu>o;��&I�Ҽ]ob0�8�5qH��c��Z��ۅ���C�9"�9�6ㆉա�V"K-Z�ܹ�Z(���X�����ތ6E�c�␫�������Ӽ��b�kh5���(F�S��-�TXë/J� K�e�ՠWV��j��/ ��L[�o�+���^�A���WJ���nۼ�r,�4��ul��uwe��EH#T������>SIxV�xWv^ݎ{��8�E�l-QE�� ��/ ����;�� �^�xʢ�U�M��U�;�xWv^ݎ�Z� ��/ �*�ʪ��K
����n��^'+ш�[=۫�BʌD�h7�<Cb�����]��el˟@��� �kQ`ۑ`]�x����W�Gd��~���t�8� v�|S��Y�����}~���wc� NJ�e�Wut۴�4�Xv�XWv^ݎ�Z� �y��WI]�,v;w�uwe���}/T�W*�m�z���]�]*w|w��n��p�>SIxV�xWv^�rI���}��3#��L�$6���v7K��`(ۈpӶ��Z� �	Y���Z�6����z�������0�QH�Ֆ12�Ec��d���/ ���4���Uq#�����m�:�uccv� ճ׀wc��¾Ք�(�"������ܓ�s��MR��]�U�������}5���Ȱ���
�+����cE;�`Mj,�r,��/ �� �����.M���t�ZJ3s���q�#u�@��+�j�,�:�y\���H�Zi��r,��/ �܋ �kQ`o6��w��,vյ�uwe竜�U$l�y`�k� �܋ �h⻠�T���w�wnE�}��X{��%���ul���T�N؄ݺC����>�dXv�XWv^*����r���b�;�E"cVX��-wi��r,��/ �܋ ���{��*s|�_�3U�Bir7f�ظ�� �ܼ0�m*Ź�<lN��67&+t4��^k�s� �܋ �5��ʮ|�e�� +�^��e��
��T���ۑ`��`[%����	�0V�7t����	�ۗ�ul����KV�^������W݂nƬI��UKn{׀j���;�"�'u8`o6���ݫmYN�n����Ix�V�x�8�ª���;�PAm�Ѷ!�s��pj���6�Xv �MS`�Q2�\��znR�m����q���x�d� k�a��k;�!��������דD�O)<vu��Ӎ�.o%�QmB8Ժ�P֑�i���B[�f��,uc0vrEM���v ��!��.?U#o/�<Jg��}����6viݮ3�;&G����뗥���������n�l,�R��}�'s�<��<�$Y�,n0�p�^Y`u�m�)�c�CbCQ��sX˸4����ĊI����5{��	�N�����v*M)e4�M�:I7x�V�xV��IxwRSE4���v��r,�v^�$�v;� �AHSV�WO�؝��������'� �=��'bp�;�"�
��+��ۤ*�-SV� ��/ �#�ݹ�v^��r��%{��6���gBM�cN)%��V�R3	IQ2Ÿ��fB)r�ѣ�A������;�"�:�e���W�5Oz�ܕ뻻���M�Չ6`[%����H�[P'�RJ��!	@F�
���$��;��{~�ٹ'�|�,�r�;98�_�h�2�c�x�=xV�x�w l��vS���m ��n�=�r��/������������v$T�H-��aWI;w�N�ܼ�d���/ �^ J�=�qôpA���F[s�W8א�p�s"k`Ս�Z$l`:��2d����d���/ �܋ ���>U­Zm��>[c�w�|���ˑ`Mr��d� ��bW�t�WE�wn�ˑ`Mr���>�r���t�l����vVt��RV���,�5l��|�e��"�	�R��嫫��v�]۳ ղ^�ݗ�v\� �;� 6*�Gt�J��3���fj�9�;xӴ-���b�1�┌/.&��:le��n��%�RK�$�r�[%�v�V����I�Wnۼ�Iy�/z����xV�x�H���[�
T�n����ۑ`�<�Ix�D"cHb-��v��r, �G�uI/9\�s�IӴ�,��7{�����~����<��� �G�{o����z��۞� �/��.�˙hZ�!\f��B�ҎMo�Y�m!0��n��\��qfv��.�fjB�E����:���wn\�v�X�G�N��e�tՎ���J��;�.^y"K�� O{� � w�R��Ʈ��i���x�ȰI�r,�K� ���'݃��j��	$xv�Xdwݹ���.��$�][V��;�"�;�.^ݹ�ܒ{��krO�� �H���$H���B�RV@��E��_i�&L���E�]�z���Ά��h@!6,L9��tZ�&v]*S6�tF`Ʊ�1v.�mf��L��*e6f�u2���t<��JH���k\��n�[`SAP�Ζd�vx��� 7L[*m���c��pYhW�W��'7ا�t&���M`X]��/5�&���]��hQ5ڎzD� ���n���Tc�Q�OWgjyn��یv��Ƹ��-�zN�L�FG�pjD��8�;J�����˷��j^v��;����9�WT��C*ݤ�ʶ�*��;��� �܋ $��ۑ`!�N�-����r, �G�wnE�vGq`��I�V۫�|��v� I#�;�"�;��Xv�X_vYwq+mRT�I��xv�Xv���;�"��<{Q���Ul�P���r��͏�_ O{� ��/ �4���7Wck�g����hR0�Yp�A�e����Ϣ��9A)��7ݰ�֫�E������Ӡ�<�r/W9_ �������7X�5�� >�ﯟӾY$��{�
� �"����`�]i'�b1$�ͩ�}�Iw\�bI-ݬ�����7L�^� ����� y���}��u�F$�[$|�]�Ef[WMr��hĒ[%O��K��#I-�?� ��{�z =��N���q0�ϾI.똌I$�H��$���x�Kd���
_�t���
p 8��g\[�N�Pj���s�N�q�Ӄr��ᄵ�ͮ�5U�>[i;hĒKd��K�\/Il�>��I)�01$��e��$��*lV����%�^$�ٵ>��I)�01$���={���I�<=��T�4c��dۖ��~;Ü�߽�[&��=_��18������T	0 ��5
��@��dܦ��ȚR�y���tY���eߘ��������޴�T~ͬ���4�1��p��Rd	�zH>�}�7��������A��J�>>�y�X?:I�'��9�b�sA����3l3M��%(�"��`J0�����b�Qw�!�A<����JB�{OH���޴�j	�G��0�3��FLnFa����8��My��3�S�lٲ��Ʌ��.#P�(K����,B�hBc���d<M���$J�7�&$�ϪX���yh�P�B!�Rah�j��� zJHɈM�l�iGg�4��6Nk�5[�~�ن�^n�h۵B`�"Nxs�r)Z�� ���`�˯9���|&�	!H�0`CR�c�^y�pʐ�B��>��6Þ���[�5+�Ѹ'����7Z��=��4�a
E	���!��6	`\$%f���0��aVЌ���#Q��b�]}�ٸ�cs�$==||A���~��<~`PU��pC4"��@_>=b�J-����6���S M $W._���-���~�ݶ����s>���p��^� ��{�: =�׾�?��ݺ�ɶ��g�}�s��E���m[��$�͏�K�{.�I%�j?� ��{ֽ ��o��Xۃc2�#-�fe�i��̚!A)�s�Z�8��T�m۔��7L�/}��M� y�׾�Iwf3ܪ��i%=<��$��)��;��ZCl�� ��'�}�Ól��M� =��� �7���߹�[�,��;�l1
,^� >��M� <��^�>�xo�7@��O�� '��gVVe��ge�����{��=���n��}���[��>	XEcP�"D #HFU.�X�G��y���ڛ~yNa6��`�{��[m��#�S}��=��g{�f�m��ﹽ�oϟm�yL#�������u͜��� �,፺�q=�8DjMn6X"������&�rY��� <�����=�= �������y��� �O�o�t�PLf/}�y�M��m���{��}� }�z���s�/�����.�MX�o@����}��M�}ͱ��O�� =����O{[J��vW���Z�{��$���^|�JI�ĒJI�$�{az:s���a0.z }�z���$������������}�_}}�@���~��=߱\U5�[ ��ڇ�����e{�E���e�R�!��d��m�^lI�th$�����y�'p���b�m飚�2�,ѵ"�uo4Cƭ�@�Y=�s��r�b�)6B�a%��k��I�Pn6(R����i
�������u��\�(���hݶ�9��Cu,�ۓ��^��{[���M��w�&Yj�n��f1�lsz��`{����zZ��"�Ur�-��]L�`���X=e���������4�~�g�Q�p���RI~���$��?�I"I��U��ﾟ=� O'�^�X,��;-�JI�z�\��{��x�I{ޯ?�I%�t޾�s�`<��Mwڹ��MCe�$O{)�I%$���+���UU�m�~��� �����7����4c�ec�oUP����u�[o���&�߾��s��I�L{�_W� �σo�vj�f���ۓ,Ē^������RJ/?�$�������2�Li�)�J�eT�%5C9X�-��òr�4tY����w�y�]V��&�L�� ��{���ۺ }�z��~�s�?~t^���~�,��vW��==}��';���,���� Ꜽ���;�r�{�wy7m��ﾽ���I���T����צ�s:Zs9�� ���������^���ͱ��|�����t {�S�t\�Ka����z�w�Y�m���u�[o��f�Vrm�����`�}���U��ͮs�@����ܒs����� }����=���� ~�I�v}ŷ[T�f�ثoZ亰"iHCAt�fbʴMu@��hUIQ�I'�S]���F���������I%$���	E&U���W+봒��������b��WvU� ��={�E@�������m�w��9m��ަ�/&�9���}�٪1�������m�߾�\���b<�X*|@Lc��J�T���J�P�d@M�Ǣ�=����n�i��Ϟ� <�kU���.c�I˻����$����ĒKd����U˹�vހ|���X�7L�^� �{2�$��r����y��$���ĒJI� ~��z:�hn#6��XĦ6�L=��[���5͹�X�������4�;���y��6m�?������|ϴ�JI�\�w��==��$��LW�uvƖ�s��=�}�NI�NNE@����s��w��7m������:�������`*��&�(t {��}����7oEP32���9m��Z��|�܆��l���e�>��96�޾N�����9m�{�}n�*(�ϔV�� �B3 
PBQCQ�$+2 �up^NG�NI!�����`o�I��4�.2��: |�z��Ӓ}�_v^��~���S���{���*�l�JV���.x�-ץ^�]�&�9��ԛ��J�,�;�'9��&ۭ��4a�b������S\��IMq�W�i%�����S���V������������~�V��?�bI%�߫��䒛3=�]�^���t�Tn�2����� ��={���I�Ӓ+���R� ~����}%�b�wl��6��{�IOz��o���$x�\�s�9�_��~�߃�w��wLAJ�t�;&V�����_�~����~� �*<k��R(����;m�#��U`o0��F�jRmm%ՙqsa�%�Q�6�b1e+p6��V"66*˱	�,[A�!�W"�mQ���&�6�@c��@����ɤށ܂�rf����r[:����&�1p�`��L-,�Uu�l�7k��]f�,i,�Smp��h�I\���a��(C���m��W5������������N�{κ�<i��B�9֩U��*�KI�0	H�-s�==Hx6��w���8�:�t@U�R�W,��~���n��	%G��s� ��e`�Y~0��+��^����{��N~�rmo�ߧ�~����H���9�$yi���ݾ+m�n���y��ᇫ�\�G��<�g� ;�Q]ܻ.�t���xO�'�T��y�nI?~��[�}�{�ܝBrrH}����|���$�vX�\ހ$���Us�磞_ {ޯ<v8`�����k-�\�eHE�\��3B�3ɠe!���h�vwlߤ��s�|I��.��m��� I*<{&W�U\��	�y���e���e�@ۻ�O~��[�����*�,#��q��T�����F�
A�Fb-�q(�a �;���UV�~ﲰޞxe�Y�UW)"x�wu~cX]�t�7����<=U\���<�{��J�J��&ۥN�7m���q)�y���, �*<s��/z{���Ҳ��;j��J�KذW+�{�����V l�����F�Ui� 1b�`�k]�0*��t��)��;%P�A��sDW����y|֋��v���m����� �\0d��'$�﷿[o��Z}>5�.��٦�	5�?Wꪪ����ߞ������z��'$�o��}�|L댍S7�m���$���빷��24 HR !���� H �X�c0DX��,\�4'��~����$���7j�(BN�eջ���\�qK������ ٮ�9�JOy����.�K��_n��Tx��ʞ���	=�6< ���1�f�{G35(Y�,��,v����m��A�u�lKVTu��I�xk]f���b�=��d� ٱ��U\����J��x�]�t���bnـul�����s�+��]��{��	����5�=ʮs��iY~��ظ��RV� '�� weG�� ?"������rO�~��=�O��lӫ�v�V�i����s��[=^x��VI<���nM��������0���&�=#�!�6�h2q&�;�6�1��C!$�I��;���;�/���������v�L˵�o ٳ+ ����s��߿_@=�ߞ weG�l�Qt^]j��I[mU��z���"�WGiG�W��lr.�Y�15�R�i�t���<Ex�ӵm1��|��^�l� �ʏܪ�����V�+�"�J�t�.��n�Se窹U\��g�� ����:�K�W9��;�/�l\wn��� 6z���2��+�ʪKT�� ��׀|�}+�ޭ�6��9����t�;�#���~��}{��nI��߳r~U� �O~�� �J�_�*�ګ����ݳ ��/ ��s�*�������	������Rz}"�,�e_,���؁�p��ޙ��ݻ��Hl]4}��M��摔�E��1�Y4B@�!Z�d�<�%5�q^'�����C!$b%!BH���Z6�`���.�"@"FPK�^�]��sG�9��%g+��y�l9P��<��H]��@y��x@�,O��'�zh��j������������Sz�jS�����喝gE��F��A�@n�BmJ�j+Y����6�1nv ��"���imK��c4��8�٠K5pd���PF��B0����s9�vcu����#�}�RdT)����'me��5f�66��g�f��H5S#���Wf��js��㴋U��fn��;�4�hۅ	y���Va#6`[hJ�f7XI[.�b��FUث�7\2��7@AUf���J�P�ɳ�aʯ(J�U�.܅��A��/J�c�NYz8Ø�Y]�q�Z�%�#����W�G�����v��M��tC�&v�~���=�;,�GEb�d�'-<��k����k�l͜7WB��z9���՚NA���4�r![[�ь Ks�A(�Ճy��IK)U��#\Sqf�iSjGk�#%p�=�.H2�]�$��Gie�cc�ZB�D��hn'����Ocm�B|��D�Kp�iW�m�Mp�A���(�X
�k��f����K�lhe��q ��'dM����]�[ٰj4e�R
�)Kv�t� �h�V��f��*J�'Ll�K���K�B�RX�q�*4�Vڲ�V�T���7G9ճBً(u�ͷ0\�0ƃVA�6��SbtW�VExv�a�i�y��/Z�0:��#�}c��q�R64t�n��k6狴Ή��iڶ�d�+T�<�!k��(�m:ۊ��/k��l�h��cl��j7U�gt����ۮ�'-��䢄�c��x���8mۤ�C�n�6K��4�pT��T�NND#lۣ�~����:���mFZ�{`eZ��u�*��F��6}�8�Z�T�Gc���7n�&�ILe�V�2�iK�:�0m����i��ɑ4�U�}���S���/7���'���d�M��䤛)��Mȁ���٣� UT�+i� [v���j�il�U�Ƈ; ݀��gg17Q ����eiIUlQ�^��Iր��d��f�=��&�f���(��z�v�����*�#�v�zu=��*"&�N/���}\_���w�->��SM�E�lU���a�eX\X4���-yt� ��+�Zh����kai��<���tlV�'��.� ۥ!�N7Yx�]�P�ܛ��$�s��v��̙G�m�Ց�n���p�k��iS:���![M����'.]u����$ĽHL���݄+a}��i�s�z�3vΎtR�
�<3�;7Y�0�j���ERnD��m�J�5n��ޓ��t�����_GU�����������=��xl8l�:�mgd�-S}�{��}��)��S������`vTxvL�r��ϐj���i�+E7WV��ݵ��Q��G�T̟w�훒}{��nI���}d�%�]����+�t�����:�K��ʮq-��, ��������ܺj�[Lm7X�r��n{׀l�y`vTx�r�ų���I^1Z�T��2��� �܋ �UUW�W��l����&��߾���4��\	`�ptn��K܊`2��)��l�a��IӼw�����ںCm|'�� �d��:������&D�,O����ND�,K9>��N����]���rwy�^Kϻ�NC���cQ!bPV��2-i Ƃ1�Ph�UG"��ȉ"� D�Pq� �"H��bfw�ͧ"X�%�����iȖ%�b}��v�9[ı<:}�@��S0�.��ND�,K��{�ND�,Kߵ�nӑ,,K�ӷiȖ%�by�{�iȖ�������o���Cgu���"X�b{����r%�bX�}���ND�,Kϻ�ND�,A�=�����Kı/���1�3Y���35v��bX�'�k�nӑ,K�|����Kı=�����Kı=�_v��B�����~�N�E�9�#n�0nq����.k��5��nǢ�qu�J{mh����e�K|P� tǝ=�н�ϻ�ND�,K��{�ND�,Kߵ�ݠr%�bX�}���ND�,Jt����ۿh�\�Z�Ο�Jt�J'���6��ؖ%����nӑ,K���t��r%�bX�����r(X�r��}�^��R��6:�����b{��۴�Kı>�];v��cP���U��5_w�6��bX�'���6��bX�'��p�˗5)��e�˚�r%�g�H������r%�bX�w��ND�,K��{�ND�,�E[߻�&�)��һM�m	l�gf7��'@��ﾽ7�A���ٴ�Kı=���ӑ,K���t��r%�bX���p�&v�	+\<s�͒�tc��3q̬�:�U�k��ٝ1su�<�ݣ<|$�:i��*��9ı,O{���9ı,O~�y��Kı>�];v�"X�%����:{z}�toB�??>"?i���]]�"X�%��~�ӐlK����v�9ı,O~�xm9ı,O{���9ı,K�l�vh�Y�,4L�m9ı,O���nӑ,K�����ӑ,ı<�۴�Kı=���ӑ,KĽzv��;�n�L�mֵnӑ,K? �\��~��r%�bX�����iȖ%�b{���ND�,��@$R @C����Ț��~�iȖ%�bw�݆~ѫ���kZ�h�r%�bX�w]��r%�bX~E߷���yı,N���[��Kı>����Kı/a;>�P��(���Ֆ7zonې�M�[q�b3����X7wo	�1+���Uo�?�X�%��u�ݧ"X�%����m�r%�bX�}���<�bX�'}�{v�oB�/B�����/�Wɑ��y�"X�%�߻�۴�Bı,O��xm9ı,N����9ı,O~��:����^B�}���m7�B��l�ջND�,K߻�ND�,K�뽻ND�����iȖ%�bw���9ı,ON�w�-�aL0�.��ND�,B���nӑ,K����iȖ%�bw���9ılO~�xm9ı,K��e˝�uf�:3W&f�ӑ,K����iȖ%�a�b?��ߥ�yı,O����"X�%��u�ݧ"X�%�4�*)D�4�ZAc	;߉	��\�Y6`U�IJ�i�)-�XU&��yˤ���HN�Rk�������C;f� �a�����q�l\�sa�_(���]n���p��9�nݸ����ri��sm���R$�."���eb0��	k�=����ks�Sb�2�������ΚL���ݓ��;v(،�.��fA.YX��y�nt���:��z�R��ץ�mӮ>-�,]���I:y;����jG�9�$@m3�h�e�7�#�s���\Nݸ�ʞq�������<�x3G.��<��t�K���|~�ND�,K߻�ͧ"X�%�ߵ�݀r%�bX����m9΅�^��O��>5�] tǝ=��%����fӑ,K����nӑ,K����iȖ%�bw�t��r�t�Jt������+nlWd���ı,N����9ı,O~��6��`��bw߷�m9ı,O~��6�:S�:S�￿�m-�SLeo�9ı�=����r%�bX�����ND�,K߻�ͧ"X�"���u�nӑ,K������55�5�n�6��bX�'~�}&ӑ,K��@� �(w���6�ı,K�u��iȖ%�b{��iȖ%�b|g���_��Rm�f�Ѕ�5�^\i_'\�rv������eA��vK}��'R�+&԰&�˚&�Ȗ%�bw���m9ı,N����9ı,O{��lDS�,K���o��r%�bX�t��mְ�L�Z�M�"X�%��u�ݧ!�
����C�����DȖ';��m9ı,N���6��bX�'�w}�ND�X �dL�oC���#����h᫏:{z�z>���ӑ,K���o��r%�(�%�����"X�%��u�ݧ"Yҝ)���C��h�M��Ο�K�������m9ı,N���ND�,K�뽻ND�,�T�=�wٴ�Kı)�Ӷ�rM]L�m�ԛND�,K��ND�,K�뽻ND�,K��}�ND�,Dr���3���G)�r����������˨��[�0���cw=Kf[49-��J�iA�E���v��y��+nlW,��ҝ,K�뽻ND�,K��}�ND�,K��$ءȖ%�b}�{�iȅ�/!y>�߬�m)l��aS�N�ı=�wٴ�?�S"dK�w�$�r%�bX����6��bX�'��ݻNEı,O;��9���SY�S0��SiȖ%�b}���ND�,K��ND��n�
��4�`F1�0
�$ %h� ����Cz�;�MD���ݧ"X�%��~�fӑ,K����L��h��asS5�6��bXb{�{�iȖ%�by�����Kı=�wٴ�K��~�I��Kı>;���˭Ra2]kZ6��bX�'�߻�ND�,K =�wٴ�Kı>����ND�,K���ͧ"X�%�>����?q_�K���r��G�ˋv��L����J�����=���lU�lg�m-�c�5���yı,O���ӑ,K��߷�m9ı,Os��6#Ȗ%�by�����Kı)�K��FkD�-�M�"X�%���o��rX�%��}��ӑ,K���w�iȖ%�b{��iȟ�A�dL�bS�O���Bj�f�nh�ND�,K��߳iȖ%�b{�wٴ�K,K��}�ND�,K�{��iȖ%:S��{�O;~R����:)҈6'��}�ND�,K��}�ND�,K�{��iȖ%���	b}�w���Kı;�N��[�WS����r%�bX�����r%�bX�����ND�,K���ͧ"X�%���fӑ,K��!��י�,�Y�3$�&�]��fBLIcK��;��)rB�cu��wC5��vhZ��>)�ı>���iȖ%�b}�w���Kı=���؇"X�%��{�ͧ"X�%�߾��2^��	m��f���Kı>ϻ��rؖ%���fӑ,K����fӑ,K�����r'� `DȖ'N�?^F]CNe,ֵ�ND�,K�o��r%�bX�����r%��%���I��Kı>ϻ��r%�bX��~�n^�˙�r�I356��bX�b{�w�iȖ%�b{�w�m9ı,O���6��bX�'��}�ND�,K�t�vh�jMa�Y�ͧ"X�%���I��KİC���ͧ"X�%���fӑ,K��>�siȖ%�bb��N�_g�����pk���5m�2�K ��h����.]f	���u%�^nݹ�F4&�'����,kFu�dˉ1���W�[������\�o�]	������. �֛�> �"�+��fm�r͎1p鲼X�6S���쾴��<i��3E���^7(�lhb礜mر�ط�t��Dyt����U[mg�n�v�ɦv��kl��z�!<�5WB�gC)��˵X7M-���;'\�ʚ`��PK��&���M<H53s:)ŉb}���6��bX�'��}�ND�,K���͡Ȗ%�b{�w�m9�)ҝ>��e<��Jݒ(�y���N,K�{�ͧ %�b{�w���Kı=���6��bX�'��{�ND�'rtoB����ϻ�[B�Lj�]��9ı,O���fӑ,K�����r%�bX����m9ı,O}��6��:S�:|�zk�߭uM��:r%�`'��}&ӑ,K��>�siȖ%�b{�wٴ�K����w���r%�bX��ٹ�%�f�%����&ӑ,K��>�siȖ%�`'��}�ND�,Kߵ�ݧ"X�%���I��Kı?!��O��Xj@�z��;/r쯝�-�d��Wf�����8���葲������?�!ı>���M�"X�%����nӑ,K�����'"X�%��}��ӓ�:S�:_�}��~h\޴@�<��%�bX�����9����	�a�BH���)�D�!�@�� �`P0`��HF0�@�%�d 1� �����I&$���! D� ����P`�$I���� �d
+#`AF$	&!JHI"AdH����B!B$k�����	�E�2%���o��r%�bX�g��fӑ,K����i�N�t�Jt����4�3M���'"X�%���I��Kı=ϻ��r%�� 9"}����ND�,K�����Kı)��ۅ;�M]L�-�iȖ%�b_~�u��Kı=����r%�bX�����9ıF�����r%�bX�?M���us5�k[ND�,K�{�ͧ"X�%�>���m9ı,O}��M�"X�%�}���ӑ,K��u/e����&QY��.h	1�ST�l�ƍ�fiƵf�)�s��l��s��ՍM5�O:)ŉb{�w���Kı=���6��bX�'��{�ȰO"dK�����6��bX�'��d�\��W53��ͧ"X�%���I��Kı=ϻ��r%�bX����m9ı,Os��6���Q�"X���o.K��Y!n���&ӑ,K��;��m9ı,O}��6��c�N!�=ݒ����z^{u$ȑ�dq�!� o� �M����o��fB;��)��i�I���	,l�!����� �z�R/��:cGo����+�F섏$B��Cm%���r�g%<�$ČB��rE�$�	�CA�sD��ˢ&�䬑	D�##5]C-iy	7��hN�8�	!'� @�co36��Á�q��W�<�đ�����s$H!��0��6�kGhڐ	�p�j9`�M�Ѭ@�e��I2��g��5�H�(M���`@�t�� =�������%�I3�Dp�@�I��X#	O`9�d9�����ְ�7���������0l��@�$\���0"�4�(oB���>T���E������D~)�} ���P�O'P�9Y�=ͧ"X�%��{��iȖ%�bz}����2e�K5�fӑ,K�=����r%�bX����m9ı,O}��M�"X�%��}��ӑ,K�/Ͼ�m?�ݨ�6O:)ҝ,Os��6��bX�!��I��Kı=ϻ��r%�bX����m9ĳ�������߆�L.� ��������t���Ce�K.���-���'�u:جцh�պ5u��yı,O�����r%�bX����m9ı,O}��6��2%�b}���6��bX�%:�����&��h�扴�Kı=ϻ��r%�bX����m9ı,Os��6��bX�'��}&ӑlK�����c�z�E�:)ҝ)����~6��bX�'��{�ND����>���iȖ%�b}���6��bX�'}�y��-%`�MvSΟ�Jt�Jt���ݧ"X�%���I��Kı=����K��'��#�	H�	lOs���r%�bX�~=��B~5ɷ��O�:S�:|��v��bX�'�w�6��bX�'���ͧ"X�%����nӑ,K���_ߐ�3YSV��*T�jF��;!����l�r��]���ة1c*�s`y�L�iȖ%�b{�{�iȖ%�b{�wٴ�Kı=�]��r%�bX�����ND�,K�����FL.B�ZѴ�Kı=����r%�bX�����9ı,O}�y&ӑ,K�����ӑ,Kľ{�Y�vk3Z�dԄ���r%�bX�����9ı,O}�y&ӑ,K�����ӑ,K����iȖ%�b}��ӹ���0�jS	sWiȖ%�b{�{�6��bX�'�w�6��bX�'��}�ND�,Kߵ�ݧ"X�%�O��{'f�5u3D�Z�iȖ%�b{�{�iȖ%�a�?}����Ȗ%�b}�~�v��bX�'����iȖ%�bx(z�'�´=(|k���pe�mm��穮�m{VeB0�fkz��=[��7a�Fj7�ђ���f{�'Ok�9���و	�έ�����\tX�gWM�&	�S`��V�\[�v�t��km�J��r�K6%a�Y��`�.ӌ'��b{��}aC��m\z�Z�s/m�lp�In� ��Yc(#���!-��C�q=�g���0l̑!�����s�Og's���a�j����#km��T�(-gR����[���m,�Ra��B�L9���|�D�,K�����Kı=�]��r%�bX����M�"X�%�����"X�%��zvp̚���j�f\�jm9ı,O~�{v��bX�'����iȖ%�b{�{�iȖ%�b{�wٴ�M#�2%����w�p��\��d�j�9ı,O=�y&ӑ,K�����ӑ,�#�2'�~���Kı>����ND�,K�Ϧ�0�3V�353Z�iȖ%�b{�{�iȖ%�b_}�u��Kı=����r%�bX����M�"X�%���Hvrk2jB�K�kFӑ,Kľ���iȖ%�`��{�iȖ%�b{�{�6��bX�'��xm9ı,O���3��iF)�a\X�v�-Ip����L�-���l�55�s��mMT�z	����r%�bX�}���r%�bX����M�"X�%��{�D�,K��{��"X�%��{'N�WD�3E2K��ND�,K�{�I��(<"�""�H�E9(�	�! 
4:(� 㨖%��{��"X�%�~���ӑ,K���}۴�Kı/�̽'n�5u3D�F���bX�'��xm9ı,K��`	bX�}��v��bX�'���6��bX�'�~��'u�\�����֍�"X�@ (؞���7�O�ϻv$�H�y�ƓpID�O;���r%�bX������2��WS3Y�k[ND�,K��ݧ"X�%���ͧ"X�%��{�ND�,K��{��"X�%�{;�f����jF�faaG��8ԍ��~m\=�
���v]t��zЉ�'t��|�i���%�o�>X�%��߿�r%�bX�����Kı/����Ȗ%�b}��۴�Kı>���f�j�Y�f�h�ӑ,K�����"X�%�}���ӑ,K���w�iȖ%�b}�zsiȶ%�bzw�;�k3T�d��kFӑ,Kľ���iȖ%�b}��۴�K�AI��&��H�﻾iȖ%�by�{�iȖ%�b_�}��~�����<��t�Jt�O~�{v��bX�'����iȖ%�b{���ӑ,K���o�iȖ%�b{��������kL�rwy�^B�����r%�bX�����Kı=����r%�bX�}���9ı,�����vGQ¸��Jaю���-��Js�������9)���l]�;F�h�扴�Kı=�{�iȖ%�bw�}۴�Kı>�]��r%�bX�����ND�,KǿM�gu�]\�CZ�kFӑ,Kľw��iȶ%�b}��۴�Kı>����ND�,K���6��bX�'}�a��e�a���|��t�Jt�O}~�t�:S��b}���6��`ؖ'��xm9ı,K�~�bX�'��xe��d�պ����r%�`؟{��M�"X�%��{�ND�,K�߻��"X�܉���fӑ,K��{w��隰�a�j��iȖ%�b{���ӑ,K��w��iȖ%�b}�wٴ�Kı>����ND�,K��{����8+2�E��1��l�vԵ�ӝB�(]Rq1f�t�q+	�+͡�u�h�r%�bX�����r%�bX�}��m9ı,O��}&��QY�L�bX�~���ӑ,Kľ�ܳ0�uu�jf���k5��"X�%����fӐ�$��,O�w���Kı>����"X�%�����ӑ?C"dK���/�Ae�P�6O:)ҝ)�﻿��r%�bX�����Kı;����r%�bX�}��m9ı,J|���N̦�պ%��m9ĳ�C"}����"X�%��>���r%�bX�}��m9İ?*�2'����r%�bX���7!��T�\�Z�h�r%�bX��_v�9ı,?�{���v�D�,K����m9ı,O{���r%�bX�OWd�I�t��d$�Ӭ�=�ol�6
�6�+���
K�rVk�k�%ޚ�ۜw6v:ZD �5�e�B���f�]�dQ%��ƶ�Ǚ�.�!�S������ь=�"�!��`�i��`�3T�%�)U�t�V�*�R�mjͥ[���N���dM��=6�kl�Y��f�J��
ƍj�ǭ�n�T�e���-tĎ35�:�.�f���^��<���C�0P��ح�3��N����r���Tk�<YW{q�9�{�T��7e���lCF˦�5J���!��K�b�M�V����N��N��_�]�"X�%���o��r%�bX�����Kı<�۴�Kı�_>'���#Wa�󧷡z�x�߷�m9ı,O{���r%�bX�w_v�9ı,O���6��bX�t��O.��f��G4ه�?���N�O{���r%�bX�g�w6��bX�'���6��bX�'����iȖ%�N��ߡ���������Ο�Jt�K����ӑ,K��;��ӑ,K��߷�m9İ?�	�;����"Y�^B�{�.���F�D1��'w��bX��}�m9ı,O=�}&ӑ,K����"X�%��{�siȅ�/!y?����K����DR��u�		�BZ.%%��6��0��q��Z�96�r�ABk��t�:S�:S�Ͼ��:r%�bX�����Kı<�~�l? șı/������bX�%??����K5tL�ԛND�,K���6���O�)��"X�&g�w6��bX�%�ﻭ�"X�%���w�m9ı,O_u�R�u��5�֍�"X�%�|���iȖ%�bw>����K �"dO{�ܓiȖ%�b~���ND�,K���p�љ,̚���ֳZ�r%�g�D����m9ı,O{�ܓiȖ%�bw���ӑ,K�2&{���ӑ,K������
�&�tnWΟ�Jt�Jt�￿���Kİ��w���Ȗ%�b_{���r%�bX����m9ı,N�d��)�=��e�舍�b�u,7L���n�t�F��Ɔ��n�Wy��K���"X�%���w�ӑ,Kľ}�u��Kı/����r%�bX�{�NND�,K�ޛ�a��XL�d��h�r%�bX��~�bX�%�w[ND�,K�{��iȖ%�b{����O�:S�:_�}�l~º&tn�:�r%�bX��{�m9ı,O;�o�"X��Y#HmD6E �bn'߻��ӑ,K��;���r0���/'���i��LZ��a^�;�bY����|6��bX�'߻��ӑ,K��=����Kı/����r%�bX�����/]B�h��]ND�,K���ND�,K����ӑ,KĿ{��iȖ%�by߻xm9ı,O����3E��&k*���ש�XDZ�-�L �%��1B#)PԬf92%�.��4*�y���N��N�7߻�ND�,K��{��"X�%��~�2l?O"dK���p�r%�bX����Y�i�f�l��rwy�^B�{��i�6%�by߻̛ND�,K���ND�,K����ӑ?S"���c��YcvSD�����/!xX����,�r%�bX�����r%��DȞ����ND�,K��ߵ���N��N�=��c�"�vŹj�Ο�X�%���w�ӑ,K��=����Kı<ϻ��r%�`]���z���D��s�ɴ�Kı=>��;�:�)2��Z6��bX�'���ͧ"X�%������m<�bX�'����6��bX�'�}�ND�н>~>|W�Lb����-��	BS���2�%�F�>���nĂ�V��j���\�m9ı,O3��6��bX�'���ɴ�Kı=����<�bX�'���ͧ"X�%��t�K�՘Mr�ֵ��Kı<���M�"ؖ%���w�ӑ,K��=����Kı/�w��r'�L��,J~���$����h��՛ND�,K����"X�%��{�siȖ-�b_>�u��Kı<���ND�,K��O�.wYanh�ֳFӑ,K��=����Kı/�w��r%�bX�w��&ӑ,K����iȖ%�bt����gF ���|���^��^�����ӑ,K��w�6��bX�'���6��bX�'���ͧ"X�%�դy�P������t̕O5&H��B�h��]>q��P!�  Qw$h\ �g ��	�x�cHb!N4G~R0�e����8K��OO1p�)w���ݦy�yÚS�7,����H�dd��w�wK=l>|�
������sN�UU�G��j��+���n6��x�A�
�b3ά9�2	� /m�UO$Ku���^$7��8����Х�F�40�]1^)Q2zA���]ۍ�#��3�����B��kw0�{>��s�l�r/��`����pF�����[��,+I�%���S\�kFa�ۑO[��TsT���2�:wq�d8�.��yL���6��x���E����+��c�nJ.�:MJu��!5�-��f#�!�lN�Io���lҲ�K�m����@l,׬Tͮ��ك�n,�7&�x� B4s�N�iPN%��Ŏ^�
� 1A5�U��TV;5wjwl��.��ȬN�]M�tlS���u��Qɴ�Z��
g�����G����$ZZR�xk�.���S��@bN�1�̡��n�k�����F$IQ���Սq�l�v�0�Jp!����^�R�C
�Lȁ3��mq�1L<'��#�{Acz�tm�t�Ƃ�4J�+S5�S��ـwu��ʤs��8v��:T8�F��6�eqN�7+=��N�s+���G/Q�r�Ze��%��c���g����Z���\]����0��c���v�m�zX�;J0�%r"r���m���Y��,l5K8��bE��
�`�Z*d0/h�tk��3̺{NY��훘!����%���=��u�&�'�{t��4AI�#����ڷkL���H�]W/F��Z��I��X;g]oL��6.�0�-f�2�Utݔ3�񴁸���Ar�ӽ�^ei���e�H��Ƙ��R�D�����5Al�;ƕZ��%��wbm�J��n��S���&�ۂ]M������q�eN�Ժ��Һ�t��6�TЬ0,�==����ܓ���^��n�C��8���N{M'9�4-�R��Iv�P��gr�UR*�UU n�W]KJ�MV�d���z-u�2�T�QUT�M��Ư%��	�P�ePCgH��+���oXfaY�f��U5E6��Dx(�UO�I6)���R;S�_��|+�TOh����`�U�A=Wߥ��9��%֦Lɘm,�l����͵ѱ:J˸�p �f3��s�[�X���6���T��ڤ\�iN#cX��s��{vKN]�n�A�2����p1ST���#`�x���T���#���v゗����i�b����	�a�p��L�x����粀�"�Ѵ�쌖ٳ����6t�z�ui庮�v�[�M��*�mҲ�ۇ�f<^U��?���Ntލ���R�a����Ŷ����llvv�Mp9�h1Nͥ�Z�p��*�::h:�r��>)ҝ)�߿�d�r%�bX�����r%�bX�g�w6�H�"X�'���ٴ�K�/'�W�d��m(e^�;���/�{�ND�,K����ӑ,K��=�siȖ%�by߻̛ND�ș����~�ka��K�f�ӑ,K��>���r%�bX���m9ı,O;�y�iȖ%�b{�wٴ�B�/B�>�����#�|���ı,Os��6��bX�'���ɴ�Kı=����K��<�~�m9:S�:S��S����Zi�cL���Kı<���M�"X�%���fӑ,K��=����Kı=����)ҝ)������ �ʰ�ň��\�Ui�z�0��w&:v���x
��qAS�x5�kYc�<��t�Jt�O~����Kı<�~�m9ı,Os�w6�Ry"X�'����6��bX���{���.Ļ -��O�:S�����Ӑ���SN�X�'ٯ��ND�,K��,�r%�bX�{��m9ı,N���f��-������f�iȖ%�b{�����Kı<���ND�,K�{�ͧ"X�%�|�ߞ�;���/!y?���N�4�2�ֳiȖ%�by�{�6��bX�'��}�ND�,K����ӑ,K��~����ҝ)ҝ=�}ğ�����3Z՛ND�,K�{�ͧ"X�%�}���iȖ%�b{�����Kı;����_�z�,I��->*�B��)t�h[v}��u�K3=��=<�n��V��I�f w��r,��2�r����7�~0�-]]�]��V���7nE��+��$wg��}�� ;ݏ?$M�ԩz�c��O�h�k ����ც�Ur���x�r, �x��WjYL���M[��8`we��"��Už'����\J��Wĭ��fd��r,�ٕ�wc��J�~�[��8��pĎ�7&�s�̝�s�;ہ�X�0��>�#��֊S �������v2��p�"엀}$��iS�Nն�!6`�̬�*�������~S���;�� �ږUKn�]�WlM�ݎ]���p�;�:��O=��؊Bm. ��[�I��w7$���f�}=�f��O�	��� ��@=;D-��ܒs�e�/�MYB|�i�� �0�S+ �0�e��RK<���V�:It���7/Mι�ۑ�:]R�&�T˞K[��'���J�0.�6ګ�w��{+ �0�e��K�	8�V���2��M5n��ឯ�g��~��߿^�T��>�h�WěHm[0�e��K�6j�Xdp�6TTț�I"�WN���R�x�^��;#���%�cJ��luN���T��=\�����<����K�/�ڭ�U����RYP(K#ʠ�:�L�kn��D.o	7��vk�(��IG��0\�n��{T@nL�۬S�@�_cc`2�g�{Is���*�CJ(��F�ԙ!�b���+�`���Mhj��M]ctĠ$��/�8j)2A�Y�Ø��99n�'���r���V.\Y���S)n�0Z:�]�e���`����WOJ� �]�M}�;�����{���\�����p�ۧ`�-���ۣ���]e�P&�I�����`���;�?[��[%�� ���X���;E>+I�f�V�x�S+ ��vZ�<�e�n�M��� ��2��8��]�x�:$p������չX�� ��/ ղ^4�j��+���V���0���[���fV!'��kwl:	h
�X�������v%���^ő$�amݠf���&ˢ��ܞd� ����fW���;�?���>Ғ��3���y绮����Ӓ���G9UE�2���E�/=��*����`c�J�i�>[M��'���\0�J.�xv�X�Բ�Kj��WV�؛�r���ql�� ��z���Xa�+ ݣhqR�||�I�fd���l��;��z��k���bl&�m]3v�ea2�!,�e���֡t�;�F��H��.�޷i���;/�Xݙf��-�xȔ��@](�����&��3���q#d~0)=x�r,i�\�����t+�f��-�x{�O�|�$5v�6Y�����rB��V��vʶ�ـE�/ �nE�Mٖ`ݙXvTXSM�J�tջ�>[%�v,���+ �v^ hnԺ|WcC�EZt	�yr��ո�<�X��l�)�r�}���퍮.��n���7utX�e�ڷ�<���̬-�x�d�{jYH�ڤ�XZ��N��̬-�x�d�nŕ�nѴ8�S�>]���u�E�/ �l��Mز��̬ ��i]Gl�(��v�n���x݋+ ������r�UB�Q�!>���nI8|_fI���Z����v,��+�U�g��='��܋ �$J�;n��خ�e<���'���6�g��z�nd�\�ۙ�:��h�S��V����t]�� �� M����X��+ ���p���m�mݳ &�x�%���dp�;�����t���V�m����N�2��� &�x�KwwV�����w������� ���{�����6׬�W�T�WB-��`#� M��d� ��e`��9��Q�Ui��0eMPe���m��W�L=d��K�Q�Q*�n��M웙��H���$8Ț�׀�=�؄.!�M���M,s��Kɦ� +)��ֶVm�ԕ7Nv��{z�\�;gs=q�c���hF�%��Mdƙ�]����S���N��y�5�6ͫ��αò/P��v�,m�tG=5�:j��6`;,[����i����Z���"&�A���o�Iffp�!A,��J�+Y`nU�X㕝���ĝuY�l.w��%��D%�֮O�~����<wf# �0��u�B|�n�o 6H����F=�� &�x�JZ_�t�Jһo �و�6G ����4�j�Ej�,vрl�7c��<wf# ��QN�|m����`ݏ 6H�	݆V�8`P%��m���h���:��K޹њ+\�іd	e��`y֕�+s��F�������cd� ��e`#� M������ ��|b��	�V}�G���ć��cd�܁&1��$a��AN"�9��ɹ$��~��d� ����ʍ�HwI�i��8`ݏ 6H�	�V�*SUN�+��nـv< �#�&�YX��wm+��N��nݦ��Ix���I��|��� ����W'}|�O/�tGh=�3I^�藫���fN7=7[nq\N0��������ц������I啀l�7c��4�j�]��:T:t+�f�0nǀ�<n̳ �y��n�l�n�7c���l�;Ir��r��Q�"Aaii���h@�̖"�b "I�JB� H��Jn�� .��. k
�t��'��D�a�@��d̹�O7⚊��D����&2b\�!�T�S�h������s<�@�`2[	$�.+N��qF���r�y��i؛�dvP�MCa��8�����# �	�UC��&mp"�E�0#�B��X^�XM����!5:�ۯt%l-�����$)Y�2�ZZ�#
��c%B-��RF訕�6�W3 &e�|%�����bA�b@�Fa K�㕱	tT!��12����)I�{�aSd,��u���� ٳ<Ko���&��r��l�OD] ��$�!���@��C�P�A�Tب�(/��_|B*₁��wvnI�k�6V�@LtZWm�����)=�zO,��8`n��>�Y�ں��v�|e�x��+ �[��vG�uhm�J�c��.���v���k�k�����ql,��{�N�Q��b��
��I;H�6:����-�x�#�'vb0ԩMT;���I�f M���9�${� ��b0��wm]�4��ʷn�o 7dx��F�0nǀ|�J�6�+��U���wf# �7c���r�ATH���L���YIV��2HF ��!�UU"L��;��V��VP��wm�#�	� n��	ݘ�I���ػbkV��vNy��I�l��0n+��i5
<a�M5����kl*�.�\� ����;��$x�.*���vڱ�m��;��$x7c�W*�;�z�L���wlo��o ��b0d� &�x�G�on]�E\��	;cm��v< �#��9�/l���%z�Msʚ�t��m��	��S���l�)�'�}���<���!�d dI�y�wn�|=��.��X*�)\��l��vt�FS+���K�f��nk�1�`�D�ĺv��K:����ilȁq<�����W1�qq�Ĵ�,n�0��"�A�q��nYs4%�Ml6fb�m��l./A���#q�+{/f�t�w-�`��i�E���D��V!r@�nyҢ%@U�B���Tc�+moK���u2��r�z� p��ٺ�����}�ӧOy���ꎭ�f�Ֆ!L��v��)�g���F:��n@�dاp��$]iC��۴���ǀN��`$��W9�|���xQ�T�'�N��,�Wm��1�2�nǀ$x��\-X41'B�h�6I��v<=��8�=�<�=���)��Eg��ݲ�6�������	��N��`6e`8\T+ U��Mݷ�6<vLF�fV N�x���W��%q��S\Xa���876��v\�<:=��c10�ۈm��i�;"�e|ߞ��<f̬ ����|���x���+�l�jEi�}���$�(pN/wHT��ER�h�Z���:��jHB$��4�� �B@�ڄ�PmY�P��6��d���XApV#a��0Q�"H�,��b d����rݏ ���mJ�k�S\t���M�X6G�6<n�F�fV }�1��HWD�9�^��������t��# ٳ+ &���) �N�Yv��vb0�2�l� �6^6@�iۧe����ؑM��k�����]�����a=�� e��U�"r,I���1]�`6e`��l�n�F�Ȁu[�j�M� M��͏ ���lٕ�NK*R����ۦ�����7f#
UP���4/�{���'������X�*����-��Mو�6l��	�< �#�7c��EJ�K�����0�e`�/Oy�=�<n�F oV�M'L��� �i�L��J�R�942UB�U�Zf�f�1D��d(���'X��+��u�dx�G�Mو�6I��wm]\�wMݻV� l��݃�6I��dx�JT�U]2��ݷ�v �&V M����S����j�$ڶǀl�+ &��d�yς�Js�U\*�	FD�l%B�рD��D�ˊ������׳f���	��[t�ݔ�n�l� 6H�	��d�X�T��K��Z��Z�N�r�6ff���6Ƀ���l,�B�w�e�#,�1J�[��o�	�y�vX�2�l� �Ie�Y��؟-�� ����;�2�l� �l���z�ȼ��R�\E�WL��X�������7w�V���j���]Z.�m� M��-��	����+ >�ں���E���j��>[%�vXwfV>�ﵹ%G���1"��C�ӖJ���f�Z�i�!5��g3K)D5 "�mfHƦ����m�6�&@!�J��mn�1 	l@��^=���d'��`<�]�H��	n�i	�61j�]Tt"5Mth\u���t=gq���{�f{Zv^ea��ucqf��Ɔ�/+&.n���ܦ�����vzg�	βn1^3���l���O �y���U���6Gj��4��`�%�7�38��K��8��j���rr&���>�Et�;l�g	�эc,t����.Uw�=���ɀwve`���/ ٩�XA����LWc���+ &����x݆V{�H�sȦ��N��M�� ==�|�K�&�2��̬r\TK�+v��6�x�*��K�=��=��+ ����	�<��QR�X툾[V� �ٕx���+ &����x�����b֔��.vƤ:�4�Mԕ��*6�n�nS0��-5`�ŉCz��9�i��;�2�wc�>[%��2����P��*t��v�n�wcª����V�*��)�GS���fV�ٕ�ݵuq�Ěh��ڶ���x�̬=\�Kd�V {g� }R�m��5C�Rlm���s���v�	�~��	ݏ �l��l�MZ�]�	����ٕ����/ �ٕ�~�Us�OW�G�YVA6-�ɉe�^�)�kv��v�N�B��Vƺ��$pY�VwP�|�x�d�wfV�ٕ�Nn𞛎��`L��m���w_����ߺ����X;#�>�Ag,�_-޵��}�lܓ�=�f���Ƃb�0C	bĕ�f0$�����i�S��C
ܘ�(%P����T�U_�?~ߞ�s��7n]�EK�Wi1�X�fV N����XݙX�ki�S���VZ�M�X;#�?W9������V�ٕ�v��t���:@�<��8m%����ݜ���v烓�g�f(z��SD��5��Hu25���l�n̬{�+��o���ԡ~��t�M��o ��+?UW=��X��� N�y��s�������˻u�{g��vG�M� ��+ ��e�Z-���|v�� N����[�}�lܐ@pMP���X��&�v�ry���ح[���m��c�&���7�2�vG�j��EZ�q�V�������G��k����4s�cl�ĨʂE��^�W&75W�������2�vG���|���<B��y��������`�2�vG��7fV{�I���^`�+-]�m� ��� 'v<?��r���e`�y��m]\��m*nݫo 'v<wfV N�x�R^�� �=JZ�E��L�ۻ����X;���ǀ�=�+M��4!Ż$4}KÜ!����$$"�<Ē7��֐�Cu���I!}<4FXFF҈��ӌhd���7��&�ѻ��fg�57|�А5HS^)π8l7��O��<�Mi�iu�S�
�{���F��F��T��a�(�PUN���*|U���_{p�r?p�dG̉��of�`@8�OHl8��h�(R� B�HZ;�uS�ul�s��/q���!�x	Ô!w�$!2��q�#	�'!�-�!1�����'-%�<~7�� KZOY�:	�0�Ü'7�sza�5�Jճ��S^!sl<��Y�D� ��%�JK��UUuPhi٪����UUWj�P���b��(�v��mڦeU��s�d��Y�Kg���멨�EJ�`�R�к�GZ.nN��Ş6��[���:;M����h�nC�:�<��:��0ӊ��vi�A�L�+¦jv�aAv��-�b�a���,�US���g뚖�h8e9t'U���F�x���>7a�q��%T�P����K����\12]��$v�]�1�pS�#&����XV�-��i���f�.���Z%����N��d\ђF�;-̪�
e!�T�.��� G`�$�6Y]ћ.����)ا\�N++���p��.�1�7Z��h-H� 2���j�9�s�n[,.W�u��1jB���2mxQ��v|2^�`<p��af�nTզ�N�ܩ��ZY�2۷f�Dx�M��V3��D�XG����P��q�g��k�)h۩;rc���f0������6mB\҃^�ٺ��&T�\2N��h�;5��w�v,W!�M3ɞ_+��m�v
P�8��1�ա��15^������
�;cˇ'57.�R�uY� ��@�X�۞r��pu1��d�hFf�	i��!-�k+TS8bs��n�jR:=[����E�n��X֬�@eU4Ԥny��tO=�`���Ռb�z@r��;u1q�mrc���Pm��^]���jp�y#q�mm�A�*N˕;;P�;
f�e@�	RjQж�+1lAs�SZW\$Xh��Ti�GQ�A%nZ+4*�ҭF�Y���͇:��O4�e�g@�镝hn�}���@Z^ћ�U*��Ms�v�:��D:3qq�8�Qoiv��u�ވ�9z�i�M��N�x��m���$q�G,��(�I]��7i�܅v���c]['l���T�u�rU\����U�Ͷ�{<ڦ��#QM�,RfmM^�r��&�����v+���-��B�#�(*�A��ޥ��k5�z��ABȋ�������߾<J�* lU��P�4|�{⧁DpVs��9�E��˨xkr��݌�bF�.̀�F��)Pe!�Ld%�u���K3M�=����е$3B���.'�#���ƹ��K���V�Y�{oDN�h�!)�vѱ��Q%.��	�cq��8vj7���o	ˇK^*crP��<�Cn�ܗl����{�i��d\3�(�ll�[`�ɳ����k����q4��x���ㅃ�p�m��`���w�Ӭ�x}�4Muuڰ!;]���i3�Ӱ�]9�oV��]��qPvs=�mh��,�GA�Wn�d� 7v< ���I2�	9L.�ۦ��C�o 7v< ���I2�	�2��ު��e�n�U���	��ٕ��������	�� �����I�|i�x��O}X��V ov< �����"[H�m7XݙX�\�qM� {}焜�߶nI�S���Iffw	JRYtHS�ĕ��S�NsOa���X*��[��3)��n��:t����m��l��	��ٕ��|��{+ =��ߩ��Zi��:��ߞ���N��sӞ�/I ��&V7fV ov<�J[j�]0�iSm�o �l��&����ǀEݗ�lԝ�w�hwI4��`�2�{��n��>�2�	�ىЂ۫�wt�7X���r��W�O_�w��X�X�A'mU�:�m��&�Omɐvg00�Tݚ�	ZYc)؂�`���D�uj6�ժ��x[���̬vL�r��W�	�� �Ċ�ʥI;mU�v��M�X�X����e��,��`��m7X�X���8W1B���$EBE�9TU�Ur�+�);x�fV+�
w��t��U��:t�[��>����>�2�	�2�wm]��+i���J��	���vL� ��~��ړ���,���k*�m1C4��RP�Y�)R%kRfi�f,�1������)�j��>�2�	�2�{������'�h��$�-��Wn�	�2�ܮr�	�� ='��ٕ�M���E+i�v���n�{��n��>�2�	�2��٤�wuj���Um6��e�Mp�'d������9�]W.9� ���QeR������w�}6e`�e`�c�"���>Zj���]��@�r�hA���Ä�3��i݁2{������wlo���b����i�+i��l�V ov<.��+ ��Йt��*�u�ݏ ��/ �l��'ve`�ڻ�5v���vҶ�����̬?%���	�� >%UK��]�ջ�>��N����ǀEݗ�l��uq%e�,.۶ـN���=�r����[=x�\0��>�%_,j1c2��J��aQ���w
�t-��dc�=�����fy,\$�,�K�[+sЎ��秞�)�:2�t���.�?���O�<�f۴�A۞�<Jyk�e��1#umfਜ਼c���#�B��-B�ȼ�m���[b���h�v�������)�.HSY���d�猬�d�&
jd��WU'��ɷ@ 7)��I�܄�V��g�a�78إ�3Ye�f���=�'m`��6#uǫ�qa�i�Xe�-Y����|�ݗ�}6e`�2��ި[tn��i����ٕ�N����ǟ��\�Gv$x�*�'m��4�x}�wfV ov<.�v;T�AiЕ�l�'veg� �<�-����փPjƅuvU�v� 7�v^��wfV�UJ��y��;I������x�]J'�K����ǉ-h�����p��$[n%-�S��[=x�\0	ݙ^�Us���=B+���V�-�w�}5�2��L"��h�aX� �VD�T��-���+Q"�P�F%C *��~��rBl� >��S�J�J��U��v�0�̬Wv^�W����������6sSB�N�i�6����/ >���{�+ �m��t���Um7x���W}3��M���5we�~��i훕��6f��ˋ���k�R��nF��9#�{�lL�,�Cs;��Q�n��>�2��̬ �����ۖPJcN�M�� ����s������	�2��kJ	�!�]]�vݺ�	� }��*���EU�`�������ο{+ ��e`�m+�C�wI���x�\K��<�=��w�2�wc��G%ua˱���N���;ݙX;��ݑ����;t]�Vĝ�Z�`&��8v�t�;f�jJb��1S+6��*��9�/v+ĕ��cV���n�e`�ǀvG�N���:�6�UCum���f N�y��s��r��}�`{g����`o;]�x�tۦ�4�Ɛ}�68`�`�ǀ}�H��(����&6����r�{g��w�� N��*�\�_*����dx�v�P�j���m7X{0vG�jݗ�Mٕ�uj��|acT��8�Bw�e(�i��K�E��[�c�k�!E��"�6����4� S�;I+�e]�����x��xݙ[��U���� ��/�Ս�M�i6�[��	�2��p�	�~�9IOQ^��G0�؝ۼ�{+ �G ����e�"Nҹi[LAv5n�`~�s���x�o��wc��\^��Vռ�ث��n��t�6`� 7v<�fV��r�ɾ������-�� �:��`�
���cl��;u�����Uκ��ճ7,�Lm��ئt�֝t�h�Wb�lYe���#�h
����ѕw]\籫��[> y�<xNI���N4�v�"�C��Vl�a�d�,ԟ�c��SHJ�x�km\��krث�7�Ӎ��v)8m��9�D���]�#<�%�j�ȕ�+u�K5bi{s�{-�t�$�t�wI��ye�9�M��Ҹ8�fb���1��e�!X�6�]�I�s��c�;�(1��#M[xRz�͙X�8*�_ʪ퇔���	�"��T��v���n�͙X�8`�%��e��UUr�"o���1؄Վ�����y��5vK���~�*����x���X�*N1�I]+*�� ���[��͙X�p�	ժ҈��T���o &��W7��W�o��`�G��X��M]&�s{l4�Dc�z�i��m��.���6`"J�Yb��s�e|�}�xdp�� 7dxȓ.���6�.s<羾�=�t!Мt�;�D�@B@? .l���&�y���͙XWy.�P�M��j�M�����ٳ+ ��mlJ������V��s����߿~x���X�� 7�<�QMEEn���i[xf̬lp�5vK�	�<�UUR�EOSuMQbQ��Ry�ɷa׸H�s��JУ��њRf�V����#[sD������ǀj엀dxf̬�*U�V�]�M���x�#�;6e`�� 'v��%[V*n��j��� �ٕ��9EN֔QA��K���9c2ZjS+���jF6!9N?y%���!Pa��<+Ȟ�YN���7��ic.�n�!20�(I��b������X[�vj�CV%`�R^,	L���ƕ�	�� i�Μ�C�(q6/�na�f���c_2иBL��P��IRVl�c�(C�P&�IIV�(�0#����bsÁ�͗�R�B���h�+)m%��xA}&i�#��A�&�y}5����0���w�@��7� ��x��p�A6�����E:@U�!�� �;W�@=>Q>C��ˮr����g{LT�xʥ���N��m��fV�8`�%���%�Wp.�SJ�nݺ�6GWd� �#�;6e`I(UytRX����Xƅ�a��V�u�i�.�"�6�LfPE.�q��ة���tuS�>ߞ��vG�vl��;#��[R"�����b�x�#�;6e`�� ��/ ��)������|V�ٳ+ ���x�G�oc���hm&[V� �0]��vG��PE�Is�}�'��S髓IZ���jـj엀�<�fV�0��E�+��$RJ�X�ݍ	��MM-��`�j`E����O�R=ny/OKH��wt��c��w�$xf̬dp�5vK�>U4VA0�T];��ٳ+=ʮr�I�~0�޼ �G��s��$Oy�w�v��`�ݺ�=�?��xz�'��o���]�WJ	�Wn�ف�K�z����ٳ+ �8`U�"0-�'V�n�I��{߻ÒN���ܓ���f��D�U�� �T,��1���d�g�ܥr���B���ݖ��eN��u�f+*^Aꚃ*�ū��gQ�^p1B�r%�t��$q���-�6%�e"�-��qV0�2�C�`�*b3��-�ۋ7!O\��b:�w%�X1�b�n��f�V��L<5rܖ�=:s�W	�ݛN9�1��WV;q`����Xc�Q�5��=u��ט��Mm:݆T|���\��5��X�wOd�7N�%e���*C����{�����P,2F�"��R�H![v��i5l!��w������	5� ��/ 6lx�;DChi:j��j�`5� ��/ 7�<�fVڕ��A�V�+.�l�5vK��G�vl��;5� 'v���W���[������|�m����\0]�����ȩ���v��6^��Wd� ��x���<�U�+��6f�cU8�Y��鴅�آ�eɖ�j���n�r����ӵjۼ���x�#�*��UW�7�<�[�]�zЛ���4����{�M�@D�3ڮY=��krO�Ȱ��mVԈ����Iձ[� ݑ���a�%���E����E9j�5|w��m�{�W?g�,~����x�#�7��"黴��2۶���j엀�<��,���J]�t @-���v&GkB`�P�\9
�+֕՚�W\mK̷_�L��P�]�l��޼ ݑ�n��;#� n�u.�b��c��w��<��$yI��7�~0�%縑�OP��]]0��Ӷ��<�z��ᇕr�\�s�r��^^}� ����j�Wp��ZV��{�U�-����׀�<-�x�%m�Zt���I[0�%�ʤl� �v^�d��>P*F����c�WhN̑V�ҷD��\��)/V]U.�-��c����0fK��ϟ}x[%�wfV�x{MEe�����E�^{�H��e`S޼ ��{�o�C7v��w�wg���K����l��v�G�M+V���7X�UR��z��<���}�������������$��e�)[E�n��j������K�>�̬-���	2�-եcWƴqb٬�h.�W+E��hq�����fs��r�F	��2r��{~��x�ϳ+ ��^ }ݏ ݃Ue��+����V���� ��/ 7dx]�x�%mPI�J�Ӣ�]�xݑ��K�g� �y��%T�3�!��ح� n��������^���dE5�e�����Eݗ�z�{�W�{c���ʮ�Q�ª�(F
B �Go�]K&kZ�5m ���ݥ�7�Q!e0Ia�V� ��p�h��A�jbL1��a�A,s�%���jÉ�X���a�����>wUS��u�ۛ���m���\l<Ԣs���u�0FR�R�Z�Ś�̬��%L�\�MnzLrB�8��.7�O7�Ξa�i�2{5m�/����p���+2m	��zj���J��ܬ�x��� A�]K$����Xk-�v�L�,�(�m�l��Jp-���ђ��w\��	��>OO�v�gM�v���ݻ�	�߲�	����I��~=��շ����C5ګ0	��=\�s��y�S޼�L� ޭ��S�+�N��&� ݑ�n��;$��'c���Qw�ut��N�o �d��L�lp�����WT�ݤ�v� ����<-��	$
��������զ��xj����;	��n,��F�ؓ)�q\���Nt&�*��Fk��=����߲<.��8`�rNƐ�um]� 7dy�es���W*���|��Mp�'u�=T��"���Cv�J��<��^68`G �#�7�,%&��Vں��ۼlp�&� �#���s� �x�]�l�e�e����p�	�<n�`c���*~����~�:����@�M�%+cC��Zh��ˎ�̪u�g��63���N�ٺ�����	��`c�k�c��m����������z`�p�	�<vYv��Mڻ�I6� �0	���9��
+�T&ȵID	χ@�Nk�krO��~X�&�a7V��;��(�dx���qz{<`��{�3�!��ڻf�$���+��x�	<�`�_O �=����R�.��ѻd�V�Vu�j�
K��a��@G.�I>�c9CX�n�aN�SV� �8`�� �8`RK�7�.�@�ج�Z��ݎ�� ��/ ��,�9č�^=�ݻ)YiYvճ ����<K�`I��ޭ��S�wE�c`�0I�I2�=T�\��UQ�y� :m��t�N�o �v^$�X�p��<�چ��'C.Ĺ%�n5R��4�^�b���s�ɵ���E��\��r�U�.�l����}�x�`������{c��XW�7E�T�&� ���G�N�d�X����8e��f l���� �&V7\0���_ v������v8`$��&��Ix{j�n�M��e�� �0	��j�^;0�ͪ+j��]��Nk�@&��S	o�i4D�p�<��'���\4ĩ�]gC���B2HI�@��ˊ�o�#4������پ��=~P�>���# ȡ=�p�0���~¡F3�����3�n�)�b�&F�'���u��!�w�\5��_|�p�6f���d]� b!�K$űv
��n��}��o�O�j�yh!,i�S! ���_<���Z��A)���9����?���@�@�bń<�3�g���Pϔ�T׾�x��.hpj@����n��H�%���w}��5�%�'	.���Uc��� _1D�-������9�0��ra��9%�o@x��C�3zu�p�q.́��2��7�l �<vnFp�ǜ|���Q0����s���`�������",b�L]#��a�iM萉��
B$T̿��˙B��e@�!CZ�~���%�Uϑ�𫒑}|�����#	YtJ^p��%�IW>�H��MXքIe�����h�C�3����sfs9�
|�k交W���u��H��t>I��c�c}����+UU�R�i檪�.��j�����X�A9j2.���ۺ�eeU���9ኖ�yݚN�F6��'��#<�Rc%M �	���K/t��3ۑdrK؎F�<A#g��㨷g
�EF~��ƅC��[[t����1�:;?O���e)n�疒��B�[�gvf��mc:7ZQ�%7Vy��I��V{��xl�x�\�l�VۗBk���C�Љ�\�B��k]��%s�U�,��@��Xh��
��:�nK�\U�ҁl&�d�v$�5	v!䖨���'[���[�i�A����ͻ8���*��f�aYS�S�"����W+�%e7�l�
 ���
^�b�G�=v�%�`���f\���f�RRXf�ԍjf:8`(B�VG	N��fXa����y�r�:ބ3L���F��n��ᰇ��Lv�r��`�M��.���֤�.�YD-�UL\\�%%��kiw$���>�5qz{U#��Q�h�\4����"ㅅ�y+k��l!�M:�H�)�mu��:Y�gs�o)�u9��T��ad�X:Ь$ؓc�n�4�H�G,�2��k� m�x��ݻNhug�X���C��t�a�l�hd{[mذe�+h�W��*Pq(�Xݢ�.�+m�0��g�)�H1�;�h|�q[Kr۝�6݆��\.݊����9�蕎�`g֑c����]cP�5U����-����ح�m���/;��#q�mW\7R�:�'g@U��]�gT�䝷���୚ngT�cq�s�ã�pu*�ԫzU��P�b�]�9��� �*�1����ۤB���i!�̨���h}��^8 �bILNF	(�J���{K��H- �k����l#L�f��u�\9�<�3����$U[e�<��[dY֍*�Y�*R�\MU�@n��+�Fgm�j���5UU6$����5U�VZ.�d�ei��5LJ�TU-T��`J��2��!Y@^���I�Az���3n�6�MO��~�b �((t��*�Q�z/�� 
�ѡA8�$��zH�I'��zC�L��+�[y�$��-��[ni�t=11N0n���6,�rV6�r/bٸB�d�F��8EB�i�ֹ�^�v�1t�l��v���*�f5h��%״��,J��v�f�EJBţ;V�r�iv�D��^#��t�׫\0,Ԗ )H�O-�cf��$KF��jk����v	��Ŧ���3��aS2���aTp���=:J�)�|��.�"R��1#�Q�f����jl�;����c+#Fm�V��J�J�c�@?H��%��e`$��
u)�;��1�&�eȰ	�2��� ��ʺ	E��N�uv�Xf̬dp�7�� �$��R�$�]�.��[u�l��p�5I/ �ٕ�sv�	�.�e�ـl�eȰ�2��� ;R���&�����t	P4s��Uа�	�Q���tk
��=JY�׋
t����v� �G�lٕ�I0��l�C�qX5W�Ҷ�߽�f����a7	؃��N(�d����7$���nI>�ߵ��UImx<lcl�-��� ���l� �c�6l��>�HC��|Uv+-�ف�R��� =���6l����g� ���+�Rc�-�ـv<f̬v8`5� >6+%��-Τ�nm���YY�sXd��Yx��N���%Gh��ST&#V���� ��f�z��|��g� ���;��˻��|I��N�z�I���<�z���=�W8�NzQa�&�c2��ܓ��]��}|�������>U!����z`���o;́��;Wl��ǀM�� ��;0�T8�ՃU|M�o ���`�� 'dxޢ�U��Q`�K��@B���,#�.ԩ�B��D�A.Y����,�[��i�6˲�cl�&�;��Ix]�x{��2;w�Wb��V�w\0�������p�5V����ۺ-�ـ|�K�"���;��}��|�h�R"��N����?-��� ������w��!@�q
�@��b#*��9Y��|�����D]��ۡ;o ����� w�<�6P��`�:�X��q�g����S7��l����\#�����Ն�m�[��>|���܋ ;���rs`bIڧV鴮ـ}�"�U$�� �����U5�5t2�������a�K���{׀obi�v��c���o �u� �0�r, �#�7��C#�|Uv+-�ـM�ݹ M���`���s�F@�+��D�>���]d���qcwc����t�\c�-����n�8�f�i]�����j� 
y����G>1P���]ṙӶS�֭q���$ڂ��v�Lp&�Px�.�lu͙p]�՚�Q�+���su��� )+g���������c�5��<�r��B$@�sQW"��FԶ�L�h��i�7�N�1uE�iN�d�w�e�5u�K��D�we��eK�}���A2oxK���Ե��F�\��XؐƱ�-����qt�-�u�#u��xB`fՊ7-k��m���ӫm�H��\0	#��/��0t����dy��#v?����܋=ĉ+ɗug�V+V��ݷ�n�� �nE�ou� ��ŀ��Z�
�I[L�[0��X�\0��x�+���0	���ڧV�I��ou� �ݗ�}��}�"�$�nՓ�.G+r^]�o2��a��ƥ�11��xB\ �%�����N����3�o��:��mȰ�fV�bj��n�7lt��m`v8f�w�U\VK�� �ٕ�M�:j)�.�1Uج�ճ �r,�ٕ��r�/K�����j�Kl�)�n�*ݖ�X{{6�Xݎۑ`*�%Ԡ��:��0	�"�=U\�w}�>���w��J�YNӻ�unڴ;����yu�n�����c:�M*:5b�c:CA��ɣ�V�t�����`nE�oob��=/�X9��K¶�V�,V�mȰ��Xۑ`Mp�7g)F&��V���k ��ŀM�
�T����B�`�T��/>�_M���;8���WH.�0	��`Mp�'nE��UU)�<`�&�z�uv�ةX˶���`�"�7�2�	��`�EI��J�@؅���,[,B�XP�ʹ�]դ
���k[��]�K�C�c-U���V[� ����m�^��*�A�G� ��)e��U���ڶ��7�eg�\�G��� ���M��� &�a�V]��&܋ ��� �r,�ٕ�l55WvDUWI�v���r��\]�g����w�����^�=|��+���u�&��OX�Z-������ �r,��lp�>�p�=ʮ߂i���t���r��wmڎ[�������%ҳB�\�qRt�we;�����`c���mȰ	�LP�*-�t�� �0��{�_ ��y`nyg�#�j���M�iR��� ��M���� �0	���Um*���l�&܋ �\0	�e`z������ +b�]z�U���ڶ��&�68`�� �r,Vs���H�d�H1A!d �;t���'���Z9m�2�	Cq�ل�m�X�[�I�Bd��7T�EXڌ,�'5���	Ѯ���%�eMpA��Q��o;������MGO8���շ/����s�]g���M���lq�k[�s�֞]#�5�ja�]��9�r쪚W�+���N��AՆV���6�dqԢJ���3cx�=f&��hxN6��h;k�L��];������{j�B�b`+pMՌ�=f�'g�ͱ
���+\�s��^9�<�Ր&�a�E�π���X�p�&܋ ����e�ĕX���J�u�N�v�X�p�&����"[�m7le�l�'nE�M�n̬v8`NN)�C�ln�k�����H�`�� ��;��)|(�]2�[f7\0	��N܋ ��+o��ڂ�iں��ۡ�wEu��t�W.�9u1l4Gu�P���n�w8Jϲp���m[J���k�I~����ݼ�S!j��Wb����ȳ��(����s��8�E$�n�g��$إ�^�j�վ6ն��G� �v^;{;r,��$m"�0����f�v�,v�X�U/l��Jv����IX[����'ob�=������`l��I�0�͋�BuNf�ù���FD&�x�&����(+4HQűq���*uh�����mȰ	�p�"�/��m�,}�R=Ŕ�;���'u� �d�v�,mȰ	�MK�*�N�ˤQm����f�y��.�ܫ�CI�pV�GI�#��"mWBh�9`)��H;!���D�"�/��4F�{���sc�
B�����)��1�����<�492��*�L��h��֜!�XbC&d�[ks*�hhVS"�MG.����EA�C- �)H]fA1�B��C^���68or�I�q	LQ.B���F:�C���b��@�� ���#4m�1�smB9�l�0c�Z7"+ ����0#~`� �1Be���p��@�⧐)PBdqIs�)<fHb:>z8��&�����d@$Y�XC�<��lP�3e)��T���	)��u�r$h�&ȁ�kq�|�5�f�H���0�ZsD!4�	L��"Eؘ&� ��S��^"
m<3b��S���r<\P�	�0�<u���n�I���XJn�jƨ��n���ۑ`5��\^��^4�)�-X�Wb��t`nE�l�-������5r�e�����E�,E������o/\��<-4��k;��{B�V�[�|m�m��&V�xv9G�\�9_ ��y`hl�,V�	5G��-���r�mȰ�p�6�Uw�����%m�ݎQ�M�ݎ[%��ږ(ݍ�n�V�рM�ݎ[%�{�|�L D#�P�D���dV�X(a�-J%�"G$��zK�����S�y���UXv8`l��wc�`nE�z�_O����f���h�ӌ�<ó���f���m�]�v������3��J�lI��!6|��� ��(�&܋��s���~0lL��]4�`��i��;��o�l�����=���ܓ���f�*)Q�<�g��e*��Mۣ ��y`��E�^ݎQ�j�6��N�[嶭��=�s��{<`S޼�� �r, ���nҫt�j�%m�]�xv9F;{ݎ*�r�ÇI�]C٦��k�Wjm)��������ܝ&v�s������.�gc�Cceֺ4c��	��b���A[&pv��PtCK9�[Zp��`M��^.�継z�v8�Tqm�F)�p��y���J#a�0�1�Ku5�����X�׍	n�v���ػvqJ�Y� ��F޴'����w�3C���_�{;K']fUgNb&%x� �A1ZWv��'{=���m$Eͳ����ܶ��c��Ya�B$�سbR:G�ϷP��ٍM�W6�vV��J��<�F;{ݎ]�x�6X�;�l�RV��'ob�;�e`we�������G}�H�2������m`=�.��� ��� ��r��`&]2�V� ��/ ��(�'ob�7c�;����n��wv� �Q�N�ŀn�.� ���Twc�'@2�]������F��d1��:#tF�]v�VFgu�r2��J��Wt�t`��`�� ��/ �Q�uWME��wN���Vۻ�{���o<1XH��H�'�� |���'�׀}#�`��`MF�e��I"Ö�� ��/ �9F&�a�W���`��+��E�J�Ӧ���$�Q�I��e`M��sv�qջl�RV��$�n�`M��N�(�=ʥ��]/;��1�M���Why(�0�1�[iw%��*WDu�Dw�az�_[;-�j���E6^;�Q�I��S�v��.�t���)��	5�0M� �\0	52�1Э�
lwv� �\� �l�4CB�`�QKs���'����=�"+]�)UةS�t`M��onE�E�/ ��(�5WM�p��V�m���{r,ܪ�����`o�����Wh��4�Ō�˘�gّ4��݄��8�2���7D�(FYE����"엀vk�`ݏ �܋ �.+��lUv�������7c�5vK�"엀ȶ��V�j�I[� &�x��x]���r���H��T�N���]���%�����
�(���ʯ�wN�%������c�ړB��p.w�E�/ �W+}3�|�<�]���N�~���!�C��]&��L���5�J�M���`e��2�.e����[���n�}��5I/ ��/�ϐE�z�	�ȤcN픪�T�ݺ0RK�7�"�6\� ��(�r��H+��K�n�[�;�x۞X�p�>�r��IxR ���eRf��)���:���w��}��DN��Nĝ1[XݎQ�uI/ �ve`�"�>���qUp��"h-*�X#He�$!%,�to��/��q�T��2ns�6��=B3�B��C�=[��"��Z�sĽcR�kZ�-��[2��*\��$��Ɏj1�������H&���&�\�<U� ��Z��;�`r�Q�˃��:�ƈ�=�b��R��'�;�-��d�bV�&x�l���3BV�W������܌cV�s΅V��n�U����H�@]m��շ�ם���m����:I�H��1��.v%���6q/4<����t�2^[�2��l�t%�;�-��m[(V����x{�+ ����(�>�m"s-�S��;��;ݙXv8`v9Fղ^��j]�WM]_�]۬�0�� ��/ �ve`�,#h�aN�V��Q�ul��ove`��w���+J���;�Fղ^��+ ���� �U��;d�Ъ��Դ�QLJ��SE��5�X%M���']rT�@�<�%�Q����ٙ�WUo������Q�}�ذ����%�1-�������Ӵ�H~��*b�I�!�bhM"�	�ECr{��ܓ�g���{�n�	[{wH�ҺZ�0�r���ŀn���>�`j��(+��ڶP�р}�ذ�̬����(�>�m"V:):�MZm`ݙX���� ���`�lQ�]�fg�u9I2�2��6Y�R��Rb�M�36�6.ړJ�r�W3��}�Q�}�ذݙX{Z�a�J�h�M�f�Q�}�ذݙX��{Hq�j��ةS�t`v��'����τ�0��0&@w��}#�`*�K)[Un��c�w�n���;�� �G(�:�K�
��\��
VQe$��ݎ�9Fղ^ n�x��%O%�W��;�T��0���[�NB�Q)A�)���s�fQfq���vݑ�A���d����|�d� ��xv8`j��(��[j�V���[%�wc�;�� �l�x�ͤ9M'J�պv;w�|����p�>]�W�ul��w����Uҧw�|�� ���ݕxV�x�2 ^Y�r��\��TH))�ZX�Mj��ٹ�D�	Vċi��jـ|��� ��/ �we���{����b��<�S-�AV��.���	S��獷:��	U�R9n��ar�̙�!(�wm�Oz��v^ݎ�v��`U��r�n��6���ݗ�wc��c�`ۑ`BTWm�+(����ݎݎ%�wnE�|����kZ��E��YM�ف��W)w�����uwe����K�]][jƩ���;�"���׳��'���{��~P@U�AU�tAU�҂��@UȂ��_�P@UȢ�	��"�T"AP�,�B AP��T �T $U$,(�T" AP��B �T �UT$AP��P�B0T"�P�AP�B0T#BAP�AP�B)P�T"AP�)B*!B
�B"
AP�
 �AP���T"T"�@T �B T"�+B�P�T 0T"��B+B	BAP��T"�B*EP��P��T �BP��P�EP�B0	B0T"AP��T ��$B
AP�T"T"�T"�P�P�B1T"�T! AdEBAb�B �$B�U
@T!BDXEaP�T$BAP�EBAP�B$�BP�AdBDX�T T!P�BEP�BAd@T$P
�������AU�

��V� *�D_���W�� *��AU�*
�� ��� �����d�Mda�P�`�f�A@��̟\�|�T�v�S���:��t��@( �"�4�� @ ��  ��=�۪���N�l�*�34��&��%IS�E
��@��� 4(�U%$��f�e( ��Y���    ����@�44Qzėx�1��=���z�:�0��%���@�ϐo{�mgOO������gs|n�9t�    ޷��n�p�=�O�e]{�!��x�z�ٮ�IOgz+�o��ګ��XZ����٫�;kU \}H�%�� ��ч܅O��N�����wW���V�}��)�z��n��z��f[}�|C��i�糭7�}�O�7g ��p  �y�{}� �B�g�w��3G}�zkﻀ��:|���{>��u��_f�l<��|�HPR��
���{�K�|��}�>�P{�p z[�砠y�ն���(��y�@��p==�: y׳Uw�p�s�O��g�   �Δ�Ɣ�{���� {��JR����R�os��/=Cf�� 9٠R�� :Q��J;��zR� uF���� m�p))� s=���(�����v�N��w�s�����{)�����$z��������< .����{���[����My�t�`-�F���	�{C�{���m�  {��E44W�t�V�Z�#��{e��;���;����{�˽`;�}�޽���wq�<�^��{��������J�À  ���O'{�)w#Ӽ�{�O��t=����{�}�!Yoxy�A���{c���\ "~�Jm�JR   ��U*T��� d��'�J���T@ j{MTSb�H  ��T���)P  ԥ4� h�OQ?�����k������y�O�ﴹ�����W��_�( *�APES�� *�저���V�"��zO������ٽ�K��7���0�Iф02��n���7,Ա��B�g��M/���[|8,��J�&g+���)�Q���_Wi��:{��|)e>P���_�{�\%���}��|vO���!c���.H�t �X2$#$F29�f������d�#"Y0�"I�̗^��=w�</����[�RI"d+	��M���q`b�=.�S9쐦����e�N��t^2�#ynRJ��$���xCe�>��L$�ЁX�13!an��3�ϒz�+\^���u�o�d&�>�1��`�IIB��B����@Je+h*A���YPR����e8��[��q"M넦kxKtM�����p�4]��乼��H^^rk{<)��xal�$5�֒<!vj\�]g�\���y�n;�r�xo^]y��/ך	Jz��<&B�L��7�|�ao�̄��&����ϒ�4����F&�I�e�d����u�Y-����ݺYe��I�F�f�I�\����1�
&A�#��$|)�� ���&���vj�F���!nh�f��˸�섺Bk%�T�3����.����ⷙ�?%�!��Vs�?�'��b�%��Ź���.�����jRI��b�����z7WTKol�
�\�v��t簉��s5f���y�ZB0��R|(��\+;��W�(��Sk���_*," H�I��57�\��o�.ȖD���7�ny���<׾�6�rVVT��������5��ٟ�2�hd�����\���ͥaj�߭2�|�R!�a�)<�FB��@�M|-�Y5�]�fI���V�$�Z��1�h��iH�	���	c#y�Ha{id��Q�Қ^^$��x�ǐ��
d�z�6�F1��Bj[�rh��ߔ�Ֆ�.X�h����LA]yԻvw�u��Pe1,��0s6BMo�xSp̖˼M���u������	F0to9!<��$(KL)R���ܵ�aYIqÕ��Md�n��\��%�����(k�=���s�1JL������N�)	8@�xa�����5�#IB�2ʑ���M����k.��e��p�h�	D�Ñ��o�����X�5���������Y��J�*�+��ۼ�e�fq.��ͣ�Ra2F�(X!d�נo����~#	a	R!YI[��B�!�Q�ܺ�3DR�di��]h��1qaH HɁ�q.j�Y�ك�B�5���¬��n���#�)�ٽ��#�$f�%ɜ!L
��.��A��u�S٣��g!t�.�|va@ӫ��d�����fc���&�����c%
|D�B$)$�Ő0�H1�	e���NRP<�XX!BZs9J��<�(dd�$�¸I=6����-V��B���Fŭ�!`Di$-!	8YM��:���*�˹n]���y�!�=�ס����^���#�eX�GO)��V$B$mZZ��Z�,�:�9E�	R��0��Bo=l8V8��7Y��f�dp8r�l����#ѻ���ڤ�V�pri��B@�0�0�	���������%��7���5C�=���Ȓe2cZ,0	q�M��Gq�����K�$כ䬲@��	����Ol)��9	��g�-�s���������9��9�@ߧ�`�Y��,��s!~y�h� O5��6����re�)��Fy7�y����7�;��9��?]�s>٨xʓ2�����E�q�5"�}��QL�����V�:!dޗ����C���g���n繨e}"��4�AM���ڼ�3=�	N���8�`]_�y��T�
�0�\Ԅ歅���#�5�0*Jh��S
����<.n��1)S������	�g��GÒ&����r�ܚ۹5^z�|w>����t[Y�۴JuG
gc�L����"���d!Ime���mc�t�Y��d��)�A(��	,�߻�s���zq��D%0� 2�B��#a	k���ޱ��:����9�ɫ�!��А�)&�~���=&�ybs��Z89����y��J{�7������O-%,�]��k[.��O_�c���*ʡ�
�ğO�}����uݠӗ��C,�f���&k0��J��b�&���R�p�˚xCD!
���ZYYa�f�]�I��#�Z��ߞy�����K�e1�L�B��0�Xf���Sa�MkL!!�i2$	g��9^k^i�M�z�5����3/.��.�硴�6q��	~W��9���S�� O'�±jF�$*�k�#�of�2N'�7��X�#cHR%�Q��e�k8��)�sW�!�ԀE�2���9�bP�NkDԺ����~C�\�B\�d�G� ��W<�4�6�B,)>X�0�,VX�H�E��Z�ā�\ap�oD)�j%a%e�K���
�J$�B0*BS{�������ύ�։H����<r����$ hufƾ~���jo�+f*��˞ZOה?�rG��=@3�{��*�h!�A��s߼���&������JjQ�4F�
o�>��n�a.���a�S���S'ľ�х���݋�9�Iy�fA/	��JCi�Aw����.�5�h�fr�r����M�qx�߳V\ן��5f���%�)V���k{�g%,��P���c`�,BA�%9�M[ B�į�����Y7
�0�aq!u�2����L	`cB���a3R`D�dq��#HR$�a��d��L2Q(1V8�HH�����1fBMfo\.�Čb]	��Vl�%��)%#!Ia�)���0%�۽�F�ސ�.B��!��a	BЙ�Ӑ�,�C� @�=% ZRS���Y���s�+EJ�@Ef*�e)�Xa	hOp��9�Cg.sH F$B.ݐ�����M��h���5Ni��xo����BOO|כٰ�p.��f�W4r%bP�a��ֳ�\5��rh�vB' I@�#d�� ����'����Om��k��39u�2f�C\$�Қ��g��֐�f�RF��n��{��^l��k͜��,�$��I%i�����Ɛ��I;�[��4�'4��SY�L�:�^G�w�F�m��S��@�B6)5�{�bX���@C��4�zMa2re�]���/7o</>��s���gǃ
�*��A,�0�R2�<n&������y
g���h!tm l���״3��A��%¸,h��*D�����#!�Im�)4Jd�B��4)	�
��p�0lK���	I"���a$�ցH�$�D�>Cʄj�=��
0.���=�9�W��:I'!�I��߿s�0v0�C��`�d*���!�	c&�9o��w黲]]��)���e!	��Mp��l�old%ނC
`.f㛾�NB0���T�	�у#_n�I)
D�g'�d�oVjxo\$�o�� C��ۡ�%#
��*D�
�����J��
�0j�>@�e��d
��6��1Ԑ��@��B!B4�c	r��#l�����	4!XR���d�HXSDK5�32��r&�ޙ�@����P��!���}�c2С�%���=\4Z�'2a���<�_}���K������+
,+-Ke���["KD��9�����hd id�4��H
}I����K�ixI�bm��d�H������O|���Ҳ� FHg�m5��G�g5<-֦hּ<f�sz�ЈBdp�I��	l�����0`c,�d�:78Mp�z!$`!��F5`P�Pw"H�l$�*8B��\��W��95�5��ap�Iw$�"H���J��4��"K.�%%�4	#R8²�\&�H�!"@���+*HE��@���,R���9�320���2g��=�2��q��4<<�4	��'5Ü��c�C�{�I�0�|�oW6�ɮ$"ܛ���ȗ�eփ^jɧ����}=��#J��(��
�B���$	0c�Vb�
����5�n{�[&��5���覌�n�f��M���L�Khw��S�jK����|e���5�3w9|��y��&�sl���wFK�f�p����w
Ra�7m]�Jfp��5���1"i�9�̔��L5�LͲ�&7�p\�y=�p�s���ޟ��D}���ц�p�.]�����|皧
�t�2��>Fg>��370�l�*�ʅJRK�殥)(@�Ɍ0��5}��_��F1J�=!�p�z� �AF�BJ22�$a,�%��5�����0���I̦��O%�"BF6$��f�$޹��ͬ5�20� I\3�����V	��򮌣��~�y�<�5�7�L�E���#p�#�����\�.�|�'�d��g$&�G�����m�UI@i�9C��)�J���l�^���=�}��g�
0$d�VP��9�3�5�x��,FI��nkZ�X5��XF%H@%d�km��R�7�������`OC)_R2�)hhJS73́�ĊA�����C4��dA����5��>�����5�b"�KJ�@ Ā2I"��HF�!dH�"@#�a�l
%޹5��$M�秄Jf�1��$,��w}��))�]�7>�B���g�p�j�s�%$HI�%&,�(�2R��F��M�0�ۓ{�����f��V���)5�{�,��2 ��l��h�#4�`Nn��!�;C�7�}���8񻎸�BB���6�3�>8B�3XL�%�l!�כ�XB�C-�{�Fo�a�Ӡ���T�e�\q.,)(q�D!�.�u��V]�aaI"H��0���4A�(L�M4�y)S�O4LC�0q��T'���������ܪ�*�ث�UUUUUUUUUUUb��(UR�UUUUUTUUUUUWUUUUUUUR�J��UUUUUUUUU�V�T�3UUUUUT�APUUzU�UU����j����UUUUUU
�����UTUUUj
���U���T�µW]Tv�U�j�)�&UƄv��g��n�%�Z�;�l��J��˷J�Oh��ABzv�����ջ�ġg��@�g� yo��1�m�
�(1[ �UV�R��R�:���Uuӭ5+��Ū��s8ĭJ�r:
�:4	E�Ү�½WQJi`��Oc70UT�N�*�mT���v!��ܫ�Q�b��sGj�^�{�}|����UUUкcvxe��eh+���Z�j���gA�*ڪ�j��jX5�7\�UT�UUmUUUZW�TNF�+h�\���U�`g��-�vNiV�V�"�Iړ#k���͊ګڵV�Jɨm-��W�<��g�M� ��qj<	ImU���Rۭ�@�B�+r�r���c�KU|�|�r�E�B���.���+�=�n@ ��قU��<��:�2�U�T�U��9c9mP����$C*����N
j�H�,go]R�q�*��@z��}w|m���*��d����᪪�=GUU!����WS�*�IB�j�
�j���I悗����2�l*�*�v
"�g�
�����
��c�X�y�p`M`r��r�q˧����Q��%7�E̦`j��2�U�]:~�����u��5*�Q�n���&
�VN�A��;�K}:�i�`�X͙	��c�������u@�����z�WA �Rk��e�T��m����_,��n����&ȸy��K�l \�'mФ��j:�n�A۝��b��W7��[��t"��a��*�T�ۊ{g��!ĖPx.o �65Fʠ�-+n�v���Y\tsю^�t6imWKVi]C��Ƙ�A�]�W���i�Ә�6-v��Qٸ�y[���7i��V��]����U����]��LS�N8���(kq�l
�X�j1�K�U�W]��ZU�����S�@�bfڲ��F���n�F[Ĝ�#j���s�-@��va�u�p��D�q��+-ml�r�� �ڪ�]>�{5S�]��:6������:� k��Z�.1¼���e�ь�^(��5��W�-�7/\r.ڣ�ӆS4�7�)�M�1��KhH�`��b�]����끷R�Ħ5��UU�L�[s1TqX�f��ə��6��� �Qq�ۍ���r��k����v����oU+¨شtlm��l
J�Eڲ��f��+q� 	:0��[��7+��$�UC�s�AU[o�C�Z���#K������G��IHp�L��������5Ð�x��bἐ\��`��U�1��#ҨV�nPyimt���Xuk���]Y�=`N�U�ՠ��K�˴mEC��Jᶍ�cn�ڹȴ����;�3�c�m�U[b�8@��o/*T�����aGq�N�@JUp���nvEn�1��L���u�>���V���$v�P����gdyKcr{EJ�媕yV��
V��rb��v��u���
+FN��Y'R��rۭ=5R���w*�(rl��r��v���n�^U�b����U/-\wo#��8���$)p�*��!0�����"�2�f"a�:ͩ�������32�u�[j���U�j��ƒ��Vՠ5���b�WZ�X;j�<��c�"��AT�rgM=�&��ʪW@tH/jv4>�U�U�eYIj�����
�m��W7�����̶��ei^9� ���;M�-J <d����eeeM��4���499�����Jq�ҭ�����[R�8ҫT�uKS�6�bF�ح�T�,����l� ��Q�T��ڌU��Iӗ�p�^�	pq�G%�n:ٹ�	V�d��m��b�v�#/n�kʵa��1��X��5\nC�=m��e�+]� �heF�c��J�Rg]Ó��CBw9���^K��.�ܼ;�sv��j���]��C�U�c�]��Yg�\�gzV��j���m]j�(4�;`�ʝ �����ƹ��yN�[QYՑ��X2f�b^�ۮ.��T�W�]O|R��R��m]M��j����UUl��*�FCJWK��̜Rq6�lU@V��6���p m���W'j�sW\�B�z�\�L�@�������h	ڪ���y�PZ �k�	7-AUUW�]]UT8�ZD�BK;	����ێ�:9�<>�x+h:��ք�6�`���u˨�s��Ũ�������g�
=��^��PJ�q�;��5�(-UW�N~G��Gmg�
��kUJ��	1t9m��X��s-N+ ��T�l1GA]
���}�~��Uyr��8B����n�C� qKU�Upm��WR�û!+*�RŞenZ��I�;%��U]UWT���Z��jک��27�_��"�X�m@/(����t�ܽ��
�W�����kQJ�UAKHt�P�樮��
�֪����#���Z���Y!�i�z
��I�xTցU���*V�Uk9j�	V��ڦ�]UG^&z���/��# ��U�Ka����@PUUUU�U��63�B���[E����|��UT�UTpUZ�Urql1�3�6�j{\^����Z����@J�P�9�,�nQ��W�������_���Xۍ�R�‪���\�KUT�&�j�Z�����lVi�1��6��A=U6�4�nKQ�cMq��5I�O!�=�UAW���J�ʵUUUv��C��-�`�
�����l�*�@-�����UUUj�
���
����������U����J�uDi*�*�*�V���kv�z��ڊ*���������
Z�����
���T*ָ�0�U����	��A�UP�]�UV�[uL�e�(�ٴTL�cj��*�V꠨\ʴ�U]UUR�qgfT
�j�����h
������
mUUUUUUUUU�S�5U5UUU����Pm���*��j�y�V���5IZ�V�ڀ�ѪM��V��畀�2��]�`��m�檪�]�Z�HZ���������U���V����(��^�kX�ɹ\q#m���@ʵUTx+�mT5@UUU\�UcM��A�6*�YZ�Ur�[@����j���!-UuFK��^��5Uu��Y����ö��AT����������*��a���Qڀm�z��@m*�UUJ�J�PQzX�ee[�X	"n����� ��6˵�9�U\�p
�l]HM��j��;q"MZP�PA5h6ն��lH��u��m\��;c�,�[U�UR�s�TUUUG�].2�uQ��Δ U�xlbڼhvZ�X
U��UWWUJ�UUT��]luf�� �2iyj�����:�UUUUUUPU*�WRqA.R����
ݺ�Y媠*��s��j�EUPqUU*Խ9`%y�nu�<�ī��Pp��8��F`f�r�5����Ty��V��6�*�T���US�ڂ���S��mUUV�X�2���H Ok��1��y�ڠ�	����UU[!sWj��i��^��T��P3i�:$�v�h٨S�iYt��
�ęB�/PR�W+$�V��UUU)ѐg���܌���V������7\GY�b��jY_*�
��n��۶��ȹT�5�{!��,��Y+�=���	�(�ݵE�骞Uc�O%̬cAE�YB٥s.^�RE��`�/\;N+�7oB�Yc\ƶUR�\*L�\��^�4�5(M",�X�Z+�N8gu\����U`xuCi��OY�nͥ9��gB��i���jn�	�aE;�\������QPbn�b�ҭV����8���P-t�R��n���I����.zrn��N�[�TR�	���j7���^^Vt�Gh�٘�[�k*b�+5]���L��G*q[5��5u�sWlԭ���Z��h��#UUqN{j*�bW��R���iIlk���[e�4�UUT2G"a�5���]�SSUT��WP;{A�U��UZ��_v�j����ݮL�UUg�mUUF;pX�l�
�U��ڭ��<5UT�@��>�����h+Q�//S�)bZ(�������Uꂸ���TUZ�u0A�PHU�f������LòdYU�*WV)��uN�t�t��+!*���;�ٱ��!�WU��ƸV��Ƹ�p��R����ө��s�&v����
�p=U@UO`�ԯ��y�U���'FުU�V����F��>�UU�j�������j�����S�q����_���[�SUR�UT��etUmk�eve٪�
�*�.�mT�۴�UR��T�UT� 4���*�UA�A2��mf���EUb����������U@6����55]E.��J��UR�5T\��HJ�UU*�T+�=8g��csd8(Z��������߶�ﾥP⪪���������)cTT�vݬuH(TSr�AU-T�����Z�
���U��
�����
�
����Z�-UT�p*�*���
�UUUUUUUU���[[V�1��U��X��U���V������X*���RU�U���e��h�PU��ХZ�V^��ەft�UTغ*�v��]v�(J�P{-�a�UUUK�=,�k���UYV�v9<��s<S�p����� �nt����>��UV��e%ڲ��DJ�M�n�0N��ɨMv9e ���pV���"�?(�W���D8 �P �j��!_�� �"HH� ABv���@�[$�!�N 	��x(`!�ljHT��^*8 ��)��!M��W�)ਞ�x�&��SN�q�6�z�x�M:0��|EO��
��#`8qJ��)�mA�#"�U=8
| �x���O��6+>� �H�`����'�WE}P�_TU7��BA�B����d+>CPҔ��!� �#�S�����4x� |��>t( �� B*�  ��PE|P�� {Q���>�	�G���P�`� ��@�ֆ*������`*�XQw��8��">�p@�z��_TW`���	� ,v�"��BE$Fߠ���'@��q4`��R&��_O�<uꀏ�G�Q`��7(�G�B
�Ͽ��G���x�	���|��B0�H�Z"x!@���.x���@��� R�TT @"�R(�b�x���|��b����1C$d �����!��L�:!�m ��+,!"���a	J"V�!�E�R�F�������#!)
BX4��A#��) �
T�FQ�@�@�$,� ���	�dnǈ��m
 �L!"H���"���x��T�^	����5*�`h���~�+CI�+��AU�W���, E���B�
�"�b��H�.�D�V
EaM��"AȥX��k�����qU\��SiV�%YPk��Z�UUKX�sv�ⵅ#�[7� V��Gi��yꑣT��g� ��xyi�khdj�cgx�A���j�΋�s;/�|���&N�Tc�y�rf�s�tPu�]�T��5�Z��xֹչ��V��Λ\QU�� k' �PL;�$�s���X�w�����z�/C'��{j����L$�Z�6 ��fC@�Q��q�w�Xy=���K���gGYႇ�Y��:ܺ4�*b��-*��!ʵGY�"e�nV9x�B-�m�¸�ύ�9��˝mɸ��eݙÀt�"�6��$W��`
���IY�i8�2kv�H6z:B
ݏm�r�%K��q�'+@ˍku=M�'�vh'G9��ͫ/��`�������=�ь�z�vzvlnV����Q���9�3�gh�0i��;(7]�
%�1݆�=#kpT�5S��yN�/{m��h�̼qd��i�T����fz{f:��Rca�ͳ��E!���l`�s�SDu�n�re\�[e�S�\�n[8ٕ�LM��
��6N���.^2��<��%��m� 9��h^jtUUJ�d�v��n̡PUB�����]���J���LTԠ-J�ڧ�ɑ� �t2���a,�[Z��e�hr���c�.�]`\"�u 5[��,�e:|7S6������`D�<v��i��v �T)p�L�mYF�b��K��Ʌ��ųI���X�F���e�y�*����']M��=��X�l��v��@n�$x��˒�kZwU�l��7�F��:������(^�f���X�&4X��f�&�bF��A��5r��U�[:x0�cb�@L��\˛�v�����l�pA�+\8<����clq�j�@�¥W8�K�t9�C�t�-U]Xs<�M����*j*��:���'64g���@�l.ŭX�j���W-9�v��rc��b�0�b�E#^6ǋ.��9��h���]8��ᯄ�T@�Q�C�ρb��x(��= �+��F�.O���م1�㱛�O8�맮��ݐ�bR$u���������t���n��+z��25k{1�0mV�^F�]vV83Mn+m����q�Z���۱��^9��n^.q�D�4iũ���{AȬث��=M�p!���{iV-C�6�� ��A��Yu)k�1��Q��e����2�K#�2��ss�jm� c˲��`�X-�rI	�D��.�L���)0�̹�e�=��x���q�.]�.��YM.��D���� ~���u��7�~0���e�N�MJ�ۼ �IJ�H�x�p�"움{�5��:R�]6^ w��x�p���r�������<�q��j�V���M�]�x�H�6��c�"����l��we�`vK�	�#�	�ݎ��\�?��<����c�m�f�.m�&Q�:��4��n;�0�6�O��K�v�-��e{� &�xv8`vK���;)���T;n�� ���g+�CS���:���o]��uM��v�xk��.զ�Ъݧm���I wjG�ݏ ݽ�]|�i.v� >� >��x��x�*�wfx�%W�{-�ZC��+�o >��x����������K�Bw�j��c��ĭ�[�<���z��vn�S��^��Iaw�8��uD9��87j��� l�x�� �dx˻R���6˺���ZBV���>�`]�x�� }�z�\�H�yQ�t�Z.�����V�׀wH��#"?@�Jʀ���w���R6n��7�۫M� ��G���� }$xݭ#�j��ۤ��� ov<�� ��< ����"��-��QI:|��ָ����w���(G�:-�v�h�N9���3�p�λ�MӤ��N��>�`�#��j< ��x{p��*�V��v�f }�<�r�����W� l�x{�y6�[��;)�m�ݕ n�x{����c�����FZ�t��RM�Wj� ����\0�#��9�E6����s����$��~.}r�jĭ]��w��I }�Q��x�O>�������*�b���^|v����-����kJ����q�Z-y)ny�͎��BWh�΀o�ߞ }�Q�����ϐn�� ��x��-��]�M� ����ݏ �u� >�<��H�֓��M� wwM� ��x��=�RGg���<wU9n���n�%V�v���T�&x��y���< ��x{p��,)Ji.v�f }�< ��G�ݏ �u� �9��Um`��I�����v�fP�M�]��n����V�3�]t�n�n�Yc���+%���Y����8��:<�aQ�#�M�*��к79i]�q��\�]�cP���r�D� *��lp�zA�\������D!�L'�ۜks�E��h�7�@`۶��d�;j謀
���wrq�CE��xǛ��5].�l�� D'��7Ne��S
SEQ���b��y'�o=�=X�w���^�M���p�N5pjŞ�����d.wZ{'<i�^��F��vjۀ�<�wc�>�p��� ���{��kL�6�/ =�޼�rlwc�����[v�;,�R��n��X���������ݭ� 7v<�b������]�`z�Uʤ��y�v�� n�xݽ� 7U|bo��i��v�< ݑ�v�, ����Us|5���7wv*��p	r���)�!���Lg]�B�ݷn8�8v}dV�R�%5](;h��{�� ���`d���s�v����m�wmդ�N�m�v�,�}Á^�8.z�E��-$�)�9h`ZB�*��!
 ���[�`���<�{����� n���o���M%®ն�}�< ����� ���`s�*^+hbl�Jշ���+��}ڞx����ob����"�m؊-ګ��o 7dx{{�R�{���Ͼx���	�܁P��)��n+�틜�����۩��=�l Ru-��e�Kfm:�ڵm���� ;$x�jG��<�b�D�˰ub�����G�v�x�#�;�ذz��[M�)[��m�ݩ n��]}IV�W*���y vH��ԦSj����o 7dx{{ vH��ԏ �vc��;Wm$!Ӵ�x{{ vH��ԏ 7dxݎN��h<�,�=Ze۫�zݝ���]<H��GB�[�f
�@C����-o�?2G�v�x�#�;�ذ�ڔ�Qn��IZ���ԏ 7dx{{ ~�z��<���1o�dʒ���闀{� �ob�� }ڑ�v3��U��e%v����;�ذ�G�'<>�[� �C�|@�	��s7Wb-B��ؕZ�cm`d� �9T���?��{׀w��`��6��c�折�LH�k>�p΢��⸇����ct��4A������:�������d���� ;$xejS)��V�b��m��K�;�ذ�G�v�x{tէi[�ۼ��� ;$x�jG�j�/ ��E�)ƒ�e�k ;$x�jG�j�/ �u� ���N0�WC��E�o >�H�[%��`d� �qr�P! F(� �)"!"�H!����wD�,���L�5nŇ�+Z��zZ殃3��v�u�6� �6Q8�n�\�75�7NR��x4��k�kRw9f'
*��Y��3�kWQ��\5�=�u��h��.���# �zNfEc��1�u���n���\R�@c6iB�V�Uu�c�|����Law&́�y�ã�gp��۞,L�Kf���kc3lv&�t���{�s���߃���{�B�i�.�O
C�v��僒��u�:�x�v��7*��6|��Kue*��Z�������\0�G�v�x݌�d�N�(Wwui��;�p�� }ڑ��K�:�"�A��V+�պ�� Nԏ ղ^7fV oUm\m�����]�M� ���d�n�`w�)#�>ډK�*.���.�鷀j�/ ���#�	ڑ�)"�CO�WB�&CN���=��[�=�׈��Qz�;v�tSW&��]�;�N ~�z�v���\��E=��"<��aK�h��L�M��V�{��~�H�# @%D��!�,��� �ξ��"�/ ���ڔ�ˡ�e"շ��#�5I/ ���G�M�K�m�Z����շ�j�^7\0��x;R<v3���6Ң��Sv�7\0	��˗��#�;��`���/�c���WtRT�,���;�Kuluvn!)��Iۮ�����:�
c�����>�{׀�#�:�f��ק ?~�ٻ�ؕ��ó�;R<�)#T���?�n{ןW)"i^Kל\�����N�`���w_M���z�~ׯ�α7�(E�J��H�ID�İH��+�ad	��WI��)��B��]���le%c[>�i�r-9���HX%�F!�A��˻�8ʒNe��0�m�c�&��t� Lc��&m޹�dԒ�^c7�Md3D��$R�t�R�e�Ս	X��SK�\@�p�4���).϶����y�޹�˛Rp�O~8|2{..Vf�0�L�bnO0���N#����R���h�M���^fQ#,�W.$�����	�HR%�`L��jHa	Ij���%{��B�~y|����>c��0�X�IFR�*B!�a��NC�!�
]!xN�1���.e�J<&P�����V1��aF,P���$HB �`Ќ`}�	ik�oX��	)_Nf�Z�&�5�<apR��}�}ᣌ�*@��$��f��RQ��b��s����	�2�(J��.9`yWA�!f�y��	M��MR�Kn@�`	���	17@Ȑ�F+t�3"R#���M=R-��{�7��%B1���O�w���S��q#B �i�ղ���u�("��V�h7���4p�)v0-�i�)�C�Da+m%!��ᐊ�Q��T 0 T������WV,�+(F)1$�!=tCc���e�����)()�x�'��\D==C�6 eUF(��tm=\"��(�B(��� ,������"��g��b;P�D"||+���8��b��}�nI=���n�;��N�[�Wm�7\0��x;R<U-�=xG��,){���f l����y�^�� ��Ӏw��eܕ�<�7.�f�M�;d2.u]uyc�W]71��6��]V�>��Ns8n;*�m��y��7\?UrO���߾��������
��a&4���z�#�?�{� &�G��U$o��U��E�ڶ����� $���$zJ��{�x˱��Wi+-6`{����< ���H�� B1�TBЅ�BE1P$@l[�Sk��O����߼��[o��>�a�X�%��oj,��ʯ�U\�~���~� ��@'����X���0���4д�!J���v.v�$���^�ٮ�w�H��smQ$4]�_ I?<v8`�<m�E�컨�N�[bT�v�x�p�	$x�ڋ $���RF�Ǭ�a^��E�v���{��=.W� I#�'c��$&[�X���Jշ�M�E�H�	�������{ަ��Wn�"�v����<�9����?}���߿?� ��z�	�EPW/�V��=����oR�+�1����r�6�/���'؃���W��sc��mچ���gt�|F����G'�Tڧ�O@A��{c�}���tqr��f�����3�u����̂M��&�lqĶ[�ST�$�p��v���� 7�����j�w`}���w�뵊w y���yyy;kcv����Q�Xń�2�,�0��M�Y7�{<���6/�����N{r������\G �3��ƹ��s��x�<��FZwM+��vށ�ߟ� �#�"�l�s��{�xW�������V�tZl��<�9�H��z�{�x�ק>�yh{헳�Y�++M�U�-�W�6<?���Uʻ������� ޑ*��H�v�Hj�ڼW9IOO<?%�ߟ� '����R���v�u�4�wm����m�c����\�~���?)���M� �n�W��C��t2g��W)�XZ�HM�1��ܸaʔ3��:-��׻��j�*���EE�> ����/ $�����zy��;�x�7t�e;�e�krO���3~�p �`�D������=���ܒ}��k����|��Y�K.pl���~��lp�ܤ�{�x�� 쳄���4�V����r��=�0����/-����{ﾽ[�lOe]i���L �G�{�\�I�K�{�x�ᅿNI'=��JX_Kt��6h��m�����F�nLA���0X�X��-��}9�s8�S��@�MZ��?����{޼lp�s�_ $�x��W�8�Jb.����=\�G�?�{� ��g��$wo�cv���IP��m�ٮ��=�}�nqv��D�� z"�)"��P)Ar�{��s���� n�� �BYJ�DS�]l��8���<�#�H�=�r��g����cuhC㳗v���� �+�����{|�`d��?s�?yl�ـ�55&��.�F�\R���/#�8��=��^�kM��n��'��sp�1�V�M� ��ߞ;0	�e{��|�����#�B��Uݫ�J�m�k�~�s�W+�g���V��;���G��T��O���M���Y�N���' �\�xz�ʤ����z?ӢڗY�f&���p>�_�?o� =����u�ܞ��%TI(�L���bM �`�h����(*2#*T��(!E��Ǩ<޹畀n�J�������j��d� �s�3��I�e`Kۗ�~�9�(�z�r:�m�9W�J8��Ƃޟ[��nӠz�x�L��t��\�E_�o���`�e`K[/� 7���"<��X/"����V��&V~�+�*��ֽ��~�����g�^�/��{-����g.�n�����<?r���]���� ����' �vn�f!�L�S-9m�ͷ�{��`��M���<�w�I9'ӏ�^��/@���a����kl2e�دI~��U�߿mn���?،I$�$v�9��r�Ik�f�;j�d��murC���J�\jt�w\F.�FKL/m��E�aM9v,{;X�[��k�:�s+�s�;���S�Yx��uv�Σ��/b�O11�h`����2m�Bra�wT���!�8Z�dt]I���g�g&=y�b3������&%��q����U�a���]��V܌�!���9��+Cl��V㉉ͬ��Ɠ��%�@�ܵ4�J��i��9����ˋ�j9:oţs��za8�kD��n{�������]���97����s��?���zIvH���W{i/+���I-��m
� !��� ��î���''�N*�}��`�����w;��Ns�b������JZ֛g^������<���/s��U���}_|�^��,Ē_k��i���.�*��rrsK�}�NI���[�����Ü�߽���ݷ��f{��\�$�<�eN�Qt+wx�KvO���ނ+ߵ;�9m����\����ٛ�7���%��,���&�ב��*w@㗮�Z��C:ʶ�"8���}�$���t��5Sg.���I/K=�x�IvH��$�����P�e�������3��ѩsYmɭ�m�Ͼ�\�I�$>�c	�hċ�Z��`X����ж��	�����3�fn�o}��9�m��>�w�S3-�Y/�����ٵ�^� �o=۠���}��s�w~�~�X�Io����$����9r�G�����9��{���|��F$�]�?�I{���7=w�$��S֝Sj�T�c3��<��z���No����RK�~��$��'���%�-2U��;�2W�m�b���X�YXj�a�<<���7��\�}�'Z㮚�ҁ�šs/`[~�{�r�=ֻ��[m���ʞy�����/@�����u�WF&w}�y�K���W�s������������1$�ײn��s�l~/��!�֖:��L����Ü�߽�kdݰ?��B@,��Q�"������֍j��F8QJŊ�ȥ]���y�/~�\��7����<�xv�v#5�l,�=�W��}W�$�����$��˼Iz��]�{���`{fu��1��2ê ~�?�I/UUW��+�$����}�IMd�2�o��Jӹ!p�̶�uk,qfC��:9l=�����G�pZK�5�k�Ğ�NNmd�N����k����y� <��;�����־�I����}�S�M}��������<��s��I$����� }��=��y�^󓓛`���7�,�V\:�6g}�{������x�򨟄ֵ�3��7m���~��[m�x��J[�f�s�m���?�I/]�]�I-�!���U�s';U«�F2B����F��V1�5�&1K
�daQ0:�C^��䟿w�|�������r:�h�G^r�~�����m��~U���������w���x���]5���.���föP�vH896.(n�v�4. 8�Wi=����t��A�5��)n��݀���o]��ً�$�vG�s��W{i/+���I.�x���i]ӦS�ݳ�JlňϽU�Z��2���뜶��?~��m�{�����Y�m�=���1��R��: �{��䒗r]�^���UZ���|�^��,���xy<)m��J�ﲟI$�qT5�{��3v�~�������}vf�O�$�_=����M~��.k5��m�}�����U?���|3�h{��}�y��m���5z��e�������pyV��h�^��,͚�kL�$<R�9r�x�3'�$��y]��k,��Iǃ	Sxxߑ�a��2,f(A����S�Ԛ��J�/�������Ӡ��C���f�M�]پ(��y��b;"�D`p��1)��>�J������Fd���܌���d�NnHi$��λ��UV*KUW*�*�lC]�UԮ�uUB�5Ɲ�7����;k����(��H'�SF��V!����v������*�syt��>�k���GI��v�2t4%m͊*yz�h�ļ���H\m�6$0�R�E���b���զI�fC��٪H�m��t=sq�m֎ɉ�NW��y��8@x���y�Q��)2]���@����9y��vx��6�n�\�1��}��i��݄�8�^`-{l�8��{M�G���+� s�J)����W�ڵƍ�qG��	�O�C�ô�EF5�]5�e,:�Ŵu�oh{p��X�/SqEb3����_[�� �eW;.O
�����9�6�x�]d�4f��fv�(sx�|�s�4p7��'V���>��xl��tn� ��"�@*��=��i�--���U�;A��:����D;[���ŝ�8e�U\��Rg�sˉ�9(��=nEw	sڇ��"��ڂ�nf�nxd�K	���z(ge�r"A��P6$=qĒs���(t�t��Z�d�:�C�+-��C�U��H�m��9J�MUR��$ҍ�ܭ�APJ�궮x���@�IɐY2�Hq��ܖ�,�84�n��-��mV��V"-V�P�#)�y.�0KE�=��u�Tn���=.�ܬ��e� ڲr����������+��5u�G�tL�Y8�S�P����;?t��<sv�U�.��M:ټ8�mLb�^��8��i����h��"Y3 Bz2����j6-��38�8�v'h������Z�0�b5ɖ���]���[��yy7>n�D6u�,��:Ғb�)�\��Aj���e�-BZF;Y+��rFf���g	ob�.t��jv�ei�a�8Iݡ��]5Ua�J�*�fuK��-ԏ	Z���F�L�+����-����W) �m�'��1mn�P;�ָ�w��1���)4hDҁ�]�8a��� bу�x�_E:��>��qP؋�m�D8+�/;�H�&�F�
�:S �R\&Nk�G���˞�:!fX��P�����݃��\�����VWcV���Fà�p���������뤟u�7k �㜻��c�MևXԻ����j8�p1��:�ĝ�<��Vv2�E68
��qɳ&��s�f���ۯ*qm�hn:�ss9PW�գy����uR��5ņr*�e��#'��7����ц�Y�ь��J� K��~6.���� n3�#]�h븬hp��2���'!��uV]2SiL�| ��~�n����=��߼��rrN���������9å�P����� ���}���9�$����~�w�IO~���$��L�=U�r��/h��TJ��������P�<���g��rNE~�|u7@�|�����ZS�4Yd�\���z*�����,�ўʼ�#ϒ^��U_��+Ē]秞��ga�cͳ{��χZ� {�s����y��%�~�I%�d3�%�ē��I���2�k��N�6�؎;�*��z�6��R����w{\1�����I�7g�I)�y��IK��x�Kvd?W9U��'��{�:���d��JO�\�;:�-��Ͼ��ET� �$FT�EB/�h�"xeQCP D�H@":�@Ң`�E�o�w~���{��w�t ������l�>���kk��ĒR{<}�IMd�1/W.�o��$���ݺ ?i��<�2SiL�������� ����`m��t���}���}�_/���v���-5ν d��K����$�����Jk&Y� �����Q�NbᶨŸάe�-�
w>�[Ьn3TnB0�����ߛW٭ ѯ�˻m��W�$�ِ�䒚ɖ}ϧ�y��=����Rnu�`�Kj�$�{2}꫻^�ňĒKw�|�<7��y�9���;nPj��ٽ����ݛ��|���_�^^�w�~������z����K�晋72�2%���s�W�=������ ����9�o�Q]w�䚶��@��V弻���$��D�IJ��>���IO{#A��x�B�v&��/�aBI�eH22��c���P(�,�JW:���.��i1��I�r�;v�Se�V[����M� ;ݏܪ����?RD�^�i۴���+f��`g�H6O<�{׀}�^���i���}��ke�\3���E�^�]�~0I�+ �.KM��i^f�e�߹�9Ϥ�>�����ߟ�rO���rz��X@z�T��S���p�矽�ܓ�����sv�lT]
��H�~�Ur��s��_�] ����vK�6�IJ򓱫)�v����۲��X5Κ��wN�.LA1v�U�.�A��|c�q2ڊGͲ�{���wc�"�/��}�� ���z�t�n�v�X��窩#�������M�Vz�""��J�ҥip��������Hᇫ�{��V I<��Su`1���w�%�����}�ܜ ���=\^�{׀M����E�4ZN�!6`I��~���r������׀}��7$63Д PO|��kXa��W-�{P�9�-0�y�r9v[��+����,l���s��uO�e-��Wk��
����|W�6��.ޫ�Bp�8�ѳ��=מ�<t֭����D��6��%��A�����6l�C��D������lC��-A���{�՝@s�m�`�H7��ktH˹�f�Z���.����� t��m=��m"j:;!,*ͭB���:�]zE|ܦ�%��f�1�p��8�'��<����m
���K[�]��Zj3�I��3��,�i�:����$���r��{���=��֛�V[.շ�E$���e`�}�Ϥ�Z~�}~�w-�F[a���}�� �L�=Uʤ�'���z��T�c.��O�v�Us�^��ՀO<)��2���W9}���w�yוӧ�L�k$�u�rI����?�2"~�����7����$�+ ;*J���x��=�e^�k�غ,���S�ss�p8۴6uES2�4o
\����k\�v�޼�0�ez���+��I��Ʒ�]������ӌ�R~�BB:S�"�EDr}�|ٹ$�ﻭ�=�}�o�?���>�g�5�p�r�N�&�߿~��ݏr���*������~0�u.�XSm����X�?"�k_w��'o�߳rN{�����EVn��?� ��}�ap.%M�^�^��f̬ ��x��j"�6y6�A،��(��[�Zf��D#:Fx���f�ii��rrN�H����6�.�ۿ����I�+ ;���W>A����7��x����6S�ݳ �fV~�+�*�Wa�{��?/��x�8g��q#ޢ�y]:m�i��7X$��;.E��@$Q�dX�� �B�H�dR	"I�"��ǉ�xG�>y��\��w�wf���l*�Yetշ���s�|��w�~0�2�=ʮRSg� wOy��h]������+��9�W����vy�l��~�W�Q�H����|m	��v�U�q�-SF��F0�]o+�4l5�h31�d�������}�' =��^��r�U�ｕ�H��WCVݧJ�n������9I[=xw���'��:�}�9������1��Z�kWX7b��?)�׀lٕ���U%��e`�y�t�D+ĩ��EۼW9T��=7$�{ݛ�O~��nLG��C}�{�܆���b��t2��0	$���ǀE$��0�[���+;)_Z7m\ۧe��u�����3n�\q;��wlL��$�!�4c���+?��?� �Ix�8z�ʯ�{��VTJ'��VYE�Wl�"�^z�\H����vnI������>�~�R��Ʃ��B-7x���+ �&V�W))#��>����?��ٻ���e�3��s�����	���"�/ �l����Y-Ҡv�aj�`�p�=��+�����{+ �fV �\��s�ԃGe�f��z��Nx�0uC���i��m�H�L��y���tI������"�2ēU�6L�NB���"5r ��i���.wF����>a���v�0�1ѬMЪm�
۩���Vz+N���x�1e���p/q0.��J��e��ݤ���ή��k6$���f\����Ye��L18l[e�Ǘe3K��5Pt���p��o�����hKbe���F
��MZ���%i-��p�4K�m]~��̼Oݺ�t�ĕ��{�� �ٕ�I�+ܮr�A7����^B�J��IQt+w�vl��W9ďI�o��.�y����W����6qҴ�`��X�8a���K�}��7��Xډ�z1ф5Xl����^��|p��}��{��lܟ�+�����v�����̗VP���`vK�=\�����������~�W�(�W^I[w�e�J��(<F�Q�1T���lam�t)0b��asZ<a �	S`�S�HE�w�=�߲�	$��6k��U_ ���xV��ձ��ˡ�乣rO�����!�Yc"A�HBKH�"F	1�X�:b5�J�*�, �'�Z�$�єBW�b3F!��(�& S���VY� Fܤ$aF,���!�a�@��b�?+��S��~�7$����ܓ�>�f��'8�_�C��9��:��Ͽlܓ���nt�"�}����?~��f��[wn�am*TЛ�)%��X�e`z�U�[��ՀwO%�+Đ݈At+w�w�� �9UU^���|ｕ�E$��JڻD�t첃����
瞭݆�t��q@�Mr�&��X��G%��NI3��c|wE��t�n������L�)%����>A��e`R����ݎ�ۤ�u�vl��"�^��+ �f� �̟X�;��,%�fkF䟯����<��nh�w����*p���!�DeH�$	��$Qc@,� Zp�HCt0�'��!$"�ن@���8�B�l�4��I��HVNi�Z)��5$��(��6z�N1)R�=�FE�����sIs�ow1�"fx�B8�C{���d^x�:��ja�BO/9�n�\0q!~(��y�n`(�"'M�F�D���<=����i�"�H1���(_�`G!�6�"@��W�<_<񔔖%"T�iM����$! 6< �4�\$��� "�B$ �f�Bz�Z��%�{�A!�E_L�3H�bNsiĊ�8��0�0�G�gI�9��+�ˈK�ߘ]���T ���a�z�B07�(ačߙ��DxI6H����gg��<�'���qTO�N��)��">����'�Ǣ.<ET��8��ES�q�/D^{�}ٹ'}�vp����ؠ�M�)����%�߾��z{+ �d��"�/ �V�wn��'@��+u�I�+ �9��{��/O^��-�{+ ���,=V��T�E�\��Z%�n�yڸ�x�^�y��`c�9�Ȇ�9FN�=�ε�t9��f�4���g�}�s�^����+�U_����~���X�~��ݺ.�[J�ݺ�"엀}$��&���7veg��$n��Е�H�b]n�����&������{+ ��z��tr����g+M������Հ{��ٹ'�Ͼ��S��$"$"F@Ā�H�,�2\�ߵ�`{=�ٻn�afUY�?{�y8��{����V6L�~��ƕ<$9n�M뗵۳��ݫ�;hF�����@M�ť��:��=�|�<�8�Uߐ?/~�x�&V6L�W+�'��i<�M��0�Ћv� �0	$��&�����Ge���t؄�]
�0{���&�����K�����?_nڃlav�ӫ�m��qzO}X����;6e`G���v��7wv��bI��"�^����S��v��ߟ� ٳ+ �Ur�s��܇���v�:�W�e���B_���X���
� 靗�t����g���V1�盰��g��.�.E�,1�nE���X�n��0�tR>z������g���ꮋ<���T/B'h��n�!�R�j^7n
�۹�sא�e�cp[�aDg�;Oh��9�\mlC��˺�6�ݔm�1yXb^׋�GJ������FN��[���\K���\tb��`�=��(�ި]���T#�����2�Kn� ������V$p�'u� �Ix�Laui�+M�$p�RG�?����'ves�O���w�}n�afU��?{�����W9��W��e`�~�Q���k�WH�X�ـE$�wfV$p��){fx�	�xm%n�%t��n�	ݙX���g����� �Ix���:#�)eU�0%����?pH�������Ʒ7T��Z��r7����n�����{�~0	�p�"�_�s� ��e`���}��ڣY��p����,E< ��� �!" $X�!�0Dbx��'o}�nI���7!$p�;]��i]�ն���6�)%��2�+�U���� ��� ��+���ۜR����~�O'���~��}�� �ތ;9\�U\s%�ͨ��˥c�0V��lp�>��E�^�ٕ�obQ%�]�t�$�t��2�n. �X��	�x��7-��1��M3m�����Vn[�Aٕr�����p�̯W9ʯ�zy��"8DGz�B��ـE�^�ٕ�M��\3ܮRA6/ ������Yi��&�e`{����F O<S�ALE��?c�j��xT$��-ҷV����$p�>��E$�R�=�`���g�3M�7ir���zp���z��=��I0�ȭN�bM^c��'�\m�#�!�c���s>�!ئ��FU��5]��s��$8o{��;�fV$p�>A���yxI^
��|IB�x�̬H�N����j8�˥V��4�`G����<��^;�+ �-�UĮ�`��nـN���	ݙX���W+�O\�Q�%jD�pV+�`RK�'ve`�� 'v< �dD4.dn��� �ۀlbM5��z�'S�ƌ=6]����lrK��#��3?;�+ ݎ;�����W�5{޼T=�-ڷJ�:���7c�z�\H;��j��x�fVz��/+��av��ڴـ���:���ove`�ק �?u閨�)fMj���~s?~�x�߲�����K��xv/W�]���Э��ٕ�{��s�{}��N��u�'����=Q>"��j�(�I`(bZ�X���$���Jl	�p����v�kH�����ܸ����v�����s:2�dc[�u��Tl�,�H�V�C
1Z&9�t�h};c����n�M��n�N�tE�KQ�\e��^�GhȄf�"f�l��*�GB����mk����XV�8af�L.���������D� =\�CZ/j�Z;Hs�3I����fp�6B;X(솵�$���Ej�����s�.�S5n�֍C1�d��(�书�0z۞n�jx����Bq���<�LЪ�2�&�����;��RK�'ve`��J����ۦݳ 'v<�Ix�̯��	<�g�#��G�����#����j��x�̬v8`~��q.�y�}���-�E;�e�w�ove`�� >��ʪ��q����;���s����3�~��N }6<�d�{�+ 삨_)Z�]�pŕy�)��n3VNpz�Xe��k�_]2��M����&p��;k������ ��/ �����s��]��������ْ�4�&�^����2y)<��$�s��ʪxI�� ݎ�����GaU�Ĭ.���v� ���0��W9�RG}<�S޼v�r�v���N�V����x��y�����*�ٞ0	K|��CWN�ݺ�v� �lx�{�_�M���;5� %mIV�X[\D,�Ib��1���۵�B��p܋��ױ�����?�q�Lkɏ.����߽x�fV�� �lx�®"�v�WJ˻w�oveg�7|�`}<���{����}��7f�6³Cfp}�7$��ߵ�(֠���=�?m���X�u\v66�6��զ�r��]��~xS߯ ���������ߙ�K�2̚�x�����6{���?������-�W���]�1�a㓞_G�-]T�k���U�#���B��i�18ͷ-���mЫ���~8�8`�c�	�9ڐƕ����t�[0	�៫��o�~x���<{�Қ��]:v�l��ǀuI/��%6{+ �����E*��R��uj��:���ove`��}�[Y!I���v��>ߙ�!�aWi�I0WJ�v� ����=�W���~:���xV�xռ�H��SO�I�U�d7J����tiד8z�֒�����	�Nk��k.�U�]l+46g ��^��6^�6^�ٕ�E�ĭݷi�6��+l�>Se�]���̬���?�y姳ߙ��[T�f����z��`�p�>Se�BX��*|t;w�}��w�� �n��:�%���XҴ���uv��{0����^�� W9�ܪ��&ʢH�p��m�|kB�`\� �%	Hy��9���|���}��'�a��C̄.fRH�6I����`����5�xk-���_�)��$}M���I�7F0�����@+額ӥ<�����L�6
s�A�=;����� A��y�������Au�G��'%��w犪�U�eU�r�R��U�UUT[@U!UT�	'Un [��	�8�骶ʒ�"�a�s�FY.����D�Ө�Ea+vYx:T�th���:��G]���� �:1Wl�.�"G3�K�B`���+��"��$&�/2�j��f[�r�UuXħV��֥�
�t<P'V܎�;����{j��=�ӆ��5���l���N��и��	۳��]EOs�1È�������=�����t��d�F�F���8�
:;9�AT=�c�Dcgp=���M=m��l�(��$��s�m�1`֑���!e��]�c68	h�r	����s�����9xg:|�]�@%.9�-����Ŗ��j,�D��6l��F� �y�^6،�=��Kn�6�� 9�^��זT��e��u�gS57R��d���v:��	yq]v�(�� (^�n���qb79�cH���	��)��[=�aܗ�{v�tc'�����&�j%�����Ec�	����!d�X��^Z��P3�r.�W(�Q���K��i#�1�*Ը�w����urPr$��,���=�)�V*^j�q����-��l�2\W�u�,i�Nܠ ��-*�IK����&^Z[j(����WAFr�g��e(�Jz�"&��ɋ��:j1ڶMEhd��9zz8��:�\pΊzi�1]��[k�z���m�`j�r�;�
+u7[Hv�O�V��E��:�A����U��[q�Ⱬ��c;]�Om���EE ��]����y��w5ѧo1=Z�� �Ån=F���8tMvsp U����3	��̛����e��r�\�x�XF�i4�����@�Qڪ[SQ���Q+oz�[����Tu�;��A�Z��NKG�h�۲-t�lúrk]J��v���+
�7b�]�T�H�7lb.��ft���6������d��.�s���ef�)F$TL�ڄ�!P�ε�g�x�҅H
��T�)��('�3jF/��*�|��B��`)؊>?<��ET�+��g3����f���4e��G��AמtZ<�;P����z�zqYsM�� ,�x��<k�j�7=<��W]
����;��⢹���5��k��E��I�Q�qY��^\�!�C��h6s
�P�:,V��|�;'At�"
 �[6]��@��7���Ĝ3*lv�ב���kY��; �:E����0��.۷�,mvN�%k$���u�oF���y� �9h�S%��F�mfCYtT�囶
Q���l�g�@������-��/T:j˧@��6�T����/ �u��UU|�}s� ��
<R�#��V� ��/ �u� 콋 �n��Ur��w|W����`�������e�X��x�����Em���huam���`۱�vK�>�p�;z{�s�����)��}��=�K�7��M�Ȣi,k��tN;���t�� u��Y*��Z�o�*�{=мNw��<�M��h���_�>����=����&��U�|�吏����a�Ri�a5���'�{���CdFzk��W17 �dxRK�%M�-b-�Ll�J���6G��^�Ix{r,x��Q��tۥe�0��x�%��Ȱ	#��ڂ��T-#��v� �l����ᄓ�>�_��,K��BMS��L��F�r+��R��j�<�g�7Z]� �ۚ�9�{Uv�h��iM�:��߃ݏv=����fӑ,K��~�fӑ,K��=�sa�Dg�2%�b~����ND���/'�}��\�ͳ�\��N�!Rı;߷ٴ�?
�G"dK�����r%�bX���fӑ,K���﷮N��y�^O3��u��k�é��Kı=�{��r%�bX�����r%����)���9���6��bX�'���ͧ"X�%���wf\�EJ�V��듻�^B������rwı,O}��6��bX�'}�}�ND�,�2'�����r%�bX�~�L��ԓL�%�k[ND�,K�{�ͧ"X�%��~�fӑ,K��=�siȖ%�b^��u��Kı=ϧ]��P�_"$3Y��6A��vl����.��D:���a��ˬ[��Q��D�,K���ͧ"X�%��{��ӑ,K��;�siȖ%�b{�wٴ�Kı>s�-�a�Mk4\���ND�,K���ͧ!��DȖ's�fӑ,K�����6��bX�'��}�ND�,K��쥹3;�Kl.Y���r%�bX�g{��r%�bX����m9��2&D����6��bX�'���ٴ�Kı/����֍�)�2�iȖ%��D����6��bX�'~���Kı=�{��r%�`~���ͥ���I'?T�[%��������?t?5������'w����/'�?x}��u��SiȖ%�b}߷ٴ�Kı=�{��r%�bX�g{��r%�bX����z��������移��
�Mj�]��V]x{=�\u��r��$v��z�lzȩ;��s�X��uS�O��O%<��{�����Kı>�����Kı=����r%�`~&D����6��bX�'�Ϻ.7����]��'w����/'���6��� �L�b}����ND�,K��o��r%�bX���m9ı,O}�{�fHg	4�a.��ND�,K�{�ͧ"X�%��{�ͧ"X�%��{��ӑ,K��;��ӑ,K9��<�Y�zQ�52-듻�^B���;��?M�"X�%��}��m9ı,O���m9İK�{�ͧ"X�%��������k4\���ND�,K���ͧ"X�%��=��߳i�Kı>���M�"X�%��{�ͧ"X�%��M�
���w�s)�Vi��hL˸�a��4�]�v���8��x��rH� ���Ѳ�f�H,i�������O\��-.Ƥ�{g�[�pi�p�@m�Վx�f�P�M�fvh�O"�ͫn7
q�����XV�n��8#7p�x��0�nM��&�=Ī�J6$y��fh&�h�'�"�z�"����!^%�������td����c.�����rBN~�9z	�݉Z:�PsZ���y�I\9;O�Y.�^�
tM��Wh��-�]��'��^B%��~�6��bX�'��}�ND�,K��}�^D�,K���ͧ"X�%�}����j�ɓ2K�m9ı,O}��6��bX�'���6��bX�'��{�ND�,K����r'�c��^B�}��������r޹;��K�����M�"X�%��{��ӑ,h�lN���n	"��vmI�>����&2ffe�&��b{�����Kı;���ND�,K�{�ͧ"X�%���}�ND�,K�ff�Z�[�L�ֳ5�ND�,K��y��Kı=����r%�bX��wٴ�Kı=�{��r%�bX���ܺ���x]+�93�ỳ���	��{;�FR�`�N{VkK��WZiQ�x
����/%�b{�wٴ�Kı;�wٴ�Kı/����~@�DȖ%����si���������:�K3���o\��%�bw��i�hA�+�� �br%���{�ND�,K���ͧ"X�%���fӑ?
��S"X�s�~r�9��L���r%�bX�g߿fӑ,K��w�ͧ"X�$2&D���iȖ%�b{��iȖ%�by�����u%�B�s5��"X�~VD���m9ı,O����iȖ%�b{�wٴ�Kı=�]��r!y�^C����]1���rwy,K����iȖ'���>����ND�,K����r%�bX����m��B����N}��4��k�[Wx=?������;n^¼X�5���^�����%ub.���S����O%<��}�?�?��Kı=�]��r%�bX�g��m9ı,O}��6��bX�'~��R�u�rF�M�����/!y����i�F9"X�����ND�,K�o��~'�2%�b}���M�"X�r�����*�1��56N�;���"X�g��m9ı,O}��6��c�������Hd	�`\��b����O"k��m9ı,N��߮ӑ,K����d�	��M6�K�fӑ,K����iȖ%�b{��iȖ%�b{�۴�K��L��w�ۮN�!y�^O<��u��f5#S#���Kı=�wٴ�Kı=�]��r%�bX�g��m9ı,O}���rwy�^B����ؖ�Z;	UN���K:�^,7�P�,�\�m�z�NU�Ӎ3D�f�BY�ٙ���Kı=�]��r%�bX�g��m9ı,O}��6��bX�'���6��bX�'��a)�w5��Y�.j�9ı,O���6��bX�'��}�ND�,K��}�ND�,K�u�ݧ"X�%�~���\��ccU��Jy)䧓�{�ͧ"X�%��{�ͧ"X�%���nӑ,K��>����Kı;��{�[�&Z˖����/!y��{�ͧ"X�%���nӑ,K��}��ӑ,K�j2(| �*���o�rm9ı,N���Y��]d5�Y3%֦ӑ,K���w�iȖ%�a�R?���ͧ�,KĿ}�����bX�'}��6��bX�'��{c�^:���5�uؤ�A��M��y�=�F�b�&�V��[�LL�Ҝn�k��Kı;�}��r%�bX��{�m9ı,N���m9ı,O}�{v��bX�'�gݒfe��M6�K�ͧ"X�%���nӑ,K���fӑ,K���w�iȖ%�bw>���O��O%<��{��'/���Dn\ݧ"X�%��{�ͧ"X�%���nӑ,K��}�siȖ%�b{�۴�Kı>s�-&t�!u�)s56��bY�D����v��bX�'��fӑ,K���w�iȖ%��r�'�y�m9ı,O�����~�h�l�˗5v��bX�'sﻛND�,K�u�ݧ"X�%��{�ͧ"X�%���nӑ,K�� =dRE�D� �)�@'��?l��s[
`0ۑ�ɉlD�y8S��,�1���F�j� ��u��Sl�k��m��bѥMq)���9t\E�K�"B���B�"�#	��W&���y6qs�����F0p�܀9�b�@ܳ����T�$�Y�m��<[:�j���x�G���G���%��dѠ���;n*�C���b9��N9Վ�Y��a�0���d���\��QT�oy��"k�Q����Lg\γ�'Uq�rOa�n�2����i�ve�,#�泉�Kı>�]��r%�bX�����r%�bX�����9ı,N���m9ı,K�߻3YtY�˩54MkWiȖ%�bw��iȖ%�b{�۴�Kı;�w���Kı=�]��r%�bX��E�̝�f��ɬ���SiȖ%�b{�۴�Kı;�w���Kı=�]��r%�bX������#��R9[��lv�M_�\�]�#�"X����fӑ,K���~�v��bX�'~��6��bX�'�뽻ND�,K���32K�)��k6��bX�'�뽻ND�,K�w}�ND�,K�u�ݧ"X�%����ͧ"X�%���gK�f��̄��}��&y�:��z^`Χn�l�]@3�/K$-&,�h⭚�*�rwy�^'~��6��bX�'�뽻ND�,K��{�ND�,K�u�ݧ"X�%���vt��jI.�E.f�ӑ,K���w�i�z	 I@�����H꣣��'�s�q=�b{�o��r%�bX�}���9ı,N��xm9ı,O3��)2wZ����˚�ND�,K��{�ND�,K�u�ݧ"X�%�߾��"X�%���o\��B�����<���*S\\.�r%�bX����m9ı,N��xm9ı,O}�{v��bX�'s��9��<��S�O%���Ք1��,�r%�bX�����r%�bX~Q��o���%�bX���߳iȖ%�b{�wٴ�Kı?�߿K�I��<��٠���y�>Zpl�v�����w\
��OW�3ӲI��:Esw���=��h�'�k���Kı;����r%�bX����l?�&D�,O�w��"[�^B�y�}�1���F���'w��bX��~�m9lK����nӑ,K��w����"dK��?w�m9ı,O����$�-䆌��f��ND�,K�u�ݧ"X�%��~��"X�|ס�B�I;GY$��@�3	�P�HdP���HIX���@��[HRRD T��%#XK|!a���%�IH^��!BU�D�c���U�1JU����嗄b�CY��	BV2��
��2I݆`�I(J�Э`K<�(p���{3�ݶf$ٛ[�'����d�J�{�P�B�䌁2BH�X���X�c<|���1�X\���2�	�!$yJCN�(d�!$̈@�&�J,V�X��U��
K�%s
%����ƹxg6����5�0#
,���"A�Z0.��,�!+-��V��ԕ�d({Mj�H�����	ea�!m���i3CBR����$�K��%�M��t6��	d1ڈ �@�Oq�*�i_�=�|��U#� O�y3߾ͧ"X�%��}�siȖ%�b}��ܝ�][�i����ND�,A�;����Kı=����r%�bX�����r%�bX�{���9ı,O={��5��BY��kFӑ,K��;�siȖ%�bw;�siȖ%�b}����r%�bX�����r%�bX��O}�
9%9�4�Df�m,5e��!��49|W���u����x8c�2Z���g��bX�'s�w6��bX�'�}�ͧ"X�%����ͧ"X�%��w�����/!y�y�ꚸ�-�L\�t��bX�'���ͧ!�c�2%���w�m9ı,Os�fӑ,K��w�w\��B��������Vku]���r%�bX�����r%�bX�g~�m9ı,N�~�m9ı,O���o\��B�����g�7�<��vƵ6��bX�'�߻�ND�,K�߻�ND�,K�~�fӑ,K"�D@$UdD$���A,ZD=�� @��DG|���~]�"X�%��gw��L�������k6��bX�'s�w6��bX�'�}�ͧ"X�%�{߻��"X�%��w��ӑ,K���z\��Me�j�Hf#��7(a�f�k���*���v��1E<oJ�.;Y�L��M�3Y��Kı>���m9ı,N�_v�9ı,O3��m9ı,N�~�m9ı,O�[ѯ�ɗ�p�듻�^B���_=6��bX�'���6��bX�'s�w6��bX�'�}�ͧ"~T2�D�?y��d]ej�'\��B�������ٴ�Kı;�����Kı=�_v�9ı,N�_v��Gșĳ���5+�6��듻�^B�?g�߳iȖ%�b{���r%�bX��۴�K��Ȟ��߳iȖ!y�{�iG&��5��rwy�ı=�_v�9ı,?G����v�D�,K�����r%�bX������Kı8k�d���2nV0�H��4���L
��I61�o<�$~�͡,)��p:R�d�L�Yyk8���+���H$
��3�<U���ւ/HNq[ac�61ìA+K��ґ�[��n�8H��h8�w]/z�E�ik�]� A.lk�������Qnt2�I����� :!��6|s�{jC=nR�k+����-��]p����!kD���+[��۝nzs7n�X+��6mj�@ m�gV���$�9�	��wn�3�h��49���&�=a���*qۘ���kO���𚂮xfY����_��%�b}����r%�bX�g��m9ı,N�{��~U�L�bX�}���ND�,K�t~�s�e3N��������r%�bX�g��m9ı,N�{��r%�bX����v��bX�'{���9ı,N�;��.���j��Ku��r%�bX������Kı=�_v�9��ș0 ~��߮�Ȗ%�b{�~��ND�,C"|����2yL��)���m9ĳ���>�}�v��bX�'�߷�m9ı,O3��6��bX�'s��m9ı,g���z����r�rwy�^B�w��fӑ,K��=�siȖ%�bw;��ӑ,K��߷ٴ�Kı;�'h}Lj�53m!��3v#c����y�6�n�\k/�OGmx�	�ݔ��\��r%�bX�g��m9ı,N�{��r%�bX����6�y"X�'�����9ı,Os��Rau4]�Y���iȖ%�bw;��Ӑ�Ĉ�$��	��P �@�dVY Q�B���pc34�	�]*m��B�FT*�#�B$�Uٝ�*���y���ɴ�Kı;߷ٴ�Kı<�{��r%�bX���լ�\�듻�^B�����\��bX�'{��m9ı,O3߻�ND�,K���6��bX�'�w�K�E�N�;���/ܜ�'$�M����6��bX�'��fӑ,K��w�ͧ"X�%����iȖ%�o'�3�{�i�.λao\��B����{�siȖ%�bw;��ӑ,K��߷ٴ�Kı;��iȖ%�o'�������R9	v�HM\��t�&��K\{p�ݝ�̸���s�5��D��Y��Kı;��siȖ%�by����r%�bX�w���r%�bX�g�w6��bX�'���'5��M��]k6��bX�'���ͧ"X�%���}�ND�,K����ӑ,K��w�ͧ"X�%���ɻou����MMkZ�ND�,K���6��bX�'��{�ND���I$bH������n'{���9ı,O~��6����/!y?~�_b�n��#�z���,K���ͧ"X�%��뽻ND�,K�~�fӑ,K��{�ͧ#�^B�o|�]�JGmL�;�bX�'{���9ı,?+��?M��,K�����M�"X�%��{��ӑ,K��5�;��R蚺������9SQm��8���)�d2��-�o\p�U�ҕT���������z�6��bX�'{��m9ı,O3��6��bX�'{���9ı,Op�ڬb��Qo\��B������]�ND�,K���ͧ"X�%��뽻ND�,K�~�fӑ,K���=��3L�vu�z��������߽�m9ı,N�]��r%�bX����6��bX�'{��m9ı,N�;�jd�s�s-�rwy�[�Id*w��nӑ,K��߷ٴ�Kı;��iȖ%���!D��E�D����K���m9ı,N�}�r�fM6م���r%�bX���y��Kı;��iȖ%�by�����Kı;�w�iȖ%�b^���b}%�e6��JX��F7�9����k��*4BM]�R�l.@�դ�̡�����%�b~���ӑ,K��=�siȖ%�bw��n¤�L�bX���y�wy�^B�~��:�̹4"�ٽrr%�bX�g��m9ı,N�{��r%�bX���y��Kı;��iȐ_قH�����0��-�4��H'����ؒ	"y�i7�?D�{�ͧ"X�%��{��ӑ,KĿ}�r�-bEBR�w\��B�����y�}'"X�%��������Ȗ%�b{�~��ND�,���6��bX�'�w��X̙�S=rwy�^B�{�{v��bX�'�뽻ND�,K���6��bX�'���l��șı4rNH���nc��y�'�Tڂc&ظ�Gn5�����\��"���,0�b������8�$��(�����i�L�=��$�8�18z�z-Wu��ڬ��9�a�An����m�t��t����v�u�`�l�l��ʆF+)�!�M6mid�6���RĤxRP7�X�Ǎv������:��>��o��G���X�c��ӸZ�=�"���NIܫN��舺�h�+�9s��{���^|۷Py��`��d���+��tR��z�5�3.�=O�X�%����۴�Kı;��siȖ%�b{����r%�bX��wٴ�Kı:{����j�u���$���r%�bX������Kı=���m9ı,N����r%�bX�{���9�TȖ'��߉˭H\4�f�Y��Kı>���6��bX�'{��m9ı,O=�{v��bX�'s��m9ı,O;;f��K�sE�SZ֦ӑ,K?@ȝ����ӑ,K���~�v��bX�'���6��bX�'���ͧ"X�%����L�亲Mk4]L�M�"X�%��{��ӑ,K��;��ӑ,K��߷ٴ�Kı=����r%�bX��$սzbۚ)�ł*�Ԅ�	��ю�b�\��l�9�7ZKtJLu���ʃO�Ȗ%�b{�w���Kı>����r%�bX����m9ı,Os��Z듻�^B����=�*�$��J��ND�,K���!���U�O"r%���}�ND�,K����[ND�,K���ͧ"X�%����WZ5�S5�ˬ��SiȖ%�bw��iȖ%�by����ӑ,,2&D����6��bX�'{��ӑ,K���;:��5î�-듻�^B��K&�������ӑ,K�����6��bX�'�w}�ND�,$N���m9ı,��~�s��1��Z
�rwy�^K��{�ND�,K﻾ͧ"X�%�߻�ͧ"X�%��{��[ND�,ay>�9�?>}�D�nM�-��\&�Y�+�7=���P�v,m�6�0K�>�nm�	u��yı,N���M�"X�%�߻�ͧ"X�%���u�ND�,K��{�ND�,K��ɻnw-չ���ֵ6��bX�'~��6��b~2�D��~���r%�bX����fӑ,K���w�iȖ%�bx���3�,�&k4au��ND�,K�u��6��bX�'s��6��c������ �X7�� 3h%>}��br'�k�.ӑ,K�����6��o!y���{�ԍ�:Z��vq�'w��g�FD�~��ND�,K�����9ı,O���6��bX�'����N�!y�^C�|��0V��Zͧ"X�%��u�ݧ"X�%������m<�bX�'~��e�r%�bX��{��r%�bX�����2f]MB���ŢJ�ư�K2 �b�F��b��X�5��dhYX��V�vq\�rwy�^KϾ��"X�%������ND�,K����Ǒ,K����nӑ,K^O|g��efѮuι;���*X��~��Ӑ�H%r&D�;���6��bX�'ߵ���r%�bX�{��듻��&95�/'��ߕQnkeM����"X�%������r%�bX��]��r%�bX�{�xm9ı,K��v�iȖ%�b|}>�9�4�j�ir��M�"X�%��}��ӑ,K����iȖ%�b_}��[ND�,� 2 l�V�D���ɴ�K^B�y?{o@L_b-n�u���/����iȖ%�b{���M�"X�%����nӑ,K����iȖy)䧓�����t1��e�[��1�N9�%r�ܘC�i�P����J�]´t��g�e�$�kS2f�m9ı,O}��ɴ�Kı>�]��r%�bX����m9ı,O{�xm9ı,O3���Cji�fkY�d�r%�bX�{���9ı,O{��m9ı,O}�xm9ı,O���ɴ�Kı/���Y�e�S�W'\��B�������o\9ı,O}�xm9��ș�w�2m9ı,O����iȖ%�b{�����%1U�g\��B�����xm9ı,O���ɴ�Kı<�]��r%�`~fD���~�ND�,ay>�3�~��uks�ι;���*X�{�y�iȖ%�by���r%�bX��]��r%�bX�{�xm9ı,Mo���L;J��\�m�
V�X�R�1�L�ͺ!̑�`a����2�/=�CM BնRFC�"A��	���m�H�s��_��8�p�0,�Z��WZ�9>m�����9�6M�@����A�<�y�85��e	%<�֠Ü
h�"H������A���Z-��CU��i��L�8g�!	1�)����&��!	!�N }��y�d<xh�HHE Ï��kӑ}�SK"}���=C��%�q7�*04���A�e�HW�D�}ѐ>����a$7�$w��&�N!5�TK�h8F8oȚB�W �����|�����@Uv�b�v�MSΖ��UUAPVڥ�\����Z�g�.[��D8x3o��Bn�Wn.�X�#�K��^��I;� e[XP�.a���y,^�f�S�4�${	�c�X:.�nqFr�5�D3Q��9J�asgI��b��k;�h:�fwO�� ���i���u�k��H��QF�^��p����v�]�%�.�J׹��'P�ۣ���#�E)2B[͸XB�P�)��W� �|�N�<Q�#��������t����A���^Z��n[)��$5n������6�H8�'1ɮ��$�jI�7gtvSC�i�rW�-��"��I�`)��۝��pek��2��;��ny���� �!�k�͝���5= s"�v�!֖J[ώ8ȏ=�m�,8��F�+�3p�燧u�ݷ�Qxֹv\�A����'n�n�c�)��n�WSF#E�cN��t89!:�Q�;�8��y{�j���<6y�@L��7=��^�f��8d��h�`5�zZ�l�v�/���d�ͱ�9� ة��\�e�-�yV��Z).�0���]��`y&��&�ݪ��\6�5�k�����4"ڰ�G*�*+Tnl l/7I�Ҡ/���Ò�%�Q�puu*�YZB�s�KR6�v[gf�cJQ�mf*��.��
)pJY���8�v15$ �+,v�=V+r��'�jD�b��ܗ�HF�+�^�+��"�ZGH,v Y:io3��Yt1��1�\n04��Gh� ;%����wo1��C�0�U��V7�ѳl
M��4l��.��Yd�I�c���EüķS�t h�t��n:vy��rT�����o>�ɷ&�%�m</ B���i�h�y
�wM�c����ӄ�+ kn�����/NM0�Q�kQ)�q��8f�yϔr5V�6��*X1n�v�K�+����q9C]0JJ�c`v` ���Yz�v����Gz��i�e�91�'l�lڣ+�gc�rNs�9$g'$�1TÇ��g��qEo�p�W�T=H0��)�� �<>QP�K��h �����aFU���;6Y�
6&3Y�9k�oI6���uǝ�/k�FS6������<���t�Aۣn��K����	ݦ��lQոΗ��@Q�����'Y'�[c�9�>�A��!�t���C��)5�И!8v<�u�����2�n���@�<��n�L�����;�ã0����Cci	v�k9�\��\�^Yǲ��w�����}k�ё8����=c'�>�Ϧ��XƸ�.W�셲,!K�cr�ܣ3j��'ǒı,N���v��bX�'��{v��bX�'���6�y"X�'~��d�r%�bX�;;����ղ��n�v��bX�'��{v��bX�'���6��bX�'���d�r%�bX�{��v��bX�'O{$ݙ-욙��5���r%�bX�����Kı>���&ӑ,(�"dO����iȖ%�b}�_�]�"X�%����L��35��]kFӑ,K��߻̛ND�,K�k��ND�,K�뽻ND�,K�w�6��bX�'��m횎�ZI35�ֲm9ı,N����9ı,? ~��߮�Ȗ%�b~���6��bX�'���d�r%�bX��s�㿡��<��4�����=���2����e�<i�
uqx�)���Wsk�E�Uoǻ�%�bX�~���iȖ%�bw���ӑ,K��߻̛șı?w_�:��������O=��p�9���Kı=����r ���&>���^D�K���ɴ�Kı;����r%�bX�����r%�bY���;�q�����/!y�{�y�iȖ%�b{����r%�bX�����r%�bX�}��m9ı����[��X�FP^�;���*X����v��bX�'���6��bX�'�w}�ND�,K�~�2m9ı,N�N���j�5�Z\��iȖ%�b{��iȖ%�a��������ؖ%�bw��̛ND�,K���ͧw����/'��=���H�J��f��:{=��Wp��=h��,.�1�&��[Grl�.ff��55�jm9ı,O=��6��bX�'���d�r%�bX��w6�y"X�'߿o��r%�bX��}=�>նܭ�sz������������r%�bX��w6��bX�'��}�ND�,K�{�ͧ"X�%���z{j��^[v��:��������=����Kı<���m9ƞh��4���	� g�$w�9��iȖ%�bx{�xm9ı,O����ݮ�(��N�!y�9 "{����r%�bX����ӑ,K������r%�bX��w6�����JO�}������:�mS�����>�ٕ�un��>�p�'kJD@�=�g��]�����U�����L(��s�����S�z���=�ܴ|�fVջ/ �u��>A��� �5j�I�I�Ք�u�un��s����ؤ~0�?ջ2��IA�Mڦ�J��ۼ���0�ve`�e� �j����;m`H�p�߶nI��߳rhE� @\U5�oq`�*R.[\)��e�0����"ݗ�}�"�'c� }R��B����x�J��%�9["<��h�u�8fs��yP�*�KuAo���m��p�}��mȰ	��v�fVy#�%=bT�t'iYm�w�v_��	��v�fV��SjX��鎓JҶ�v8`�ٕ��='��=��}�S�-�%c�Nĭ6`V���	6<�ٕ���L�z���ět�Ue$�`���Wd����~0�n��7�F��.��r��q*�2>g^�u�Busۍڡx�!�m�@p�G.n}�x�,5�nm��	y���퍷DmSI@��r�:J,������--�2��`�:ņ��夫�����w��n$W4����c��#	�6�m�=��y��a�ȼ,�o��}o����Y��7(��Nck¢]�9�᪭�Ge�3se�mV̀��Iy'=�9�:�z�d�$s���:��2�=塛	��vJ�K�E���(Q��<���m�ڧ���+ �\0�n��"�/ �Q$˖퍖�Sl�$��[%�� ��~�*�I��)m�6�nճ �)�^ N���Us�.�7\0DR����L�wCn�nǞ��$n�� ����>��/ �%���`�v7v� �u� ��Ի���e��W*�T�As��j���*��&�ܜu�4�{t+QYu����x�85����L<�h���˭�s��ߟ��/�{�7c�*�������=.�~)Sn�c�Z�n]jnI���ٸ>qh�		"T�B$�H�+Z�R0�*	X��HJ9ʣ���Q�W*�0�>xv8`�� ��CMSN��*e]ۼ ���w\0�U�ܻ�??��{�x֒PlJ�bT�J��;�� ��˲/ ;�xC�Y�l���T�k�����������X]+h���]��6K.D��`��ë�s�z���m�9�-˹�M=n/;�j�㪆>�F�I��X�� �$��|7u`���x$�=ĉ����y��>[#xZ�ʴSe�]+�[����X����W?R��Q\9\��1C?+�T/��_7�x��������uc�iZN���\��{<`S��H��p�7n�iһ�v$[fˏ $���2��p�'a)��Wm$��9v�q�s'�0P817#������/2'�yy���g/����~�2��p�"�q��%�ĩ���ĭ��&VJ�W*�Wf��0<����{�=�γ�m��K+8��-� wv<�0�I�wl�;f�U\�/\�����<��}7' ��"����M�<��8��v7m�wc�;�� �c�ˏ ����u-��4&���?Uo�]��b��r�Y:܅�&EL�8���Uq�NNp�u���b�e�����תlp�"�q�+���y�V�͡�Ɔ��ݺ�7�� �eǀ� ��{����KO}��sY�+�.S�yO_� odxvL��\0	*�M���&�^��o}��{߾��;5��9K�=~x��z��bT�IQb��ݓ+ԗ}��z��{׀I:z�Z�5mm�`�Z��OH�'Wcv�v$@�t�lz㷎�44���T4{q�4``ؘ;TvJ��84���C��Kv����z�LD�m�/��&�Qc=�A��7�V����z!;nCDQ�W94Ã
\��bt,Y�s���F�r�ʔ��Y�i�^HLlU"����XLF�����c��^T��[t�nG-QAؚVm3Rs�����rC������V���\)����@���gk[�W��n�#j�t��m��b�m+�@�m�@�k�E�������$�?��{��N�����h|�e��Gd�"�q�����X�\3�9�RGTJU%�E��Wcv��^ݎ{������������F���M�J�hm[��0�p�"��5vK�5V�V�1�h����0�p�=ʪ��y���}��>��}���>�ԕ �� y��U����L��u�D��Ťu�#c��`�.c�H�=a�`l���%�lp�;5� �u��d�V X�*�o��sI���@@�0# I!C�Pء�:N��O�����)#xt������m%E�v� �d��&����������Ӯ�K�
��O'*��g��{��we�l�X�Y9-��Sm��[0�F�����L�w\0s��iz����[��z�6�
���ۘ�J��ԥ�lFљ�'��&�In�v��-p��ԻW��{��?�l��'u� ��7�DE��)�b�|�[M�����&�v7��<Un��X���V�v+u�M�	��ߵ�͜�|V��̘�@�!		�hL�[����r����!���]BB��R���vC2�A�!*K%�����m!��i�5���4�cBHI=����>ޤ��Y���˂a�LM�	�p�l0�f�͘H͏�ľ{�4J\k�� ���EܮnT�II502�BHJR�Q[���D(2v��y� �T8�_U�يq� �#�G�U����:|*���<P��~��V��D<�}�}��9�l�KO�:���#v��5�N��~^��/ ��e`u� ���Jղ���"�m���<�+ ��["���{t��P� l1#���nt��؞�����!��BX͆�,3clP3m[i*,Wm�M�X�`M����y��LU��-�J�4�`�ឪH���� {g���+ �lb��C
m�ݫf�� ���M�X�p�q#V�*����Ӵ+�����'� ��v8`r�]�J��S则7�}�nI��_~5`ݱR�Z�w�}�2�	��E������=��f�cj��؋tķ���� ��ݸ$�nF�Yʒ4ee�t�^0�4�d��Y�t4դ]ڷ_���E��"�/ ��2���Jq[����զ�.�o?s��s�IS޼��e`c�{���->�u���í4M�x׿}xݓ+ �0�cx�d�ZM�V�J�Iۼ�ɕ�I0�cxSe�MLT��Ī�ջu�I����z�� {�� �l��)r�}l��Ԁ纛�[�j��֡M	V�0ɎT.a�R�t�Z�uq9��NwzU��eƭn�@*.k���;
p����<86˦����=���r�<Ӷ��.+��Aj�>^z�+�>I�;F�	��s���k�+J�J���P�Gn!-�v p�dY�Ǭχ��#�O
� X��gһ�i�s�(����]�9}j�m@�)��P{fF�&��m��(؋����XkR�K��5�d�WN��W$pg�5nO]��"p�9�uu�Tι=��ߗ��x�\0	5� ��[�(�:-݊�m��lx�\0	5� �lo ��ڻ*;bE�]�ݷ�}5� �\0���vG�j�K��5MU���f�r�zL�yzy� ���Mp��r����K�V�c�h�i� ���x;#�>��M�)"�7L���`(�]��H( ^����up��<�d6X��zc9�n�G�j� ���Mp�&뇹�s�������$�g���b�m%E���T8*�s��U>s��᙮�lo &�x�T�)�hL��v� ��Scx7c�>�2��e9i�+ubv��m��� I��M�X��uu-�B�LV+������̬dp�"��|���⋥t�m!`�K-�j(�S%��l��[��z��!�3LF��b.Ku<�\��~��r��� �lo �$�V�KmX1�j�U�v� �3ԑ��y�)=x�8g�����n�V;���m�$��{�nI��߳s籌���
&�Xߌ}��6���l��nЩ�m���r�T��� ��`H�E$^�l�cWCd�T����zp�G)#x��xkvR���n�X8qr��E����#p�v��Q�z|\-n��)v&�[c�����?�צ�� ����p�;��ګ�V'n���0��窒	�� ����$ujR�%�Պ�m���� �I��l�)#x��˲����9v[�oܮ.����	��`_��Zܚ�� �`��G�r��krZE-�alJ�ګJ���\0���fǀvI��I�R	Avs(���`]`{m�^!�թ��A��y�N��b���0.�|3slq��������c�;$��$�mG�lt:m!U�n��	6<M�X��|���	�����.ؕ+m��2�	�ᇪ���_� zO<n�0�5t:vP�m��N�����	��Jk�X�ѣ��]�Z�c�`]��\����g� ���+��$O$���@�C�5F�����+:�K���C+=Z{s�P-�M(M�1{w.���/ˌ�KV8F�z�������V�x��	�/3�l�hzB)��U�vӔd�`v� ��d6;k�x��>M��F0C������"ƨ�ƭ�x#�%6������h�����8�N-�#Rtݎ�*���i�9���,c��Sp�:�T<f8�7\]��%�NNN��é���Rn���7�� nq�@�V�Ѫ�2��PE�<�з^�'T���-��ݷ���� ��/ ���U��W���F��_=wC���m��E$��r�#����z��I��R�LI�wVݶ�	#� wb� $�����H��m*vZ-� ;�G�lx�#�|RnC �Tp�V�:M�;V�x&ǀ�&�`�.<�[�2]�w��#m��OYź�b��f
R�i�n�R[Slo
��s�$�6�3��c�$�.�ǀ�<n��T�1؟j�w�M����\�9_Us�XZ͸��#�;�س�T�9��&�6U��[� ��~x;#�;�ذ	��j5m.�pmX��� ��x{r,������#}V������Z-+o ��"�>��jݸ�wc�=UU��W��U��P�����˥�	���/nѦ.(�rY�ל��,M�f��Ɇ�	����V���������uH�c�ZumU�Z-ـ|���]�����ݭ�˻e�ۺ��&�V��f��G�D�P���M��g;�����d�Wv�N�j��ۼ)%�H�|����*��=x�@i/Sj�.��i�X�8`�W+����)=x�r,-*R-$�AceM�Bl�b+��f�[���br��$q��W4.ֳTڬ�����w^�v^;r,�0DS���ڱ]��Wv^;r,�˾��y%����'�h8<�5���?�\0��x����$��J�'v��M�R&�`M���{�nN��OE?~�3;��'��h����-���E��0��x���\0������ӳ$���Q�in�z0����r�=���H���c����=�VD.��am�]�v���/ �������>�w|���K�le��\3��~0-������	[�)M�ڻ�M&ـ}5� ����5we��p�7��M�iڱ��;feǀj���;��}5� �5mQr�pmX���Wv^���]��|�YTQ�E{���jɽ�>OO��$�/��������Y�����$p9�jl�Y�ȑ�H��
T�!���%�9�9,�C�Zy��o��n�~s8�R5%|#LׇT�+�y�o������$My��� ��q��%�h�h����`�VQ��/��3�	�zfh�sS5�+
8:����׾W��eMs4���P"�����]x�y���!xq���7����C�cO��=ܼ`h`FV��!		�u A�t��!���4�ˣCki���&	�)<����і]��Hi�ϔ����l��P7O˓ �S-y�קƴ��=5�Yx�8hxʔ�0�B$b�8�}���@�1$2*xӥ&�%�<�f�d%�}�y�=�P�����>��6nց�R��tw�`Be���y��n��n����!�B$a	yp� F!h�^��{a^C ��o��H�I��(fs]֪��C*�UʌUV�TqUR��V���G8�.����q��o#FTQ��`�h����]&�I��qB򬹢�ڧ�j�yz9z
v��^�b�6k(&�n�I�c9��N��f�#(F���c�v�)2m��� �n�f9%�OR�ݦ��)�mS����tK��Ϟ��]y7nC��<�$�qr�;�ۏ]���n�ݴ@��rg�s�2�,�KT34���fi��8��1��CxЄ���	'CMqq�ɹ�3vbsgt�0�:�XW�^���������x��V�"Zm�8��Ɏ3��7y�dV�s�X�z5т��a���t��^{P/W�	���k4�S��j\�/n8�62�'�����R��=�9��ȼ��:�&�TI����д�ʳg�yy��KxP�R4�������B��]6#�[8��OC��r�=7�\R郆4�h\�N�i�� x�Maw'+"dݮ���&9��B�:6%�d�-ΰ3Z��Zsǭ����j���>��q�7G#՞E���$'Q6��v
H#�مI�tk���f�w��{���e�jA��;�X��Y��0ª0�3�s��H�8-)���J�%���_Q�<`�k�:z۪*-,�ö���*��j���vueI���<�p
+� rհU=e�(�B!As ɺ���0Z
ǭU;D�ʲu��}�!�	�O�P��WvՐ
��lp ��F�#�[��ͅ�1�<9L�7;td�R tT�]��t����(�p-�!-Ds,��3�c��V��:T%㱂�tf���8��{v<��9<�[o�x���J[�`]���ܘ}W4+s�n�v���䀋ۖB�Q��&p
���X6�]�uE���6���u����gi�$����� j���+1�9�:Z�ؕ��X�ʣUO<Z�,J�Ź�Ss/i*�\p���	mi���4��@6�YV��m����B�q���Bۭ���ݱj\�r]f�f���'=OC�ب�"!��>AA����|*��L"�c��v��|���u�u�a������r0<��..��9���;�x�;9I۶���爻�^)�Ɨ<����s���X6�q��9駂	zmc�h�)�u�d���N�0����n�
�t�9�LU�v�4�p���+8��d�h!1ŀ��g93qc��<LK�n{s��mzxrI9N�V�Ў��]u����Uc�t.���	����$擓��/aCw06���4�3:��آ���x%g^س�d��
yX�Q,(�lGDq������~���Ȱ�.<w\0]�]�[I0N�X��k �\� ����7��wob��G��Kʋh���-���<���n�Ke�,��y`V�y���-��s��{�N���o �G.ˏ ��RPV館tݳ ��ŀ}#�eǀn���pמ��0�`����Gy'�t2�\��p3�)-�n���X�8`M���p�;/b�;�ڊ&�-���[� �mǓ�;B\�O�J�B1:�b�OE�OȦ�*y����ܓ�s��'>�_M�AFKOi����n.�r���� 콋 �G)��WvT��줁]���qo���;�?Sn<W�y`^��Ym$Щ�ĭ�X�8`E����`/b�5l�J�����K��Vᕪt��ɻv��^��1#�)sp:�n�oXpрEǀn�ŀl����W�;�?�N��L�-�D�� ��^��y<���\��;�?D����RF��ޠՉ�iP�f�\��>�����>�H$,Q`���W�5|_~x������V��m4ժi�m��0�����%��z��.�F�К��bm`,�x��x�ذ�p�;(R
�B`��e̐7��nz�k�&���'CX1@"�#���"K��&+[�gb�
�����^�y|�� �B<��*��]ݫT�]ۼ�{�\0��Se���V��;Bi+�m`5� >�� �6^ݽ� ��-TU�1����q/o���� �ݗ�^��*����ҫ�!�D� ��E矼��ܓ�O�\٩�K.����i�T�x��f�`{z��~��Aeeܳ2�A�n��M܈�\۞ě�%724�-f6RYL�ca(�Qt[w�j���6k� w�G�j�/ %mij�-;+��m��6k�~�r��n�y�zz�]�xx�wBj�n��l���Se����	5� �M��Q5���WM��)��]�x��`݄xQ]�j�]5I��$v� �ݗ�I{��~��'��~��>:0 ",� ��y;����4#��K�j��9Fԧ"q���Ÿ�B܅�hq䞈@�ۻ�`�k�Wq���v�a�trk,���nJ�[��_|��Ck�C��v��t(�%9R.���KO�5���#��nB��Ct� �d#%̥I8ۜș�R���]�۩E��;\�'v{*Q7�%4e].i KWC�v�Q�zvh����#4�l�WJr�UL��s�y9�=]U�V��y1̚�h�S	r5pD�Ӧ���댂�2�&1Wp<��1�^7<���$0v��
�m7����E�j������:���wn��*�M�4:���5wb���T�����5{޼Kس��q �Θ�J��)SV��^���Ix��j��x�qAҤ��:aE�m��$�Mp�5wb�UW8�~�� ���U�����-ۼMp�5wb�)���%��3I�<i��zU��3>�G6R�Ν�;Sݔ���0��h�ϑ
�����3o�߱݊����:�����j$�W�h3[�o}�����Hyy�.;5{�^����+�:��WR�v+�ݻ�5I/ �\0���RQl���׀m�wL-�W��Vջ�$�Wv+�"�/ �^ݺZ��q�����f����Us����}�<Mp�>]د���BN�mxo�e��1�6���\�\�:�6o=<Lr]�m�u���6�,vM�;{�w �{��&�`�ax�P�T�l��bv� �^&�`�axSe�mu(����M2ݻ�$�V����=��b�B�#��`����sꪪ��s�{�j����`��t�un�t�� ջ�$��Ix�\��L�E½�~��Z@���x��j�/ �\0]�� ��=���ݺ$�\��m�u/8۲>�0]��N(co7�ǈ��7��p�����5M��I���_��ϐ{������)ҷe.b���%�Y��$E�=x��e�Xv�j��q���C�m�Wa/ �\0���$��-����<���!QwV��$������Rz�	/b��(8�9����r� x!�w�����_gZ]35�$��]��"ݗ�l�� �E#�5M��I��!�L��;�BFJn��v��d(���{s��d�7��.���gW]�M;k �{�G�j�/ �{�v�m���[�Zk �E#�5M����<�	�Y��F��W����	&�M+o ��׀M�� �{�G�uݱ]Gn�
�,.��6�,e�X�)�\��O^�e��)ҶX��[��	/b�>QH�	5ɹ'��]�>06@E �@$	~��	����}乔�ffkS�4\k\��M�m�;�����]r߳���Ƚ�9X����=��s��j�@�"�O�/nj�9�;�I��a^1�ms.έ��뜭ւ�秦�6����m��A���l,�v�J%�P��KE]M(줏p��<�v)k ú}c-��v�<W��xaxx�K7��N-����x��L]A6�h�s3�伶xI��fK�|BSK	�e�p�Ktk.��na
d�"��E,�b�؞� �*َ���i5E[�)�ƇV�^�/~x��M���ϐ{�<�����IҶ*T����$�v�,Kذ�<V��*�Qm�ƭ���X��`�$x���D@��U�E4�v���, ��� ٮ��Xy�8[n�T�Z� >�#�6k��{�\0JlE)E�I�C�Gl��uӨCs�={,q��q�&݊�w#��"��.b@��t��ﻢ��u`�рen��:��u.��%a,���ܓ�s߮�4AS�j�~�ʪ�W��}0�{� �6^~�$yzo�#6n�g7�w� ���� �6^ݽ� ��-TU�e1�4]�ـV��Se��ذ=ʥ=3� ~�I�bmYti
�������?m�X�p��dxȢJ��`S0��3H k3f�Z�b1���DG�n�ĝ0@{+��Wh���U����������BG�j엀��DQJ��4Qv���;5�W9ă�H�]��	��b�H�.�+m��;i��l��#�5vK�N:�ʮ%T���
��V���>�O9lY	B�k!J� N[40�r�4$Q�j����-��P��)�L &�B@�tb&�LŅ�8���I��J�j0�lZ$a_4��P�4�3A��V�U!�F�@�]Z
y�T���8&���y�`l�˾eƧ$��%��o�0 2��3V�z�FFCG��X���iC�20�p��|���ҿ4|lq�t�����ɐa�� �=JD����R��Ԟ�jc4�7@g� a���y��h��Sc�"�	2�3P���µ�7@FMe+2��f 8z�َ�G�	N]��)�I�)��, ����A�00X�r��]8�.x��#�`n7.��6!���y�A���� 8�C� b�"� }D؇=U�
(�T���"� �����m@C�}'�AJ0�{�3�_�r��|���¥|W�SC�ݢ���*���x��,�\0=�Uq.������+�;j�Z��w�M�� �� �<Wd���J��e M�Um��)�#7*�h;4Z�������>5�j�琨uN��b��ݵ�M� �<.�~�W9U�K�_|�K�QQ~E�V�J��0��y�vK�7ob�&� ?���fnκgΎ^�����{7\0�����m;N�; n�7xv�,n�{���=�q�@�N�8��$$``aP0�eU�.s���nI;=/�QJ�e.��X�p��dx]����X�s���Q~�ISWwT�b�H�d�	�^�Uَ����Bݚ�֞^@�`��vU%�ji\���~������;��z��s���\~0��T����������"엞�s�<�`��`t�窹U�H�T����5av*H�n�����\0�H�]��	{�v��1f��i�����׿^ l=��<�8`�J�TwJګt�wV�X�$x;#�;#�6����w�I N���-�8v�:[��r�.�٭��ňNܛ�p��wm�j/Z�cp[��V챀��I�7�5p���f�u:�'��ln�qڰq���م�ב9��c�9z�y8�W:��U� �v�,������Uv��[,���`n��'�����&�[#�_��;��}WI�չM �!ӀVn,��]F�$a�`ι�y�T��-��ͩ�=W���&�?�� �"
o|�5�Z��95h�W��f� ����fC�N;{��9��vq���f��C+2�����vG��/�|����{���ݧiݻ�v&��0�p�5mIx��窹Ĉ�H�)x,8]�ـo��jڒ�{#�;�� �M�-7o���;��`[R^ odxv8`��}5�]���6X�un�{#�;�� �� �ԏ �Ը'�ࡹ��[pCj���Q9z�cQ����,�ܠr�x�WYKX�nHx�Ep)[���ٮݩ odxSj+�R�]!�b����\2�9�P@A�d$ �*��S{��< ��xdp�?��ҩ^�]���ݖ����< ����ᇼ����׀�l��vm�f^ odxdp�;5� 7jG�N�x[���*�M��8`��`�Q��G�{���'��H�V#�UZ �Gv/C�{U�Gp��z -��H#��z҅n�v�!�cE����m���� nԏ 7�<�8`U6�����;�v� ݩ odxdp�;5� �Tj��Gj���WV� odxg��n|}S��)��~��������:��mڍ5t]������n�p����	��K�|V;J˫��n�`�Q�� �0����EӦ�M7-(�ܦD�F\��7$�^��ɞ1���n�8�N�����M�fe.�e8�{:�vG�l��p��U��Ch��M�� �0	��%G�ou8�c�i6�&��8`u� 6J� 'dxWiV�J��i�`u� 6J� 'dx��r��	 ����<�y�뿺p�w�ݕ���,�' 6J� ��/o��{��7\0UUy>��|lF��hd�*k���Wj��¬f��L�d�����{GG����۵m+�� ��� �0	���U|�/z�x��QZ�M]Z��+J��6Gn�`��x;#�s�H�/]մ��v��Wm��~0d���RG��x���V���j�[E'uvف�q)�W� {}�l��p�����Em:o 'dx��M� �*<��TW(+�Qb*��9!e$������Wm(��SA�;���E���T;�(� \+d�77^z�3�Ӻ�L�����p�~�|qê�q� ܐG`9Ө��w.gc��NN'�;i��c����N����9�;tdWk�n�9� ����[)��`-��Ĥq� ����L�X��[���tC��S�����j�%��\y�l\�z۸�����a�BTf�����*�M	��_�I�&䜒]&�G�us��E��Wە`w��s�m�p�6�iwA+'n�I��MSE@ε_�w�_�6�, �*< ���~[{J����.�l�I�%G�lx��v�m9i�M���jڒ�M� �&ǀ}*5wr�;�C�������0M� յ%�G"�j4�t�Qe�����lx��/ $��UW�����q�Ё��οaB�-aj��'-q�̜j7XrHu�(�����Z�:vF)������RT� �c�6G�EZ���)4���x����W9��ҩ-5��.ErA O�5'ny���&ǀ���N�4����� $���� $��[R^�/T��]6�T�;o �&ǀjڒ�M� ��U�R�:�8]�ـlx��/ $����N�ӿK��f�4I����mO#nhFw![����`�m�w
��=�ͪeh������W�x&ǀvG �}��?�:ݷt��6%���	6<�8`��jK�:�E�����"ի����lx.R���`H�@��u>�;��������÷6�t6�l� ;6<Vԗ�lxdp�:�Rڍ]��C�Cm���� �c�;#� I#�?Us�ۭ��gen��r
 ]�ƣ=Tvy�H��H�v���`�pL"�9�
�;�����צ I#�5mIx��ܦ�][`��v���vG� >�< �< ���]���R�WcG��0�#��#��q#uǀvG�Sjcn�aĕ�o ;�� 7��01�D�F�3�k�(��f�����B�@5�rVD�H� 9�5�$���+��I�*)���V���ǀI0��a#�=T�%/]]��P>E�݇���ܧ78N��qC9�nɼY��l���)��e����p�����G��պ���umұ]]]�`�=�H6��< ��x�p�:�R�2�&��-���#�	��0vG����N��mҡ��m�{��q/I�I�� 'dx�w�x����8ڙB�gW/ �c���r�����z�����9U�_�� *��T_�( *�AU�@�
��P@U���������(�2 �F�
�H
�b�B�
��� �" ��� H�"�b( �@_�P@U���W�
�P@Ux� *��AU�J
��P@Uʂ���_�U�U���
�2�Δ��
�������9�>���>��h�Ӡi�X�� R��h �

H�H �čk#��3��x��� @t 
U�� t+m��:t���4
  ��Ҁ(�ӻI@�
 �@  �AB�     Z

�{3J���mtz[��>��>��;�}���w����O�n��w��`9���Sx�u�݇    W���;ءxt���fϠo0�7��x�{��{�ִYޣ����0=�8Z;������� ��lcZ(5@�w: �� d�{���璉�}����_X%�_T*Z��c����֪�h�>빗]��k�0>���   ��`����t��ٕ��{� ná�}�b�r�E|������� � �R�^��>�Exǻ5�O�{��-�$�hӀNށ�t�罠_[|����<  �m=��=u��\���:>��O�����L��@�X}����� �3 ��>΀�[���l}zǾg�>� .�Zכy��� :S��
S�� 鱃@�#�f�)�w �� @ [�Ҕi�g@�z��' L@��Gs:P)���@���s��R�����Δ�����P��A@  ��CO@�5�](���r�C{��� i���u�t���w{6�u����z�:w��{{٩����Ϡ{�p  �������k��}����������`�>��k�=�|A�ǡ���� "~�Jm�IUC#����R�G�T�Q� ��eJ�==R d ���E<J�  ���U!�J�  D�5) �5=D���?��u���d�O����s��U�5��DWJ
��W�_�@@U`��*���Y���?�T��$�e��!%$�a)j��g�h�.o9<�xM��(t!���| �0'�d��Q�\�2�	��9��B�$	Ą�>t�&%�FB\HB�7υ���,%�!8���χ��︼�,�R��y/�Y����6�K�׻�l�P�$��g�In3̴��fg0e֦�8&�\��3����7��)	�o�{O<�����������y��>��>We�ϳ� Nn��y噝6�!q.n�C�K	�/gs�]��ܦ����d�%�ۼ�����&��o=��k�0��&2��dp���L�m�f�B.�M�S4x�|Ŗۋ���7���MBB#Nk8e�|�J����	 � E��p��(`D�Y�\�8KM���{�X��Z֥Mf��B�!)���sw��&�yw+�'�5���#7���)�4�!f�X<HCP'�m�%&��_y}����e�3[���[&��<�hO�i���H;6��M_:b��B�/��(�(���b7i�s��Ϸ��(H�B�%�4CY���D��WWSzܸˮ��!w������s[$��7���|���5i�H7�%�/}�u�c��T�a	`ZJA�u$L\;0̈́
BBj�&�¯5��)�r��i�$2\9)B��X� Y)`�%��xRQ�HR5��b|�K�)
``�+M�>��I���!�zIL���S�cC,��'��fsF��7��}��/F�j����dCn�$	�2�eK�1�	���|�4y���f얄 �I�P�Hnm#�շ�nS�wN�ם>btI��5u�xJ�6��s�o�^s���	����2Z��	r��}���g�F��s�}�O�yFUP���V�9�tq]P�>���j�:/�>[����o��˭����8���k)�F�i�!������5�BB��%֘m�e0�>5�y�vf��ĀK��a��.34N���މ����̳�o^;(I��	�slM�26����fp�0!�ĕ5�h���l�|�!zo'�88�N%�g�dn$a>�a&����	PHf����*B�RB)&��YV�-�Y	#$!�ϣxoi��sS>���h�
I��qs�7wބ��>BB��@b;W]���9EPfe�Q]VӬ;���.-���B�Ɔ�O�ђF,JHo.��{��n�吅�	+�`��f��B4y�6��>�%�BaB1��ex�����H\!s�S4¹�P�א՘�zB�R�
<5���C{�
�՞7�a�i)$�Yr����p�KyTgݣ��_P����T[��Y����^p�	��K�]y�L���P�"I ��R�))�K�^yu�Ĕ�HHJr��k�3E����!l�\��"��|���3.��m䬚=>���8,"a��^�y���K3^������.y�W�۫��HնR�<挓ӄ�P�N�r\e��h�H$`��W�'�]��6�}�f���r���ybC��l���uK��)a侱=�5X�OV����j�5�1�8�Ë��L	s��S3�$ɶotc
e%6K��r�����%�"\��]���YI���ri�.r����,����2Dܦ8)��P���CB=]��=���ȠY��YFM6�૖��u�Y!	��y��.0�5�5�ځ�]�!$����	-�o7���rY�T��!��a�	9�{���|	KВ����B])s'ބ�}����P,XH���K�}43E)��H$ �2�
��j����	 F2��E�����:�-9s
��ݼ�-����Rnh4S� �I ńH��k�����'5��|�I�b�'���J��IIx�BSt$Ё���[ IU�0�$#˚a��lљ5�n�i��JFRF6R�v�7n셒��>Eo��V�C�Lh���3�>�4}|�pԸi�!sy˯L�d�	r�n��5<���D!�lq���K�4�,� B0�	d	"�a��2��B���!��ae�HL��+� +�*Ő!&��6���dI:%Գ{w������3i�o���)²����R6o��o�p�^}��H�}��$4q�L�:�����ђ��xrE"�Ʋ�-��`E�53Z!0�J$��x��)�K4��:�y���2$H���.�.��o3�	�+��\&k��	�����K�����29)ɚ'����T <8�!�~s\	��3�aHҘ��nf�}�<��<*B]>uy�>|�JC�Eb�J��лOK�隮����ONa�	�������9�]C��+
�み5I.Mo$�8��%Xf\���)�nG���[����Zj�	u�ua��ˣt�ԙ���{�0$HDi$#0��淲GE��!�`K�}�xn�����K��,��v����Ü�L'>�>$�M�S�)�d��ZֳW�ل���㹮iY �$	r�[���.�l�ÄpƦA����<�ܐ�<�k9��U���_8`FN'<9��%p�.L�'9�0��RZoD)y�]/�N}$=�ͺ��B$X$H�.zk�����u#5�� I�����(B9��Wh�����[橚��d��d�J,
@4�a�� M=��zA��)�p����"D�$��)�,,��$�H�܁X��7�a��4��kRA��a1%&rs7p�i����
B��
"b�˱��	�34;�������>I�Vr���y\�x�˸�6�����X]�:��a����jf�9���I���y���sS9���%ֈC�@��f��bF+����KOk�H$"b���A�ɸx�H�v�Jy{5�#p��.�����L�0��	��Q>���0��B74Yn� �vY��)�O��++�,dHO7���Np��&�M0Ht$	��4XU�o��~�ύ����H��Z2�}=��[�l�I�Ys���S|)7�p��xF��즋�	cc!���a��	+�6B��,d�*1�5��;�#aB#`@��2Fx�	��x���Bg�I�y}�p%��s��%�Z��8F�줘�{�k�!o��L�g5���?����Ysd7=�$�3�4��K�<�G�z|�ƵJm#`T��sWp�A�IHJ���I�[�[��Y��A`�	'�ө�<s2��,7ʲ��9�a5tr����c�����p�٩�WG.�)�"2�=)-[�!5�j4�60���>_B� `����˯|�6h!�"��p%���5�����PbcB�%!�K��-l��h��7u�o5�2g��ȗ|�*B��I˿�\�0�{������0�
B�͞H}Y�{L\4r0����VtJ�C!�k��6�a
�5����y��٬,�K�t�H»��|1��s�nl%�_u�k͛8�{o���z���f�	�.�	�j;��f�q�#G�!$�{	�'������i�B\���:�?x��;lʀ%����|t����wE�$l��n\4cH�0���_35�7�!��.��l3/��^!�^�Ny�!��.Cf�D��tn�W$�BYb�4�u�)��c��K �!)�H�(F���BA�%�ᰇ��% ㎁ �)�eg7��B����0�jD
�A�,�!�#I�'��4�\'C�]$.�A��aL��P
l�r%50wo<��Ɖ#a�#�{�E���f���|�ɚ�.�7ݷ�	�H[��I�M�{���6K��|����M3JC X@#m�0�`a!�|%���߉�H��$$���=�#=�k��$���H�?1(	mc��.�q0�FA�� �
� �\!dF"Ї�x�,d,S���㊷#���T}��.�eV��
��U0#H�-leJ'�m`����|�
�\'	�U�)k]���U+��;[�y	��}�9���Y7'�~|	sSfP�hh��d�����| �p��X�	B3=�rH��\�7���2q�c�0�
�,�Jd`D�aq8�|�8�$�8��R����w2�^.���Kz��7m>����%�{Ô�!RP�$�!R,B1�Xg�� C�P��6��f��]���f���436;���
�����q�Mp\U­���ٙuAʢ��z�}ﳅ���!L(ə}�19�K�}�k��qv7w�:ɚ�0�-��aJ��	q�_�,�ךg:�3� �K���\�Ů�Հ.tv���L�*��?�U�
�;�e��!��������<ѭ�����
��w�e����G��B�3g���ޓY!3���C��ܻ+������[����Kl-e�B��M	2Y	�1a$.$"X�3��kb�-��a����HӁ.V�a0�����G0��S|����[���N�:�M�[ڷYWxÏ��w�֙���4�v�)MM[�7M��U�	cP��"V�g��~|�%�ĸ��م��	d*GD�7ҷ��~��u%!v>����G��*W+t���E�s��t������7y�*(
�e��I=�k� �%��m�S�%���u��0�K	�x��)�}̘}����˚�g'3y�9��ѽ���7	w�e�e\ۧ1���	,Kr�6h�`���M����w6�?������K����}�k<�,1��̛Û%��:�Џ�ǎec���[��c��
�\!/����!&�	I�.K��B�({sa3�w���2nn܄�b��\��}� K'�q8�s�й�X:�=8��<��	�o���36�|'�\�P��C�|UUUUUUV���������U�U�j��U���U�����������������UUUUUU���������*��������UUX���Z*������UUuUUUUUU@J�LUX����A��3j��G���+gsV��^@���kmj��A,���(Ȗ�X/K�J���$0;tV�j��M�kc(ю���īr�*�[s��T��+`��U@��Uj�VI���+�U}UUUUJ������������V��%[TZڌ�5[UUUUTs� U!u��UUUUm�Bj������X)	������j�z��vh8���v�UUUU��[<���U��%�]��U�6�;l�c"�J�UQF2����.�f���<�5����Q��A%�j�:�p駐���[�5���Y�Ф�����s����4q�����1��,i�Kr[�S�q2��mS�v�*ʮ�l�bƯ"�1�Z�
������h)j��l� �*��V
��U1	�]���glr��;qAN�;Vͧ����,�ĮZu�T�V�Uc1�+]�����U�����Kq\k��T�p�
���ɸ�VquYm�^�9����lݳ�Y��3�@V���R�n�@UDt� �[muUjڗ�~5*�[&Yqڗ�l�j��ӣj������*���@U�Uj�@�J�*���X
��5�:�e��TZ���Gq�{l�媪���e�۫�]<�GZ�TU��t�� tp�L��jB�*���NU��m��M�ܐ�ei�4T5u����gS�҃ u�gpv��ʌ;��z'�($���p502�F��f�[D� ���v��
��݃p.�r�2�LMpA��Q :���(��`�kll;u�U@T�VR���Z�������U*�U�{�����U@UG	�H@4mUUr��ƀ�[V&�v*� ���� ���t�Ի 5 QTS�M�T�T b�f�*�SUJ�UT����WUUUU�UT��UU�V^M��UUT�VP�evU�\	�P:�/eP/+UmUuVC�T�u,�UZ��@T	�b:c�ER���U]Ue[��U� �b��XCf���:0ҩ���U�W@.Q�V�U�U*�ii`�mB��.U]�����V�֥��ʫUUJ�*�����TĹX�A��R��cUҬ���Ԅ��nGuHZ�����U\�@�h���� Ұ ��nSk���ڥU\jUYIm�V����
A�q�,��BM�ڪ5���uJ���̩S��R�"���WR[!�n��u���V��Z�մ� R�����&v,bXU��-fݝi�H(���E�֬Z�'ǌ�%��U:A�Դ��'�.Kj�ۇ�@�{U������R��m\����mq5�q�[���%��c3��v#v-xE̕�S���DjR��$t��H�6�J����a�VJ]FW���[`Y�t��8.��#D�4�F�M���������,�O�<춆t���=Fz��c����!m<ph��K��KM�,-���W��W�;�lO[nG�������N�Z��z�\�=���	 �5s(�2��5BX�Y��/�nv�I�Wm���d\�N�c����n ��	e
�m^V�(�m�j����=q�mKQTd%�z祐����>9:�um�tU�Uԯ4��#GL������s��ҵ�8
[�gj�CǮ$s҅p!��&F�j��ٌn�J�A�"�.�9L��m�U~�����;q�eX/Q����5���֡���HF춳���U�@l�-�Vl䁲��TR�:�(��n]��:�#��]FFVu����՜�E3����˖ݚ�K[m�Ul��^�K����g��l�5R�Q��8�m�m��Vܳ0�h��%+Ҫ�l�) ��mU)!�O;L"m�ܣv���=���L�U[������l�ZX	k������=;g=<��Cm���$,���We4�*���`p9
�vϘ�],84m�
��bр0.A�*�ἶchxU�bG �A)f{j��
�%�N��Y$����TZ�D�V[5l�n	@�A�D�i`ј�
o���&����@p�qe�/[e!m]ր�f�2�
�Xm��e��+�5z�R[�$�.c��僈��@��M:'�
{"Y�<l��d3�h��qo�"N�-T�R:ѪyZ��@畮�"��
�E���g�Ų*�Z@�@�+�Md���Uqgm�4�8 9�}�R��nVH���[;^����#��h�hg�Bj�i9j�^u`��TN�N
9[���=����juЭ��3:�V23%�*U�\��� ���P �u�UUUq�UU��Q�x
�í�h*�Ym��j�P-[A�Ҭ���᪭R�j��$��k�Ǜ��ʧRsm���f�
C���7�T	3njy��Ojq�� m<���:����e�n��Uu۞���٠*�z-�x�YZ�a��j�8ۀ�y�YJ*��;)��QV�κ'r�qn�����/Ò�z������Ԫ�Ȼ+ �uP%�M*A���V�Rl�iμ�8�V�m*P=����}�x��
����+.�9�� ��j�*�3 8��A�z�J�;�*��S�p�U"a��v���7@
��*��B�[@�	s������_O�|D���b�� ]���%[�m��+��<��a٩�.�m��W���W�tHQ���U+��ù� &����z�\5�U���k\H�S��WY�i���۶������l��\�h��1u�0�b�%��6Ӹ�F�u ���l�j��9��7�R^��=5[A�����[�a�1@
�U�tM-F8]nq�K������wJ��xɪ\��!ۊP 6�l�kC�W:8��jԇf:ٕF��@- V��j�j�e���[�d����d��r��MH�
Z4���0-5Uu4��U*�ŖS�P#-Qs�pdQ�\�۞�mUUWUT��\h�B5J�S�WktT�U.ϘrҭU{l��[Un������+T�$�l���`n��n5�6�t���g�%,Q�UUUUUUUUUUT5T�eiV�mV�
���!�vļ�on�zGy�S����(L����2�!*�7lUUiV���~ �����a`������ۗ ��c��A��1�v����r��s]�Ru�M['lHM�>�s�i���lMi*��(5m�[}�{ء��ڼ�
����ܨ(�eZ�Tg��[H�N6��յUUO.�j�ȵ��v�cSKh�d�5��\�X�%��ҭUU���UUU�T�U���
��+�W[UUUUUuU�j�Z��
딖��Z�j���Sj��y7J�UV*�Uj�*�2�4�6|Վ�T���mUU[S�y�P�Zڪ�Mc�����M��^���ñ,U������h
���*ڐUU[U�����Eͫb����6vO��7ݴ�W:*���UWi�,X�� Z�b��U!5S�kko+�T9WeRU$7=uUC�uMJ�U@r�^�MIUP<s�k����m]m�&2[-U�UUUUUPlUV�J�U6ej���������j�iV���j����Z���Z���>����ꫴ놠6����r������\6xp[��UR����1|�m�Uj��f��]�fƳmE��UX�\��@S%PUU*�����UPUX��nvB�j���Pbf�UUAv�2�;���SUR�qUQ������
�A�d���v����\a�hq��n�UJ�UR�ԾX)٪��*���kj�
����T�������
��,U�k���*�Z��5T� 7���y.̫�+Um�["c���duLb��=����]! U@�U^��٨b�Z���P��T
�i�n��ŗ7�K��Ԫ���v�[U.�YIN1���Um���PU��U*�
�UR�f��q��t��[I'Y����';T���:����Td%���*�N@�ӡ�g
� �U*U��cAT��2*� �-�ي�D�)6�U[uF�x��V ��T�V�u<��h�P�t��la��YP*�h�O�`ls�+*�;���oIё<����gB������z87P
`��JZp����[�$)���s
�6��X��Q1\��D���i����=*sԹ����m"sQ��JJ[R���! �N��	�m����-T�)��k�K�6���Z��c�p:x7������X��ʵty�N0�J��S(�F�)�h�j1�Q&{m���_W�UR��Y�V���k��ؙ"�,��E2��Z����������m;,�X+oI�#ok[X�Z�WX��̊��]�z��H/  �\�=�rX�]�f�
��6��U	���i�`�/	�4��)AuV[B�V6�rUUU�F�/`j���һA �T��` A��k�(��n������ʵUUU,��|pm���UJ�V��#v�UuSuR�%Xծ� ��UUUU@UJ��������UD�H�*�����@Ѳ��5J�UV�UUT�-����9�55J��UUUV�UUR�*�PTUV�WUH
�[UUUUV�m*�J�UUUUPT�����WʨQUW`���5sUUU[U�@U*� ʵUUUUUUT�UUUV�ԫU[TUUU�T�
vF�
������,�J��-U �Cl�B�alU�0 �	�.ٵ�EUA�UPm �2)-mUUUmUT���9j��X-�ڥP ⊨ ^Q̻;[N��-�U���B<���+��� _��������k��
�~�Q)�QxD�*��Ё@����"� 	 �#� �!$}D���dP5�Tڏ�Ea���Ď��	�<\ �>��6!�S�T_D�"�Om�.�^ �s$��*���O��8'�H�Bx# ~QS@�Q@���� M���x��CJ���=��"�B
B � $��x��z!�Q���'�'�GԒD�0 I"1!	!>C�x.�v�`�_�v�| x!���������@	�R��|__Qqz�eE�P<E�
z���fi ��������OS``��+È|�DGh. � Ҡ);Y �!�qA��D��
�!�6�R:AS�0��> �AS�C�(= U���`�{ w�|�~�Q��4�P�@	b���|�1"%P�H,�A 0D 1
 Q
 # Mi�� �b��8J
c�B����	�=" �R1 �[T�H%�d�#B��%�1��T�
�
E$�e��%�	E�$%e �Fԍ��ĄĤ�$�İ+@$H�h�6B��
H@aP�d�dbFX!(XK!D$���.��@Z!=pX:DC�`�)�0��4@>�A��`@h� �A� 6���
���@"PZд��0���T�JB�B$"#b� �b H2 B	�f��;�kZ֥ ��V�UUh��T��R�1R��٩�Z�R�f!yv�<��}��$JڪY�brCjUjtW]�P�R�ls�lwclS��&�ֱ��*�vE���⨌Y �@�z�����x8%� -A�֋+��U�,5X8,4#bL�)�Tx(��wm-E�<k���	ݩ�F�g�̯><9;O�/c!b�!`&�odu����p����uR��a��Bi�IJ`��X��<q�ZM�=f�G&ZV]�-�x8\��l�6����{k;P�@6�؍698N^wg�ܛ�:]O���2�e�8YW:0(f6�܃��5�:9^��
'�=	ڬj�sc�ȝ�z�8��)+��Ԡ�Hu3�b"zƤ�4�	��.���U\gS�Ȧ뵻�d�j�2ݻp��C��
��e��K�`*ٔ���m��@����&�WSZL%�e#K\eA��̓I�^4��*;p������&��� �%3 -֬�H%���[cK�Z�V}� �ʍ����s��[�v'p:x�%�e�hd\ի,."�!0t0����x�NǱm�����=&���fn����lE;9�'���o��1�d��&�cZ�DB֌��=�/;���.ּ�:ݵQ&.�e#\�6n� \"5ka��: '8��݌����s�Ͷ�@	�e7\<Vy��3��8���l�{v��ʨ�ҷV����6�KW)=���4�W��8zcѦ��hj��vv�K�l��f6ε=���A۝hBC�٤v5�4U�xRv�3tJg�5�ݠqъ�8M̠�m���֮͐�n �5ЩK�!3��c��F�� �e�i��a�4R��H���Xݰ#̜�;�<��j8�,��i���p�P4 ���k,s.�%*�@��F����19�N�8��A ���U�+#�"4�,sq�[��VۣP�!���e�ڻjVU��Uc[L� �=RY�$��.��� �炎M�m��u�! lE�Y9�sNI�I��<�hW���T�.iG�ASB����
 |��> �h��h�X�{55��њ��.d�@�/[�W\m�(�t�,cA6JYo
�v����;7X�i��B��Xؖ�RZ�+��������Y3����2.9�y8�Ӭl�՝4�u���p�W:5k�H%����p�Pk)��֙�W��ś�d`)��T �;%l�S�1�Y������[��
!�k����A��e��j��,���{�zw)N(�&�/�ܖ�-˙�r��p�<m��<��������U�-]�VWv���v��;�e`�m�w{� 6lx��]	[mP[ݻn�M�:�l��vG�lٕ�}�5|H,J$��i��6< �����r�)�� ��<Kĉ,�V��V�o 'v<f̬ ���fǀ}ڂ&U�Lb���x͙X]�x�c�	ݏ �9�W+��z��Mqk���恓X�[�qX�F/��1 A��4�6�Z�Ԯ�E�"j�gvߖ�^ l����x͙X��R��EC��Wx��޾|�O�C�;������y������s���rOo����i�Je����v�o �M��lٕ�j����$j5�al�����7�eg�"-�� �O<s��qw�y`�~�*��in�]�xٱ�Kذ�X�t�*�r�eLXbӜ��6�C�
�M(ۓ0e5
�0V^](���q��K<c��}C?���O<�{�fV��/ ��q"K)U�iն��>��`6e`���fǞ�W+���U��i��v���'���7$���ٹ��]��+`��yUU�oӯ �{ }�"ն�-�jƕ��5we��#�>��`ݙX��R����n�n�x�����XwfV��/ �h(����I�V�H!eBmՍ�,�fm(�9����1�[!�74�&��66VV
l��>�o��wve`�����c#\��Wti]��wveg�s�T��^ vO<�{���I;�hCHi]��5we��Ǉ��Iw�<����&��ZJRw|m[� �v<�{����r|+�8����k�ܓ�Og�de�M�V���}/b�>ݙX��{��^��I����-ݰ����f]��e��JƠA�ӌ�v�c��q��A���"��	ۺw`�m|d�V��/ >ݏӒN����um�y����.a�����5we�۱�Kذ�fV |t��E�n�n�x��x��,=U\K�{+ �g� 4�'t��ڻo�UK�s� ���5we�۱�c,�۠m+���fV��/ 7���� Uʧ\�*��r��?i���+���l.�+�B��MVK� ��(�2�o�G�*fRʉif���kgY���jC9m����Iˡ�;n[Lm�3�7a���
�vݞ�ƕɲ�#�����e�U�rm;�N�������/@L���b�ٰ�;���5�vD��+Z���r�E�¶�0#Ga�F�(���k�u��%����5�2\��=5�v��wt�9�����;ゑ������:%�C�;O`ӻ�Ω�Nkul��=���t�cA�պ�5M���c�"ݗ�}6e`�5h�J�R�VSJ���c�"ݗ�}6e`vK�Ĉ��)�:i����x[���̬.�x��������`E�&�ewV�����>��-�� ;ݏ �v^�����Z�wm[x]������e�ݑ��s��K�R�~�*؄ E�]!��:�[[΁��H�2��]�v�5"V`C��Bh����vq;�m���� �v^ }��Uϐyo�x���ۧWMИ7����_}�7ߤ��>k�E�Q�L��"FOE9�/;�nI�����'<��ԑ��b�&�:j�2ջ���E�/ >ݏ �v^��-*;�hCHnݷ���W�}����Eݗ�nǀwb(Ui%���V� >ݏ ��/ >ݏ ��/ �JD�YU�.�^�����.�cf�d
�gp�J3#c�M�c�]�i�����5���]�x��x]�x��x݉q'����Wm� }�v^ }�v^��	K���iSWn�.� ��xeÕ�r�Uw�x���㠶��t�b��m� w�v^ }�v^ |wI��ա�!ӻ�o �v^ }�d� �v> |>�Ƈ��ͤ[]�����XL�ƖT��h�U�=�M8��nj:�]d��	��� }�d� �v<-�x�9t�&_���x]������e�۱�$�(Ui�*��V� ;'�� �v<.�x�Ҥp�WV��Iݷ�E�/	'=��nI���rm ?'�Aw��|�;�aM���ۼ �lx��{�_�g���5А�/f��I`:75�we��Ŧ�t��Tm��\�gV��P3�,lQ�[�V�|���x���������Am*�m�V;Vۼ ��x]�x]�x]�x��V�:I���v�v^v^v^ N�x�1S:wwn��Ywn�������wc�"���>�2�R��.�Гj�.� ������wc�%w��2"D�2,�2�F(�"@��bȠ���L��]�$�3�@ٵGn$+��	�K��l�G��2Wl�c�;q�V�c,ڨ�W�l;.8k"� �D
Җ-���J�k�ln��kEe�v�8u�� ���q�tJ�"R��n�f�����6<�'�#�(Hl�.�� �"����jy:\�(RJ�H1 �˪]�*�y'�J&��eh�hٛ�^��hVWF�QZ��@M�^J�����,�������r�j�mPFJJ���gM�r�Ng]QrOd�����S[M�E��!���{��@Eݗ�M� �v^����v�$�.�x�dx[������%I'w/�j�v��� >�� ��xSe���%wV�ZM]���"�/ ;ݏ �l� �lx�m�Jtմ՗m� ov<)����M��}$��4�j��Q����x�w[��3ٮ
�i�:�4�uX0����053�0�Ç/V�Ov^ }6<)��r���6y��/bi�f����ߤ��������υbR�	n�0�J4!�\�όOݼ ������>�2�R���즄��������ǀE�/ >�݈N����Wj�ݻ��ǀE�/ >� ��/ �ZT�D�U�Nݤ���Eݗ�vG�Eݗ�� V��)�-:,I"ݵV�F��օ�my�)+
Wf8�и[n� !�k-ġ��&+�]�x���we�fǀwc�>��,I2ڲ�.�m�.� �����x�����A����i��X�w���wc�V�@�aD�a>8�bi����3D��h!�2S��2h4��nyd�̈́ᗜ5VRD�8�"e���JC�LH�],
��14Gt���5�^��6s&�o^
$�LD!� ���iD֪a������.bɜ_)�$�!N_��<�.ZbJ{��I��$׆���X�VA����Vk�0�'Õ�M K�J�+�(`�$a��,
H!te0#�@�S��PtF%H4�YdBE�l�c7����p7�k�D @&�Q���B!I@˓zK��h�(��cb�� ��!JP�"I��{��h6[�K��ZÙ�3L�h��,7��n�*r܁�G&bT<T��<9�䤛L5N*u�_�tU�%����!0��eP�P��2��h�����CN����yo�Ä=�|7ﻄ�E14s�W5���J�B'(��)|��'0�6l�, �U0\%B	! �D")IeH��%$!13_y��󇖞3.BF�1�10t
���Z��ֳ(Ĉ��9��Ѕ�����g5� ���޵��|ۓ�Ҍ�Dd��h�G0��q���u��3�I��e���|�<]�[<�p.	e%Hx� |�� 8!�G�|!�C@x���P�+@UIP�@�S���:�|� ��"b��X ������;{�srI��e�:I�n�;V���%ݞx7�x˻�����}�շ߾>�i͜��0� ;������G�wc�5l�{���V��&k^���%Pܶ�[��M��ey�`�ݴjd��J� )��v^ w�< �v?W9ϐ���=�諻y��S�n��c��c�� �vK�ԑ�"�y:Ut��e�m�����R][�^ o���H�Hpe&�Zj�oܤ���y}�srI����ɲb/�ЬP�EHE@��EkHE�UU�'����krN�}��we��\��v�o �vK�;_�ʯ��9T�{��g�< ��3��lE�B-Z�AM-�����f@�[�>|ԻF��r9�Q�0�������Hci7v&�����< �� od~�U|��g� :I�E�$��Ҷ� }ݏ=I�y�Rz���=z�$�_>�~�X.qW�ojzy�V�^ l����x�j�L�un�	��o �we�͏ >�ǁ�)��OD;���̤�;�w�6<�UU~����߽��-�x�����븙�jG&2�*S]�rX�k��t�O4��uy�f�U��\KkNa�ó͸v��Mo�Ŧ�n�<�:q�N��`Hu�n5t�պZ|�F\_K[�m�{.Kh���f��3��1�Wi�
�H��Gcر�t�=\Ǒ��5i�êf��+���@
�Қ�(6\x����/�ì�������^
,�:�e���%i����g���'XKf�5�
�!Bi��80���p��+�c�5E���q�gbX��?Q��zM.�ͽ ��� 6lx�v_�@OO<��T�SJ�eݻo 6ly�RGT�� ��x��y��9Ď��yX�V�)2�o �׀6<?�_�����پ����� :hK	bJ�v�V+n�=��*�)���� 6lx�+��'� :l�&�ۤ�mZ����{�������ߟ@��߯ ;�< ��E6������u:����9���dGu��n{/C�Ʀ|M�0!dO�',z:ꋬa��%�m���x�l� ���UU�l��$���
�n��ա�n��>Se���k1 <C��C��f��$;�� ;�<�UU��U\�?~���/̤�;�w�߿<{�]{���'����׀N�.j�諤��-[o��9�6g� ��x�l�W9UIOO<��T�SJ�e�M��c�=ʮs����zy��p�?r��Uvz��9J+�k,٩1�K((i�e�Ǵ�Ĥ]�^�!�5]6��;�I�*Zy��I�b�m�_���fǀove{�U�|���x�U(~��I[M��� OO<�U\�D�� ��x�l��*��<���Щ�V�.��&�e`͏"���<!	�X��2�E-"H�9 ��֫�ŝ��}�<�"�Jݪt�[����u���RS}�uzz��c��Ur��� ��®�2��L���o �M��z���}<�l�V odx�Uz����;YF��Dc��Hɪ����9�.άa&Ԭ��y�=�|K@�oq��n��~��ove`�G�r��^���`��^tr�[�Z���ٕ���ܪ��Oߞ���^�엞�r��H�<�ו4�Al�j�`���>Se��UW8�V�׀M���>��I%��YN�m�r������:�޼{�+ �R$� ��*ShE�� $Q`������Җ 0R Q�\�\��UUk�w� !��G��+i�i	�x�Ix��l����� �M��o������u��Eԃ�cF��$>�kz�c�kl�x�	4��5-�5��'(��G3!յj�V�z{�V n�x�l�W�:��^����U�wN���4�۬ �������9vj��׀j����ݙY��'�����mӺV;e�xW�� �I/�U���.�=�+ =�~x��tvRR���n��{�I{}�M���	����g���ٹ'~�+{�?��.�x�fV��r�W�������x;#���<���7�Gj�b���T��b��(ܜ�g�݌�K��4�hYS(䗝��T.V�h�vNڵ�Б�z�����'l6�vX��YRVH�ng��q�ԜM���le�&��[�ma���Y����G�F�F���'���]�Y{Xљ��˱��l���3=�NWW�^���8ݝ[�=�+KRvf8R��CLy.]e����#-�śMq� '~3�����Mf���6��/��R1srE��.�34a.xJ�Iv��C~����[�胔��fyhw��<�/ 7�?s���d�V�߾�l�R�]EW�og�{��'$�9�a����7�����z��� ��^��_.�Uv��w�}�}�2��W*�#}<��=x�� ��:Iմ]�f��?�	� M{���ܒw���ܓ��~���T߽�u�'�N����f����i�v� ;6<ܮs����z� ��<{�+ &�j�WMX�i
��.ގx��or�X'vr�]b\�P�lb1�s�I8��J�e��SV[wv��uzz�{#�7�2�ʪ��^�� ���]�B��9�������{!:��'$%��B#	"��#b��cVHX�B�X�`ȉHQ D�b!�'A95���rO��� �M����q#}`��үr���[��6{+ �Ixz�T�W�� =�y��J��]'m�����R��z�[=x6G��qw}�0�<�,����Jۼ��/ �s�����w|�`I/ �v�uw؄ M��'���IMzwg���v5ƱE�V[4#��f�s�	N��]̭���p����o����"�_��s��z����IU�J�j�����}�៿W*�����E=���#�r��7�x�U�ۤ��U�k57$�}�u�'�g�]� �RD��B0R�
�@�H, �_�4b �#B�A(Db��E& bH��GW
�����Uߎ�ߞ=���;#�
4V5�l�[��'<}�������c���U%$��;�aJ�P����wm`� �Us��g��='���ŀM�V+���[�$�;��CfD�pՈ_Bw7���Kxt&�%nC`���a&��'wx�x��Ut��Zm������	�����UUs���x�ԒMZ�n�HV� ����r�\�ܮUU]�_�, �߿<���9ʪ�Gd� �X%V;�[m��<��#��W+���s�\�������<�Z��D]4ƕ�&���9��W��M���ݏܥ�t����P�ME"�CDY]R4]f���馌X����DtOB��Tߝ矵�$�~�wE��h˫�&f[������7$�(~@S;��ג��� >�< ��K�1�[�J�Ymɬf��
ny;x3u���:,��݀,ny��c�8���:ya�瘙Y]��s���}�| ���vG�W9ϐ{g���~�*LM�)ڶ�� ٱ���9UK�����{��e`fǟ�U�W)#ވu|Wj���m� ��<�&V��9\��������'l�Q*��Ui��?
��TL�~�ܒ}����$�߾�����ܒI&�}��շ�����ߨe��[� ��x�Us�+��U�~������{��7$�+�COEjJiH���}��q�"��<�_|{�lg�V�(�3����I0ס��E�x� �@<iU<L��xF4�D�W8�l$!Ϸ����;���xN6q�����̹���a�FE NNB��+7���A4�[�FF�l��yXXB�i�t��Uk\*
�����UAUUV)UHu�l�uC�:3���E�j�Vv2UV�A�*������kv�K��9�p�=^}�>~�Ң'n�.��P[�mB���J@�`��q�v�ˏ�����y2��#F����32�d�u��5I��BW��7	�-�3�P��["�%�.+��,'�����%���T��g��v���H�D�Ҁ��S�����Y7�"���#r�UZ�+X�Êz]�"�pv�r���h�a��OVø�8��n�kk�� �c�ĳQ�p��r��rj�q��sf100I��*�v�i��T��+0����|?��t�+��؛��n:P��@uݭ�5� n�dt�̻$ڍA ��5���,�5
�k&��8ڲ���c��.��M�vAE��d��Ә��gѮ��0pNxZΞ�1<x�ؾҖ\�{K�j�e�ZYC6b-�mx�.����]1���uq��g�6�\�t�y����s��[v�m4-�s��6*�y.�r�c`��\��Q�Uϊp���[T�J�6��1�hc��(f� Ҥ�L\��H�³� �m��GhT\F��C/kq+Zfn։-��!���睎�`)�7�˙p$**V�8�nz��u6h0+B�kZjؑ`]�ݢ��o�q���X#��6hF\:[�E��a0nVzvN�	�����G.��ňYK���C����V�m�e�s�dN���V-P�].��V�@���\��c"����\В���`��h9:O*�ݶ3t�x�{��1��"�vps;b��7e7/�c�π1�����Z��h�sm���@���:����Yd:�:��lr4��� j�*1�m��hrֵn"G�.��\-�.Պ�1u����8�4u����Rn֌�5�F�gF��X�E���Y��F��iV�iP�T��U�e��	����MK	��Y��j����@���V�l�ö2��N@~44�D�����C�j��P�> ��:>�@7�zN�zI���O��Rʨ�狦6rD��\��"q�4��;��mv*@9��jc=��3�mf�m��1ۊՄ�!���N���OlF��,�{	;b�yi}�`��2�+z;N�	�qq�ٕ��F�����VuZ�i4F��[�(��dy�m���kH�t������� (��K�S{kX�ޅ�e�Qø��;&䤐Ѩ�V���S����;v�sw����C��p)Lͩ]
52>$�͒=��բ�.*㷉�&���^�K�����ޗ҉^U�Uc��ݷ�������2�\�r�@l�x�j��+��m�o >�Us�9UUvO~�������#�r��IM��
ڧcMݥm�=� ��xz���$l�� v{� �h�e�v��ګl����W)-�� 6{� >����R��}X��ք��c
v���o ;�<ܪ�qv{��6{�X����8e��˻i3��[�V�=�9a1>�wi՞[�ɪ�
&0ux��w{����W�v�,�J�� v{� �ɕ�ݏ�*�����l	�ߞ�X���*?��f���<��oJ'Ċr ȋF,D�@ah�"� ��R�1!���TR$T*D��اE|�N��5�$��w[����ׯ��������y���:�l�xݑ��q#��x�{+ �t%!+ʰJ�N��o�Kg��g���X�%��x�j��+��m�o ;�<���}_ o���'�}���H��&XmX�QӴ�K��f�[�P�������5����h�N�]ح����� ;�< ���_ $���D=�U�t;�j����#�U$=�{� ;�<�r�7�~��Mڢ���v� l�� n���J�q*�w���u�$��w[�|{��1���ƕ��?W?s�w�~��g�< ���%{�\���[��Ĉ��"�V�wm�+����� ��<�vG��{�w�e�eԘ�b�)��Hj��R����G vp�` Յ������ޜ�еL�w`�|�����t y#�;�I-��y���-�����Vڡ�*�� y��t y�}���]� {�}���i��u�L�S�$�����]���/]��{��Il~k �?���FZ8f�je�?s�䟸����t ����������d���]��=|מk���r�{�/�u��evMQ2���}{��s�������RI/{����$�{�I-ةD��^�=�U��Ճ��GM��"m��t&`TI�i[UF�7%�Ut!ʋ�c��/}����$�[�?�I-�r׾�I-����߮����O�-2� ����ߪ�Ը�kI-����]�5���K� _O�B���+�`�_�� y�}�Nm�>~�� y��=��I�cB�L�:�m���� ���V�	$��?�Iz�~s=kIvC�B_2�ɭe^� ���� �?NG߿~|�����]�m�߾��[n��8F�N����߸]J�A32m�D��2�Ŭ���Q ��ׅ�v:�t'kJ��*���[@��m���gX��%+�RKF��@�m�^�]`��d�+Mgh�K��� 6�4�@��N���α�"�����ʖ�Xe�p��[O�]0�KS��-j�U�\J�m�ا8b%�yiɢ�.P�wT=s�K)X�5�����UgX��\D���ؿ$��s�7=�c2nZ������i�L�Ϳ����չ�m�A��fv�f�8� q�F#[pL1�� �����`�q�����9?��>�}:�@?��ߝ�\c0����`�q����=���}�}��u���}{��'&����EuX�a^UqВ[=��Jm��X����ݭ�������t y�^��U���]��������.��~�u�[o��˻oUC3�߾����e����Y����}���m�*~_��~����~�r�|�G�t w��tu���4K
���0Q
j�	��$�l�"�]���KJ@���$��X4��H]�0�������O���g9m�zf����̶�~�u�[o�alI��uШ�+�����w}��$$���v�>�蠩�r��Z��|���9m�_u�����
kZ��ݿ�B�����˻�ߢ���ݑ���s�ʮ]��~��$��|�[u�R�gQ�^32ӪI9�ͷ����i%�?�!.�>Imz�\�S�Y�K ���>�:�l�S/]�?�n�I%ݑ��Iwi��$�]��$��)I��i-4"U�v��Z�%��7M."Z-� ּ]�"
h0��$o�Iӊ���,e�[�v��$���?�I.���$�vGꪮW{i-Q��I%���Cm;Ab�e�����NN~�r*�~������ �=�￹�ɶ=��e�ħ�#x�8� <��� �<}�����%�2 H�`.�F5`# �#*Z H�"�	�Q�og�w��`|��t {=iy��Se^���M����� <��� ��Ov��$�y��=��:|E�,F�[� �=��Nr}�ry�]m�	)=���%ծ�$�UW;���]�
�:.��j6��Q���bY���sH���0�m�����PJ��������T�^$�]��K�\/�9U��In���J�R�:��֑�C� ���׾��f_o����m����9m�zk_[��*~NqP�O~��-��a�2������$�����+����ߒĒJOy��H��ފ걆ʰ�>��m���?�I-�7�$�����%���W���w��� ��z�RR�GkK���`���X�Iwd|�F���$%ݑ��I~��������C�������@����e�ѹ.�-ʒ1�i���rN�1մ��۾SCe�I%=��ϒIm�OBRlrN`<�W� ?��!o�!w*aW��7�����rm�{�=���~�@ߞ����I$��''=�)+���.�79G��}����u}�A�9�6��}��e���� ���@��(4��w�I9&�����P߾�ﲁ�#�I%��_�$�����yN��L�Q�C� ���^� �s��|=�O7�}���b�N����<��$6�ٱk�0j���,jX��B��Np�U�����3I�lA��ږb�m��s-�$��X�{[�$q��L�:�"h�*ٴj��qIc\+l@'msk���[��g:`���sٖ;GR����z(T��V*![m��1���St�dθ`%Z�5Ev��r�e7GT����B�|i�GD����)Y��fR�P�2��B1dXA�;aa����}δ:�LM/(M	�B���v��j����u�2��K1n�)��y�Ι�ZV2����}� �}�� vG��%���z���Io��$����fX�Ua��� ��={��m�~���s��?~���e���u��6���}�	K�qH�u�~��t=�׾��m�� ��~z��,�,6�=˹-:�ͷ�{��`��� y��s��~��g�t ~��B~��d-�o�Im��I{����}�IOZ|n���}{����-��ka��T��B���XJ���D�GC4"�aiJlcT�f��؂ּ�ge݀�{��`-��W�$��G��������;Ē]���t�єv^� �ܞ��Ig�� ��B��� ���$Vh�dg�)�	�!�!D$Hń1+	�@�ģ�� �DH�#"��I� @!!P�V��J���FV�Bz��5'7���$���ܒvly�s�I��Ez����L�47x7�xv�X~��~�UU]���<z�/׀n�]v�
�]��n܋ 6lxv◁�Us�OO<ގ��C��7m�t��X�c�=�W+c���=<�ۑ`�JZ���V�V�v�%�y�8�j�r9.]��C�ǩ��5u��4c/�rH�]`�61�Rawv�=��V�M� �܋�W*�r�����߯ �*��(V�/ͻ�4[� �c�;�"�"��nI�}���U���?�R�����Z�*��	���E6^��/��0�\0���MB�{���Y6F$	���t�HA�p�-X�4�OU S�"��$����Yq}!�s��<�"&�v�6��l�U��z��(hTpÃ ���&�I6B�@ �iD�M�CF��H�����1>H@��A! dD �$A��Pk̉J�b�oF�BX0�WD�+��!	�D�IW���c	Kd���%�Z��B0`�WQl$$0�EZHmy����A!	�B'ރ��lƆC*_���� �	��qh�p��%�����zf>�@p��f)�u�t���0C�>�3�l�Y(��_CL�� ��B���Br�!W$�a��!�AHd������JX���+�f`����`��Q4��?!������0�_��,p�^ ����
] ��_�J�j�W�7�s'�^ I<���Tmڥr��6��f��^�O^���x&ǀn��ȅ�um�Cշ�wn)x�U�L��y��	6<�T�T���R�t��Ml���O]..�c��v�\nx���N#�O'�f��c��}������I�� �6_���a=�����|�wJĭ��ȰSe�ۊ^ l��ܤ�z:������v�;m`zz��j,?W�=�ߞ�_�� �&X�J������7x���x�I�~�$����<]�� �bH�F$b��0�@� %�/\�x�*��h�w�t�0fǀ{���/O^ݨ�wu9E��6�X�1���z�p�J`����Øۑe+������}OE�]��e��U~e�� �6^ݨ���=<���Qg�v�ջ��Se�ڎ;#�;�"�W;�x�m�6�V�g�� 'dxz���<�H�`��T��e���M���%���%�,n�`l0M�`]:nՊ�˶��ذUI3��vzk�rIϾ�[�*����8L���PKV�]R�P�Vt�]U�ru��f	�{fNz�v7u'��Ͷ�ۗ��۶D���x�h�]b7iaT��XR�S�Z��.�q�j�pXgOg�7ZU��8&���,�f�$p,�6n�ٺ�P��B�4���h��əW�b�/h�����5ՎvM�E&ED��dm��O��,F0�r�ۇeάL��m�3n X�_�~���ho�z�ù��M�Fm7�.�,%��:#�ԡN�)�2�G��h��R��EY�wզ�?� �dx��XvL�P6]2�HM� �`�6<v�,f̬��Ү]J�#�|��fղ^�{��9T���Xg�� ږ$)rЩ7Vm��7ob�7ve`mG�$��.�j��۠-�v��7ve`mG�$��{���x�R�=.�mθ��]`��x{1�����ݸv�Ҏ���!V�Y���Sv� �j8`[%��ذ�X�
*�)��&�T�l�:�Lލ �,! $@�E�DR1Y �@	�"�C�|K�� �ٕ�}�0���+�@��I_.��ݽ� ��?R]�~��5Oz�	��]EM��l����6���.{<0;*��un����{��e�(i���$�� �j�Xݑ��ذ�Ȱ{�R�j����;TG�1���% k�WSKLzsrVf� r(^1?��r����q�N� ����{6�^�s� �/^+�	O;N݁I���{&�`m�/ 'dy�RGt�U�y۷@[V�z}���=/����\x@S�z��׳� ݹ�}�e]'n�S0�v������� �{�H�'�x��˴�j�'n��#�=<��I~��6��x�N}e�+t]�-�ڎ�����Uc(�ʑ�ͼ���+;v1MX,��-�0je����N��y�Xқ/ ;$x{u�Qq���M�mݳ ݹ������OG� ��eZE6]1]$����6^��{��&���7ob�;�\����D�2�;�x;#�7�� �{�W9ڲ����.�`��|�N�m�XQ6< ����%�c=�B���d���b�[�}g�;������m� p��k�M��n�0�o��r,iM��d~�*���	�~0��,����*m5E;m`�6^{��$���	��`I���$I�^(���]�+V�;w������I&V����"�袴�ۦ�����U"��zg�����6��x�*��{� ݺ��q�6��j��l�7d��=�W6�����y�m�X�W9ӕ��R�`�P�B��Z)����熩j���	�<��㨬��;V�ۋ�����zn��p�
����V9ض�q(����&�����%h%�
���T�b���l�a�9���<�=�B$a�m�%cڄ"R�Ī�@C�r��`:�傗ZlM��h������c�gJ��2�	�5��(<3Ó��jJX4��^Ҽ�4��d��35[	#�	Y�QF8���u�d����*}�|a���ܓ:ŊYr����v����	��s�`F,�,BF��hA�Ҵ���>QO< �H���,wfV�����W�wL�v�� �H���,wfV��c�6X�K��SI�m�� �ٕ�j���?r��%����ZW����m'v�7fV��c�	����.�<���e�I�b��TSM����������,�+ 7kB:i[�R.Ӧ�֦ahUDZ�I�W��^��(-5�ȱF:����[]6��uG4ƪ��o���շ�7�`lp��W+�mO^�[�n�Qy�R�,�k[�{�{�� h�~��&�Ȱ��/ ;���)�-�I��Ҷ���X���U\����� �s� �ɖ�P��ڢ�$���'ml� ��x��,R�~��=�.YEݔ�RLe4ջ�ݏ ��ŀ}.E�N��xyU�Q��:wC���&�vS%c�s��f�Fz�5����fir���E���b�Ɵ,Wv���� �Gv���ݏ �m$H�[��:N���>�� ����wc�7��`��wMX�I�*��v���ݏUUUVs����w�<����R����v�	X�V�ܪJI�g����E]��軦�WB�m��c�>�� ����wc����J��)R��)�v��ș^�V�����#��Ac�c,��$l4�*M�b��V���0	�[/ 7dx���	�ab���tBJ�v���� 7�ݹ{�I�,���^��I5n�}�< ��xz�Ĥ�y`�S׀j��m�*\��o 7�%Ȱ��/ �\�Q�G	N�OA=Cbk_o|��y���pn�>
��K�`�9�h�����{��n�:�!Yc���`��d��n�
�L����^٣�v�"T5h�j�E;wut�J��X$� 'v<K�`mK⻬C��B,t;w�H�wc�$�)we��r�<�`�wIһ�hWB.��l��$�)we��<��ZJ���"ݫm�.E�J]�x�#�:���$�U�(6�]E!]��m.�x�#�:���;.E�w�u�V
�U0}4�%������"�`�v��3�P���/��+��ų�	�܌ � Ӛp�̥�Q D�GnH��"B��0�tSz�@�tM�a�l`@���/����D�..�Y~R$"@���9# ă	s��!��8{0���t�L_aT���$
���S���餄�����<�U[\�)u[UUU�-���ڪ�d.y�pG�➳��+A[
�6QC-�e�40���-΢n�T��)eB����f��
���s �<φM:V��d�f�^��b���wkH9����$�c6����HSUF�/j/SB
.���
�0�)�t��`�!��3���r�i+c��wX��Kٷ�0\�,\�k`M���+b)ඁƜ\zs�`�S�NvN�Z��\����(����2�x��Y�f"���԰�iA
�uOC����<j9��Jws��+����>8l�b�tH-ͮ0�$����Ç��y�j��8I�֙�u�<�\��#�n,�._[r�'�x�/Nؓ�ɭ�մ��Éy���3��l�����<aئ��ÔL�Yf%,ps۴)e�����L�����k�א�A���Չ��Y�lFv�R]�h���B)r.�*vu���բ��j.��7�.��!j���4ᦰT	�[1j����)K	��x�F%r�R����x��F��ǣmٟ)=�Q�,`8w#��y�7r���N��O�KGn���#��s���5�&��m�jt�1��5��FZ�B=�6��M,ul�i�"��w�F'9Ǟ1�V��;�I�i��X�]l�*�n�ض�%{Q	�I��"��K����\�
{eY��"��-/Z�-��']u[F�m�eM�3��1�;u�,lUC�z�U�8�Ix�Lum��Jֶy:Z��6:��e�.x3=*�N�Ḗڤ �\��qʝX���rU0r�������ՠ��=VC.�Xv7bn��i��5��s�Cy�]�	{u��������^[��h3�SJ���ݦ[<`�oM�*�h6�Vє���0��� ��:y�4k-�\���)�[��m��GM5Ӣ4�\�c��ڥTUj��ѵ@@O(*��U@[�q�[��.�c�B��ܫ�;,PM��u�,e�'wI	:2^�� hW�ڈ�A}~�~OM�Q����"��m<Cj�P� {9&O]h���ܶp���wWYl�<q�h�r�n�)P�ڕ�8��IƵ�j�eu&�mb�7r ����6a��E(j��3Y[�B&z���Ob�97���]9ȧm�m��p��-�c�((lM.�$��^{=<�3ݺ��1�JrqShL�ڈ���B˲�ȥ��$�jGx��G]�
�8�Q�W�m��!(a����^N�k��v-@ذ�(��C6��Ì�4(�5v�U�+4��l0�N�.�i�n�T2������xdp�Us� �[�^��\!~J��e�m�]����v��x�#�W9Ď��*���aB�n�O?iM��dx����e,e6�M��;m`Jl� �#�5M��M���/�Xe;��:w�H�Se�\� �]���!��JVY�7�m���vae4��)��\�$Dab�.�3���6�L��Se��O^$p�6�d����>@{���:�aj�cjۻue���$�W*��UW)�*�+����� 'dx�d�MeZ�v˴����`��X6G�|�K�&�v�ڰVU�CV���m`���/ �0��,e���.4�bM��|�K�7c��^ŀ�<{����
�ʼ��Pw6#�B�G���o:m��o-q˰�ɜ�ڤ��E�v�B��x�p�7Kذ�#�9ʪ��:��x}�#m*i�lv��� �/b�r��W) �{� ����� �ڗĮ�����؛X�#�>[%��
�U�EUVe��wmIx��mEƋT�Ю��d�lp�7K�`z�T����*��]Z��۷e[nۼ�8`�#��ղ^ HR��i��$Z���w����.�z��$�'.uA�G�k��(�[jNI��.�J�Jـ�� 7dxV�xdp�7h��eZ�I�t+-� �#�r��H�=��'��`�#�6X�ipB�vYI���$�H��G�H�	.��J��pV�M����g� �{� $��<��D�WP��=�9�g~�����������0�H�I�$�H�z��u�g�m�/,uy!Rڜ]���3�kM*7B����4 j
%[6�thۙi��7���<�Ix�L� �<U@ڋ����J�E�xT����$w��V$l=�'�wj;�cv�۲��ۼ�+ ;�� �we�RK�;5���U�
�wn�=Il=�ul��RK�>�̬t/j�Ui(m�IYm�.���*��ݞ���G�g8Us��*���+��e�u�M��e�t�X9��#˕ѽ��l�����5��5��Ԙ��5�K&��<$\݃2�y���:
ʝ��F��7co=w=�̈́��ҵ\l�/h�3z���#���2c�s�����Nz��	rV�ru�g�ɜ����mG3ʹ��ڇ݆�=WM��<Z�$�w���m>�q��j�ɬ���tݰoWmu����S�����a
�QGg<ȕ�7�YG�{q�s�#�)@8va:�7ny�#���N�b�VP��������+ 7I����$�J�*������wfV n�<�ݗ�ul������F[L�j�6Ֆ��	y�.�'8���ٕ�w�����J�Uһa��Kwc�5Oz���X�H����.:V"�+�Z����,������x���BK����"��g�u�y�P����u�֒C�X��;]y�Q�R��,nmv�#+���������?��T�� �0���ݰ�%$�57$��=�[��v*q(;��ǀE�/ �3��9\�	�󤕶��t;-� �����/
�� 7M� �V�*��m�+m�r��W).�y��~0t��d� ��Ց+i��'H����8a�$l'� O{� >�<���,J��4���Յ���ul�QD�6�2��5��
P��i�E�R:7M�uO��<�d� >�<H�weK��UۥvS���	$yꪪH;�y���� � W�PB�-*j�t+V� }$x��	��z�G8�GUS��*�*���� {��E]ڔ�����T��H��ǀH������hT$���lx�G�l� �0{�U-����:�B\BW.չ�zXb��n��`�s�S�"]�(���
��g�9���< �dx��j7c�6U��Z.���T����#�s�g���'� l��j�tڷe��o �0F�x�G�Iޒ"�1�$���`���d�$�����&	��@U� m׿?��w���]�S,l����x�G�{�T�'��Oy��>F�x�%"�yny�v�z_+��Z�h�V��%X�d��5��td�`{L���ۮ��|���d� �]ڈi]��m��t���6G�nǀ$x�v^��(-F����$�`#v< �#�>[���e`�J��mI��Lv�����վ���e`{�\g/Y�� ��]z�ul��J�o �vK�7d��:��x���ܓ�@�T�$EVN�I?���Z���c�c8m�J���rL���k�e`[tڑ��@��m�e�B�:�s��Z"9�:��x�z�Yul��v�YsM
jjza�<(�E�r`��N]����3�`z�@g�kbչa7ck\�.\���%��qg���`;j�q���A�DpΎ�vZKuH��l���t�0nl��]�gA���V�����EZ-��S���s�y�N���W�xh�@]t�)��Н�FuZ�7uGiM�䰠P̠[�Ke��]�	�nݕi𴛿��ɕ�u��l� �M��w��^:)�t��X[�X�� M��)��	�e`**D��YM��L.��	�<�6^$�X�� W�J�ӵB.����>Se�$����x�G�j��D4��ۻn�:M��6I��]��d� �M��l�f"��ؒ�b9���h:s2U�7��R � �E3
��4��!#Q�PZ�� [�u�]��d� �M��l�+ >�*�*Wc�WwCj�o 6H�ʡp(UT�Pp���Ѓ�HF 
���R}u�f�ɕ�]��ʵ�\,.���]+m��6^�&V mwc��%괢�mۤ��;w�nɕ�]���G�|���;�D^:)�t��X[�X�ݏ �+�[�y�W�� ��ާV߹'$=��O��qxU�
	v�n.�ٛ.f0�ß�=�ك�S�u�gf����ԩ��_2�����} ��~x�l�vL� ��ǀ|�ԤL�-ݔ�]%v��^$�X�l�@{���<�ey+�6&�S���$�X�lx|�8l����IJ[
JIK`�6D�F�c�ݷ0�Xdpd�ce$h@��,-%% �RH�XFJ�&9Dr��"G�e��-2��F��1�Hq!
@!
�!iP�H�B1�0HĔ�hJ$���i�܉v��
A!GE���pߊ��7��7n�	�]l"VQ��[�a)�����	����#%���̄2�HJ�J��P��32P�cRQR��)
K!.\*��Dn�hV�	)KJW�V$`JBp���LH �)8�	r\R�*��Q<GC�k�MU7v����o0���&`�&���b�u���������Ռ	e%��� 6g ��$�'3�I�0�*�sa�&�hT�,��G����H!��Z� M���/�3�T�
'���� `	>���U]�G�6^���I+��@X�V�u����y��������e`�u+�|�&�x�G�{��{����V wI�d*���fz&�D<qA�m.|V(�k���6�g8��-�-FX�Mxr`�Gi�ʾ����6I���G�$xˊҊ�ݶ*�m��L���$y���uI/ �H�x�n�m�4�� wM� ;6<�$��+ ��HNe2���:�����-���7'�>�H`�b�b
��"��a �(�(�Y$����O��������j��x�d�{&V wkc�͏ !���Y�iJ���vv"���v��1q	j�K���Md�9��4fv� �ɕ�����c�>[%�v4RT��]!�e�� ;���fǀ|�K�7�eg�\�A"��MRt��ӷt��I�|���	�2�����{�k��Ņ�ӻ�����:�޼{&V w���z��K}<�	�hK���@ݕi+w�od��=UKv���'���ܓ�Ͼ��<|�*�l4&J�	@����"!~��&M7U9n�8�m���+��8�� W)���jMYJ������7=� 7������zW��6�uِ�U�1�����sq9ZdݪA�Hk2��[1m!��f���8�ln����(�A�$>s�㩂��c��WЅũ��<�kgBn^36�)���y,j3�W�Ø�4����4A��ąK��S؀�R�Mѹ�����e��f[��5͓/4d�����!�;w`]����]��EV�j�4��,{K��֛Q�sq��U> ~�=���c�>]��ʪ�+�}����L�t�N�o ;6<��/ �ɕ�t���V�e�n��*��m�.�x�L�=\�$�t� o��wj;T]]۫��t���yM��� �� &�x˲^�u���Wq�T�U��� ����ݏ �we��y< �������hcd��f]���C��:��tc�l�ӱ����L�����\�v��m� ���.�vL�s�ϐ��x�V�/yU�Ճ�b���_}�7�&�#��@�H �! }��XE�@��1D�`�U��a�bT�\	$cS%�2!�><G�'>߻7$��{��	�!{ah���n�v� ��+ >�c�	��/ �$��Z����\��wI��߾��> I�|���'d��>���2�M���v[x7c�>Se��e`�lxQ�U���ի)�HƆ�-��e�,;z-��h^z�)6!5�#ݻzNݶ)q��YE]]���uzz�	�2��ݏ &�x���J���]�c���;&V }�-�ݏ �^�u���Wq�C)ZI���e� �����@�[ �(k^_��nI���rCz��p��iZNݶ� M���%�I2���o �V��˫�V5e����:���~����� �<� n�}[|�y-B�4�0�%s����1n�n�RJ^B�iqfKr;R�����;g�lݖ"����+ ��fV n�x�v^�H��m�U�݈-۬��2�wc�>RK�>�e`MT�XL��Wc�M� n������2����;��Um��*��[x���r^�&V }�������K�U]�W � H}�Nk9�nI�<���ff���t���;$���Tx�#�>RK�=�r�{�/~.���Tĭpv���n������`�	���qH9�x�h����w˱&��ȼ�vG�|���M�+ 7�H�][
iZN���	6<�$�M�X��<�s�vy=�J�]���W���7��w��}��K��*�F!�I�n�	6e`۪< �c�>RK�>����m��n�Zv� >�Q���^�����,�	�jD��E��[�;�a�3f�j`��Б�u��`����k�nV��=��\��ljoi�Ӈ1�+��>Bv�鶰.K�vy�,=��Kd�u����zS�`�Ed��m*��T]S��s�C�.�V�M#C��ܥk���E�0l�Uf���̮��ƈU�E����C��3v�4Q;��e���#�-�+YZ(L�e���,�5�
Rޓ�{��%�d��J�i�� �eI�i-�h�īi*7T��7��D9��J�RWMcN��wi��{�<�$�{��� �7eت��uwm��$�{��� >�y#ʷ�k�`���v�t�w�M�� }����ǀ|���}�®�|��N��6�UUs����� ;��|���ou� 7�H�]7E4�'V���c�>RK�7��j��r��g瑗U��X����x�K�o<��4���8�����ݺ��y<�<���3��O^��V�/ >� �_�K�}Lѵ�2� �����I���UW+9U�jzK�� �M��I�t���+v jـj�%�ݑ��K��׀n�� �4A*��2�uv!�W������ վ���`NU%�bxUݖ�e�-QWWm��uvK�;�p�������Ur����g��D�{pQrE�,�<�#M ��V���i5��-ϫ�Q���r\�9���_�n�� ;���#�:�%�wXU��"j�\Hf wv'�vG�uwe��`ڔ"E�t4��ui�o >� �������(�g>�U�p�%E�4Ԅ	0�̪9ʦ���������\JEautӴ+M���/ �u� 7�-�ݑ��z%V��hi4!ۼ���Sg������ݗ�M����8���\��yx�k���=�״�H�K�eq��Z�uu��s�uh���πM� ����7��l��J�1���]��m��c�r�\H�'� �����s�H�@l��Yn��Wv��5Oz��`.�o >�l�R����V:Wn��`.�zܒs�~�����$D�
��w��w�a˫�y4��Hf������[%��p��hPm�M[q]�NurQ��;�Σ�����ҝlsa����C��xM��T1V�&"�um���T:�K�7���U|�v����q/�]]7v
ݷ�~���_�M���ܗx���	к����MV� ����R��*�;��E����J�,��ui��`g�� ;ݏ �v^�T���w�T�"�YL�!�[x����e��p�>R���$CO�O$�!`�h�]u-N�����0��!�j;����{�bB%�ZK�3�4@|	bnԳ���u9d�]Z0�
�ik�p���.p���sz=�$I���x�D �� �C��X᳂p�Ԑ6�!kVԟSv�+��%05�k�9q&$%��� ������:�CA�(q<��a#2>��X�E<��
S��H>)�9	���!lDMk��3�"C���DMV`hsQ��˼&���F�L).�v�������!=g� T�e�,��ݻ��<��U[V������mmUYv ��Z�	��m��]�\7,�F�#�S��0�FG�mz�jUU��&���a���K��`�\6�gXѮ���Kc`ȍYn{F��eV�4�]����lT�Y
����ɺ�˸,%u�]�*4��[ m�,��\u%�d�gzM:A7%�nd���Ѡ���Cq.	v�M�]���-m�V��p�:�J���[U��sͰ���m m�����`�N��MyJt���vˇs�(j+�7&��!q���6��ۀ3L�ihA�%��4!��f;K�E!%.PiFPZ�\�U�p@���1]�J�ZM,�ņm�iH*�$����}�vgyC8��3k���Z��c�X!�n6�.U�xZ�^��04�#A0�1m����{R����q�Bw,�c�;!�/m�E�t����FW<���s�q���%�"�Yv��:|�o`��;�U1pt�M�s���G17��<\�nl	v�k��*�f�1ջ%]�F��r��>��Wk&�B�#ͺ�ã��Cs2v�l�p�8)ډ�nJݞz�	2ьcf!��هK{K(��6����0U�����{`������jA�ǖ���:��]N���&����g��vyzX���s�A��8��{p�X�˳f�(Y�;n��b��R˶��s�e��'�x���մAl�r����`�8��k����s�������ͫN�@ke7>� �m�j�)��i��LDBе�)���T���p���R���Ӳ����i`�nݸ`�vs""�k���-˅�L�C�	��bm��4�\vx��-E4����Ī`R�U���h�vfZeq( 5v��SZL"C0��;�;DZq�	ײ�k��,�Oh����v{k�-���1�;n­���n	j����n@B� ��j�ڠ7SҎ���P,��T�j��PxT��U@A�q�i�q͹�wmq�Z���6ڶ��:���Z֦hָ�#H#�i��UCo����.����D@!M�&"T	����Ns�O99�N��MWl\-MأeRv�C��|[n�#��Yc��X�nW�n�.�WjD���+B�B#.�eZ�-��;p�ͬ d�n�^z���e��ymm�����]m9m
Z�2n�!�C�Nbݓ�L<F����<o�:Gu��fr���$('d�%�+��v[r��l63�i��3t
Z�ƛ��Ak,�����W&�F�����Ӹ���3c���bK<� 8��۪5�IE�3k��%�EV4F�Ζؚ����o�:���ou� �Iq��c�>U%*���iS�v� ������ǀE6^��]�P�i����`-� }6<=UU�J/O^6?�Q%t�� �Ю� ��<Wd��� ��G�}*��Q+����Zm��%��r��og����< ��<��*�{�R���bGi\7E9�v��nl�]�����,�е�� Z����n
�h��2�j������ݑ��U�[=x���y1��C �� }�}��O��k�_W9J���;��v^�ݗ�vj�D]�ۺբ�&� }���/ �������Tu@�CV�Ҷ��:����� �I }����Yt��)ZT�&� ����=ʮ-�� n�� ����;���وww8"��G�4&���lv부����kŌjf�MtL��-5]�ߧ��]����s�U_ ���j��<+���ҧV����%�]�x�ذ�$x�V���D���v�[zܓ��f�_��7�!��)kIB�s�qp��ͮU6-2< ݑ�hx�i�ɒ�qn]տs��s�<�ߞ����{#�:�%���z��Uc˄�I%�Z�ӑ,K��=��bX�%���[ND�,K���ͧ"X�%�}���ӑ,KľzvN�ԬƬ���n��E��̈́DØىR�tH�ex�Z�g�f�5&\CVܯ�}�Kı/���m9ı,Os߻�ND�,K��{���DȖ%��}~����N��N�����M������Kı/��u��?șľ������bX�'����m9ı,K�w[ND�,K���δ�j�̙)�sZ�ӑ,Kľ{��iȖ%�b{�}��ӑ,Kľ��u��Kı/����r%�bX�w��\���l�m�u�m9ı,Osﳺ�r%�bX��~�bX�%�w[ND�,��z �������iȖ%�c>������A6�a���O�Jt�K����ӑ,Kľw��iȖ%�b_=�u��Kı/��{��"X�!y<��ۻY�;[[�e��6��k�9ݛ\�����m.<B6uXN�Gkv��<@�[�e���ӑ,Kľ}�u��Kı/����r%�bX��~��ӑ,Kľ��u��Kı<�v�L�;���5u2��ֶ��bX�%���[ND�,K��׺�r%�bX��~�bX�%�ﻭ�"X�%�߾�NfkL�˫$�Y�m9ı,K�^�iȖ%�b_}���r%�bX�Ͼ�bX�%���[ND�,K�~���9��ԗ�ՙ�m9ı,K�w[ND�,K���[ND�,K���[ND�,K���u��Kı>�I���2��J�z�������<�;�bX��c����[O"X�%�~���[ND�,K����ӑ,K��|�}���#���&���H�2Zm���1JA(�̗CU�d�	����mn�|C���=��![��ri����q�m�I��ۆ${/��5M�`8k��[9 ��Y�t�LFa���ue@�m�u$�[J��t�tƵ���y[I�.'[���B�#�]� d71*�p�Df	�F�ň	F��te$�ٝ�g�Xj�*���+5m���l5�h8�bN���$��d��v&��i�iaMle0lh��1b6/YK�R8���8��
�o5#�:
��{ı,K����ӑ,KĿ};�m9ı,K��w[ND�,K��~z���������޾Ĺƛ%o�m9ı,Kߧ{��"X�%�~���iȖ%�b_���iȖ%�b_;��iȟ� ʙ�������h��1ї&���"X�%�{���ӑ,KĿw��ӑ,~Ea�2%���bX�%�g{��"X�%��MV���榦K35��"X�%���{�NC�r&D�/�����"X�%�z~��[ND�,K��w[ND�,K�Ϯ��7���.듻�^B����~z��%�bX���bX�%�~�bX�'���6��bX�'��߿�k����+�TXlg�N�,�ـq�ZI�F)֕�-��������8��lk��Kı/O߿kiȖ%�b^���iȖ%�b}��sa�A��2%�b_߻�[ND�,K�~����k35%̒�5��"X�%�{߻��!�'�� bn���4 R"�%�Q�� �a *�"�JA RB�HR	N�` �y�,N���m9ı,K����r%�bX���bX�'L$��ve-��	�f���Kı>�����Kı/{�u��K���/O߿kiȖ%�b_߻�[ND�,K�=�c�m��
�듻�^B���ﻭ�"X�%��N���r%�bX���u��Kı>�����Kı<��}�V�+xr����/!y������r%�bX�{�m9ı,N���m9ı,K�{�m9ı,K����������i�s04b��n�͝�^{j�Rn1�ƥ���en�a��ֶ��bX�%���bX�'s��m9ı,K�{�m9ı,O����ӑ,K��U�L;n9�S%���ӑ,K��w�ͧ"%�b_���iȖ%�b}���bX�%���bX�'�O�a�^殉�Z��f��ND�,K���[ND�,K���u��K��VP(��J�cb�\ꨏ�0W��ı/��[ND�,K�{���r%��Jt���y���k,2vWΟ�K,O�;�m9ı,K����r%�bX������Kı;��siȔ�N�����)�M��!v
�/�>,KĽ�{��"X�%��}��ӑ,KĽ�{��"X�%�����ND/!y�����m՛i��,��ӹ��ls6Dv�s�U��#��Ċ��)3%��rrXK7M2[��K��f���%�bX�����ND�,K���bX�'�{�m9ı,K����r%�bX���Kfw1Se�rwy�^B�}�u�� U�$ON��M�$w��H����M��K���ْkVe֦]cm�f�iȖ%�bzw��ӑ,KĽ���ӑ,K��>�siȖ%�bw;�siȖ%�b{�N��.%���r%�b��%�~�bX�'s��m9ı,N�~�m9İ>W�"�f�f�{�y��ҝ)ҝ?��O�nδ��_�,K��w�ͧ"X�%����ͧ"X�%��v���r%�bX����듻�^B���~�:�X�]��ιe���.l�� ̱��v6���t���Z`D.�wt|v��"��.�å:S����ͧ"X�%��v���r%�bX�����g�2%�b~�߿fӑ,K����o��2���$33WiȖ%�b}���bX�%���bX�'s��m9ı,O����9�y�^O|�����l�����'u,KĿw��ӑ,K��;��ӑ,K����nӑ,K��'{�m9ı,OL$��;���e��ֳiȖ%������m9ı,Oߵ���r%�bX�d�{��"X�(X������Kı=3ߌ�M[��3NY�ֵ�m9ı,N�]��r%��*dO�?~���"X�%��?~��ND�,K���[ND�,K�z�S��ɓMp�3�� Ji�\ctC�xC]nۇ�v݂��e���ĵQ���&�fQ�,��w<*.�y ck�nCm��m��\�ð�<�Qe&�Wm+(kH�J�lD�R&f��m"1�uȞ��)�˒1Ɏ���
LrUԻ;E�fWU�Ԃ�X�X]���\��6on4�X_v�Ԭ2�n��J��f��gF�bwU��J$c/i1�ԙ�&�S,�
��"!rm7��[B�j�]��Ĕ��q6;TKִ��&E �)8��u��5+j|�u��{ı,O2w��m9ı,N�{��r%�bX��w����2%�b~��߮ӑ,K������K����!�jf���"X�%���{�ND�,K���[ND�,K��{v��bX�'s���iȟ�@ʙ���j��?�fK2kZ�fӑ,KĽ����r%�bX��۴�K�Dș�v����"X�%��?~��ND�,K߁��a��-l�_:|:S�:S��u�ݧ"X�%����u��Kı;��siȖ%�b^���ӑ,K�������:c+0M�|���N��N>���[ND�,K �w�ͧ"X�%�{�{��"X�%��뽻ND�,Ky<�ޥ�1~���$��Uafp�i-��1`�門�i�6 Yc�P��c X4�UDXitԷ5��"X�%���{�ND�,K���[ND�,K��{v��bX�'����iȖ%�bza'����ZY�L-�k6��bX�%����� D �F�"D�U��OP��Eڲ'"X��]��9ı,O��osiȖ%�bw;��ӑ?9S"X�������9��4��rwy�^B�~���u��Kı<���ݧ"X�%���{�ND�,K����ӑ,K��]�˫��Y\%֮ӑ,K? �2'��'��Kı?g�߳iȖ%�b_>���r%�bX��۴�Kı=Ϥ�v�i�̦��j]�"X�%���{�ND�,K����ӑ,K��u�ݧ"X�%������9ı-��9'�~���L�4r���8b����4�SG"��\ڋ2�au`�,6�4�9BٓZ�k8�D�,K����ӑ,K��u�ݧ"X�%������9ı,N�{��r%�bX�{5I���]R�Z�ӑ,K��{�ͧ"X�%������9ı,N�{��r%�bX��{�m9 �,K�^�/52u0ђ����Kı=�_v]�"X�%���{�ND��|�arE���"�I1�#B���ZY�k,��[Ie�l~E��H�%�@4�Yk!(�����HZ`NІ�q�C���&08E0aȟ<���˒��H���#I�d$�3
D�[)
H1bF$#���p hѐ�-�%���Y�, �!A��ٺX!�^�l�)<<�"��Y
f�s�t��1"��H�¨�&b�|��[�萌]2�
�R�t&㭅��M��� '�3��*���>��F��|�!�@�ڞ � !��<Ap(!�����z��m9ı,N�]��r%�bX����9�f�f���̺ԻND�,K���6��bX�%�ﻭ�"X�%��뽻ND�,K���˴�Kı=�'����Z]Z\-�k6��bX�%�ﻭ�"X�%��뽻ND�,K���˴�Kı;��siȖ%�b}���d�5rMk��P�k4�p��ڊU�P�r�@�{! �0�tjV��")���ez�����bw��nӑ,K��}��m9ı,N�{��r%�bX����m9ħJt����S�PF(|���N�%������r�9"X����ٴ�Kı/��[ND�,K��{v��N��N�����lU�ba�ü���ı,N�{��r%�bX����m9ı,N�]��r%�bX�Ͼ�ͧ'Jt�Jt��M��s�L+��O�K��2&{�����Kı?~���iȖ%�b}���ͧ"X�ReB�� ��N��m9ı,O>���|�+j�W�N�!y�^O�~��9ı,N���siȖ%�bw;�siȖ%�b_;�u��Kı>�W�z��5��k<��r�snRFZ��X������K	��I�SF`�m]�"X�%�����6��bX�'s�w6��bX�%�w[ND�,K�׿rwy�^B�}�g���m��n��iȖ%�bw;�si�~A�DȖ%��kiȖ%�b~����ND�,K�k���r'�L��,O�O���2��V�s5�ND�,K������Kı;�}۴�Kı;��ٛND�,K�߻�ND�,K�w�}��Y�C+�'w����/'�>��9ı,N�vfӑ,K��w��ӑ,KĽ���iȖ%�b{ߎ���5��5%듻�^B����ݙ��Kİ�*G��w�m<�bX�%����ӑ,K��u�ݧ"X�%���`�#BO���y��L��]�R��F�}Y�&L�zɋ���~>�{�[l���=��l�b2ֶ�N]V8��-�XF�Xܤ��q[�h�BּP,
�¸aA�З+0m
�1{�U�%�"�m��n�n��qͧ����r㛝�e�'`^�b]k�Q���%�f�5��r\�*q��%�"L�99�u�2��[j�,��LbA�S.�	:O��7wt����F:��xj��]���i���K`���:1��D89���:�{1Θ{Y�v%�bX����6��bX�%�w[ND�,K��{v��bX�%��ӑ,K��f�;1��R�&���m9ı,K�~�bX�'{��v��bX�%��ӑ,K��w��ӑ,K������MR���Z�ӑ,K��u�nӑ,K��=��m9ı,O���v��bX�%�w[ND�,K�O��un]L4d�f�v��bY�D���~ͧ"X�%��?w�m9ı,K�~�bX�'{��v��bX�!�=���/����j\�u���/!y��~��듑,Kľ���iȖ%�bw���iȖ%�b}��ٛND�,K��ׂ��u̡<9#frY�%�`�ɺ!|NV�g)ũ�Z���k>��܉bX�%��w[ND�,K��ݻND�,K�����~ U�DȖ%��?w�m9ı,O�}�g�֋�h�[��ֵ��"X�%����ݧ!�0��<PӸ��bw7��m9ı,Os��m9ı,K�~�c�^O�:/�ԉV�RS'\��B��bw>�w6��bX�'s�w6��c�P�Dȗ�����"X�%������å:S�:~����qz�{9p��,K��w��ӑ,KĽ���iȖ%�bw���iȖ%�bw>�w:�����������~4CMJ�vӑ,KĽ���iȖ%�bw;�siȖ%�b^���bX�'s�w6~��2%�bw��2��5�$�ːՙu�H��mlG��]��;�s��l	��ԡ,��j	�e�7g�U�å:S�:���ٴ�Kı/~�w[ND�,K���ͧ"X�%�{���ӑ,K������!���l�rwy�^B����m9ı,N��w6��bX�%�w[ND�,K��{�ND�eL�^O>���ܨ��k��'w���K�w��iȖ%�b^��u��K���ꇪ�Cg�<����iȖ%�b_��~�ӑ,K�����)uiq�5��r%�g���3�����"X�%��?w�m9ı,Kߏ���"X�%����ͧ"X�%��=�eu��g*�rwy�^B�}���\�Ա,K���u��Kı;�����Kı/��u��Kı;�v^�j��[v	hWiM��WAe6�hs-��PR��%#-�2���.a5%2uÑ,KĿ|}�m9ı,N�~�m9ı,K�{�m9ı,N�_v�å:S�:~���6�����f]�"X�%����ͧ"X�%�|�{��"X�%����ݧ"X�%�}�}׮N�'�rk�^C����?h�MJ�siȖ%�b_~���"X�%����ݧ"X�%�}�}�m9ı,N�~�m9ı,O�����;�a�ֵ֤��"X�~��?~�]�"X�%�{ӿ���Kı;�����K���T	I	Cb�[�~�<z������������!��ٳ���Kı/�w[ND�,K�߻�ND�,K���[ND�,K��ݻND�,K��~;�.j��hԹX�t�뎍�g��v���[=.:(M�6�laHh��`�Ω1M`�{�����/!y?o���ND�,K���[ND�,K��ݻND�,K����iȖ%�by�~�w!iuiq�3Y��Kı/}�u��Kı;�w�iȖ%�b^�}�m9ı,N�{��r%�bX�3�o�9��fA�\��B����}���9ı,Kߏ���"X�"~�߿fӑ,KĿ���[ND�,K��w{p�Ӣ�).j�9ı,Kߏ���"X�%���{�ND�,K���[ND�,�2'�����9�/!y=��o�PY�L��z�����bw;��ӑ,K�������yı,Oߵ���r%�bX��ϻ��"X�%��L�BтD��5��Uٹ��Bq;sv#"5z7c1�����F�;]�x�`M4��,t��WJ�>-YO� {���gB�k��vH@��!�n#Le�*v�:�pKW<�Ji�������]���K��p[26��6��`'Uұl��W:_�q�҄���A�5h� Ǫ�.�J��7 ��f��d�I��^z�,m�������^��i��t����6}a�V�[[$�l��9v��r�;�.�ђy��uY���9 ��n��b��}���N��N��~���"X�%����ݧ"X�%�{��u��O"dK�����6��b[�^O���k)?8��+������/%�bw;�si�~c�2%��:w�m9ı,O����iȖ%�b^���iȞ9S"X��읳���]MB浛ND�,K���siȖ%�bw;�siȖ%�b^���iȖ%�bw;�s�N�!y�^O�=�����1MD��iȖ%�bw;�siȖ%�b_;��iȖ%�bw���iȖ%�b}���ͧ"X�%���}܅�ե��ֳiȖ%�b_;�u��Kı;�}۴�Kı>�_^�ӑ,K��w��ӑ,KĽ����sV�c�`�a6�Q���ިݱ�2c��As�K�<q����.L�W�+�O�Jt�Jt��~��r%�bX�}��siȖ%�bw;�siȖ%�b_;��iȖ%�by�N�Ʃ��n���:�������<=���r
k� Cn�n%����m9ı,K��w[ND�,K�׿rwy?Lrk�^O?�vҫ1�˅�kiȖ%�b~����r%�bX�����r%�bX����r%�bX����[ND�,K����Xw]K2k.kiȖ%�b{�{�iȖ%�bw���iȖ%�b{�߻��"X�%����m9ı,N��n2���4I�ֵ�h�r%�bX�w���r%�bX�����iȖ%�b}���ӑ,K�����ӑ,K�����L�h�rS&]k\A�j�MaH7Q��H��{��f\�����e�.�Q��۬� *|���N��N������r%�bX����ӑ,K�����ÈA�I���M�$�~��\��@p\ ����t��޽<:,K�{�ND�,K��}�ND�,Kܞ���r%�bX�a��r�V���m9ı,O}�xm9ı,N���m9���y*Ā��&�}�|�bX�'s��m��B����k|��MGQ���9ı,N��m9ı,Or{��iȖ%�bw>����K��̉�߿xm9ı,O���eɫ��֮.L���r%�bX�����ӑ,K����f�Ȗ%�b{���6��bX�'s��6��bX�%���fgtkZ���bһAW1lx/xc�Y�F���&jq6d��GU6*�l �k��J��>)ҝ,N��w6��bX�'���6��bX�'s��6��bX�'�=���r%�c)��ѳ��<X���\�:|:S�:X�{���r%�bX��{��r%�bX�����iȖ%�bw>����O�ef:S��=���Y�R��r��:|:S����~��ND�,Kܞ���r%�bX�Ͼ�m9ı,O}�xm9ı,O}�;m�fR��$.���r%�d�b{���[ND�,K���ͧ"X�%����"X�!�ء������6��bX�'���2�2�	.�rh��fӑ,K��}�siȖ%�by�{�iȖ%�bw=�siȖ%�bzg�w6��bX�'��l��U0�m�+�y{&8����a��eJV���k�	�����H���,��˼���N�%����"X�%����ͧ"X�%�����~'�2%�b~���m;���/!y<����2:a(��uÑ,K��{��ӑ,K���~�m9ı,N��w6��bX�'���7���/!y����|j��hS\gt��bX�'�����r%�bX�Ͼ�m9ı,O=��6��bX�'s��6��bX�'�N�����hˁ���5��"X�%�����ӑ,K��߻�iȖ%�bw=�siȖ%�bzg�}������������a>B8�]��r%�bX�{���r%�bX��{��r%�bX����ͧ"X�%�����ӑ,K����	3��د�&t�c��IHB~�7unR���Ӈ����(8D&{��C��#��'6�-�� ���<ѧ	�xa�&�4�w�6�7�e�xJN!�qH��W@�)��6A������J�� �g3Q	�\$ᗄ��5�q�'��G�(o<���
��h(x�kmY�'���
[׸���>8�Zu(�) �������n}������e������^���)'���<sZ$GWP|�$�"�R��6R0�F�'��8�x�
�ደ�Q�$��wf�		���<����3�P�u�燜�<4��:�Q�Mm,�	����،ĂE"l��6�.�{9��d���M�p��3�u�6����#�u��)v[����9�pNq&Ͳ�&9���9�=�pa}>ִ2
FA�����Ͼ%��Fͬ� ����	�� ��Y���
����&&�z�ݛZ��2�s��"�l-�Ba�m[�No0sɯ8fx�bH���H�`�W9�j�p�>>��8g.%$�G���̽��_$;�</��������h�j�������O����En��Z���V`E��
��[��R�n
P"��:��A��
�T�qH;U'9w*e�� :7	3ژ3H2�Rh(ó6�����1�9��ly�f�-�)v��[�z�@꣣W�Z&1ے�M���c��1�biQ��#`Ğ^ݬ��x�e;YJd��k�3.l�:XA�y\�b�:3Ketc��Tٷ�ir]�nءm���%9�kV0Q.D�EZ�{=O��v�n�8*ų�)����3�� 6�W��D�O<6�hʊ���y٠8M�ۑ�v�S�mk�Hd
GtjX7G��:{�0&X X��D9�������j�(d�=�M�;q�����ulcF#���wòc��K�\GS��=+���ͫ�}Tr�<]��I��os갸��%+��`CC�tH�^�Q�h�5�:��]��'*��V�	+]�(�)�v��4	��&9-���Sl�up�K=�;���7n9�n҆���L-#��3����q��ۇ���6G5�Y�#�X�ue��zf�Z�m\�+kW�R�J;�K�b(�۞�m6��B�ˈ-Ae�lj�&�I;h{<��uz6���7�����a7(y5�ԵgLk-�]�2�/k�ev�hOL�C`�X- ��Ι1Hʆ��"�K�!���t�R�9+����	����fNXpn�Nl��7�evw]'dS#-7eb�����s��V�Խ�.�fy�,�W#]VT�M9�T����b����"�I��m��ka(�5e�a���:�U�jf �hW�{Ҍ�<Tf-�.���wZ�r���P� ��jM��=�^���SU��vw)q�X�)s���g&@9�n6��r��-��0y6=�c���c]lr�kA�'9���������y�.�i�
6-�m���}�����y��S�,MT,��Ar\�Tr���*Bc�1���U@����T�+��԰*��ç)4�۸d�����sh[�%�;���+�§t�SE�����@ ���*��/�� < �v;DC���rG�q�ġ߶c.��j`6�|�9X��vͳ�۷dm�%;�j�}��G��j-�`��e��d-�b$ŷ<vЭ�$ ��9nw��g����̩$&Nwe�Ԝ�U�&@�;��s��0�kܘ�n�ѡ�'bg�#����N��gj���v5����5�Y8��>����s��W,m3#rb:�֤�	쩔X9,nM�BP�0���i�ԉ|��,b�l�������L��&�2&�9���u���3ٞ�/�э�E��f����ı,N���ND�,K�=����Kı;�}��r%�bX�{���r%�bX��vv��5�&jI�k6��bX�'�{�siȖ%�bw>����Kı<����Kı;�����Kı<��2��˩&h�&���m9ı,N��w6��bX�'���6��c�!�2'�����r%�bX��fӑ,K���{gd��B�nkY��Kı<����Kı/}�u��Kı=3߻�ND�,K���ͧ"X�%��I�� ���u��rwy�^B�y��\9ı,O����ӑ,K��}�siȖ%�by߻�iȖ%�b_������dy���-��`����\���v��Bk�9D���M6��T<aA���Kı>=�{v��bX�'sﻛND�,K���ND�,K���[ND�,K߻�R�L����&����Kı;�}��r�XA�*��Z�4P?`r&�X��p�r%�bX��߿fӑ,K���{��r'�Q\��,O��?e�?j�YrkZ�fӑ,K���߸m9ı,N��m9ı,K��{��"X�%�����ӑ,K����S�c)��	�5��kZ8�D�,�����6��bX�%����m9ı,N��w6��bX�dO����iȖ%�b}�R��ظKl�rwy�^B�O>��9ı,N��w6��bX�'���6��bX�'s��6��bX�'��d�9�\q��
i�u��N�qH�a�^�
���v[� ;��c X0n
�hf��t�Kı;�}��r%�bX�����r%�bX��{��~I�L�bX���ߵ��Kı=������B�nkY��Kı=����?r&D�?g߿fӑ,KĿ��[ND�,K���ͧ"~ʙ��Iޟ���fk&j��L�h�r%�bX���߳iȖ%�b_O{�m9���az�OXdM����y�ND�,K����"X�%:{��Ȥb�J\k��O�Jt�%����ӑ,K��}�siȖ?�dL��߿p�r%�bX���߳iȖ0����߾�n�3W^�W�N�!Rı;�}��r%�bXt��w�ӑ,K��{��ӑ,Kľ����wy�^B�}��p�9E�4n�iKҵzư�%��]�܍a���Xh�	b��	f��F�̹5�f�iȖ%�by�{�iȖ%�bw=�siȖ%�b_O~�bX�'sﻛND�,K���jO���\���N�!y�^O��}��Ȗ%�b_O~�bX�'sﻛND�,K�{�ND�,K�{�B߉մ�|���N��N������Kı;�}��r%�bX�{���r%�bX�����r%�bX�w�;u��d�`k�듻�^B�o��ul�߻�rI�������Q�hs�U�P�D1�uT8�R���� ��UG��j|Jۼ�ٕ�lx�vG�E6^�e�,��.C���	v۞Ru�Ѕ�q^!z�̻7Ze��c+żʍ�tSG9�n�����z����x�v^7GR�E7CeՊ�+o >����+�Rz��<�vG�N�b���)�����x[������ >���KTT�%R����ݻ��c�>�"���<V�e�qK*"�Z�o �\� ����e�{#�;U�Dm��`2I��,��螲��J+�r���ӷ&c�ۍVZ�2t�����m���dWf��6���o�]`Kvr�a�����ʦ,h��A9t��KK7c�[����l�y�Z�K����'l�+)�`�
�1������k��Z�T�4&�Z4�	s�9֬���4D
�8jy� �hB�*����kT�\�V<�,��F�[��5K&�33SFO�� q��ƀ���trv�mi��ME4Yn�9J�HY��E�%ۘѤ,-��i�`[�+e� F��������e�� �\� �P�Ќ�h��+;o ջ/?��I�<�~��:��縑��\<�M�+�V�����>�"�:����e� ݲX;e�����6��Ȱ�dx��x�s�l���/4�������lx��x���K�`fР�۶��c�i0�n���Yw"��RQ��]���Eښj{��V�`�[c��Ym�V� ����Ȱ�lx�j�P��S�+v� ody���;ʪ��߼���� ;6<m��T��Z�j��7�"�:��x~�W7�� ;���>��������S����ǀ�< ��<v8`"TY�m�%cm�d� �W9�����Is� �;����{�S0+����6F(ӑ��ů&��+pga��l������-���6����x�dx��XQݏ >�<�*�Ig��n�ڵm[��	.y`��x����c�7��F�t:��.��Qݏ ;6<%er�QYu\���DK?4�@/9=��������7�at*M7m�
��xٱ�ݑ�ۑ`~��-�g���T�IW����o >� �܋ �;��fǀvl�^S�$�ݔ�S��f��v�'������	��\4ZB�Z��{]i�H.��v�{r,��ǀ�������<��P���5WV��k �;��T�o�� w}�onE�nĔT^+L-:J���͏ >� �܋ �;��.ur!D�!_m�W+��U%�O<-��Qݏr|x��)D�����O�~s��������jݶ�j�ڷm��K�5���G�M� �Ej�W�m*��ۉ���E�.G�BŔ��Qn.�iA�BR0$j#xQ���x�}���d� >� �$����;wM�v5c��d� >� �$���ǟ���j�^)*��B�����RK�:��x�G�I`�d��]����$xQ� l��{�\�]���6�I�����m ��xQ��U)�y���< ݑ��TMĄ��	$آX��8�N�=<�˾6��.�rep-��h����˻[nݦ�kO�&a�*��p��Tu�(Ey�Y�
�hlP�;3v4�E�	��fB%���Qg>1��8B��Ѣ4[�+,�T�����5��@����7q6hSf�<�[�s�4�qm���ɬ3�1��9�H�:+�[��
Y��n9��擭���́�F7�� �<[�-m��%�F ��;�Ns��I��څ���f��F��)�.�Ac���	5�ΰ7kcܦ+q���ְ�N�%�\0m�?O� >� n���v<�Ϊ	D@�BWĮ���G��<�ݏ ;$x�v�JVն�J�ݦ�ղ^�nǀ� }�<{������Ywb���v< ��x������]	۶6��X�x������#�:�߽|��=���f;`)4�)�������؆����&�k���n�uM�4���0�4%��6R��n���[ ����t�>���7lH�]�q]�ݴ�� �ϵ��@<G�T���͛�I����G��I
�;�^h�WM��o ړ�Xݑ��#���!EE���B��m� vH�����\�ړ�V�P�A�MS�]�]��l� 7dxkve`fǀ|�P��]Z��j��(��ݕ�D ,�k����� ��'/�l݃�.^��inݫ�j�o 7�<��2��c�*��g��{��6��Z*˻J��;[�+UU$� }$x����$od��M�c��(j�n�nǀ�ﵹ뵉�fn]>>�4��
I�@9"1���@��T����dM+�k	�Mo˒����Zy ���	�٭��đ`�����M����66ᘛN h2�F����j�D�)a%��^͵�����	h���S[�.�E��"WDu��䄂���[1׸���P�M�HD�}6��
#"�ر�<"h�D�C�j'�=0�Đ��W����f��6�[}A�s8�
l�)���Z�eə�O9�<��`��ͬ_7p��-))��!�8���i�`�1��	a��>`pAh��4g��p7!0%e�	J�b�i�1M�@�Y�p��:�E�n���t&)��"�8blPO���&ß(�� Wo=jx��~@ !�G�f�E�*�� �؂���u39�~�߻�f�xh)"ļ�X�շ�I vlx�̬s����� ��#»���Wm�����c�7ve`�G�I&�n�U���i���$軇pme��P+�9_p��:�4��q�l\�vA���*�X��m��2�����G�s��ޞx����wWc��m�� �l� �dx&ǀwve`*"�	�Ӻt+���x���fǀw�2�Se����[jݴ��V�x&ǀw�2�����4�s���U�ʲ�L �ХV�%�1# �
uP�>�]��ﺳ;�MS��e݊��;ݙXSe�ݑ����-��n�U��n��ML��!HѤ@њ;��WIɧ;KY<r��c5�ɴ�v&�i�u�^�� ��< �c�r�ʯ�n�e`���+���X�;w�ݏ=�RA�O<����"�/���9$�ڟb]��l]���z����}6e`����ǀI���qS�MՈ,m�Ur�}=�`��x���fǀn�D�N���	��۬ ���{#�	�ٳ+ ��:C��~Hk凌QssԲ��P�����{�.�W%���sx�\��^�6�mj�x����{5�:Y7,��+�h�W�Y1�;-B�Y���D��.�a�A���/R���]q"kJ��.�م%q��X��r3:���l���q�c�=��s��qZ�&���)���1a�w�`7r�x��Je�H�`�Zj�:��Փ�7R�yɮ��t2���]�K��5�ML-�%���̸&���V��e#	� �ifc@�hSF�������t�
�V����� &�xf̯�|���� !%y��M��ڶ� I#�;6e`�< ٱ竕\H���kΝ�M5�.�M�o����< ����G�l�-m6�j�E۬ ݑ�fǀ�<{&V&�pV$�e&�5m�fǀ�<{&V n�����r�mӦ����	KY�^3�d�4���t�1ó�N0gf%�J�fٛXl�U_ >�﯀~�X�#��G�w�Rڅ&��S$�\ַ$�Ͼٸ�$��X,R,Y��"�$�k�l���d� �씗����];��|'���c�	�<<��{+ �DR�RN�Ю�n��͏ &���2�l� 4ݢS�t�e��v�o &���2�l� 6lx�N�~�����:e5���rk�=���к���bjcI%X�:�)����˻I����X6G�6< �#�6I�$5m�5N��V� &��fǀ�<f̬�H��;�#)5I�o 6lx�#���UQQP>A�U@�5���nI?y���K%��wr��n��m�jJH��X�G�����8�-�2�ڶ��X�G��< �#�ޞ����ݫe!R��b\Hί����� j�����1�:��5�d�ݙQ`
WWcwn�d� ;$x�G�nɕ�!�DP��:��ݷ�� l���2�vG�uV��]�6X;�i���G�od��� vlx����0���؛x͙X�#�:�K�u_QT9�
�*��'x�z������ܓ��ݘR;mX�:�[� ݑ���m�z� ���wd��=ʮs������l��M2�a�5���C��f���3Y���f#��/k�Wi]�!��T���T�� $���2�Uϐ���z�]X]�Uڢ��)�� $���2�Iղ^z�#wʐ?4����abm�=� �G���=��{�x;�Kv��um�uv�n�=UUI{���5Oz�M� �ɕ�|�D����[����d� �c�;�e`���T$�$�$9@�$a ��DlI�}/��4�XFf��ՙ�m������[a�L��5nɵ�OJ�dC����oG�lma9��j�S���bR��@��)l�i���܊Ev���Q���ѝk�mp�D�V����;]�s���#`�����{l�Z�� 8�&ص����թ����-��4б�cV�ݍjTt�� ݊�el�a�`�案�U���E/+��3c~wԝ�:Y��#}���-n��W�hA��Dgt���'mIAٸ��q�Wp�훬X�,�ui����<�L� �c�5l��I�Z�v��v�o �ɕ�lxV�x&ǀwve]*����E۬ �c�5l��lxd�X�Rw��J3�շ�oob�	6<�+ $��	�K��eڢ����M� �l��	6<{{�����s�Z}��وV�L�6�T�m5%����r�Li�����m���ZdK��ab������	6<{{ I���"��tݍ��պ�	=�[���!
$'@!���+BBŕ�AȣZU(@�c!��TH'O}�^��nI;�ߵ�'>�� �Am��t����jݗ��<�&V M����)�5n��իw��<�&V M���ذ	#V(�4;9eݫm�l�X7c�;��`�ǀj쎮�4��V]�3U�!�RP��úџe�i��
�����i`�(�ks< ���_ ��ŀ�<�+ �D��At(�[V�ݽ� 'dx�&V M��	,�V]ڈ�T���k 'dx=�훜@���T-��JDTUs����v_���PAN�M;�MXYv�ݓ+ &�xv�X;#�	�Em��wb�&� &�xv�X;#�;�e`���^��+�)5Gan�0���'�n��L#��&s����d�kK���GDr�o�?)�^ N���X�ذU�JLwt�X6�7x&ǚ��&V%�XV�x��!V��:�.�6��&V%�X���M� ��ʺT7n��۶� �l��d� �ﵹ5��IcI�eD���Dm$�kT1,�`��!V65�U5<�;��<��Wab^C��ջ�5l��H��2����~�W'��V/��N��|T�hv�x֑7b\�ӷ<v��[Go�������9]WWl)X�����{�xd�XRK�5l��}ڂ*���7abm��2����6< �G�n�5ui�i��cI��"�^ l��I�fV i���Eӻ��x���Jzy���<f̬)%�����v�v��m� �c��'���I'~�jI<��u�'�U�����U���P_� �������W���(��DX�DX�`A`�DT *
�E��Q �`�DX0DX�`0DXc P�PUD������tW�^� *�U� ������P_�@@U�U�(
�� ��� �����e5���u :0Ř� �s2}p�<�@�.��v��*�  ݀5Au�����waJ4:   tm�b���7Y���lQ�v�SC|U 
 R�����P�	(R�5� PPV�J@ 	 P��F�h�  
.     ���l�hh@	$
��@ܝ)J;�)M��(�g@lΟ��F��O'��p�>��q�p>)��9<�;>� �� E��O'y�|4�Q�Y�>����� p��p+�%�]u�����gP'�6�м �ͭ(Q@ ���j^k^�r5{��`�A^7�_{����!���ݏC�z=���;��<���>�  y�����x�6��x��ް����=�>�KO ݀;a����@d�7��%���� �H)�k��^�g��j��g�`;���kx�l�u��]������Gl�{���À �oo����^{«����7�|09�3�=R��ws����篡��p`�� :�%#@4 ��GN�/ �jC���� ==�������`���[Ѣ����n�����9҅��� ��Ȗ��s�	��ǶM�����T�>>������D   �����4��V�	�wek-�����;�8�v��)J1��;ft 73�h-�Ӡ4�� t۹�O@oW�R���Jm���٠   :i4���� .�I�GOM7��4۸��zz��F�*̀ �·M)��̥ t��O@ ?I�6ԥ*  Ob�J�����  �d�*{iU(�  E?h��)U4��=�R�  "$#IH� )��T������?�?���۟�ZI%R�9��_��E\?耪*�(*�쀪*��TU�
��PES����?��Ѳ��?�M��}ּ�L�����'���g	!D�2[�;�g	L5��?�ߡ!���;�}(���Zr��L꿕8%T�t_3�N[�v���/����(��9UP�@��׼����)-#�l�������5��ӄHd��8��!-פ�����X�Pw�=g�/�7i<�ba%�.Fjn����Rd��2�����FC�=;��h�5�]p���	IK-
_3��\&]H��uOd���nR�%f��',������nj$OO,��
B��5��6���B4������X���i���L4H@�#.h�lp�:#�@n��s[8�L!��6%X0��__BO|!HB!.Cl�Z��\�\�R�"���p 1�"K�˚�yu�f�y����X�氂iϋ����Iz|�n�O�.�|��J�Ba5�e X�b��B]@�&@��}��tVII�xo'sDR��e���w< :�sOl�cqzhD����0��b�:Ժ���Nxi
��H�a��a��y�<��D�
�	4B��C�fA�!lJ��n�v���{�!���<�31�uEV^�F�uB��> �`h\96�2 �,;�0�R��q��NY��{��!uM灳C�fSE���RoP���RII�ݠc����!�pLї��%��a3\!�u��1�F�n�i�w/*q�y��5���C��uBZ�%0�#�á��fxVd�3�kN���%�ćn:�I|����.�������$<�۾k��</����ޟ3P��f<IsE�C�`���_ ;�+>��U�利w���_ ǅ����8���$%�t�)L��]{�<�=���:���K�|�\�"c�r�/cCr���ܥC�bh���y�l��k!9sS[�)HH����P�I���}y�Ȕ��98� �'<�	���}C~�#;��n2���<<<���9I5���5�-f����Y� �Z@�J@):�r�5�s���a|���|���y�9���$��H�
rT�[���y��.�szܘ�D�Np̈́��S�,�����:��'R��##1���7�����<�/!%e�	M��,�HRߓ�~��τo�=L2��,X`�u��L0�)u�k\}����ֵ���ܘ�]���V]%ܪ�w)S���N|��
¤K���1�H>>Y�o�s7�s4˚aL�7�*�$�'��ɼ��O7����G�!I� F���$`�3t�ht3�����5��l4r&ر HXb�1�B"A D�a��o��wܞ��l�J0�(\�Y��a<Ǟ<���k/��ׁ5����$Q�����&�T�0��F�		<��;9���^p�0��!���ɯOc��[�5
i�ӎ���<ْ�M��C�s���H�1 Hɛw�YtA&�=����M���w5n�8�p�5�\6�S��P��� -y��Cn��� �# ��%3Z��58@��#,B�1�H$,"a@+$l5�f��/q!	�;���y��$��xV:*��*��(��Tu*�O�~u�<&�OW��������R���ަfzl3��1њ�՛�e�!J��%p��b�k�<��\7Ēf��8�<���$���9���@V99��tdBᣇxw&F9�Ď�3f�挜�wԁH	���39��BX_f��Χ��Y}�q׾Be��[d��֯���$&����hҗ��f]�;�Ԓ@�HIHYF�$��t�F�a��B�����{�y�g�����0!fK'�a=2y`���,e}0���ߩ�%ى�$D;��0ü�l��\��k�0��i��7��5!06Luu�y�o�{ͽ8P(��%,���,�yL�����HW�5��#X�n0e��T�c/�~i�_�&�i5�
t��o�R"�$�S�N\��ծ&Gf|�ɥ���e��<�O8�U�3�J��Ghl���
��l.�s[�2*Snp䒘CN��BŐH�l����e���T�Ť��5�k����gK�!�a�k�!!x�q=��L9���|�|��#<����s�7͞g@Iu�漞�I��&k}ݾ�T�Y��0�0l������*��7t+g�K�\BA���iI���Ԥ �8���_Eqp�����}�_7�}�Y\��J�!��}W33�R������K��.g��\�6��@b¦C��#H�F�l�R���߮��β�C�� |Hę�a�� �M	�}y=��<l���,�ۿs=���l�0���@tz���F���d}&�ԛ��r�A
aM][�R:8�"`A��~}�h�	Iw��N����xl��F\�'C�XHy��.�]Ns�M:��ܧ�rv��;M�;��,!=�3�g���g�h M��=��^��{���C0� Bg/�������ĨI������=�35�Аk����)ۡ?�����a�_k�Sʡ}[��׭��m�h/���c�m>BX�#0�%<���;��0�+��5�����63y���͜���N���#���ٞsz�IK8s�qh{�����I�s�=�L;�B���*0�s&�R�y7�Md)�#糼��k��.�$��y�]j#��36��<��n�o��7�@��0b��o_g�4��<�Hp�^��7T�h��ۚ3.��{�$�}e%�<���ٯ4iӼF%Bx��B<����{����ְ�I�l�[������wV2�)�{�v����s�s�H$�JFL�ִCXC1!\�aaT��P��i��~�'���k|cpb��J�J�)�M�����ѳ��g\�I!ʥW�+�|�#:�^^�+R�|D!KuIJc��
�ĂPF-H�� !Y	Ie�k������t����4�HP��0`�L�}Ӛ$�2�°�
B��:euS+{�	�}!��4"1d�f��rH:�4�XD�cX�HD�w�����xlpcR1 Ą$"�0b�c��FCX�Y�(��j
B�)
F�X� �0�#a �|�<3�7˗�4H�sd�kd3W��=�ͲO�����֣!4�!aR#��jT��"�,�2Vc�a!f$!���A,1���!==������$D�8ݖ��B��p�����y�J`K��5y�K%�6aŅ`nva�\6r]�i��"B�X�Cwz)&�, c
�]$�؄�9�'!Ö�u/����Bx�6��F�r��B�$R)��"F6$
�@��D�)�ŀB �4��!4�F������I$d��k��%H���n�s��ot�L��̇-�#G�i�N�OF�=���_��f�fz�$���
e��<�w�)���A)$׷͹��dFa4�
CP�$H���(B�BYJj\$ �D�8R��8��Wyw�v������A��<M)�Wܐ#��<t�&s[������w��(��)��&s�}�8Ǔ~�ܹ��$��f�'�=����|Ϟ�pY������D�2���c&;��Ⱦ�_*̬��jy��l�����"I�q8r���\��9	(K�a��)���0� �m��FB�/0��a2���%
���V[�(\�y���&�?����Txy�m���Rs��[��Mk�:��%	t]�jM\��f����]��b�fߦ0� ҵ���mWy���v`��>K�S�'���˹��K��<�a���		wYa�W@��x���7˽u��!�����xI!	!������Ѩy5��O3i̏F2!��sZ&ah��B�u^M�$�		/e={�p��aph�ǫ.�0�f����W�~:Wo0��e�.!��K}�8�y�Ӱ���9��[�[�[u\�s��}��K�ݮ��5�xy��˭3�D'��y��������;���G=2g�.1"J$*B�j�fzʐ!�+�n<�6�=h͸��g��!.a�OK	����u��T>�T9R��Un\>�7�tw���}��2�ue-̅�i�,�dp�HF�Ѣ�3�9��l�'5�5�ynT�V4%	l�IH4�T�(^,���,'VIr4�eJ�F���%l�&�]{�$$B�^a.�!�w��<m٠�C!LŅWC.:I���6�����]i�,�ĳqf�SZ܁�K��݅a��$a	IB^�۩zS���]��J�R0�,��\��r/���!p�&�:���0ю�cM�J�@>�<�D����hF��)��`��A�0�c����&�	tKz'l�,H�a}e���kC���m�0o��$���XD�y AH�
`Ȓ�!hA�7u���Gu��XFRu>-�5���Z�0��:�y�7s�ˡ�2K��0,�f��<a���Ly����<������+�aćJt���欹F�p�8�C��A�B\H�=!�apjD�o�<�l!��2)a2@`R$#D����GF�37�N�!$;�k����{�<5�$@�1rYJ�#+!(2�"����&�������%RմQ)D�]Huvv�;��Bz��� P��&���'�_9���g�,Ӹ��:$RA�,X��z�}(��hSq&�xw��q�	BA.��S5ė7�Y��_}�|4\װ��Є��V�
�!L4Ja�L�Z��@�"2B�bF�L,��C�I��,��HZ��)a$�N�^�����uѐ�����$��}�׋de�L�S{#L�JbB�c)!��h�5˸i#B		�����oʯ��1�qR���RUPq�+~� ə�nFw�s��a��I)HZD����7�Op�<�h��� cB0��}��&S����72�vFI��O$�������M�C:�c߯p���ЖC����+UUUU�UR�UUUUUUuUUUUUUU@UUUUU++Uf�ﾪ�����UUUUUTUUUm�UUU,UUUUUT�������������YW���������U���������������*�����^Z���궫��j���V�U������n���w��b؍fɒ�u���j^� `�]��φ��B�E��k"bb�*+t�0��K�U�����Te\����J�I�R����G5J��3UR�NR:Z�v����6��iTw*����U&�%Y�J�UU>�Ի 4�+�j�����t��9Uv�D����@�H���jsx�u�n�+s�xлsU*�}���P�h�+�ŵ�2��eUUK�2�@B+�Y��[p%l��k�<��R�R���T��M��`T3eª�z\��963�ۨv�8x��VݗfWj���⛠��C0v�1UUe�F�ܱA²��UU�U�U,TUJj�w����5����� JU��BR����6����p�/G4��Gs����ayu���м�[�vTM�k��O=V��'j������՘�
��Q��
V[+f8�N��7��]����R��s�m[� �]�[�-+m�$ D+jt�R��:=U^S��ևe�tW0�ٴ͞V��ڝ�_�}��UUU� ��Ò�6
����ܨ]]\�U�TJKT�j��>��x�ʪKUB8J|���UUJ�]�f9X���A[j�ҭ �V�UUHC�ڪ��q�`�@u�����UZ(j�` ۳�75㡖����(�Wf���@Rղ��j�;X*WLU���ڇ-laK�Ĭr�b�V��M��Z��U]��h%9��J�����W4�R�A��T���jX*U�T�+�[Us8��[��T A���sR������mS�=@K˰rF����kfjV��6��j�$Tu=[���V 6)w<�G(,���k�ڇ5�8����u��l�s�Mv%��
�]]GU���T�p[�V���a@j�VS)�21�j�A��1�y���<-F�I�6�뀹Z=��y�o��!�Q�)i�-��lS��4lѪ�軶[7n�R]Sۊ�{9�}գ��9��CuY#�(����,-�q�Gm�Ƀ@�i��=����5Ep�
�j��b�kl����9�ۜ*���ޠ�xc����+����ƶ9Z�n�
�*�֨�lݗ�unԤ��ZR�Gh�XR�X�IKv��[�������+vB*�S.%3Uf�ʰeDE!E��UUUb�KUWA>�şX啇�89NG��;���wj�K��eqΞ��ͤ
���ۜ�yf�L��f�˪];)2����b�E�5�7�	;��vh���lfż���L��Jz�}
%� Y�Pr,]ښ�&I���Y��0kj��>�@(���Z ����o�ӱr�f�ldFYvIx��D��m�SA�tCrͶ�=������q�*�ܭ��7;�R�sUUUmP#lc���ЅV��^*�͕W�*�j��3�%�<�j�v�kk`݋���j�wm�:H:� ��U�D谑���B�r���*��iUUH�u�`�<ҶR���1.�+���6(A�2�a7a�+]����ߕ�ݷi���P'��r�B�խ��A4�#�79��S����7&�n�Vݵ[J��.^6��^YV�s[���8����������[���W�����:Z���@օ���r�y� B�q��r� �x'p�ZG|�}��ʮ�+/��Ut؊3G#X�6����mnwuc]-K�cUU�������[N���g6�������#@{��"�U[[W]C.��r
���R%�
�cI@R�U��*�); �d:d6�m��x3R��K�����Jݩ� ��Wt��)g��8+���\�
k���I���n�ͫE6��e%�]���څ����i����K[%v]u���v��Bj��y�[Mm�UU�WT<��[s���Sl���y�����r��J�PI�'����6�];xz�����RY��/<��n��!u*�TUU�)�CT��M�Bʺ�������İ�V�P�[�N�N�K�{T�� �u�Aut N���+�[pUUmU9�zN���������[�����#�j�(�dz��c�n;B����A
z�WT��l�ƥ���]C
��P����
Ꮋ�:�*����¸�j9ݹ�r��+s8m�7�-�rմ%�N�6��M�n]�7�c͞7,��f�
8�nx��֫7`۲�AД�]b
���fLm�S�.P����6PV*����J��`�L�٘q�gI���v����(�iUIaXdnY J
��p �v����$��ȫ��]�#��,��� �G )��;0qT�[t�8��������x���UZ4�նzt�v!���a�DwF�-89�댁�n��+K���l�^��������w,�W*���u�UU:� �6z�l�f�Z��EUU[K�-:6۠�ݪ�Z��UMX����@/YN��U�����f3�u�;:2ĉ5�{m=�t:֒5K+�b���R��I�vKi6D2qA�� �BF�`�`�Ӟ��D8W�7k�umR��2���9J�:�\�h��	���m���'��`)��Mq��uQH5#- R�U�UA���q6��Q[+B��Ebi�����C#Ui[����R�=.0�Y�Z�
NwU�U@UmN'P�`�6շWWV�pA�H<����UUU��J��d�U�򴤻T�i{-U�U�
��+e���pe��/C������lUU6^Z������[�j����收�ۈ
���
wf���Fv���^Z�V��3�16j�G5uWUUUUU����vb�l��m@b� �+�lR�r���˻���ZKj�:Uꪮ�y�j���Xyf��S]@[mmUUT���U��Y���y�P�m����k��*�vV���3VZ۪���U����7��UAKa�V�5��Jʀ�UR�UJ�UUuUJ�]A�
�Y�����WT�Ä��[UӖ� ��U_����Uj����
����ڪ���Z���V���H�j+N���Dx7n�/�UU�Q�����=��=ۮ%��kv�Wm�'5P�9��������F��-gAUUV����
ꪪm�[P*��������3U����+�h�ir�u��ꪂ���CB���.��ʺ6�5UUU\�+����٪���ڮXv���j�����������j�
�+j�����M*�c�k������k+eX퍠;j��XA����j���V�ݪ������j����4v���PUUUV*����P��m��[PUPԫA��QvVW�c!-@T�����궭��S����*�UF5�� ��Ptʪ
���٢�UUX��]�UUPUe�����UUT�N���ʽ�ʴ�v^�"n�`����Q��/6���i�P
KUJ�T�U�F���������UUZ��U�UUUR����U*�Ί���V���YNU���C̬U�
���������h
�*�U���'����U�����ZU�j�V�V���4�Z���4�I��u[�d�N��<�\ JH��n�3@�j�b�U��mV��P ʮR�9�)vY]�ڭ��^�j��ـ������^Y	 :e��n�*����ݴL�Udz��U9J�s���Q�hΎ�1�&Uƨ��G�Rڱ�40���aW���j/W:����vQ�v�$�k�Jpʡ�TAX�m���m+�X�@V���o9٨z�R��v�"���������v��O;�����$%6���ke&�0�C�(�<��"����vP��vCDp���O[lF���ڵͶ�(n��@��ۣ<I���/������vR��r�n�Ĝ&TBFGqձ,��l���0s�u��xܘ�-mJ�+�p��Dҽ����pƳ�X�(�D2TaQ��m,����vZ����/Z� �DJ�,�x.j8�<9���N���M'X3v'��`�y�q��C�8v��ݘ�.1�Uꫫv�Sa�φ�+�1�V��e�`*2�fS��cv�P�dr�P���l۩��9���kԯ����r[�WM�Vd]U��Q4�P8k�����$Ʈ�
۝R��R�/n�����ۑ���V�����7vZ�m��n݋B�UM����X*5���T��AS�5]U���%g��dn�]"�'D�[�j���P���%��������߻�S��~ ��ؓp�nR��Tڄ������ڪ]����md���y�`�r�us�	v@���U�UUX��pi�-�UvV.v�UUU+�Q\/T��U)�L�yJD�U�V�ت�+n��������j����~���V�j���V����������PYU�Z������*�V�`��R�a�UUUmTUUUU@*�+,�U]UUU�Ys�W+�Un1J�WUQ����HRҭ@[TT@UUUUUU�UUUTU.�UUUmJ�mUUUUUP@KUu[�Q��UWf����ڕoUUWUUU@R��ˌ2��UuUUAKU@uT�s���-j�  ���宻�j��m���mU�M�/P�7�YW,��U���6�Ejj)��ZU�cWU*�UMS:*�m�eZݠ�*����V�Z��i�kj��:����fQ������Vr�����]s������a�r5�e�v��[�X�WIVx�nrY��x�B":�Ɔy�B�9��r����}(T[���n�������,2k��g�S���'w'� ��
!��Q��A��J?�]��RE�d��H2X���D	��M n(b�8&�"���!��n�W�� ��x ���h�.
�Ah��!��>��QM�tD7�' �S��U �U�"���h��Q"��X	�����z:4�����E��>�`����*���H$P��"!$H�/��B &�ΆЌ������Eu��!��1���� � H�J��= �j9�Q	�Q��#����q$E0pڜP@�`��}��P�6U���)��;Tب`M*
;��	R�`n1���2&�S�P��C�`��BiUU=�_ ��0���$��+�M(�@��v(�xt�_Ύ�����I"J���:����F1,-��"�*D�
��D(@�m����Qv4F��4.�}z�*i���-!F��B�%��ZV�D�RB���FE�k%�ZR%-�i@
F,�J0Jư�B��B�,�	T"�P�R B YX�B����x������. =6�4�H���@� +� B���`:�(�D�!���z8�W�ڧ�PE^�1"��$`�!�(PGHZ��ԩS ���D
PJ�hԁ+��U���	�BF�D�wY$������ʂ��P��UJXhUUUb(6�eUUPX�B�fج&eU��y%u����&x��;�΍��p�U&�VUJ���g�v7$�q
(���@��f���d8��b�X��zlk�VC����,
Ͷ���d"]i��VF��F�*���p]�g�yy����x��ś<Cvfu���;�R����h^�z�-N�\��&�e�e �o\lF$�V6a� �K+`���saM�56��Z*嶺j���#������Q�,� c]@ά]#m֘�:T�Q�t���.�Wf0v�v�@ �V`�RWRk*F(p�f���-�T����1K�X11�kv�{$m!��*6\��`:�n��[Y��.��Ã\� f�s��z^qmb$s)v�����ݧEv�*�S�E�+]�ǋ:�� .gtsВ+��{:���TSL���DPb���W\qŬ�w���n�Bf�v�ɬs�9У���1��w7 �/qnW�.յ�t�"�k�d{n[�\���������4Cm�9��7��u
 vυ��T(�n2�p��k��r�U��Mm��\�#s�63���mq��r- %f(�����uP�Y��k��I��)#JA��C Vv]ts�lh���9h�a��x��QT�f`����h�i�\[s7;�� �"br`ʰ].�b��s��M�i�s�4P��+���y�/bs4�++s�\�UfH�4�c��%N����b�NJ鱷Y�X�<J�#��<H�!#ŗ�!����ࣛ-)SFm�+�LL�ۉh���|�R�|!�f�=�p�m�����'hR3�,)��m��m3@�r��phM�LK��QҀċ�A���l�`�Җ�k�WkD�2��ګ�t��;�ɱ�OJYx��r�J�Z�����o�b��Ш<U�:�X*��� �VD�h���Zq��qe�փ�AT���5(�;Q���{;4�/\Nx�m�ov�b.��H��� p �AU���*�z�A� ��}8"h@�5 � ��7��D\v�h��ȅ�nzg;��k5J#3HW[v�CS��5i��b�R�č(�y���,�-��>�Lu��D��MJ.����� �	�P�n��B�\G3��T۝͞9�!F66�u��ĨC�ݨ�;��,yEn5�!���ڢ����%w5�o�s]�M�N�t��\F8�#n\[ 6��V�3V/�� *�Q8 ]�o̅��d2[iHalT�Ԗ%
���0�m��%�S�Ѣ�/�����������$D߾{��A$��Iؖ%�b{��ӑ,K��@�~�|�ҋS-f��ҝ)ҝ9�wٴ� ��,K�;�i7ı,O|���r%�bX������K�S����k��˚[���:z:S�8�,�֓q,K���{ͧ"X��B"w��ى��%�by����r%:S�:_�%�IT�k��U���ı,O|���r%�bX������Kı9�{۴�K��dL��z�nt�Jt�K��ϴ�-XhS4��OGKı=��ى��%�bs;�siȖ%�bY�{�&�X�%����ND�,K�	��2ɟL�t��1x���؇T:9�� �ksp
�VX�ai�KB\��K��HQ�G��нн?�߿fӑ,Kĳ��ZMı,K�=�6��bX�'{{�17ı,O3��fdѣ	�j\-ֳiȖ%�bY�{�&��������@}Q�"y��~�ӑ,K����l��Kı9�����Kı,|�;���R������N��N�=���y��Kı=��ى��%�bs;�siȖ%�bY�{�&�X�%����;#nvW]��Ξ���N�����|����#�2%��}߳iȖ%�bY��kI��%���ȝ��xm9ı)�����/�](��2�n�)ҝ,Ng}�m9ı,K�{�D�Kı=����r%�bX���vT�K���ӿ������51�A�`�u���[5�AX]��/\c�Ǆ�l�7MpT��2��w��Δ�N��~~��O�%�b{���Kı=��6T�Kı9�����Kı=���k5a�W7l�O��N����Ͼ��=X�%��ɲ��X�%���ͧ"X�%�|�u����eL�b_=��h�́����Ξ���N�����6T�Kı/|���r%��	� RـH
$["_;�j&�X�%��{�ND�,K��鄖h����㙓EMı,K��{��"X�%�|�u���bX�'|��6��bX�'��&ʛ�bX�'��ץ�Bi�J�U󧣥:S�:_~���bX�'}��6��bX�'��&ʛ�bX�%��bX�����L�������댶w^�h� �W�[���Sc�Փ��͡�ow�,K����ӑ,K�����Sq,KĽ��ӑ,Kľ{�j'�Jt�Jt���P�ur�v��g�9ı,O=�6T�>Q9"X��~�[ND�,K�ߵ���bX�'}��6��bX�'���ɼ�p�5�u,��EMı,K���[ND�,K���Q7��R"}���iȖ%�bw��eMı,K���5k�4k%ї.\�kiȖ%�b_;�j&�X�%��{�ND�,K�oM�7İ:�M)�#D7}�y��"X�t�O�#>��76�n�N�(�%��{�ND�,K�{�eMı,K���[ND�,K���Q7ı,O�=�xK�>2CF�L$֦���v⃴�a����Q�XZ��IJB`d-�L4^�4Vz���N��N�~�ǒ��X�%�}�{��"X�%�|�u� ��2%�bw���Kı>��c-n�0����^��^/��u��Kı/��q,K�����"X�%��{�eM��L��)��R����]&&��yU��c�6I����O{�+ '���W
�b�wcI]�oܮqI�}X����I }$x�\�ƕ�vڷt�&� �"��	6< �H�	6e`\�N�,<�����!>�!
"��9�c�璸s���e�ݺ�m�]l��YKP���P�FXum��!�D����^;n�۬u�l� ͕�U�їq��n�c/�x�m�&�q�1سĻ�:,�7���O�W��᱆cicQ�x�֬�c6k
�uq�pZ�,%���j4x�'\�[���鍸3�0�v�y!Ku�k���tmIB&Ms1i�_���'�k�&򋢆J�P*�IR�%t��s�&8
���c�^1��\�WZ��uaG��J��N���< �H�	�2��,���1��t�؝����x���U$N���'dYX;���ăn�!n���m�wm��2��,� ����#��"���Eҫhm��U)�y}X�x���ve`���Ɔ4�_i� N�x���	ݙXd�+ �UUs���}@��=��	�;�Y�ej�\�m��P�]c���qk���fni.�����b�ͱ��<wfV�"��UW�l����i]�ƒ��o �ٕ��z��
Ր��0bR2V�����a Z�`+���(�g~�l܁��< �H��\���?S���ڶ�RM��{ו�� }$x�̬��<��c(N@���%ꪪ�f��}�<w\0	$���ݘ�)�6[�V�]�� }$x�`��_�i%��N$�_ki&�ZS��$�:�@��&\rY�v�K�GGFJS�Ѐ{2�[�lv�[m]�x�`IyX;���G�t����N����V�I/+ 'v< �H�	�p�5ul��%WAwn�nǀI��B�.�5���ٹ'}�sf�ީPV��v��o >�<vL�I/+ &�x�up�CWm�M]��Nɕ�l�e`ݏ >�< �NH�%M:(?]�!e��(.�Vq(�L�K�H
WlT� E7��	���*���=x����2�nǀI;&V�ᬨ;J�c�T�� M���#�'d��7d2��$v�����mݗj�ݶ���� N���� �#��(B݅�v�mڻ��l� �{ٳrI�{�nM�� hy�O�����$��nӟ�m���K�!��z�K���=��	�<{�Ǟ�����@�v']��9�N�X;a.�0C ����s�b������� 'v<�^ N�xvC+ ��+�n�$>	�V���/ 'dx�V M����
�����!ݻ�	��!��v<�$��9O����I��˶��� ���)%�� ���T�|�ݪ�� &�x�]�{����x�E�� �"ELkT��T�Q�ā 2
H!��t�^��}���i(�2מyu�Kty�B� U�y|ku��E//c�]E������ИɃnP�]���ul��v�]��z9��y�L̅N:_ݫl�0h����Z�;=n!�[m���B��L%��؅�(�4`6���S)m֖R�V�C?�K���aFN�����/uω�=O�Q`�ey��Y��*�n&��:6���܇v��O�����-�	u͑�wn���x]M��c�n�^۰�',=Z�Z��ށ��K�	� l�< ���[���v[���wwv� 'dx�D�wc�>RK����>m+*ݫV� l�< ������wc�5wn'��C.+�h���e����	�yUIJ��)
WN�`��&+�xSe��ǀ�� ��/ ��Qr躻����V `v�]5�6.��3Q����$�*��-���
a�ۦZC�w�v< �$x]���Uϐw��,W��]�v%n�6�(���~��S���x�&aC�0P������瓗_y��y�H������S���;�E]&������6^ wkc�>��%��l�wv�v��܋ �/ ;���ۑ`.�(S��uce�v�uM����ǀonE�}�"�5m�>�����-�v��-��:��G���B���ڜ<��%�kC��p�ڏ �܋ ��"�:���:�F>	Z�q]1�o ��ŀ}ۑ`nk�^��3kӗU@�x��7ħ�*L������ �M���f��b�ɸs��9����;.�L	�f\fe%�FXR\}:f�iK����MbG#ŉ
#��9����K�a�eIYX�B�'p�b�4©�1,e1�BZ�B�FVY������i�����l�C6n��[Ip%�#�h�)Ӽ�5˩yq�<a�)M^e�p<,����_N�9�o �//�l����.��o�e$Ĕ��	[T#�(8�
B��R>�i
�=���<��Bj����A�1���
� �V�P�R���m�4SB��ݗ �{��R�keEѡ��[����琞���|�N��b���r�`ҕ���a.%��;H9���-��;����NtΜ8q��`LH��A㸘�^�d�F����RRRYYg������hp�]zK��L�6�k+b�=�ZB�pV	H)IMF�1`�)
�eR�`�!RPH1b)H�$�3[�F4�IHP%e	HP�YF�2goCa�f�_Jo[#`�R5�`Д@��P�h��ĕ�x��	K����i���D����͙<����sz�sYvf�s=I�g��`�nN�Y�%����|�nH`��B>��Ȥ,��<�E<9�y
�i�|�
�����x�Ǆ�K�qb��זj�����f��z�|ߔ�� �M�@:8@t:D<j+�b�KT�PH@X>���Q1B%Q�C��vx�T�4!O�� ��}9��<��������A�����d>�d���j�֮ܺ�A��@�A�>�ٱ�A�A�A�A����lA�lll{��؃� � �(~ �}��~�y�Y�qgI��߼���n[G��y�O���A������b �`�`�`��u߮�A�[|�w�ܗ߾�����e�9G6�A�f�;K���a	uc�6�5������Ӽ�o'�MwQ�TU���<�~�x��j�_��+�I?������ym��~�?��Y�A��ឮU$E�z�|{� �܋=�P,=�<��')��N8�����ėTR<=\�[#�zy��vEi�YI�+�x�r��ߗ�����&�ٹ4~�FAka���"(�2-�D=P�/�<�}���yO�i�$7`���i��wu� �~�9���9_�}������[�l�G�H�ɗ��lm���%un�w
8Lh\@pM/B�ޝݯ��5��KBV5��	�?�������������O7i��%i� ղ^z�#W����?��Y��_�͟�����.��ݦ� �9����o��`we�d� �j��qU����Eݷ��l�x�<���vG��/����Vʿ61�Swv�V�-�x�UU-����/� �� ��r���Kj	��ն��jˠ�r��m��g�#4�����������ss$ {@�Y���$�ۚ�a��8)f�te��.:��V6q�	`��?��6>��nۖ��ۏ&:F.]�zM��2͠m�hK�Au�:&=AE���g3�q`�h�Wr�6�R�c�c&XD׬��<�P�ėPMЀ^�pf�6pk����v�c�[3���/���%��y�ǶY�q�@Ŵ�R��ۮ˘G]���i��U���'�����ۆ�u#�٧���z~x����U|��O^ C���YM��v��x��{�I�~0K�X�����RGT��uJۻ�W�t��o ���M����UU�=�� =����>QE[whS�lV�UUqz����"{ߞ {����\�����OZ���I;n��������O�������"ݗ�J��J�cm�$s�v5���{h×j4q���-�؃�B�������t�\jl٫M��������0�e��@l�xv��W�Ywj�CWkrO|�6� |J�R+r��c�	�G���UW�U]�����[�6�n��+f�O~� ����W���ω-�O.$��kg�����6��ʤ��� =����p��9ʥ���Ǽz���5e'j����=U\������ �����s������k?.6��.y��J��8�JV0ŁR.l-��hRДߺN�w��d�y]&������ �ٕ���ʪ��K��?r�o�=��Ӳ�T�n��|�{+?Us��y��/<{3ܤ��4	�T�1��'v� 7�� ;أ�Mb�֔ABaV0E�9��@"��S�v��ϵ�ܓ�{�+�+��[JI�)�&��^�1�_�7��;&V����y�*��x����*���7�� �r��{�W���uIq����שk�IݵV,�E�$Y����Wt�dЎ-���N��:�-����;[�V61��@����߲��c����s� ��� �W�-��[�t۫v� ;6<�\�\�������=??��L��Ur� ���𱃵Iڻm�{�/ ��=��U%==����j�6�'n�Ut��v���UR�����lܒy�{���h��P��%J>�*i!��0��3D��T��
1A�q2"��:�'>��|�7$�������-�ݳ ٳ+ ;6<T���f�$�W�wV�+�G�� )�����峞ѻY����K.ę7��e-:��Nc�:wM�I	��d��5I�>��lٕ�}�w nݤ�mU�Wm�e�,�s���`��V ody�s�|�;��i[hT[ٮ�2��s�H��<z煀o�[�X鍵v�V��{���o����X��\�ӣ���?_-�OOg���U�ʹM����G�~�~�{�{�����6I���ԝ�H!����n�b�lQ��M�x�75V����'n��I���'X�<����ܓN��+��!�T�m٥K���H�ܪ��I7\Tٚ�5,�f��*�ۛJn���ܽ7!����P�m�ˑۮȸ"*��a��Kv�XZiW68ݞ�]lM���#�f��*D�vZ�]F����z�1�d�#J-��m�FK�mNJ���]:{�
i�5�n��*�n#f�T�4E)���2B(�-��e�P��!l*_�*y<�l�j���M����^&�`�ez����O<V�6�'n�V%W�헀I������U��~����{��:����[;}��a	����ִnI���� ݑ��W9�K}s��7��V v�K��kfu��O-��I?wt��~�ZO����;$���Ur��JO{��=�w�"��&�ʾ������N�$�����O{+ 7dx�:�؆ۧJ�hK4�uɯ4���5c�MNLw9irp�mnwkWE�N�::O/������r_@|�����nɕ�$~�UU|�}s��'�+�e;����i[�vL���h*�W(�X>�%��`@%�VH$daF$����	iVD$���|�{�s�u�'~��.�$��UW8�Iϖۤ�4�ۢ۬ ����6��UIO{�X��V H�j��2�i;o��%��=�e`�e`z��J{�x�����Awv�����e`�T������������P��@ `��n�c�<�Y��1���kn�B�m�bƌ��b\�~��u]�T�ڻm��~�W�����������ܮs���V V�ү/;��m*5n�d�?U~�9Wd_���߿~��7veg�UI�;�ݡ�e]�v���}��]�=�{�s?EdI)@��0X"� �1�L���� 24 "�� �A�Q"�a*'�w�/����e`�x�VV�(-�V�VŁ�r����� �{+ 6H�=��8��<,R�/Y�c�n�i�n�ݙX�U\�~���;��L� ��(6����kL�]���3�A��U9��Վ-�=�軝�XbYls?I$�;���n�cn��|^�� �^�`$��r�\���X<��V�-P�;�x�����>�����>�߶nI��{��C�I�'�k�n�����ݱ`��V{�ٹ�QO�(f}~��7$����f��=ɇfc9��Zѹ>AP���pܓ��}��r�����B�����1r���k5�&GC���b��0��ͳI�����$
M�5
$:���U��~�ܒ���s�)�cE	Rv� ղ^��U���s��~�_@��~��7�2��7�&��ab�
̢��%i+	���٘���ȉh6����coQ�Lְ.ߺN�O+3)��i���v�j���x��j���s��W�<�=xv�)�j���@;e�l��s��9�_�^S߯ ����`)!y�����F��%�=i0��`zz�	/b���s��Q{�/ ����wB;)�V��t�Ҷ�	�S��~��f�_߿Lܓ���7'�'O��'s�����o��ț����46�rOo}雒~U?
���߼<�}}�7$����0��Mk1	L�r֖-	���@{�� ��0�tu�NytoC�M
s�.l��߁�E�G\�xE4l����7�b�f� ��8B!�$g7��Sl�B>{��A�1�hw�wOD�)�j����8Y����%IRQ\)��J��[aP42�MH&��k�o��id���R-H����MV��9�<ֳZ�*��Z9T�v�UUhe���ݪ�v�d�U׊^�]#P�je��L���۪q�!� 6]����nvg^��0n2E�!0w3v���;X�n�ss�9.��s����E�����?87��=s�I�AQ�V��݄�eJ˹y�e���t�:��/S������Ha�1(52Fmİ���A�f��Kډ����K,�Yn%�9��*F�V1��-�(�,�F�2ʦR�[@B�NZ�l���Bk��d�%	pc�q:\���u�(ͫ	A֓v�^o����u`��I�3�6 �����*F��&
����8��v�::�u��e�m;�)e�R�mm�Gv�8�sA��AգN}��N�q(볍�^�f��f�{-(��@�ٌ����݃C���
�/;�!B�Î�����A����+F$��)(G�L�1�(�hL]G.�Ԓ�]�8����n�V]Ԇ:�h٬[K��!�[u�3I�@�j���SS[��$dl��XF��ݦ���u��Mǫ�;�w�=��prd���st� 6܅�W]6�h':q�]a8p��Y޹�cj�UM���i
�v�+Qt3Plj��I=�H��$�О�@���[�®�õ��_|
����/k��ڹ�jk'E�^"nؖ��p�N��(�'.�j�Sq���-�2��,�n�lYK��(ш�����]���5�}[�C�v�_n�hx����˹�"%�.35��'պ=M��'8+P�j���.�>퓭��5GF�=�6�ĽWdR�n����$��o0X��zzc�Z�-��<!���A�<;m�M)s�5�z�8
E,��ϯV�Wna���<��r	Bq����\�[���pDb��n�1��Q�B �0�D��W�um-�V��.�:��6�<�|�̒�I�U��BV�����a���)�5uJ�Ev��[
���a �ܻ��Bg.�ժ���Z��)H9����A3Eڦj�*��I>� ��)���׉�W�R���A":��8/�!��O<���2k�wZ)6h�:tu$�E�ժ���s6xv���l��3ӎ��V���x��EK�.6�k���;�776N�gdP��]��c���42�5t���B�["���9n�눌5��	���:���EƊӹ�@v�j�G�Q�w֫d�r&�I�YUL�������I���ؙ!��l�����=��l-U����l`�:4Rkr�=N�?��$�'�I�q$�.]�S�@9�]rg�r�`O���Kp6v���1fk�����<|�x�R�q������e`���"�/��r�����=r��¾uO����5M���W��+�v~_����~��&�g�\�$��"�_6��ջ�<�=xT��9ʤ���`^�� ���ud�+�n�[�m��������� ���E6^��\���z�	,�������B��Mp�=\�Us����/O^��� z���S#.�ٶ��Vt�pѶ�q��8M-RlƲ[��<֬�Ӥ�\��Z���ݥm���� �l��r�UT���'��������J������;|�s{U`#��=�-�>*4��PXE���Ti"4R,� R!00�_�9��3�����x�����RG���V�!X�L��-���ݏW)(��^�?x�K(��C�JPM�:���^��%�<��=x�p��W��+�7�*�]�XS
��v��l�����<|S�W�v<�ϻ�.���<F.��iq&���TM���HT�4�iT�[��v׫��Q����lo�4����XRB�n����=�Xv�XX�i�؛��E�XRB��T�n�� ���Xf̬�9I�qz��Bc�@^jf䓾���$�s���=��`�|�Ͼ����<���v�,%��v+V]����_�������,~��)����Ӥ���� �~��es�tk���n�`NW9.l/���Ir,�l	�m~ą�MT���4U�ǔ��nQ� �cW&�]-�4`k���9|��Mt\��;g�yzx�{r,K�z�_ ���z���5�0�JՊ��^�܋=T��_���~0�����*�]XXS��[X�~��;5�R^^�/ �~��
�	j_-�V*hk�*������䟯�Lܓ��{��? A �X���f@�(� z��_�~��;w$��d���Y��,�j�{"x��s�_�9���~�ߖٳ������֋2Siv
f��ssU��������-pc,�jӴ��I��T����<��e�)�(���@�^��X{&W�_ &����tz˯X�!�ۺ��xˑg�#w���	��xWd��$��[nڻݖ]��n��X��oq-[�^=~��:�"��]�lwE��u��R]���V�׀l��Kw�� �/{ʹ����v��]��UT����n����Kx�.�M.������5uL)��f�nKs��k�r�ً��A�;D^�,h��\G;�+bX��i�D��(�_ax�������51�#5��,&�&NE�lu�oY��X�B�F9ۄK2��v%(�k\�(����/!@��Im�"F3��83��KRFӊ�oe��W�pcd0�m�ҕbk�o49��]n����͎9+�[�X��3ar-��Sk�D������1cԈxc3 ��DRhj*���e3jMD�б��Y��u��X����!<,�7�m2�߀�럖�� �ȝ�=�r��վ����֘վZ�`�X{0{"xWd�eȳܪ�Ge_�,T�諶�	5l�	��x��x{��))������6��YR����(����UUJ^�׀O_���p��'wu�~~�_ ��~��ƌs�����X󜪪�UU�r~�ߎ�{�� ӻ��+��X�:J)#:�>o���]u�,�Nf�oIa�Х�تj�c`��wwNg�cE�Jӷm�e�_��� l�<Wd�UUs������ վ�E�I�hְ��f����ٛ؎��;P<#��N���nI��~��y�uٿȿ��:r�����Jn�qW���O��>��Xz��\�%���E�z� ڛEvS$7�Hf��f�r~b~ �߹�� ��ߖ�IW�ꪪ�R�޼ �4��.��[m`Se���x��xˑ`ݥ,�cm����Ҥ*��R[�i�\6��J!��T���mq�;@���t�%ٚkK�	���ew�>~�����Ȱ�"�r����=x����z����]�-�������I߻��o��ߌ~�ߖ�܎���r�7n����Ӷ��ۺWm`��,��X]W�+�
BBY���� � H��El�p!������x�~��
�Ce:mէhm�˶�=��R�{<`��;�7nE��UW����g��ui�i�'Wm��܎��Ur�ʪ��.��y`�e`�5~���Ov�R��͙�[�C��h��sN@��6���ķ&6�	Y�t�t[-x`S����,eȰ�2�s��|�������+��Q�[��Ir,�9�RF����:��7�n܋?r�ʪ�U\��J!�~e�`��C���	����$oUr����� ���X{f�i�$[wBvպ��r�K�~����Ir,!!'>y��o���G�:��.���ݷx�� ��X�e`K�����jR2ו%M;�������r�.�WJں�2�ͻ3����f)h�s����<�>]Z�[�n�[:�����$��ԗꪮ|����h��M��v�*���	$��W*����V%�� �{���wI��N��>�?�5˕�Հo����r,=U��^�<���V��K�j�t��,V�ܪ�[��K�XvL��I��v������Tq��m`��`�Ul�����=��<�;۹"���P� ��l�.�\v�cIT�:�Ӡ����l<��ʥ��u�x��-��hv�2�#�TN�=��k	SBY�w%�K��V���^�*��GP뱬��m����(6�n��7m�J��,,��Aɵ�F�Kt�Z{��%ɲR1�j�}�%=@�Z�.:$��p��{���`ݗ�ˡ�w��ti���.+��E�Ls֎ѱ��V��+�j��gFy.�Ц����]��9Rعk�k4>�MQ-.�.�e���W+t���X˴�[n��V�Z���X���;�"�r�A=s� �~Ai�E�k�v;u�}��Y��6_���ϐO���g��W=T��o�0�����J�JK���{�������;{+ �K��)�r��ۡ�q/U}Fz{�Y�{+ �e`~�W�s�~�~��ҏ߇M�n��+.��;$��=ʪ�=��$�y`��`��=X���T'ip�oa�ݒ6�i�؎�Άكw�-�hu�5k��7e�]�%n����X�Ȱ��~�s� �{�X�I릕'`:B.e��rO}�����*���R1�a B
4 �#4�3BA��"�QK��R\1L����ӨH@D��b�E��		$b@�.�Aa�H��$B1a��H�$D�R!�$����Y��}���rw�ߧ�. �m�߫ꯛa^�*^O�cJ�qG�}7��[�u�ٻ"�Mf�����|���~��ݠK�di�c�$.��yG E�uv cݏ�z�����s|]�{\a�rE��q� �m���爵�z; 7�|]�c��\ �E>}�����lYcol8�ԗ����hG�$���.�nJ;[��/�����1�k�R˂J�@~�| 3fiv�7�~��}��v@3ߏ�W`����LjD�6�ۉ� ͙��<�5��n�]�t���~�N��;���O~����i�˝A��v���k��ݺ�9�j��\T���.X;3!$H���)�a�V���8h0��P0ДU㍰�E+�L�FK��3��8Bk+Cd^;u��st�
��8h�2,�˱<ٞR�M̲+�r�w�j�����6�\$�XD\ 2^I�7��]+�}с������5GQ��6c�,F!�Ha tA6`���@#��F�!<yWi����=�36&�U8��!8l�&�N5��t��� UX��C�]EI	y<0M$�w�B�$P�iE9���	$1#MƑ�R9I'������RL2��31	���m�4FH��,@�`9��D �	Ŝ[BB�"Hˀz����iH�G� .�$�"�b�;ǀM# ��:�Q0n��Hk��3*'BU<�QO@E(� =X���D� =B��J� ��8���-@}%}�UUVM��i� �Ox� �1m�#JFG��� ��W��W�ڻ ���� �������3J�!��I	�hr��0٩� ��V{�� ��q�ꯩ��^���~߽�*EX�q՝��u0)�X����ƍVu�����4̶b\�I���]�<��D*��o�+���~;�~�g Żu꯫�Uf@�O�p 2��#�R���$�$.�1�� �v��f�S�vf�~m�6RL�F��/��nFp �z��nMS����UI7�������� ʩ�I�Ԅ�CD�v�������~�~���=�r����A�!�d��B	,,1@�� B&�系��-��fޭ�L��A���S�vf�`��7�e���]]�.��8 U~[���N��M�M�k�Β)�r�5R
��������1ԧ,&,�9�ʸ�s�I*A�8�p� ���� �v��wf���=7��ѫ��GDppt9��n�]�.��8 wfiv �w���a�M��GI*7*�k����f�g��m��r� ��]]�*�I-�� �E"' ��S}�7����O��ͺ� X�I� �n���mI�L�� �f����uo�]����;�{y�m��`�Q��i���kG!�2�m�݄�����1e�&�;yç�'���|ky�k,^պ���9jA`�`e�C��W͐��l"6!ZE�Gh�Zř�%]kL1!5ֹ�%T5�D�#M���:5�SG�����u�cJ�d�'+��:�uXc�QXeWlX��Um�]�c�\@Z����S�z�$�G=�˞W\t\��WFa�ve�̙3�:�j���;�|�3���iPR��g��<��cJF�/gG�p�rlGCOey�v]˧/IL�cp�$��� ?mo�]]�c{�� ���؃�� ʩ��n����Su�����a�M�v������۫��3�T�9m��> �4� �f���_U6�+}uv���� ��[�I*A�8�p� �sQ���۫�ou�������u׎N:D%*D��;Y�W`���� w�|]�fɡ��������� ���AN%�R������S1�u�����ى��c0b��7Mʻ Ff���f�`�4=_}m��[뫰��J���\*�M]k5�m����i���(���B��$*��E�$��"E=O�|�k\�v�~�߸s�fk� ���
djH'"c��vM ��uvg����"o�����v�ԒkcCnO�H���;���\����I!I�x�K���INUUU�s� 7"�|�n�"���J� X�I��7K�� ;�v�������x�i�#F�[Ë0�Z�omp��v��ͩv4>]$f������^υ1���!: o���� ��[�W`<�� gin���
�L��]�w\�p �-۫�l| ;�t� �Jӑ����J�"8 w����o��u��6�i�@�pG>������� �sQ�_pkU!8�'CC�v c͏�vf�`�5 /�����J��"��E�G��3K�뚎 �v���o�>���N���7*�b����J�\˖zӭ2��q�[�D�������6�J�q��$H�!ހf9��x�n��1��� wfiv�e$���Crq�� /���7�� ��?w���(��^򡺄�$DD�v����3K���Q��n�]�w'��"B���6�H� ��.�;�yG �ݺ��}N���L��> �[��"�����7�����n�]�`�G��3K������c@��C�X��؄	����G����.����S��u�����f�;4 �ݺ�c�8��<��W�UU�vG� ��w^(E7I"��V����Ş��q#e�,����2��\H+�
<XR� r�M��l��}�p�7�&V�ob��K#j���m��Zm`z��vg�mOe`���=\����'���ם��ۤ&�]��okfV��.������ob�
\��8��,Jx��
���z�����	ta�GZJ��u����k YD匱��ó�&���i�����*#�aiL�Wb�m7b,&�F+gl\R�:�@#�Z��;r�=>g��6�X���]+��mr�-vw�Q���	]��n���H�לk��i(�֥n�AA��*�gy%��v�\�����sc.)�q�0�d�I���a���])T1�y� ���$[VѴ=w���^�z��^�4��ebR�U9A.I��:x;) ����ܽ�Y���Xޭ���bT�	'���� ��"�7��+ ��K�&�;��.��Ȱ�d�v�e`{���Hci��[I��[k �vK�7ve���x�U\[�<��ybj��[h������,��c�:���=\�R�x�<���B)�I]]ݻ0]�xWv^�c����0���V)C�qvՃ��@%nZ(֐���]{k�0c�Y�����X敺8YaJ�"�v��]�xݎ��O��r�A�g� %o�y�M��ۧI�M���\�s��U>Sa����v^�ݗ�Ip��[��mح���o �ݗ����r��������}�8�R�:jؗ۷�jݗ�uwe�Kذ=T��z��s׈M�v�컴;w�j���;.E��-��K�;\�7����۶+n�X{r����^�RN��F,��F�R�R�k[86i���V�N��;.E���[%��e�ݘ[�Ֆ�"ۢ����Kx�{�v^�܋ �e�B�St�(�v���;��`�e�� �"�Ԏ��~���'{�s[�N��᥅*�Q�i6����=xg�������Xڛq[�n���`���� �d��wob�5n������>�m�Q������� �������{[��n�Jd�&�u�_�n/�6 �if��۱�|��[�5vK�5n��;5É+2����8��G�K5�Ibݗ�oc� w�[���Gvs׈M�:vЮ�M�)=x�8a�$n�����,�	17lb�l�wm��� w�[�7ob�\�:(�J*�����*��򾪯��� �Ʌ�N�ui7E'm`�Kx�U���I�}#���o�]�b�t�HhvSL���	��!b���-�e6��֐�4!(�Ih:�쐤]!p�v���7ob�ݏ �G ��'��\4��
�bm� ����p��"x��Y��W�KK̤��n�m���V }��7��`�ǀM��&���n�ݺ��"x��, �����X�VR5ղؗ���7ob�ݏ �I������39����Z�j-�"�t�P%(��XJh�9=gh�r�}��R(̈́"hu�L���
���� t8DO"��$��Cf@$a�R����Ovxin�����B���"�!�}��!^�q������'�؁�Y;ܾ���	��~�*
�������R�UUeB)j���8.��a��k\��"K��s��a����ij���*�6�u���ϳ���u���[�#�؃5�#q6(�LJ��0&���7ZҪ�}ю��IJln�m�	�6a�v�׍��⹸�W��=�5�ey�W˥)�h$��=�� � <˖�h۴nxۇ�k6Uu�[N)�]U[Yr�i�L
Xc�)ˊ�m��1���nf#e��m�����՞\s\.8�Z�m�v�6�@x�u�l�v))��������l��A���2�w+5�/F�q�kI���-6w5]g�i�w]���2cr�M0�1)�� ���e]f+[�dV�4�t�Gc�u6+ώ��96z��D$�/jj��]�َݬ]��.F	�#Xb0���
PD�eL
���Ґ��-�h�%���-�҃��@���רm4�`�+)W2ѡ*��,�K�k!Âj��g<xJu�m�ݲ��&��kcV��d���O�.�+��y��srk��gOSͱ�t��&�x,�/ns:.^��Le�f���z�+�6&����\ f�kZ�Hד�v� 5��ky���-z����3P�7�*�9��R��P��`N-�[��T��p�G]Q���؃�������T�ֆ��sPOR-��4��E��3��`��U�v�8�bL���;Xr�A#��=���r�&�N�NB��`D=�Շ���S�u����镪�v��[��g��	.�֥����{]*Њ���7v&{�e!��$�"���%��Z4���6uq���g�L���;���'��T\��.�WVium`)	�D3.�)�-4B\v*�M�%��Ț*K�������tk��ܥE�sq�!��3!�۲�qUl�: /"a����D:*��s�j4��t/�Ch�4����$9���(�#F�F���Ju���7<k�0"Pm�+���tnu��س6�f�j��MMqDM:�Qt�u\Wb� O����!�X�T�P�;E�>#�D|@����殮��q�nkC�zcK��d�%=�dKK<5�v�\���8�\����)3!-�Ļ��½�
��S+��8��K����0��WM-�#@)`�0&�$�"fk�ٚ���[!�*�@���!q���5raGNɬ�Xz9��3p�Mv9+-� &-���6���!��=�/g��vu��á�뮦ᶌȽ��W8X�Û�{R��<ͮ�ŬV��=ܝ�<<h陴%�ж���@����%!Lp��z����m�De���M�:vЮ��k@;ݏ �I����~�Ur�A%�,��{v�]�J�һm�I2���o ݽ� ;�{�č��$���M�M[� ݞ��n�ŀݏ �I��E[.�BE$R�v���7ob�ݏ �d���Kx	K��� 8�w��������o ��ŀ}6�D-=���ֶ8�a���X2�l!��RU�����zSc�ert�[��ڷ�k�l�X��o ����r�ϐO<ʥ{ä���Mݎ�`{%�ʮW��C ��Ҧ�=�k�rI�;�nI�{2��e-IX�llK�m��;��`wc�>�e`{%�����lM���m`�c�>�e`�Kx��XݢLv�v�!�����}#� w�[�7ob��c��AJ��ذm�PVf\똱{v.X�F��f��j�SE��9a�I�lr�lm-V�
��{%��{ }��ʮU|����j�߶�B�Ii.�W>������t�$�;'��s� $�o !)pQR���E�`�c�&�Ń�9|(��;%췀M� J�iF!ҷBv���H�l��N�U%�xZSä�i��wi7X�e�w\0wc�'ve`�QR!���KHҝ�d�fvج
�K.n3$փ5K�(< �)+�E�[�W>��������	ݙX�����R����
��6�]�y��G�{+ &���	�ذ��1۶�6�.ƅm�;�+ ;�-��U%��O<�ax�1�n|	�\K�U�f{�q%�{�I��[��v�#JJю�]Y�r�KYJN���_<�{��:������*+�6ǀN�ŀ�;&V ov �sk��֨��A��{&�s�3�JԀ���k"��8C��rg��1sX���l��YdL������;&V }����� myDy�t��I��o ��+=�q �q/K�X�=xU� ��wv�m[� ��6�,�l�vL�t��ڸ[�ĸ��	��`Se��e`�`��8��V�ƅwv�XT�x�\����W�g��uvKܓ`x>z	�0�;i�]\5�\��
�-�H��7�Z��̷�����iԏe�ۍ�^yw����qɪ'sY�W[��F��:�6M$�;	��7k7+خ�D�̃j͍�p����	t��n�2�$:�e�0�,l��T�RݩA�74��gmH�J�v���+���2�1sZ����ϊ��m%��Z��Gq���kd1`�!Ur��{������i|�CCY]�<��z�'`��r̽���:Qy���XФƎe6v��m*�XЭ��&ɕ���:�%�*�A��׀I=��ҷeZ��� n�O?U$j�z�^����+=S�-����ХΔ�����o���ϔ:���UR[�� �؞ t8t������������X��<��^ v�Ѝ*t����n��fV n�O �vK�:�%�졖KCN��o�2y���`�N�,oL(�mNz��eܺ��cU�U�L�[���wn� �<��엀uvK�r��A��e`�Y^���7M��]j�rO/��oh ֥�w��wd������ʪ�r�;�Ez��CcNݡ�x��� �d���7v[�5l��}�6c�ui�Ue�Э���W+�T�}� 6O[�:�%�]��ݘ;�M���b�X����s�j�z���� �d��=R��%]�렻h8�0.v��F`È��Z5��&G1�d��r�E�p�G��,�V:�}����`v�X{&V N췀�\KJT��*����v�,�s��H�����=o �엀�h\E:V�N�5j��O<�vnI9�{u���~ɘ�H���,����'o�XUmH:eՎն�V� >��:�%�v�,��+ �*��7���A�q%ӻ��+��Xݓ+ >��>ݜ���R�J��n2���%�Z�)(�fr �eq��ፕ��ά,���Ct��n�v���>��Xݓ+ >��:����D����T�cM[k ��eg��a#��[=xݹ���h��o�%n���xWv^�$��ɕ�j����IRt�n��ݗ�uI/ ���UU�z@`!�wz��'}���m.KK�����$�ܪ����=�xWv^�c)P�.ʺ|
ݤB��2Ʒ �a2�j�Y,
�A�P�P��Ye���f�t��Uj݉��>�p������d�����;V�ڶյn��%<��/ ��/ ��e`gJ�L�j�M��:��������+ ;�S�;�D�V�-�Nݡ�x��=��;��Xݒ���ʤ��� ���c�am5L�ۼ��������xV�xj���*��S
�@��j�U �"���}�g��\v3�U�K�SG.���*3�����8�Iv.4��	�Jh�ś��Z�38�M��05́�̵$�.�Yj»X]��Y۶�@@�Pcێ7V�^����ά���c�ڞ^������wKvl�a�7$Jm�s��bY����s�.9:�C���Oa��<�.-�rQ�ܳ��Wh���n%����	$��4f�[�Z����Tb M��o&	�� �a���Pt�P>3��3�n^�C�6��N:�W+������7�n�ٲ� }ݏ ��/ �ve`6Y�Mۺ,*���x��x����fV lڏ +��|�U۶�Se�n̬ ��� >ݏ %��Wv�V�؛��ٕ����۱�we�U�*:wN�mZv� 'kc��c�	ݏ �d��>������m5�wj@�n�{,e^��d�nB7Fٷl��WR�_5�%ؘ���x����'� N�x�&V N�ǀn�%c�]6;wI��wcϪsh�	���\�����d���W*UUf��+ >���wc�6Q%�[�.ƒ�o �d��	������we��1��[v�v]�(�u�����c�"���>�e`Se^pi��]���x��������������	���r�\�4T�J�#�SM*B�5�m���^IR����ˣ����-Ʈ%�?�,�Χ�M/���Z��?����>�e`�lx����aj:.��+v&� �d��r�ă�S� 6O?��-��*���'t�6յn�v�< ��x}�]Uʢ���!	}e.и`��Co�i���Bi�.�e��R�!Fh�bG.�a	�0����[��)i!�T�P��I)[�@+�3�dN�<t�fУ�]ԠBFN9��e��qZ�d2��)��KY	c�F��/0�%(.l�a!�����XP������,%)4<7��ޣ{��h�	�T��!8��D���-�6@���1!@�Z:�����{#
�2�#� �h@�+))���-e	iY+*�S0#�!鄚�H,d�$��+CA>)Ф�Y%ز�m'B�JP����F��R�4
ҤF0�-R2�]e		r��e	IJRI3jof�	�L	�2ku 6�P�:�dAH�H�
&��&�C�=4��Т��p��G�	T^f_}�6�2���*�T�-ڻ�V�x�-��yl��vL��ǀ}�D�,wc�lv�m�we�vL��ǀ�ǀE!Wr�v���9wb�f���I�{%��(^-X���ci7 �4X.�ݖݍ��|i�	ۼ����>Qlx���$��k�K35�e8�q1����>Qly��I[=x��^7fV�6V2���Uۻ���"엀Eݗ�Mٕ�|�����D���
�q�m�v^6L��ǁ��UUh �(���QA� B0�.�"&ED�bD��
H*�w�o7$�'��zI��RM؛�l�X�-� �d��s_Wݢ5�I!L���Pr9J��x�����nJ�k�Ȇ��VRk��5��'�0���i�V�u�^S� �d�.�I2�iȪ1��j�Zm�I/ ��/ �L��ǟ��\H��S��c�`���g� �L��ǀE$�e^Xج�7l�'n�	$��>QlxRK���g� ���)�۔H�G+�+ǯ_^����z�/O^$�X�IQ�+�V���p�(Z'����n@c�,J*Y�:I�K���0���5���2��G#��k2�ȴ¡\Û�ja��-���Ռ���fYBVl�ط3�2��d�Ad4����������\�
t�9��[c.��af��%�CHK�%1�ЇXݗ��,��3H70V�L��nb�V�-�iUPU�ժ�6�.ҩ��Dk��u��V�`�q[��:ALt����[�v>��t��<ͬ�X+��h.��:�������kK(���BQ�K*ns�H�]�.���un��5M��I&W���9��������]U�˖���w�j�/ �L��r����GvҔh���7x�e`ir,=��|}��y�Ko�W�I,���lPqұ۬R�~��<�=xV�M�X4�Uq;�v���m`M��{���=�Oe`mȰ�m#H���Y(XP%��ʥ������B�����[�|��E`�i�X�ܙ�ૼ�����'d��>ۑz���A�'� ��z��6�i\� ����'���:I�&�$C0Lv�Z⒎�`5F��"W-I#�8#bqR�H�HA"o0 ��H0����6��e�����"˵V�ݺJ��u�|���"�/ �ݗ�I�+ ٲ��4St[eݷx�*��s�����"���$��6^ Vʥ�TR��e0v�����	5� �M��E6^�F��.�"�0�s�y�4��+�Ψ:xN��l����}	�첹4��4&�I4�7x��|���$�� >�ǀ|�EQГ�M7t�m�˻/ ��, ��$p��Ȫ�!��m]�+n�	.E�wc�UUddR@!" �w��f�_=�`ݥ),�v��l��m`���	#�����$�%^[M*\�nēV�$p�=�r�{=�_����x��)Y�'h����M7���Sp�66k�d�eb�M�!5�
X�U��e�l�e� �we�\� >�ǀI0�i�(h�O�[eݷx�"����G��/ 6U*P�R�R��;n����	#��엀E$� Ӳ�j��	4�;ok��8`Kذ����亪�+�#��ީD0���
k�\2$�B�O�xV�D��wHcwJ�۬�{v^ ov<wfV��W{�'��K�IB�@�C�Y��������7HPҩ��.Pz���厅���8�m�l���c�'ve_1[���ږ)���E��&� 'dx�̬ ���we��6Q�����I+�`N���ݶ����H��K˵Vӻ`��)]��	$x]�x$� ��+ ��p�l������.�xRK�&� �G�s���7*�����|�~�B����/U!H�bYI��ʭ��
��Hu4I]�(��5f���p���g�ڭ��Eki";"��׆�e[[F�5 ���|�{+�/g6Qx3\0(�/f��op�mCtR�ݦ	�
�YBAi��Pa
��e�
�;R���g��2랤��6i��6���X\U�vv嵁�gp�`�ѭؖ�*�,�wI��L�!>����Gn�T���zK��c�������X�5��K.8�l��eW@���c� I#�&܋ ��n	�:.�BV���X�2�wc�&܋ �\� ޗ@l$�I�ڱ۬ ���	ۑ`K�`�2�˽�O�k�k���|�'I%�����}~��'ve`�ǀw�ԺK)�b�˻��k �\� �ٕ��;{������=�V�jR�˥c{{]7gL�\Prl�s��3H1�	�-�fX9%��6Ī���l�V�ݗ�N�ŀ}��`lV��ӻ`��)+u�|�e�r����/wS;���I�s���=���`��RO���.ջ�>��`m�X�fV�ݗ��J��J�T��Zm�s�K��� �{׀wob��-Ǻq%�`�\*S��rF�8��d��{%Ȱ��X�\�+������E�U��[�/_X����m�s@�(�M�i�2�6��&��"�ŋR+W�'�ߖ&�`mȰ�%�K\�WM]�˾	[��\0�Iv\��Zg����3_WՔjTq(�nـ}��`�%�u��WNg+��U_<#DQڛh)Hd�0(h���*���¹���/ �c�M�a��J�&Z��kܪ���'� ��� �ob�'vZY�i�t;��I� �n��=���<|e�,�ٕ�v����~�b5���.*7Y�)i���s��e��ff��cv�&z�I�[�a����Q�����n̬� +zqR�R�TYL���vL��W9I�������9T��"��][���n�`=�m�Xdp�'d��>�])n��C�i7X�ذ	�� ��+s9GWk��*�>� }�j�*wuAv�68`�e`c�6�,{���T�e�ݪ������k����=�u�V�TV��X������K��N�`�t��NـNɕ�M�+ �{�A�y��=(�1�B�c(��;u�~�W��}_�s� �8`�e`�MSI�M�cUj�`ob�6G=�K��e`��V���E`4Qm�]����R�2ݙX�2�<���
�8�W�^���e�l�'d��6I��M�� �0U)}UM�H�1�|��#N�Ňx���$3�6��:���l�C��4I<�]!������k[=�|7��xl��r�}��_s�A7�Y��M%����Kt�6�I��B�'�y��	�r�h����4��xā#����)�r��Q�0�q�*u�$��i�	�|0l�R��"B\vxj��6S�hw�xM	2�7�_ �L�ͅ�Y����9�K�:�L�9�}�%xz�6E�	�/P�!��b˽��n�n$�F�������*���V[UU�M�����3pUU]U*�ٷ>��l�[���!�mK�F��M�,D��ki�a0+;m]����ٜ��ݲ;d��G1�:�:(�۰6s�E����!A�|<W��%��D����<�N�,p��v�s��s���[�m0���;9��X�rV��b�����0�,�:�e����r�V&�-w-
)��u4/J��*�O�[��d&��5��lp���a(k=k8�k�o1�.�&�f�݆��a"`v�R4�7Y�l�;�q�%��E�K����0d�sdɵ;Y���3��@`� ��Z�%hE�h�M��ء4j7)�uZ�b^�P�zŷ`X��d@�+C�g�kؕ�Ҙ�������1C6��+K��ۑ��hق#ū�rV��G	[�I��j����^!�G�mt�J�\$����T.kP@�Z�;��6U���i^���kƵ�t��,��.ࡕ�.az��1g�T�99g��m\�vrcu9lrv�M�]�\;m�2pt+Ptt�j���zlຼ���4sZ�2<8���oC�� yt/�`y�!��m[�V�U���`PAt� N�]j����"m�v�F8m���6WB˱��E��7`)�)8��M�l�NZ%��Bm=K��.2D�u5]�o�W�,7'R�[ml[U;�p����f��r���h��0�� ��f�sV�K������Z;���X�E<8&V�6v��KЗW��˴�lM7��� �.ֲ�+i�Lmj$�����d��]q5�۠B����۷6\�șʚ�WU�J�,JeM���U����uu��BP�WR���ŗ"0�A�ґ�x���58� �XѠ�����l9,��Z7a�t�b�j7rg�����3���УG
H*���FS�iV�y��Sl1*�j.�t�A��ե��Y�a�Lj�"��nxv��(G����J�C��t��L��5�)u���hCC��4�lN����z��t��mS�����mSD����UC=A4� ���au�e��\B۬���P��mu�#wev�
�M��b�s�>�۷m�v\�cv�/-ږ�Յ�K�c����E�,�P�Li%���؞)S��m7���ag�G�͐��t�uҪ�9�s�8��r	�\��T��0i��뢈�=d�T�]	�*����l�{����=[�Y	�i�(7����'Z�9��Ak�I�I9<����3j]�"g;��KJb�Y`��E��]5s��p^6gq��V�-ή��vݺ�;�2�	��`#�;&V��J[�*�Lwj�n�	��`GvL�I2��8R���⫻�-[�H�Nɕ���R^����yI��;�Ҕ��m��M]���X�2��e�*�r�6����1۬M�X����z�z�ޏ�;�+ �+��j�)w�i��iT����(Jc[��j�ͷ��^�2,�l;h#�(�����׀I��̯r��A�Oe`���!��@�;gx߿���I�:{���r�r��	�̬�ٕ�Eݗ�:R��B�J�]�`�2�	�2��e��� �VܻL�W`��n�`ve`n��'c�;&V�yu�Kt�v�6էn�	��`����<|����&���>�k9n�B,�t��c�P�Q�,b}	�F�q����e��A�>�J��`�Uw|��z?�X͙_���W�=.y`���Yv�`��Wm+k ��+ ٳ+ �v^��m�!Sg.����;�2�	}���\e��Y�r�yU\O�0�2�݋@�n�M��ݺ��9��r�����;<�`I2��̬T�
(U`�-��m`lp�>�e`ݙX��Xe��@���M)ncs+i%]B�c.�]�����T�yI`53a)nxi`�SZ���k�}$��7ve`��`H�E�n]�SE�t�m۷X�Y��9II��7�~0��X���J[�V2�ڴ�� �����}�e`�e`�
%��I�uw|����0�f��<��ٹ4 �C�P���w�nI�5�e��v���Nـ}�2��2�����p�7og.Ӵˤ;���8H(�΃�]v^�B�Kݶz��V΋��av[b6r�&�`�2����0��+ ��Ɓ���6��������r�7�~0�{+ ݓ+ �#�*�`��[��8`vL�vL���/ *j\�g�.;k �l��7d��5we��"�"�Q�e4]'I�6�u�nɕ�{�ʗ�����^�ٕ�wHL��+G��F�q[]�H�Z9z3���*ށ�X���*��Ț:m�b�0q[1X�S�(��3�v��8�zϱ�tY.`^3#��#;n��9���9]T�l�����&�]�g��+Vw95K�p�DDl�\hLPż�+�+H���f��:³�2�(�R2����H2�4Cs

�l�aՒo^�լ�IӾt����x���)��ji�0��YD!�c.qK���f�&�j���o�y׈�]*���ZM�@�O^�$��+ �ٕ��*����n�����̬wfV��/?r��I�v��[�Bn˴�������n���yU\I-�x�Ixj�I��*��X�̬�)#�g� ���x�ٕ�n�q�clt+�X˻/ �I/ ��2�ݙX���*y�]�������K5�"F=����H�������P�n�(�(T�g<B��Q�;��o�X�ٕ�wve{�_��j��x^�s��e�&R�̺�ܓ�{ݛ����Y,X,�!
�A�@P(H�B�R��k+�@�U+��E�D5����7$ջ/ �[�!�M�����7d��>]�x~�K}�� ��e`mXD�t�_�E�� �we��� ��2��2�y(��RN���Z�xeȰ�ݞ��g���|����|��}]5�-��з��(YZ�r�X�� ��"\�aX�!Z �WfmIx{ʣV��ve`�2��v^ݹچ�CM�ҴSm�ݓ+=Ď���T�� �ve`[����E�j�� �n��:����H��qU��"�R4&J��tD�R
�q
���Ogr�wfV+vg
�U�
-��[��\]�y`��X�fV�ݗ��EmՔ(�q��X۳+ ����>[����XГ(�V�7��I�j���m�;�c���태ō�n��M����t�]��Uі,#b����>��`[����`l�X���IGH�t�jէn���y+ܪ����}~��V����7n����]�V� ��� ��2��fV����>�e��t&���'l��+��R���V�=��_=�nN��"
@׽�97$����i�m�]+E;n���+ ����>�`vL� ��)Y
Wv���3�����ڝ�-�a���Ψ馰vX� (���:O#�|cGf������}�p�>�̯�ʯ�wg��V��V(�˵n����ٕ�}ݙX˻/?r�IwQ�vp^T����=��}�2��v^�� w�an�]7E4��n�?s��'���g� �ob���U.��Հv��<%�I+Tƭ7v� �we���.˞Xv{+ �vd�I��C�Or��c\��lG4.q�V�У�lj�9n�;�����h�U�Z^��#ixn��g�T�K�N@;^��nڭ��c�A�fa8,�&�z��k+l&օ�?�1��-ƙ�+pF�]����\q�6۶�*�v���K�'0�ˬt�6�gs� �����L�0DtqRƴ,i���43��(���0ֳ�]���[s˯/^�֦�Q����5a��T�jH[,�e C�PȆjFmj�+��� �-�j�R]��@����6�Lq�%���W���$}�2�W+����l5{߯ �?S��.ڴ��uv�m`n̬�ٕ�|�e�m�Y���I^'�[�i�t�m��&�e`-�x{�+�{���`�~��;]�pe6�h��j��X�v^��� �ve`�2����$X:�ݫw�}.E�{�U�=�|��X�v^�w�����+t��lE������Ya72��0I�)��.�a����Wv�q�������7ve`-�x��Xٻ��tf�l\����>}�y륒��H H��H�����T>S\�S��m�,�ٕ�}]������Tƚ����ݗ�}.E�}�2��̞ {�-�d���w�x���'���ߖ����ٕ�|�e��)��vջ�B���k �ve`ݙX�v^�܋ ��r�+����AWH�v�B�HYu�%!.ST�q��Je0B�1z��K@���M<�b�lv�&���t	=�+ 7��nE�}6e`��8Sl.��[j�`�c�>�Ȱ�̬�ٕ����yc(���*Uv�v�ݿy`M�Y6yHZA齥�ғ���*$cM��N2e�����-.�@�u9���[�����8�ޙ����|�$���^���z�sDf�]�)$���^�Il:X��J�Av1�B�R`%��٫B-���{�8�)lO.��`y=��m8���G{`$�@��mp���びl)[RIe�|��c2:
�x���^��S�4<�å��tC��%�H�$C�0ǚ)��L1nP�B�S��IS��Í&J���׮��R��ᇦ�Wl�@:/��� ����H�
�Ӿ/�x'��U��S����y����rI���o��{c����cm`�{+ �ve`{��v�X�ەv;�Wmm�;u�w�2�����r,�ɕ�}��b���{��n�x!��Sh�f�^�j��vᓴ���8z��c��E�S�o̓vy�v�,�ɕ�}�p����ӱ�7|�[xݽ� ��e`�2����Ԕ�p�j�ۡU�I��}�2�	6e`{��^ş�UI�O
�7t�N���n�>���}X�<�$�s����g+-R�.���䞞Jp�6��L@����	.E�}6e`G���Z�#����T�Ӆ!͈�s�Z� 9#i�ñx�]<j�e�˅:�Uv�v�$p�>�2�	#� ov< �).�	`�\v[f�ٕ��+���D��� �<���=UU�q �/�v�ӥc�6�i� ��� ov<�8`M�X�ں�t%j�ի��x�����}6e`�K��h�li�X���8`�r����� ��x���[ʨ
�"�H����o�.�#u,z�.)n�t��#MmY��bL�����J86�Fͬڣ`�(�2KV��&�"�L�&��yQ8�\�5ō��!��3e��v)t��[0��IN5��n��r�Vgv��ٮ:L�k�68���[h�NݮZ��������S�:�V�,Q%�e%m�Ԅ�֌lf�g�Sc��c�7\�0c@�a��v��zH����|� K�80��5kd-�LH1��R��*`q�#t(R,tt��f���mk��|����� n�xv8`�6$ؓ
c�h�m� wdx����p�>�2��v�q��V�n�M[x�\0�Ȱ�̬ ��x�S�N�VRV���s�K��, �x��xۮ�Ur���)x�=WT����� �n��>�p�>�p�"�E �O����[r�k)M�����5�&�]5%د��Vq�6����\�Q}���ذ��ۮ�*��_ ;�� �ھ�^�.�e4;m���ܮQ�8r�P�UUϫ��7.|�{���p�55*Q�����+f�� �������ݧs��V;uj��m� }ݏ ���u� �d��;P�m]Ӫn�H-��wu� ���}�e`������)jUؐ���f�Cr+��9�v����b3����"�n��GE"*�+]U<׿���>�̬ �����"�t	ؘR-;� ��eg����7c�}�p�RA[�.�=W�.;�����'�{����t#�b>y�5�M�=��|� {��}�n��KUkU�?wN����wc�}�2��������tʷc�ـ}��}�2���x{���RW��[L��WV���oc8����e5�V�qrBm�2�KI��ci�� M���[�j�P��g��X�v<������1�.�bv骻J۬ ��~�����;���>�2�ԑ��?'m���lm ���?��=UĻ=� �x��dT��lUl����UR�� �������>�B0A!�&���n���ݚ ���v�V��+ >�ݽ� ��%���Ue��ҥ��0YLIZڹ�+�;Z�n�˃mC��)��;O�������`۱��ذ�\0�̬�l�ۻ]7Bn�m��}/b�>�p�7�"��c�;J�A���j�n��}��onE��I�� �\���jT�c�wM_
� ��ŀwc�>��`ywfx�7|���0�(�0$8�W���+ǚq%�}�f��=�ܓ�_���(�!�2��t"ą�Asn�K����<��\8��e۵έ���c�`6,
�I�,Ќ�1iX��tNm�ۡ�Դ��]��7#�w�Z�Gf�#���$`���D�7v9x��Ξ9�f=dcx�ֺ,,K��5��K[���6�O.�Q��3�&����3������v`��k��36f���b6�a6�ͅ�ݩl�f[���=Q�[(V��&��-��IӼ�xO$z{l�p������ˊQ�ڸ���uN5���#���b���+R�gE�>��o� �\���;.y{�Uϐ�� ���*cbn��w�}�ឮr�#�� vO<�/;ʤ��S�2S
n48���y�J�6q%ff��� ���]��*e����c�>[���\0��,�l����];�6ڦ�x�v^�u� ��ŀwc�>�Iԫv����wLl#�g�9�-��ө�KD�!����&����<�,eںe[����v?��X�v< ����jT�4�Li�[0	��W�U��W9�*���>{ w��u�?RD�?YEؘ�m]4+�`vy�� ���Mٕ�w���-�]��T�o 'dxۮݙX�K�y�����;v�T���>�p�&����c�	�����/�C���1�ͷ,��4V�PY�jY���B$�qJb�M-Y�rA�|��V }6< ������T��J0�*��n���`���;�p�&��vS,:wBwo�6�l� �u��9L�rʪTR�
F@X
@�uC.�]�f��;�.�Z�;���݅ݷ��Gu� �0���=UĽ=�vY^���ͻI�>�`�� �W+��<� ��x�� �j+b�t> I" !&��i�+nf�V��+I˵m����9 �Wf��x�bn��I;f }ݏ ;�<��ݎzA8[�-ݷcim�vG�}�p�;�� >�{�T��'�դ�BT�m�c�n�.�x�#�쉰���.4[b�`mR�&Vd��d�����WyUO��� *xKUؒ�)
��v� ��^ղ^7\0�XГ;c�.Nq�Н!X���W`8���ks��a��:3����J�p���	n5O�:�K�&�ݎ�W>A�׀v�mU�av�U�%v� ���U$I~��<�޼�Ix�-]�n�I�>�`�"�"���;#�;��S�V
�t�b�BV�v^�0	�p�7nE�w�ʷt[m�;I$���� ��v�X]�{�D5�����<&zjsqf�_P� �7�M���B�Á3
И�5�o�]y�ܼ׾k�w�މwhG����$�)�'��a*��ztt��a6�N#"��ySxzf���9>�_6'��_>�3L�8�f�4!R/9�g���.���>���_ie�H�f��	�Ė}	��.�V�9u�>(�(2�k�����z����@SPY�>�$�~nk}�'����;�!y�񑺠I`Ro�R�HkI��5��B��Ow���@�)bIȞ��ϔw��z��ַ��$7*�d� ��!��R%��f�w��w�E�MkZ�%�]"I5ӈxA�Bt�&{GC3<}%Û����g�3y��~o�H�4ɧ� Hkr�d��;��x��dta	�e��]DZ��Clg6���Пvw�o�>����S�p�> l �d����d!��$4ith�b�Ȥ$�H�\� B���+"��#�kc�e����V�c�**B̙~<:/��!����]w��xx���
!�vU+	��D��N�4I��������g�a�qg�7��[j�
�U����r��R��UWU@]������k�ƒ�v5�L�Qs���vy��"�F�T�	��cCd"ز����1lZ�si ���Ǟy]j ��,6y&��pd�	Ba���lv�:(�l�9+[���m�k��)&X�`�����cmv�ٜ�g��$�p��Fbk$73��f�H]rVH�W
$�[N�YÞ}�J���j݌{uu�F�g��@-�|^m�c�����ҚQ&�B��,Fr���
���U�-���k+rh���CQ��3U��Z�c����1�g��U��4�2�T���l/$���91�E�ݶ�wl<��X�����T�M,m�;B `,	���z�΀��os�t�����*�j�@%�e�6[XY���*�e&�v����6U������4O��ƞ�0Vv���` �t�����P� N�;�b��+�q����y�[Uǋ���Ø^u.t���k��r獭g�2Q�.!yu�|�-3H�95�Ƨ��qñ��h�ֱ��hd��\���-��±ja�ed%%�ek��4��6��˃{9^�����[6Yu��6�
J�)����O]���P�
��#��` �k���Ë��3Ϯ�Sh��U��q���aɺ-�
;%I@�eٵf�,-]&�N�rc��*t/<1�UU1N�m�cT�J�.A*bCZ\���'jю�%��Jjޝ�`8�H2�)��0ѥ
V�AmCdj�T�viҦЗ��X4�p7J��i-5Z�ݜܨr�ۅn6C�2�-Jtt��be0��/��r����o��{v�^�3��m(�a���ėA,�V���X6�ݺYʻJRX4��Pp�Q1)1���-E����1�!Y�u�c�R<kG��ƥd&�\�;�����s������KÛhףZU�U���5U�ں�S��@S�Z��e�t�+��$�۴񍸲�q��̻�"(el���5�Yq�l1�P��Q\�h[�=I�;��s�=P�E�� �P|�<}���=\18���Q� �t����¹�"����-u�ʖ�Uc��s����]�	Y�g��S��m�͐u�T�(7&��[�+���ST�i�K1f"�4e(4Z��d4mkk#vˈ�5N2� tA�J:�y�[�q��gh1�ҫ�m���v����܅�m<������L�c�P�=f[�m̈́��q�VWGfu���0�mF1r�E�#�(�۲��0�c�N�xi���ȘM�� ��gCj{�vV�],˩j�^(sZ:��b-�A�8
��6k�n܋ ��/ �0�6v1.��[0	�"�"���&�w\0�Q]�W �U���.�x�p��^���=#�uM�i]6��+m�!�x�p�&� N������[�"t[t�.ճ �� �������p�	Gy�hʊ�P�
J3c<-YC4P-����� P�z�18|Uy(����o�� ��/ 콋 ���ܫ.��M6*�Cm�we���UYH�%>0������>KS��� ���j엟�����F��{*�Э�t]��n���,w\0]���%���yg�6��@4���H�`�%�vK����X���e&>;�WVح�]���%�ob�&���`*�WhwV+I������]4��{�l��{H�G\V����Scc� N7$�KN�$�ŀM�UW>@{}�j��Ҷ�:J�wHm�6�,�W+���� ��� ��/=\�RD�(!��v�!�����>���nI=����z����ל�0�s� ��R�F�ؚi�� 7�<.�?r�ķ�<��?�Z�AwM�I��o �ݗ�w���`���7gx5t��J�M�G �zz�x;v�teM����#2�LL�b��%��V���ӱi	6��ذ	�p�� 'v<���cj�N�����N� wdx;#�;�"��l�U�m.Z�M�ـ� N�x�Ȱ	�p�
������M�����>9?w���r%�bX�}��]�"X�%�����iȖ%������ eR�AJ$t $PO"y�{����/B�/C߾���el�kiȖ%�bw���iȖ%�b}�w��r%�bX�Ͼ�[ND�,K��>t�t�Jt�O_� ~c�����ۥ�K%�.bne�,n�`����M���ȔR�Ξ���N�����?t�Kı/�}����bX�%��[ND�,K��~�ND�,K���:�WVCd󧣥:S�:_�~|��~ #�2%�~�ߵ��Kı;���v��bX�'�wM�"X�%���|���ge4l�/�=)ҝ)��߾�ӑ,K�����iȖ%�b{�w��r%�bX�������bX�'�����9vɭ6���:z:S�:S���~�ND�,Kϻ��ӑ,Kľwﵴ�Kı;����r%�bX�>}��L���eV���ҝ)ҝ>���m9ı,K��}��"X�%��{�ٴ�Kı;�w��Kı?#��V�_��]]]�՗Tմe�[�X7dN�j�g�j�p�"��BW>A.�t�oDJ��d�v� 4��p ͤl0�t�%�-�s�Ea�/x;Fx�����[ Yv���Tc�0.ֲ�0�!MH؎�&�k��m�v��Y톫jە�#�;�mv�YɺuJ����jb܂g!3z���I�l�L7Rn����P,l�����Џ����j��k�'T\ H+�b-@_<���c�Vc�4����q�tۈQ��l�E�Ŏ�#/2�=c�#�a���%�b_w���"X�%��{߳iȖ%�b}�w��Kı>�������^��^����%�b����[ND�,K���fӐ�$r&D�>�_~�ND�,K�~���Kı/�}�����\��,J~���5�XKsZ�Y��m9ı,O��߮ӑ,K������Kı/�}����bX�'��~ͧ"X�%�|;d�O����ԳE�֮ӑ,K������Kı/�}����bX�'��~ͧ"X��Y�;���v��bX�'L��f~�Yu�u��a	����Kı/���m9ı,O�߾ͧ"X�%��u߮ӑ,K�����iȖ%�b{�~d�֋� ��{&Pӻ�B�s�^��#�K72��j���`�X��T%�3�Y��/�=(�%��{�ٴ�Kı=���r%�bX�w��m9ı,K�~�[ND��z����=�ܹ��  �Ο/B%�b{�w��D�$T�D`:���'�oM�"X�%�}�ﵴ�Kı;����r%�bX���f}Mfd�	�-�Z��r%�bX�}��6��bX�%���ӑ,0ș��߳iȖ%�b}���v��bX�%�O��p�!�ܞt�t�Jt�K���ϝ9ı,N��6��bX�'{��v��bX�'�wM�"X�%�N�o���>5f\i��ֶ��bX�%�}��"X�%��@��o��i�Kı;���6��bX�%���ӑ,K�����:�f�j�I��tWV�o/l��SF�0�EN�*N㱴��zxfx8jx�kiȖ%�bw���iȖ%�b{�w��r%�bX�Ͼ�[ND�,K�߽�t�z~�:7�z�����4�ƹ�Z�ND�,K�����Kı/�}����bX�'����ND�,K�_���=)ҝ)���ߧ휘R�n�3SiȖ%�b_>��m9ı,Os߾ͧ"X�w�J55��4Ӥ`ba����Q(�'"k����Kı;����Kı=��y�����)����ӑ,K��=���r%�bX����r%�bX�����ND�,ʓ"g��~�ӑ,K���~���t\ ��ϝ>^��^�������Kı=���6��bX�%���ӑ,K��=���r%�bX��e��a�Y�m��G	�z�f�1B���`��n ,�	�ab��1ұ�hT|��bX�'����ӑ,Kľ}���r%�bX��}���&D�,O}��<���/B�/C���f����%�M�"X�%�|�ﵴ�?#��,N�~ͧ"X�%������r%�bX�����ND�,K��߭˖|h�1��kZ�r%�bX��}�ND�,K��~�ND�,K�~��iȖ%�b_;���r%�bX��ߟ����6��̓Y��r%�g�U�o��iȖ%�bw���m9ı,K�~�[ND�,����b�B[4�PB~@��bk����r%�bX���~U��mV���ҝ)ҝ>|���ӑ,KĽ�ﵴ�Kı=�~�6��bX�'�k�]�"X�%���=�c�m%`�X<�#�awd����⎎һ�茱����=����4ڱ4=��O"X�%�~����r%�bX��}�ND�,K��~�ӑ,K��߷��OGJt�Jt������1��Y��v�iȖ%�b{���m9ı,K�{����bX�'����ӑ,K��>ﯝ>^���:7�z}���?�4p�V�iȖ%�b_߾���"X�%��o��Kı>ϻ�m9ı,M���9_�r��G*x~,���tPؖ�kZ�r%�bX�����ND�,K���fӑ,K��=���r%�`~	�?k�߳iȖ%�b_{���N��$�K��ND�,K���fӑ,K��뿿f�Ȗ%�b}�_~�ND�,K�~��iȖ%�bT4�(����> ���2�EI3��}���ZF�Xܤ��a5l0����2򏮃�V���[9�%�ŷ�="���o���e���h�A9�&-L�5VF)Ӟ�Փ�/Hj��a�14�@�Fh������
�1ǚЄPbP9L�(��лEH�v�3�s� nĦ
:b`�R��%��4F�]�����a�H����\)g�#����������j)e�}�:wH�/�	f4����r���#�H�F�9ڔj��!��-	s�#��k��;|���/B�by�}�6��bX�'~���r%�bX������O"dK��?}�6��b�z3���%q�J�m�|���/K�����ND�,K�~��iȖ%�bw>�ٴ�Kı=�~�6��bS�:_s����j�[v|���N�K�~��iȖ%�bw>�ٴ�Kı=�~�6��bX�'���m9ı���~��2詜�Cd󧣥:S����fӑ,K��=���r%�bX��ﹴ�Kı=���6��bX���������2�Z;Ξ���N,Os߾ͧ"X�%��~��ND�,K�~��iȖ%�b{����r%�b��?���)��MC�clD�`��,��dX[mZr���9�æ宰�2^tam��5�A$O{��M�$�;�͉"���M��%�b{���m9ޅ�^�}�Ԟ�0e�y���^,K�~��i�x�
'Qx����9��o�3iȖ%�by���m9ı,Os�ͧ"X�%�|��jZ$�YL5�sSiȖ%�bw;�ٴ�Kı=�~�6��bX�'���fӑ,K��߷��r%�bX�a߭�\���R��ϝ>^��^����{��O�,K��>���r%�bX�����ND�,�̉����6��bX�'�~�����+ns�O��z�z{���9ı,?G����i�Kı/�~���"X�%��{�ٴ�Kı<��|��8jKYja�k���&Ԩ�H�YZ��T&9\���n����.�8�1��%�bX�����ND�,K��}��"X�%�}�ﵰ� O"dK��~�����^��^���َ˜�356��bX�%�{����(�șľ����r%�bX�g�}�ND�,K�~��iȚPʙ�������L̚�х��ֶ��bX�%�߾�ӑ,K��;�ٴ�K���E�g������/2�b�̄.b�B�dF�$�k0������Rm�քޮ���%	a�F��F`a�W$cLS*�NÄ�ۄ	.�7byqS"Tߏ&���I��'���7��p��bp�@@�2S��]5�C'X�a @���D�ON}�d��'��zO��q�$�%��Z9X�XA�L}��H�$�WF�͙MD0�X�!(J�8�cCHyM��W�b�b��ק�e	8��3IF[�BI�&�I�w���4>��	e0%2��t�;�5}`fQ�"� �k �]L-��a+�%P!bP��z�P�SX�$B��=i�v�!�K��xs�<���wA�����(�
҆g\̈́�(��@ �M�a�b�Q�CФ`�P�!�	A���Jh8��U��*tD�HhM t@80D����EC��p���>UC�9�����O"dKĿ��߿��yı)��~��_�.�K����󧣥:S��2'�����r%�bX����6��bX�'�;��"X��dL���kl�z�z����c_͍ڙ`���9ı,O}���ND�,Kޝ��ӑ,Kľ{���r%�bX�g~�7���^��^�}�޴k�mnR���K��B荰05�YjP0riBVˤ����.Ir:�-��SΞ���N�������ӑ,Kľ{���r%�bX�g~�6�y"X�'{��M�"X�!z~g���M�h��X:y���^�K���kiȖ%�by߷��r%�bX����6��bX�'�;��"X��/O�����`:��o:|�Љby�}��r%�bX����6��bX�'�;��"X�%�|�ﵴ�K�)�����������Ξ���bX����6��bX�'�;���ʙı/���[ND�,9ĪV5!V�JU�D�E~iȝ�?~�ND�,K�k��sZ�5��f�%�M�"X�%��{>��Kı/������bX�'���fӑ,K������Kı?�=�����x�^��;�XF)t�F2�#H30]KV<ٚ����i���V�MM���{:X�%�}����r%�bX�g�}�ND�,K�{���� șı;�����OGJt�Jt��_ؿ�r	���v���Kı<�~�6���X�L�bw�o��r%�bX�����ӑ,Kľ{���r'� ��,N���?h�]�SZ�f�iȖ%�bw�o��r%�bX����ND�,K��~�ӑ,K��=���r%�bX�ߎ���S$�Jk%֦ӑ,K��ޟp�r%�bX��{����bX�'���fӑ,K������Kı)��>.EɅ2a�6��bX�%�����"X�%��{�ٴ�Kı<���m9ı,O}���"X�%�M	#�{�����-�ˉ34�K��vh�f2�hsvG��Z�o��y�p�H8�gB\!�r�CMĉ��\�t���uԽ'�����ێ2���������Ʊr{��t�b���ۮt+ef�0 ̙骏X6��2�J�umv��A���[
���'�6�s��D��Y���Һ堑�PP�
��!1��c=�ڏO<��U+�t��)B�d^����n����'N�����z�,��׵�:�6�.�z���=�7nǴ�h�k��k��37O�WK�WZ��ؖ%�bw=��6��bX�'��M�"X�%��>��K�G)wg�r�9H�#��Wl�T�Lcn�fkZ�m9ı,O=���ND�,K����ӑ,Kľw�kiȖ%�by���m9��S"X����CR�2�ɣs<���N��N��~�ާ�=	bX�%�{����bX�%�����"X�%���}�iȖ%�b}�[n�Ԋ�:16�t�z�z����:|�bX�%�����"X�%���}�iȖ%�b}�o�6��bX�%���K�eю�Ԧ��OGJt�Jt�?}���"X�%��~��ӑ,K�����6��bX�%��}��"X�%�N���K=A���mj㭚gd���^�{[���bܮ�E���ք k�(���l�ꯉȖ%�b{߾��Kı>�wM�"X�%�}��kiȖ%�b^�ߵ��Kı/~>��R�WM�L�ND�,K�����=t�	� �� ! ��(�M`�ND�K�y��"X�%�~��kiȖ%�b{߾��Kı?!��X~�?��YJK�N'�,KĽ���m9ı,K��[ND�,K����"Y���2'�~���Kĳ�����Q�A���m�O��z�R��~�ӑ,K���}�iȖ%�b{�f��ND�,K�߾�ӑ,K�>��߭Ds`f�|���N��b{߾��Kı=��M�"X�%�}�~�ӑ,Kľwﵴ�K���������b�\�Ҁh[Bf^.4�@�2�.n�1J���+��'�j��Xi�kY��L&�GȖ%�bw���6��bX�%���[ND�,K���kiȖ%�by߾��Kı<��Xn_����[sS56��bX�%��}��"X�%�|��kiȖ%�b{߾��Kı=��M�"u��,K�ۼ��:mJ�|���/B�/C�����Kı=��m9��n1$*Q��%F�ȝ���ӑ,K��>���r%�bX��5�)��g[�i����ҝ)�>~���r%�bX��wM�"X�%���~ͧ"X�%�|�ﵴ�Kı/���R�Vi�K�6��bX�'����iȖ%�bw;߳iȖ%�b_=��m9ı,O>��ND�,K��>�n�����`S��c��)!�l/�� �H�Z�9��cH�:	eSA.B����r%�bX��~��Kı/������bX�'�}��"X�%���=�t�z�z����{Fm��.��iȖ%�b_=��m9ı,O>��ND�,K�N���Kı;'���|r��G)����$�;j��u��ӑ,K�����Kı=����ND�,K�~��iȖ%�c/���>t�t�Jt�O������&Y�iȖ%�b{���6��bX�'����ӑ,Kľ{���r%�`i��d�	p�p� �pP��y]�}6��bX�'��K���5���f�ӑ,K��߷��r%�bX~H���[O"X�%�����iȖ%�b{���6��bX�'�~���+�\5���ΚXF��M��7F�Q)��.�lq�5x��V��`�%�&���5���%�bX������"X�%��}�iȖ%�b{���6��DȖ%���o��r%�bX����\��3Y��ԙ��ӑ,K��}�iȖ%�b{���6��bX�'�wM�"X�%�|�ﵴ�O�&TȖ%�����R�,��YsFӑ,K��~��6��bX�'����ӑ,Kľwﵴ�Kı=��m9ı,J{���_�˫��1�kSiȖ%��H����iȖ%�b_~��[ND�,K�~��ӑ,K�����6��bX�'�����v�b:�_:|�н��>��bX�'}��ND�,K�{7��r%�bX����6��bX�&?�	h��# �!!���#�����;6Yv��j��Rm`D,qVa�J��m�7���[�ra�n�	te�&�X�l5��sԦ�)f�k�3$����6��m�-������Uḷ�Dn���	�<�s�9z�0���F�8ȍH�FMƗ��-AM�s�Y�0;S���[��7/�g�y=wj�N�',m`x�Y����u�I2��.��t�ֵ<BEU�pW��t��[hAb������d`@���6���k����Ѹ��K�޸����c���ި�a&j�5�'bX�%��߿p�r%�bX��ٿ�ӑ,K������Kı/���m9ı,N���	�Lֵ��fja5�6��bX�'��o��Kı=���m9ı,K�~�[ND�,K����"X�%�罐���,̺�)��jm9ı,O~���ND�,K�߾�ӑ,K��}�iȖ%�b{�f��ND�,K��w%>�5�F�չK�jm9ı,K�~�[ND�,K����"X�%�｛�m9ı,O~���ND�,K��~�}�&j���$�k[ND�,K����"X�%�｛�m9ı,O}�M�"X�%�|��kiȖ%�b����ʟ�sK"me�Wj�fDء�:,k(��J\xy�.�8��'/�ZX�[��^�7~'�,K��~��6��bX�'����ӑ,Kľwﵴ�Kı=��y��ҝ)ҝ/��t����80n�Y��Kı=���6���F��R�5K�b�M�@:g � j����%�߹��"X�%��}�iȖ%�b{�f��ND�н?�O{ڷMQ�u|���/Kľwﵴ�Kı=��m9ı,O}���iȖ%�by���m9�S�:_�O�߿6;.��r���ҝ,K�{��"X�%�｛�m9ı,O=�M�"X�%�|��kiȖ2�)������+�\�g�=)ŉb{�f��ND�,K�~��iȖ%�b_;���r%�bX��߸m9΅�^��{�?[
GRU&�:�P�ٶ,��i�9�@�T٫�m��`�(��kC0�Z&K3S58�D�,K�����Kı/~��m9ı,O}��6��bX�'{���iȖ%�bx{��~�1�Tm�2�t�t�Jt�K���ϝ=D�,K�{��"X�%��~��m9ı,O=�M�"X�%�|��B�@�5��t�t�Jt�O�>��<�Ȗ%�bwߦ��ND�� �,�D�������m9ı,K���[ND�,K���f��R&]d�Ѵ�Kı;��M�"X�%�����iȖ%�b^����r%�bX���p�r%�bX���K>.��HSf�6��bX�'�wM�"X�%�{�~�ӑ,K����ӑ,K��M�6��bX�'�>���S/�oPӤ��7j]�����C[aK�D�MLH]�q@���דL�l#�����ҜX�'���ٴ�Kı;�~��Kı=����ND�,Kϻ��ӑ,�N��~q>����U�J.w�=(�%��{��!���,L����ND�,Kϻ��ӑ,K��=���rt�Jt�O���F��X9�t�%�bX��wM�"X�%�����iȖ>�2&D�5�ٴ�Kı;�~��Kı=�!���0��)����r%�bX�}��6��bX�'���fӑ,K����ӑ,K���6G2!B*X��.T�����Ba���(�cT"E�­���UM�E_���}��rm9ı,O{��c��6 L��t�z�z���{��O�,K����ND�,K�N���Kı<���6��bX�'��_O���Q�V�0ͬ�:�S��5��]��v�v��Y"�Q��Vۧ*��g��Kı>����r%�bX�w�NND�,KϾ��iȖ%�b_{��󧣥:S�:_�?~�D��iL�/�r%�bX���NND�,KϾ��iȖ%�b_}���r%�bX��~�ӑ,KĽ�L$�|j�d�LneѴ�Kı<�_}v��bX�%�߾�ӑ,K��{�6��bX�'��׆�|�н������t�eVQǉȖ%��D����m9ı,O���6��bX�'��׆ӑ,Kƻ�<����G)�r��Ҋ�����浚�ӑ,K����ND�,K�J��_� �'�����A'�w�ؒ	"E_��*��� �*��TU�
���@U�����QW���P@����F"�0R��"�B"�0Q`�� �"( ���(� Ĉ�@��D"("("�0B
�1X� �b("(��QW��
���@U~@Uj���TU�
���@U����PE_�*�h
���
����PVI��sݷ����w�@�����d/���3��� >ٳZ�)���n:�v7ckP��wuYN�� ���{� U@(U*���@*�����FB�
�@ E 5 G����>>U�@h�><��va���t
v	�:�}'���  �@ ���|;SZ�C�u�}��vzuMj�Ux}UG�kAU��uy�Miɦ��u\z�F�kF��Wǳ�ܠ���}5馺=���!���t����Tm-%K�p
��$ozxW�M:k����½{�V�3���c}���^G��(o:k��C��=�<��T���V����Z�MpW��M�{=+�^�C��s�փ�>8h(PQ�p��P���{�
{>U 
P����AOMѽ��C ���{���zn��$3�-�ׅz:kA���
�{ۧ�Zr"H�    �i�FI*Jh�B��i�S��T�h�       ��R�G�)�4�ɉ�ML�42 O"�TԌ       D��CA4����OȚ=SOP��S�MR"���@ 4   �> �>Ч��?y�
n/��ҿ(������k�� ��PU>�UE_�� ���?����-�Hf,a ���EXT����*� �***Ț�����}�_��_w9������{�vw�����{�@ �@���7��g��m����ym��g�p[l�X7��m��<�ެ�m����[l�@����[m�,���u yya�����o o-�w<��P�7�-���6��  DD�� @���ݭ��w9/fffg3fcm�fffffffffffffffff`��������������33333333330fffVfd�fw�x�^e�fffffffVfd�f<��������������ŏ��3333333331ff^gs)�fffgp�f<�����̬����������������ř�����3333333333332�3'3333333333fffff������Y���μÙ�^5/1�ff^ffffffffffffffffffff����X[y������Y������������3fffgpfffVfd�b��'39���33/ffffwffNffVffNffV���������b8�332�1�fgp�wfffg3��̼�y�3;�_����p�qo�̹�e���W����_>�U'�F�"�6<�cK�h��l� l9��<Vp9��M�a�y�+���w���!�(s8�\���ڛm]�G-8't��XT)A���X�P�r۴.,L�<�3m�ְb��c8�f�v��l2�pC�1�kZ�00N4�6�Ć���RM�\��8���+��b0ĺ�[e����L̙`��&��O(���qiɬ�]�P��G�6Z\��%8*��E�uV��s(��L�Q���AH�c#�k���U�Ē�Tˣ�=ĞO>x�؄̃��l!3n�1@	�J"�\�E��P�Th�jG��qdu�8&�`��C&��GR�g2ޘRJPP`�MȢ�p��5�6�`!��Ԑ�ta̱fϸ=l���N 1
��8������C�
������7�C����� gRYI��IY֡Yæ�3�0`\޲n��53,B,d	��ޔ	3�<7���K�!<�K,�Nztϩ���n'���$'D�����NN�0a���ё�(�F�*�Q���^$z�D&��Z؟g��sS��]�Yf���_>��d$O��t��p�v�
��骂+�LJ:E>B%��\�1؁x$%�d)l����A�v#+���x72;I��w��6ɽO8�}E�o=S$,Q�۱�˸*Jm
�-��dA�y��1!�@�Û	<g�H"t.B���dӡ�%���l��Qz%Z]�ګ�\���4
r8�S\��\���|��N)�ZÉE�J A�!d!��U�ff�{37�[�<n$��`F�L��71�//��HV�����*`�xp�B� (Lpؾ)Ȼ$o~�y��tK+�6���h��Y1.��|��y=���	�p:>K�k����8#d�ܝnruw��oW�]	n�i�0��6���=C��z��2�d)���6���ɼ���A���
�B�L�c;����ˌH����ᎂ�VV
�yЌ�e��d�i1,�E�[y�x��e�{t������֬�X� P
��NE"�*B")	��5�&�Ca��0-$� @�o��7�S+$��C�$j5}Nf��[,�M%�T*�R^�%������zS�g@eT���Ȩ��-Wë횼��*��#$\�*B0ʩxӳ�e�PA�@�IK`PF��7�L0��s=;'�6�B�$l$�N��q8�����s���E�Yn�E��|�ܰu~p� ��e�t,`�=+y�@�V�����Qm�e�a(�Ǒo�{Y��|e����܎��($�!Dh�Ti�Ɗ�a(#�H0���w0;��q\�ݤ�4�h�B@�����_P]�F�,��$+�/frk4�l�+X�R%g ��]�t#.����r5������u�b�[��G6�c
��R�0��$�|!  I=��4%�s�o�{��wH&-'*fOA�*�yfh6f�����%+T&��9�
	`� �0C�A��7p@!��fC��0_%𹺜k*�s$���˙H���Y�g.�23�HQk����e�y!,#t���@�HBF��p�a�I �ňU�:�F$`�FY���}�vh��Ғ��H�E���Pi,F��;!#�,峍%��喏n��"����X��xw�1!@�mH�1$���fp�Zf��,��l���֠��no��^��HXbIRh�RE�\�"I*ˊ%����+����Ynk�լ������N!i�,���'ʓ�Y.Z֎�nqZqrE�N.m-MB��9m�r�k��$B-��K75�[i����Z�U��4a"x�#!#���āy������e�6[	U�8x"Ib�,<�K��q�s��kH���KZ֖��ֵ��-ih����kKZZ�ֵ�����ikKD���XU�\�|�M�n����Y4�SKt�ԥ�]oR �v��h�[q7X`�l��wXPB��K�s"ؚ�"��Rf�e�h�h���Tږ0��3Qw�*X��N�m�=km�rऎ��I����z��/\�=�'�7�Ό��Q��Ϟq-�*V[�s),+�ĥW��M��:z�p�wc�b������=\{���V�FX^2����z���`�]l��2��RP�Y��n��(�LZ;Bɞ�7v	�ݒ��1	�N���$.�\Ө�;Y/qī����V������R~�C.
&�åݖ	 �����d��ff[neL�&f_     [@              �C�                                                                          �庬��Ͷe��i�cm& �kj�i㚎 #��T8n��Stj�i�m���U�e�ʀ���͊�ЯJ�R6 $-���A��mU)Ӝ*���;�;N�%��%��b@ж��@�`��A��6Z      l��`���cm�-�   �C�      ��    $	l ٶH�` 8:ڭ��vv�f�i �lm�HI��lBt����@p6ؗ�}�dHE�lImkdbEc�h�@d��%ۡ�9�j�����8lp�U`��@�Z�Z�We����        �I� S��i\�ҍG 5cl� ��ւJR�UgU�v��6��jBNq��Y"�2Zgk�HM�.��i�m���Zl �j��]�b��u��.;[���G��^��ntۦ"Әݣ�5m�  ;n@�Z�6�	��[@H$�I����i�A�6�ij[Qg�o2��h�M�p���׶Ԁ�J�UP#��U�U�������2ܭ�����fͣ�imK�\ו�q�.����+UWR��H5���q"d�K�1m$ �ꕘ1E���[x�=�'���vy�C��u�v�����,�������-+�>�*�8��b'�	y �^���
�n����U�����,�V�@�����ꀕl�*��*�T�Q�KU\���.�x5̈́�[%4R��eyuN1�UUQ���3ly&-�.�8<,sM�冪��mŸ8L��� �j���U�6�n
�f��)e��6<��-��,v)^�`�n�8��:wa���ke�4. �	�V�p�h����\My�Շ$t.t$l�I�����ݎ�gA�/Z�Xvb@�Ja�i&�a"����;,���Xl$l&� �`.�&q���$���] �!6 q�mf��.�ҙZ�(�,��}{N�uΝz�g�� [@X;l�^v�&�8Z�P�mTnlF
���A=ۓ<�KPZ6��f��6j�W�GF�K��e�+���k��h�W1�0*�hE�UU*��U\���K��o�7����t!tc=Ls�D8{gD�%�&F��`C���,�첮G��v�`��N�RZ�vg,�vTegh����6�.0L��6[��CX��R-�t��QB�V1j�Z� ��~=���YyP�[l�ip���aB�a�:�T�i����@@U[@�C�0e@2�T0e@2���2�*e��h�.*�ClSR���`���`�ʀ`�Pl�l�$[y"���#i�*�N�[�{랶^j�����U��kI��f����c��	���-Ս����rGdkkr���)Ӽ')6��Md�bnv,$�i�Y�])�s�%˶r«�5Źl��1��(��a�6�x΁� �Z��X���MW�B��$7]nrC�pw��h`,�݃�\�<��Iz�6�u�=&�Z����ûlf,��^�jۖ�����D8;=�.y3L��<��Kz7Ra�;
���l<pP�J��UP<UQ[Y .���6�4F��I5oD�)-������bFn�p��y�[vy���ۮ�������b�K�o Hm��n��4��4�&��ܛ	ͻKl���:ʝ� r�H�X�Pn�^����.jƲ`b�kb�2����t@�n���+��T�<��y��/[�x�tAf�6z�j�j�8����e9#�=y���=��#ݝ��NI��$��zy��]�� Q�ێVTK�-�-RɍqÞ����RX8���$��U������͕��&��D�j�[L5U���q��[bNqɆ�3���`��hx탇c{ʷ[M���1L�g����2O:k�rݸ�d��u�}&xs��3*�F:��v��m���쉹�����cvp9�Jv��z�q[Q�ے+��t�]ҵK6�Gn� �V�R���ԨR���5´����6��$�V��\Z���+i7$qm,4�8q��"@�{ﾤ���ַ�k�l#�@�ʵm+��F����j�W7A�l��p�%�n�pkm�Cm�$m��o6A�%���)Sy��^e�	�:�2��0X�eh�;^�ciUڭ�YЯ0��-]�iδ���{޾�_�"���ٵ@A �(�_������y�Z��:q[���9RR+S��R����uӪ��bi%'rtN���#,�HH�d�'��Dt88�É���6���A���B���+ZU)"JH��$��)"JH��$���H���R��T�UIeU$RI�E$�I$RI�E$��J��H��)$�I"�H��)U"�R)U"�RU)TR�E*�R�E*�R���jI�&���U)TԓRMI5$ԓRMImI5$ԕR�[RMI5$ԖRVڪRKj�Ij�$�e�(�`}B�6(>�h��)��:��&�j������3jQhF<�H�u6I�5k���6��e9�L�t�hi,CN�b�p�&UX��Dm�
d��/J�2B �����R�M �����f���(��p��b�6=@(h����D��X�A�:�t� �P-ѥ:ة} N ҡ[\�cf��ҔAС`��Tw�&�Қ� �7��i2��,P88"�Dx�0z���N*���`�fZ��z*R���4��[X�����@�BBH&^��[-�s�����Z�r4B!b�SC�F��p�]�-���ȉA��I!��Fe"��<��@0ٕT���w��S�U]��^U�^U�^U�^U�^C�/*�*�*�*�*�
�"�*�*�*�ex�yW�y^���)κ�JR��)H�� @�������>�EXD������9񛻩5UUUT�uSF����Uz���US����u�j��kֵ{_b�(�wBRȊޑ'���=��N�\h��Z8`�v8*Kz�� N:��J@���'Q�J�!��M4 ���H	'��|��o����  �              �b��L���l�jvT�D�rmB��R�J��m� EZ�w[��\hj	z��7bg�`�� ���kmVa`#��8Uۮ�cAJ`ǝ�m�u�ڧ��!�Lu̎��l��4���z{5;q����W@g!��@9�w49#�V��n�	Yu f��Xfً�Fk,��z��ctj��Gp֊� �әњ��z�v�	v�wԶ�7nRZ�:�wD��������Ց�B�gM��p�ꦪ ns�;l� <�r\�ֶ'�'�!q�-�q��Sp�b�%r+�;	z؟O8Sut�y22�a���7�]���|����![���]07=X�vZ����n�9��g���\l\�k�� ����	�96�Z�����\�quλ=�(l����g`Q�l��t$n܆#DE�e���5�3�
�Lkɵm�v��)���C
��O���L�|6�(J`��y�.��  -�&ˋm+ie*U%��i	��j�-HX��S��I���������l�[���cvm�;6��ɺ�QY�Z��a����q�Ԛ��i���w�����ʀ��<��϶�a��U��:bGHn�\O?�ݓI��3ʁ6�w_�v��(�d*��Y���b"a��P�-�K��n�̖;�y��Ys2����31� @�k{=�W][�V�\��Xܞ]��"dș`��I��[��b�LWn��*��U@1�Zq�3�=еH�Ef08c1� '���찤��� �_N% Y�^{�&��ɏx��CIݲ|;��^�f6;v��vf�(��.�Z���]E|������@�P�V�dIJ31��.���we�2ڮ�����( B���]�m!��(�Q�� t�UTc�AUꋮ0:E���˔�R��%�d�gC`�U�F�1����5��(��3c�������)
J�0��!��̼�y�d�N(2c��_�1>>N3P����)�u�/�2�5{ZF';F�u|j�b�����r=�y�:ww|�>�~k����u�U�B�!�Ą�̵&[Wb�Ő�31���YhHdI�&m�fk\��/��iS�iQI�o
��|���@�w5<���K��<�]�_<�vR.9�Q%�+�YE�T�3�T�<��]*���;z�1�c  ��fu�R��j^��8�+{$��DJd���v�v�T��u9J�;`�۴��v�^���I�MkpbR�J�C0�	�f����t�"�+Ij-�^��[�?7{����K��aŉ30��1T���3͙�N�^G:Ղ��m{3T�k�6]�D��%�Sv���R��;z*]���^s��s��q�Q���w��/c��ʇ�N�\�{�T���l��v�AE;�Q����`�`/�)�����ą�Lb��X�m�7\��:��t�{X�iG�(Z݂�D�����T�.ʰ_<���!�r�K`��� y�(�b�]�]yX�J�/".uJ<��J��{�13W��� ��@��@���� �W�L�󔋭��yy�Q�9�+��U]U��%�jm�]�gK����؜u/T���u{�Q�(��|�c�d�Aus�DI��9`���ܪ�P��j���;ڴ^��oZ԰�����u��/ /9H��jw$��*H��;� .ո���Ü�
\��l�(��ej��ѭL�\�:8|�����G��^s��{�L��@_<��|��E���W����2��P.���(���D̮ފ�,��
���]@^��9B�n�A�P.��]��WW�^DA��@� w��w�'w��~�lW`�f�:P�+&�tpEg@e�5��wߴ)؛��NڥA���e������|�]@u 9�EN֨�bʴ^���P/{J8�@���W\�V%d�:�r�y�Z�y���W���O*�0C����}�^�^���
H�(�+��c�0  �],�v���t�ٸ$��u��9v��/쎗ۚ��A�a���<	��-���j۫Y7hm2��C`�M1;V޹w����7��Λ�;���>e55(�l���C@b���k�۠����=��wz���sy�Q�+��LK��b�{���*H�ҏy@��+{�(�bb�ȋ�R�9@� w�����ʢ��P�E�y�-GS��y�"t�$�9�rYw��)"s��.�����㽽�<b�qsv��:li�b��+������"����T�b$�"���.�^*�L�q'a��{�n�n���7|"����/{@��e������|<��|�����W�Qxd�/9H���R��󔣹�ޮ���^��"����P.�SsZ�*�V-=��uFوy#:��T�J��1�Q�x�`�/;B��(�����y�]��V���(�T`{��iODb���y�S�ʏ�P.�����Ыk��wwj��n�ffn��]��݋�����ww7v.���Ϝ�9�O9�?�� ��f�7+NY��5*�H���@�sb5�Z%^X�A�s=Op��4�!�ܑ�c3�,�ؓ�c�۱(� ^�)HĄ`C(�L!�NQ���1�d�д�%j�0(kF39�.�IAd�G�]���c�/�������>� "q���?#@� |0T�����h^��J=Q��
}���JӚJ��7IQ	B�y���g�.L[-3pN�yi���6r)�y�ͺ������HHȒ.w���`�"�j�w2�S��F���9�E>����S)��el�S.\el�S)�__]��e2�L�)��e2�L����&S)����8�e2��:}��_��&��k�dˑ��.CD�t��7�|�7Y���N��e2�[)��2�[)��e2�L��e2�L�y�]2�L�S$�e2�[)��el�]�e2�[)��e2�L���l���e2�L���d�L�S)��e2�L��e2�L����e2�O��ɒel�S)�s��S)��2�S)��e2�L�y�L�V�e2�L�S$�e2�L�V�e2�&S)��g���=|�u�W���S)��d�L�S)��e2�L�)��e2�S+e2���L�S)��el�V�d�L�S)��e2�L�)���L�������e2�&S)��e2�L���2�L�S)��e2�}q�S)��e2�L�V�2�L�S)��e2�&S)��g׾�e2�L�I��e2�L�S)��2�L���e2�L�w�﷊�*�]�A$A$A$2�L��e2�L�S)��e2L�S+e3�<ｔ�e2�&S)��e2�L�S/WL�S)��e2�L���۽��e2�L�S)��l��je2�L�V�d�L�S)�y�L�S)��L�S)��e2�L�Ke2�L�S)��e3���l�S)���L�S)�e2�L�S)��e2L��	 �	��\�&&1x�hI�I�_WL�S)��el�S%��L���e2�L�y�L�S)��e2�L�)��el�S+e2�&S)��g��]2�L�S%��L�S)��e2�&Q���e2�L�S<�L���e2�L�S)�e2�L�S)��l}�^6���q|��{f��2�L�S9�߾�L�S)��e2�L�S)��e2�L�S)��e2������t�=8�2�L�S)��e2�L�S)��e2�L�S)��e3���S)��e2�L�S)��e2�L�S)��ebm��p6���6Ͼ{�� �
!�W�f��^*]U�1f�s�s�k=y��������S�]w9�S)��e2�L�S;�L�S)��e2�L�S)��g��]2�L�S>y�S)��e2�L�S)��e2�L�S)�ϟ}��)��e3�e2�L�V�n#�g���~���$/�V$O;��y�(G��=@"�S�LUe�Aw<�<� �ﶝ�v)︖��9��b�PX��JA�����(H=�=��l�x$2����
z)�{h>D<����y~��   ֦M�ĵO*�T�v틌tݘ��S�Gm�5o�uۑlNz b[q�͝��svn�����4��`��8��ݨ�1-���&���#�Ua�w�h�z�8�hZ�D��k��qs5@�y���n \��*vv���XʏHT� ��(��� �{�0( �g�N]U��(�
Q��W���R>�틈��♬���#w�������bj v"P1{�纞`�Y,�<�O!;��kʴL��hNg[�L�PV�s�/��������ѩ2U�1N�81` ��q��!9�����t�� ���y��?�" D����S�(���_8�` �<A���.Z\& �;��1�lr c��.t�S,�t0�r �[9�3;���~|���ػ	q��4ҽ�� �i��4޻����<��w��ٝ���pw�}w��w	^�4{�z��O��1G��S2�#wS�>G��RDz�hϴ��5.��&%d��|���H�����K�q����È��#v 0�ܤY�,˙Lf�a��Ȏ#.�-a��I,�Q%���Q��fH�TD#1	�7�T�1uO�y/��D��^�ﵩ�+�F���vT�3%M��¦ D sfc��{�X�I�8	'|���>y����Bр00x� 긧����^b:�0=�1�,t׶SEJ-�%��HÎ|W�trW�ܿ|w�������������2����L0��TGwX��A�âN��G� P��1:�/o��܄kF�ޱ�����P�^�%�J=�1�uǼ�>~o�;Ϟ�ޟm�   ���Kj�ԠI �6h�W�甜b��i�*Ρ}���7l�Ӟ2�㮼���e���<�\��>֢�o�����|��d��r����[L&]{N�-d}���	�y㫗��.ܥ��2��=~��>UE�3"[=��d5,{�� !�-���Yl3u�-F�t����A%d��3�Q� v�b �3
��["qw(��x��=���\��6���p��G$�F��9 @��b��Y�ߟ5�r�A�5,eɶ2��l	D��FhD�.��2a���&F�لpg�p���U੝N���@�IKj
z&u3�:\�׽����"��� �B���)	r��������⻜}l93-����'1� �xkz&_KI4�n�ë����0�j�%r�X�6�X��6����v�&[%NNi0�HV<�xG{�i��7x�׋dL�X�-k��!t�=�'u� ������Ĭ��tW�8 _]D�$K[<kgX��7!ϑ���0��97߇C����(��:  ��o+���#As2E��|둆3��}~?�\�m&��@سk�Yl��&T������ԑ*BK��ّ��Cu���H�����p�e:�>� N
�F�G|���<� =���.U\������ P� /v��v4�&�0�$VM�	��|�^���G(]�I��l�� �}���\w>x}� 4D��(�D@w��,�.e$�ʝi��җ�{���x�!|3*�����@�Gs��t:)�LhհEf�O�y��T_w��R��*�gG1E��� ��;�nRܶ�� :���y1�]�Q��0�����+�n��F�؀9]���v�#�ҵ����m���wv��ffn�����ٻ����ww�kZ�ֵ��o{��{�&����8�`�d��,���kd�)ѹ%D���v@u�%�k�Ī[�s��E��ݤ+kBZ,Yp�l'�vTBIpJ�QiTr�Z*[��N����WQ�f�             �@  ���h�[�-cu]ݘ�!��ƮvMaZT m�'m���  �.=�T��C-T���;��Ƴ��,�[�� �PR�	xd\:����AN��m	$-�ٮKr�b t{S���I���Km�.�M�g��V��U�����C�9Zں�a,v5�瘠O- �8ɘ6�K{t�W&�;�B[�j�bJ+���9r܄��ՙ����Ǻ�;	�k��p�ۦ�R�1b��<XOkiiM��%����m]d��<�E�,I� ���YUV�[W`x��Gr�e���#q�_-,�o�����O[h��ݪ�u� �����*�����3z7;/Y,���m�:ڬ�w.}[wU�ʉt�rrɺ�����톢v�l�]t E��gU���ɹ�47B���N0p"�ѥ҉��ke� �46l�:��l�R֖g2KlK��̥ �rR�#�����h���"�B�@6�:B���G �t8@��h)�G>�����   KYlA{6Ȳ�	v�S���1W'n�/n�9Ӻ<�;^ʻ��O|���'���.ӭ�;�x��W#3můe�{;6�8��=V�+;��%n����Ɲ%޽zټ85
�m���"m��]%Gy'k6�K�w��(������Hi��/��Y
f���� B��4�+u�#�k��\n�f9҃ �y�|� ���	/������Ƶ�3T�s(s7�h�L{P�_g���}���k6*]��i�f��QZԗ)T��@ �T	nB63|c��0��C5{���!%���B :R b$�0�w��/u�L��\�D���0�Z�:;������[,4��X��*���aP��s�1�H�k��,)������H�p��k+۝<�%qWkߗ�������gd�ʪ#[C7\fv���=0d�J�C�e����FԴ �_L�iw��K�̵C���=�zE|��  
��s_\�%�J7P���gϏ|����Z�v3��krS,1��9����;�m|�[�o�����hwu��#85���MiB*2s$#�4��l��s3f;�cOLn� @)ט1�%��r���19}����PD@6;>�4g}>�ʱÄI� ��Q��7��n�|��Ԣ$L̴$2iH��K���u7�o��4�7��y�/���x�cw9�\�J�b�/����C-o%KZ@n�1��w�9]B��rf[�����;�o�e�#�}\�{�I��#":@ �y;t���������O��   �q�ܴ�L`�E�u�y��[r3�N��*+;b���Jō�ۗc���C��I�l��+@-źh�(�ɭ�n_cK��\��L*YLE�����6��RN�$�ow������0��k�\�P�&S����!�r�X?c����ǃ�����dL�S���E���7V�I{�S֛eTa*���Ɍ�b�}�8�R,��5�r������w����J�b ���@�r�HGu{ϓ(�,�M/nE�%-��sb��v�v ff�KCJ7u�,� 1��w��]x����� ' ����X��(�v�5O�yPkㇷ}�a���- A���M����'�� f8�:�8G �r4�1�̦��b���B�uG.��NQLʔ��S%'=D���y��}����~^�����+1ɼ��*��&=��DD`\�?}��(��y�K�)*����t_�=�1)� �I�s�;�{�Vr���k��pf8�qs���S.kH�"�s�7B�7u���d���Jg����k�v��U۞&��ys�3�z`H��3u}N4s�ĄS{��ý�AWg����*�tG��"����35���΂�L�� r�uyE�q ��c���(�2I��C��<O��g��6�k��*d4,2<DE�2�u;�������eJ�(�Т�N4�����/pɖ�r%�4n�� #�#��b�@� C3Wp��$���Q\C� ���r<#�[� ��C4 t!u�3w  �T�al��2
�fs3�P#DD������̀ -�[4�)m��R�^I\7 ��O���v���S�t�=�at;%��^����u!P�5�|�vrˎ��ӺŎFt�i�d¨�����!�{�i��	�����c��G,�d [�N~���H�`���|���7FN+�i�u|� v�v���#�Q�꿀���fw.��\�%.,ɫ���c{���%	a����E�w2�Ѣ x��n���Q�Em-ǵ��H2����I�Wo�� �~���\�sϏ?#7x}֊��Y��-i)�Ŗ}��	U�6܊�Z�YBi���V���D����@}����rN
����O\�wyv9�`#���N�Hr�>���;���]��I2��
 ��ffO+wW����8��=��%EY�`\I�K�"��X�b��g�s���3s{΂\�)n������@q��fYa�hv��s���O�6�nn���������݋�����wv���ݻ�����wwsv�����&�uݮ��m��ե�JZ`�
b�ҥcٖфd$c�:y,�4H=Ӡ�u����$M��|��{w��pֱ(w ͢lC8Qu�p��n"�N�*Ʋ8V�ǄeĐ�j�\՚5E��B���
���P m<GHQF�O"���uKUٕJ�z+Վ�`�|#�Ǟϳ�#�Ù�������~��|�������~���6Q312\����3&Ar
n2�Re����92�ѵW���>�C�&X^���gz��������V̬�y�ƉF�G۹��m�$�D���%H��p�������6�o%���4�u�4�g9z����Ȕ�r�`ʽݬ�ӆ�2��M�s��s0���O!�̻��{3ʆ;2��j��39s�kdL�{��� �}���������;�����`  )�`�g)Ul���ܫ �����E]n��y��_���Yep���Mb%�wU�;i�j�b���.d[����Ä'u�8�r��=:��|��YmT�{��p�B�l�E`2��'��mN����eI\�U�ޜ̮��D�YC�~���y|��{5y�D����^�%6��{o����ӗ�eJmf�0=��y���6o�iZͰ�eÑs�ܸP���ۘjd:������G�#*}��9JaO}*������՛�ɇ,��9:tf̲^%�| fs�� fewtO�T�+޷;�;>." e/�jS��jͫ���ܤ��A�n -�C�)fM��ȋ�%Vo&\șkwv��Fe�Μ���N�;<��3�ګ�
 =�c��O7{�J����s4��g*�ǊB�les1�v�4�{$&ãS&�å:+nj�fAnJT�Nd���+v�'�D�2���f_3?�T3���%����HFφe�s��i)�R�e_��4L ���eKd����Ә+��즊S&T�,$&e��E��^�¸��u��?�,p��� $n�}Ѿ{L��Y���=�8�Bk�%�	���W���8bg��a���F���q�:���N�L�����{��}��#���yg�'O��w��<�_�  �+͢\
�d�Ya��*Z&g.��7���`�Lɮ�6�cZ������9N��k��N��8,�n(�B=wm�l��6h;�6�K-ڹ��!Ӻl�qd��2ts=k6�Fv�M�e�eUD�����|aR���f!���[r(�3�q���m�R\�C3�ΥHh#�� w�Ys!)q�Qg�J���������a�xźrs���=���߽]-Ku]�cv+t�H����i��Y���g�<��Fg��19�>�eJ@׏��� �6"�T>yǽ����-�1E�� ���&/��$�M47#�w�'���1]�"Rh���]1�1aÌ�[+$լ`�k��������	�Ӕ��)��cw\WTi���\�3%�m�z����\9����}��`��!ٽן(� ���.�j�>-ƾ,ν��Hr�#�A�P��&33���D����9�vcH`@K2S�T�JCNfnvn�Z6�%���ݞ��zF�Dp�g����d�*��.�V~+�z����:����#u
��t(����R\�]�1�L�;�A?�Gx ��}����{9&<�^+x���τA�s|���_9�ْĂS%�Eɜ�.��ʜR���]�/=v�-Ჱ!X�����D��+u��n��� �ףdI��wu�)Fڎ�G&�Lu�%L{3dI�n���ȼ��'ʕ)i_��;J���I9�LN~��^�n����������ػ�������wwwwf���n����Y���� �B� �#Zkd��U5���.{g_{�I�H�x����Hw9�T˔q�c0��֮���(5�vD�ӭ�3��)>o��G���8��|�uκ:���@Q�R�h����獻mm�                 �.�UP��=�!˶�N�tgk���56mm 5���`   ��u�jN�
�I�&G�u�����[� ���e����������9\u��s��͝�S7�-�=��;�jM�d �6�\�p�9�ڣ��9{v:�wk
�<�T�qZ��b�!�q�d����&����r؄q�
�ik7h�.2:v�^c��.��.�h	� 3��IP���;p��d��
�U��E�`�dX���r�t��VtJ�6�pm���� ��2d��vYocls��=���Q���h�[4�i	]D�X[���l��ƶ�mR����U���7$<�u�2�U&�BX��a��&�.�a�D�భYn��j���h���8js�R*tL@��Y�����@��hZ�s��w5����s�Ύ�r蒨�Ţ%Bx ��B�8XW i����Gw�HB�BI���
 �(?D�4*Dx�%���aG�iU�H6��P�"�I�P7� -8}@<��;ϧ��|��;���  !g^�Z��4-F�.�+��Snηc+�`R�Mwa�Tq�n��.�w7�[�*;P���E���3ɮ��R���z�;Z,Y"��9wf���w?E�PP�p�U�&�L$��td�jd3!4������{�ӈ�1�2o�JRі�n����=���ιh���q������&=C��0�0����w�9�r��w��qި�L�J`�L�azΞm�c���[5�Ys)L���hfcy��0�@:�) Rw�If�L�j�y�|#c�#���Zo�a�O��4H�G�F�����Nc����r	D��c�/�|"���c�;r����Cw\_:Ɲ1����[2�F�Ω6�v�I`��":�`e9D92T�7L!�� �g� 1��3��	2ąQ�-"�cg��������gX��}?�E���i�s�L���gt1��G��Q�d�2S��y�cC0`q�������R
 ��hi��35��^��y�����������7U���H)���\�  ��q��Lf׬�R2����qΨ�c�9#�Ļ%��J_ONf���"@�qB< ^����u����4�vt��߱�wN�����[��;l��ۊ�eWK��l5 w߬�ע�z��2@6�-�,0���^{���<`���I��9�7�rGH����8����>5%�����+�NH�A�;䆋��{��� u�L9��#��>�'w۾>�   [p�e�Zlր[��M��m�M�̵ck�҈EF-�g�*а�@��[�d;-<�G�C��:�x�N�jf��SM��N0Y�ct
�Y������,����^�L�v�)�ݼOvj2~}~��s�⸼F���-!����dYs�㍱��0�I�*4��<��Y�U(0�$Y�B�f$F[�Y"e�Zwu�=�&3�̞Ja�%�N[AvG��ed:� x�q uh�҆�n���+y��|Qe]��H��=X�Q�^Y�k��fr��V�t�ANB&7Jv������{_T�$�k�< @��zc��0��UɆ�KM�zV8F�wP����w�����e�N���۫����p^�p����J�H�����rذ �8�$�~ �\n�{N+׫��á���g���)���:!/�y�s�J������7u�7���5Eʛ�#�ձ�{��*�Z	7)$�4ړ-7*g
�).lj7hk�P�~����3c�[r��-P[�#��ukCLf�ܭjHnT��s���NfH'x3M��d��k6w��>��"@gu������X� }���;#�<������,*���Κ;vF��q!�"P����	l*��2���s5��	��e8�CH�Dn���+���|j�7���:�{τf����-�D����}��6�à�m󒐗)*�㔡���*DC�T�$@"-J���  %e���-��m�8X8*��=��;<�7\<Z�uY�����j��7���e3m����=��mV�p^�Eɋ��ֳ�'�:�I%嘮����8�$:t��I||�5#��G�5��3'd���T+sr�\��]#��4;޾��q���x�1�7F���ݜLd�*�� wm��^�[!9��|���q�3G�@��K)��/�;�����n�
�q�b�6zg��g9֖ܤ`�+�Q�j�60��9�+l8�P���	w�*@�9*a�ʥ�DH�Vc��Y�̝�%ɖ�g1�/�0��B�ԝÙ��dt�����faq��!6Q����75�b�Ms�Ԧ�s=j�VG�Ŷ&�=�u˓�,�c1x�{�|#mj�d0��}#�Q�؁�1G��1�*J����<#�q# �z?m*mUUUP�m���UUUUۻ�wUUUUUUVn���������AM=0�����\��h�ӎ)���Na� ��$��x�ӊJ)e-$*�� Z����ID�
�?	�d*ȍU�o�(��ی9��Λ�o^�H���	�,T+=��(	fVK�L7H$�kV�ğ?��$�~��U�$�
������0DVT! q��z�tu5rx���D!��,��!�&�i��i��1���Ye���餘v;�C�����!B�!�t=A��!ǡ�z�c���z�!p=C��g��}��P��}~����G��TP�ާ�JQ�����;���fs����CΡ����⻐Cr;����>=�I��_���ci����d�{�2�t܁Pp��n�ݘ�PΑ��;$��JM�b�k����Tm�׀&�xzE��q��g�E�1	r�kR�sV|)��+ �9PG`Z����s�'0cV�{���{������>��I�(;]7]L��t:�n�ͺCo|����|�z�{��'MH!�iա����<��H32��J3ǜ��q����%̖뚎��t� �C���S��q�ny���r��ʜ�t�,'q��1�c  m�`��m�ö�	5\;��<�m�����g�#J.Q�@x�g����nN^q�(8����,��^�Z5t�k��d�p���S�қs:w!�7-ۿgN&�w�����ݝ���\4��K]ՠ�wÿ}���k�  �B�x�
d�c1
�q���15�6a�
�wu®v|  H>1����E�r�����qΨ��������RI|��GÝc���wu�����*[���8{\���Dn�J�f��d��]ӌ�0�FMܤ�HP����K�bб�0�@wEBÛ�w�G~W�����4Ԥ����#��i;["N�n��9�R��D |c���}�H�^�c��2$�c7^��_H��c��rRI��bZ�V%�{'d�w.QΎ��Άf8��	�j��)6eIc32} ���Cw^�{�z'MI%�i�/�_��tŁ?��)���<�� ��Hʢ=�����q���;vAQ.RT7��~��Lx����O�?ݮ��f��)��@"�I`��$%.`�%7��Q����x7^ ���Il����q�l]��ɖA1��ݱ�wX��V-�İ�tn���:����@���hx���RX�M��!��C3|" n�ƲQ����fVZhgԬ�N	�ү⦍Q�>(����߿	�7s$sVd�.Q �j�C�c�F�LoV�t��	-�#����{1��C�5��)L�fc�3��q��!&�'D�1v��q���_;�{�3��ω��`  i[BmD2�J��J�� l�р�$װ]�#T2����3�.���0a|ܕ�U`�^��c�V���g�Չv̑�JGMci)�k;��o���V��Dr]������n�*L��D_�weƌ�|C���D̅Cs\_{ɍ1�|�ҥ&Jq��x�=�1[�ww���&m�w� c��q��{ޑ7��2�D���+��'u�������[�s#�kF��KR.	R$�RH̕C3���Ƙ�C�5���f�DDG"7�Ř�!^��3���B��]:b�� {�;�Ls�>L$�v㹅�� �#���Y"B��_{��8��z" �Dn��d��ZvW�b.��v�{���]�3*Z��1��1��+s�D�3�
7�x��{�I�צ�H&fQ&H�B���67��  �)q��2RS2���|��1��s_!�%7�Ǣ��??��C���v[sv�ڻ���4YpZGs�ue�Dl�y?Oý�g��wv��3��d��θ����[|#�D�*hwu�+���c����K)�f8�;�},�\w���D��
�#��C}�x�[ԓRE�2�N�n��i�\fd�Ln�5l3��������JA)������35��[s_!�%7ov�����\>烉�>c�Kdʗ]#���Xn���Lw���A'"R�{�W8��dƘ�� Հ�\���ΛUUUUF�n����UMU]�ػ�������wwwb��D�C���
&1�e�Eʡd�*�ۗg�q�3��w�wjB(U�|eð�P&�B�ʹ�cUP���葰�
K��]b& �pJ
�3�"P�PLJ��2H*��
�7.)�.���P��`� 'nd� t��C��zRs ��_.��v-�                 .�%a��<s�f^��j�nI�]Rً�5���Ͱ ��4N�OF��Tt��D���ݖ�nN�,� �3��) �p����P�+���-\���Ta�iq�a-�-��8�M��P�]Gf�=���R��bx�I�r�Xx����v�e��t�$rG{`;RTt9�hu��r���f�vn&�2/N]�O�ۓ�\�����.��Y�(	�Ǎ��-��+������ǤܕҒ�r��v�MT�k$�zM�d,�y:��v���hS8��E��U�M��3]C�j��[���Qj�D��=7 v.�3�\��$� :g���M�vt�nW�a<�{��hI���}�Π�x�g$u�i�v|����x�8���݃ќk���l׈b�t�b�j�s�E��c;��qs3�ȫz�n�g2^��0QW�]�]K�����YI�M�`�tO�|.��0(���
�@�U"�)Cf ~T��z��   [M[����S���+�]�&|�b�F���U�3�-Ηq{&��3��3̻"F�Ї\@�
����;��`n֘�a�z�Z�10��2�^���z�깅�7G���B������FNm�(o�y�H�q�(��&2��c$�qw�3�@f!�LQ<��tH��
���.���@>�1��&��!',�J7P�����M��IL���7�� n�LpǼ�z ���M�r��L�7"ḼH-���#km҃p��o{>����{�����ؒ�h�p��& �1��A׽>#1����.A1��]�0��æ&r��J��nko�}�4�%I0  soJ��Է1��|�Ǽ�}�8��y9�R�N�ڞ����qs2���&i�V�<b�,{� �y�ߞd�����yY�o�n�`�1�Wr���'An����@� �&���������:��)�M��@�{��c��q�a�2I%6[����;�6��7X�"��%�s7K�� ���v��S\ə2��飺�8i�I"g-l�RQ�������F��y��2K���n�bOn��5�����bg�.=�}�ϕ aS!�_�����g���SR1������V�&4�o��S%�Y�go4fn�r��c�$��I)��swf;ьp�1�|��5�2S�M�2����1�!����}����y�7u�wu�<�E�$�����n�Ɯ"`@�Y�!IT7u��>g��~�<﷞w�v�o�  ����-*ճ�,�/�PY6���v�7Uʤ���ٌcXs��?��	�}���=��N�#p3�WB^��m���ŧ1�S8�gR2���7��<����R\Xj��x�v����)�r�e&K(���N8c�C1a��� �:�Wb��a���7���S�I���b��`���.4�;���)H�K���� ����<Fy��wL��q[�6GN�kz��6zG�����K�I,9,����H�A��.�]r�;&
[��q	�{ �GwS�X���K��_.�`1:��P*���K��6w�d�U4}"T�CF��v~G�{�C� [>E�����Ln�d^��$N �ǌU��~#{�2�Ϲ.k��B&��͉m��)#-��KfA&9�b��Y��Y�쾢��sCww��F�G5�fj��<���|���#���Ԋ��@＂��E�O�	)���.��s\nn��@'��Xr$��Ѕ�'w^W�3�>~f�V�sz���l�m3.2�)̹IRU�8�u�mk��Ƴ&J��k�� ���҃�q;��$J�L��i�����kX�\�܄N�"�g{��<���*�d��|�p�"��t9����CLn�9 �ճ.QJ���Nn���q�^z�{8�d������n���z�w�b}�Ώy�E0�ǌ]�wu�f=#��aH&7P���Ɲ15����C���Q��$x���+"�BL�)��p�v�n돣��y���[��  j����V�l���=�����4­s=l�c�2�ζ�� ��B�]�LLq��MI�#u�z�uʸۀ:��MI���.��dK��F�J���e�I�'��K��jF��o��,�`�&t��#�T$H�@����Ag������^��CEĄL`�&��f)�>�g}ξ���b���g=�z����þ|������y��;ź�V�# p=}[�[�����c�1��&P.I2̂��\��yܑ(�rL���K��f�vFf8�{L�-IT31�(� �I �@�Q��'��==�R;���EIN9�\p�e���.��D��@��@ �����(��޾�)���B��n�"τo-oPR��3�Y�òK:؋�n�˹�g(�r����\x��9�����Z5���7u�lf>�&\��t�<�:�]��;N�UUUUT�n����U:�ۻ�7USUUUUv.������" ;H!`���"w΂JtX��3�	
�S(�Wd�3��3n������H�n�Z�UU_�_vA%�����t|e�]���%�`�"# ���T�����3��度�Mc��� �<^��"hx��C��/KSE R�= ��}q�ۋ����c5	�c�wX���'��!P���\a�K����Y^�v�����vQ2�H9L'&T����1�P�����%�CPJ�G�_��ɍ�L^��AmHD���/�ck�Ti�>���H�ʚ���|{9>Ot u{�j�|gX4����6�G;�sbҽCL��w�	���Ong\ۈ�ղz���m�$�%V����]^�n닱���ct/�>��`Ͻ��� ����XU��y��1�R�����R�q��4��R| ��9���D��q��� �\fc~�  �A����8�������� ��s�l��`]�eZ�a!��ngi]u�, ��u�b@�u����Ӭ/m`'5��L�3���n�3��3��J�c4S�+p�	�KM2S\�Cmӿ${���ƹ�ݰ;Rm�Ѣ��̐�ƣv�n���-vo�������|e�2]�zI���H���p澤�-�*\V��H&7B{�Q�ǀ4�	P��Q��<lyG��= ��zr1��ո���;8���G�PU�\�ƽ=�ĉ�2K��q|�f0�D@|g�3��-��N=�;�0"FșP��m���Dϐi�<@�C��Q��O��{ �,�cu
�}=;���Fm����t7�\s�q�#��Wq��ܳ2%H��Isё��ն��8Q[�[�ㅑ��f<#9�/�)��F-���fH������)F����� `O��x�s�� ��tGwL�;�Ƒ��(��)�H4�nhh��p`C&�v�#��n�rZ�G*/p�ky����	BQ)\h:E���A��"�w�
r	��|o��wXcv����.�f1��c���w��e9�,nD/?8�g\{� 1 Q󮑙ì�Ґ\�Y��Øޑ��-�]�)�S2\�Hm�p�p��=�lWV�����V�;�0�sՒ&K
�f8�����iݰ��!�����t�yo��w�tH������7E8�̑��NHI�G�Q��[�[���� !����<���wN��   $��-� 9j�jI,�P��U��G6���T�S�;;��q����u�P�Χ41���d��瞭k�K���f��M���l��Ad�Xl��EV	��^������#r���;�c��;����� ��RY�w��
�mt�=�<}���s*Z#wS��0�=�=�z�/v���,�Z�F��\;��w^��󦐙Q�������ƘNql�!�Cw\_z�f!�1S�S))�T�-�A�*Zg��"����͒0����4i��%f����=�@���j""�< ;�>y��?�{�{�
bA)E�V���N��Q��t��&[47���t�ޱ�5���s3./u��`�2�Ǣ �������ru���I.D�%���%1c���9Ln�#)Y�63���Zj31�A$c��c�V3W8� � D;/Ӻ����FXE����7P��߸Ӵ�B�1���X��n���(�$�fR-��"Sƌ��ԡ2:۴��??|}�1�\a�ӎ��L̤hf.�����Df/:wϡ$���h�l��9�;|8�%��1v��\lq�t���ÐLf!t��N$�&k����rI*XM1�,nmgGn�h��]�i�����q��_���O����<#uQʹ���=�@�|b������&���r V�f��tk�<#�\�	r5g129ޖ�(t?��|�ԵUUUUM�ꪪ��R�����uU5U��9ֵ5�kY֦�D�@bH���"5�R�ɵ�G��q!i<їw�tB
*�Ѡ�)4ר����(%���"�(`p��`�zNPd���ଙ�@����d��n������F���U�h�ԡ��R�@A&�S>^Su�NU�##Dc�0�:΋l	��8�԰�X���o6sl��L��u:����Q�d�#z�-�x�ib��H��L
���+�ܓY��X2aA�$zV�$N�\�:�q������RJK�5m�rΧ]t��,�����z-�                 :d]wM��h�"^j*@{4�B�9x����ڶ���V��Z� l�&W,cI,͊PN�	R�ٶ��%˲k0�� �\��Sa]P1B���ZFwcu��vV�핰`E����ƪ��j��л�9+�]��4[�Zݶ2;����jP��U 1{�4�.��=��~y�<�V�;�G�����L������ֳ.��Z!m��dZ�\Kڬ�h[u���i ��k�k�[���X\Jv��s�x6���\9�vlj�R�U+�r� 	��n��*���2�c�Z��z���ݵ�zz^��ۯc��z��V9z�{B3�	t�q��h9MHaMc'W`��N8;6M��T*j��z-u���rʘw��κ�q���l7*�&�Wi9r
$�]�3q�c�h�D��Ln��1�F!y�$�Ѩ8݌'1��=u]Z���cV�4�X���-!��s����x0((0���X�x<@2;Q�Y>6�	�d�~c�1�  1u�Y(m��i!5@�-O Z�Ur�������R��,&�����ם� u�@TI�
���P��.���q�a�I��-�ҩm�[�t�����n2<i�Ά;y��SfD���I9iF���1�!���ӏ�Yh58C�1���-H�G�e��U����g��7��s��:�f!=Y����q�Z`�;���b?��}��-��Y���d�ed�A�H���o�N�s����W; �$"�n�ۀb@ �����c� �M_	32�����z�Lf!�<͂S���@<�َ�E�r�z�$&It/�ڣ1aި{�P���3-��21�4-��w�m�1mɅ%*T�`����ww�1�k	�*Ӛ�G3��O�!! b�q������r]�"�{�l��mo��Hqϐ��Tm���'� ��2cwX� �dݐ��#n��#2�r�:��5ۃ�����m���hf(�8�w��b�c��%�sJ6u���s�u�Hl�YΨ}�J;��F��T�cy� ���1�D�0 �@t�&�CJ�SX!Ɍ�uE�Ux�Y�3��s6F��A��y,"���e9kŌ�8�a�r���b��MLn�1��z���̤WG�8�ݷ$��97kݐ[��1��o���(�es�)S.���=�j0Ylf-|��U�o�0��n����A	�A��y��;���v��_�  m;Y:��Z�"S<!*:-��qr%]����](;PV<9�w6�v��u�w��C�ZƤؗUb�6	�sF��O�u5�b��x�fV����n�j[�'~t�;���z޽l�sn��	�n���f$�$Sh&��i���b����Uw&6�5�܂Gmn�Y�_H���'0BE�'��F��Z�w�7�t������d���j3��q]���� �Wb���fbig��R܉�T�feU.K���b��]��n�eX��|#��9��I�僖@��� D ���$��Tt���jB	A�ܡ��}}E
�q����m��t�ɑ���ң*��Ѹ�RZ��}�v������}z�%���ٴ��6�ֆms.�m4�h]��~�>�{��&	�ű ����,��sS�1�y��9�:RK�F��Fz8� Y�2 �"" ~�ӆ�K���[��1�V��8��H�!/bdo��K���7`��;ً��ā���mL��,ːCRܣ!�۝j���r���lcߏ��Ř����;�;C���M�i�� |+��S ���ԩ�*�fc8QYi��#C� ���ɒ4�����b����5\�����\���yn����Ͽ^����1�+]��,t��`�\�!CNW�AĪ����i�J����Y"�{�Ȕ1��,qQ�~6w{Β��@���0���c3�f/7�Bs%5�q\XF�= 
��;��2Jl�^�:ΰs��=μ��
.���H�����  `�[���T%��Ʃ�ȓ
�kB�4�u���7P�A�mٶ�������jݖ´(�O�i`�l�����]ك��Ң�Ŵ�k#�{�݈���U#p��K��a�1��;M��h������Nl�cH�{�4C)=��<�!�t��8����8��{2q����Hò�W�{ɑު>�N�Z����"ct!t�3t��s��L̡(�j
��,�qB�u�0*�L�la��$a�����D� ����S� �G�(���a�g��
���u�;�3ޡ���bO��[-�$Q�C��svG��]o�hn��tgr�I??�t�ߏ���+��e�K���1a���HF�`��� �������o����A����dk�RB�ƌDZC�48y�"�}� �$"c��#�Bk��ުu-UUUUSl�����T��n���U:�����7wwWv��
�  Q��%�g&�zc��F�Г�k7�
�AjZ!VYQc 4E�Zj��@N@�S"b��Z�ݖk���-�|�z���6u�Z�n�5�ͬX	T`��OHBQ#���p�tߧ�t�S�H7�����<Q�M�J�(w 0P1�w�&^G��{���#1�O}n;�`d[u	�gϨ�婙�{�8cw]����W�rRi'0e	�l�I0�8�L�4]t[t�_;���Q�� #w\z�|�iH �y��c�
"��0�h^c�빌1��Z�cUW�k�-�)��=T�D���A(=:gN�w��k���z}�����1��A�>ː[�fT�@��.d�8m.,ŦPҪim��~~{(�(9��c3��)9FK43 G{�zA�|� �é���s2�G��&0ǩp�(�wBm��пZc�C-Ff8��(��C��y�[~yoc��K��+��   �9Ibm"�R�[<���ϸ皰�5u��uB���������eV���"�-읂V�T��g��q ����q����x���ظoC��k�N��ԓ��_^z�2�Yn�PI����\�TP�c�uE�ƟR�H�<��Jh����n�ޯ@�>.��Y��WO���!^��bq}�7!�U�#w\��39���A���Q��bN�(a�ճ.IE�������v�qnd�J=v'�q2ڍ�q��w�����=	�32,Y�.G$�WhB,�"l5�ku��щ��f7���R	��*�fq�YVXl�(�1�<�\i��>�k|��d����1�M��Q�U�����Bf��I�a\�k���3)�<�����>w�><��Fw�_�$�$"�����Fc1� P�<�)9$�.��"D@��Z&5<���v�{�V&%V᙮8ct!�����S3-��`#��C1GϿK>�z��GUt�9�ΤK�*̑�R�P�ND�2іA1��Z��xt��8����(��XG;����3�5ȖJ��qf3Ә�3�s$�mR��4����g� �0$H�6" �-V�z��-5 �wC�w�/��Ƙ�ɥ�H�°��k��m�,��p'!�$��HV7Tr��;�rt�"��'�qd#�u���FwWq�32���6Ak�1FVdǬsZ*A#" �/�75�ʠ�d�F��8�:��s����C�t󧳺N��m��m��` �-��Z��H��Y�c�iD�#�ӍFR�g�m��ۍ�D�1��ݓ�vk�"�s�gkqE��ś!�c>%��A���3bµ�L�R���[��䓡�ԝ������r.պ�t��l���b�-�Y9�zu��1W�!��C1a߸�-�)q�XY�P�U�1gdU��Ii���Aݸ��+U�\n�i)9 ��a�z�Eܖ0���r�q��1��b����o�)���.���˪6��K�ױdwN%�2ԙ�*oON��JK@F��8N���=��,=���9dB?@��#"���h�|>���3?T��[%�|q���$HFS�ӯC���CqAw��%�d��1�q1X�k2z~���ӫjI֒a:Xh���]y���u-�+n�;��=x���俢p�s9�d��l_q�9���C���Ub�WO<��gvy�p�_"H�Z�/J����&[T��Xsfu�ݝl���kH��G�����(�8��,�O�GlN�bDȐS4fJ67T_&4�{�GM��"T�|�n���߸���)%+�#�|C�Q���X��d�̂H��ѬS����E+Ib��S��OBE�)
�.�ӄ3���3K�+0��.ܝ��0v�D�b��&�naKRQ�k����L��5�,�����n����P��YA9cw����3�n$����p�H*���7\r�����&|�"fBq����/�y}�<��������)T��6۔X*�/�}�,i��) A�#3_������9�`���(:����a�`��0�g�1�m�m�dbm�b٣lŃm�RY�L�c4� �X(��Ĉ�:`2$Cpi"�AV�+�3*�RF(���*b(\ �^E�-�l#6�6Kc��0ۉ���=6��7y_�`��c��dE� ,�`j���mg��^ !���OmE?�#� 7���َ�m��a���6��ُ���� ~� ]���|����w�������V�`��o~���@���F�TB��QE_�'~����A?��r�����8�AU�B�����o������R�x"?�O��������W���m�#�g�6m���������ae+@R�����|p�$g�F����Q�Z��p�;ۍAQ�}?���MC���D��~�g��&4� �F�A!�U+m�1#0���V�6m�6����f+Z�[jm�b�fQ�jVج�٥�ڀV�jd��̈́�lն̖mkQkSm��m���$ٴ�i1[j)L�Sel��նKm�clP�
V�$�VfV͙,0��!Y�mM[
�*�C
֭IiR��/�͙�&jҥ%F���Z�����V	SSd��m��V5m��6��
�7v����lZm���X[k-2-�2,�bͦ�m5��?T��
��W!Ɍc�����C������U _JCp�Q��?/��?���?p�=��&ކ�B�����?�g����O�AE]������~������������caCFA�����Fq��a��O�������_�}����(���AA��k����	?��?����u;�(��I��*�'�"(��S�?�$>���?��O����G��_����*�*��H�$���ϰQV��?e)�o���QUQO��*p8����!��D6iQW~?����QW����?���QP����������,_��*������d����'�����E�C���A� �*��D�'�~������O����4�0BЏ���A�.w��8����1�?f>��ɿ�h"����/�����~Y?/���&�Gp���^��e?i��)��O��"�E_�`~���_ڜ��¢1�wJ"��S��?/ʃ8�j�������+��'�B#��w���H�
$i�`