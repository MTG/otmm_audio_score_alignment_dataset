BZh91AY&SY��e���_�pp��b� ����ap� �@�P�$�E B
�EU(@ D P�(EDTB�P���U� x�P��P�QD���$T�*��"%T���B��JR�TUH���BR�BPR��
���R�A .    1�    � 
b��L�)e��\�]k�R��= 4}��>��,�f��qiK =ip,�����  ���B��R�� �*��P�&�U��:�VZ�T` 6�
��U*�R�LڕAVXU(�� �     � w[��S��W�;��q��w��]�()gr��j�6�z��;ٯx�8s���*�w�e�b� �yΒ��7�Ь޽�ݼ{W����q:U� ����u]�n�͝o]�]�[��
   �� g� �o�Yss�[�w����z�p �c�������9�����{W� ���������� }o��/3����x h��뛯y��������6�� a��Zr��^����x�vU8 ��     �� )x}8���g�������e�n�8��Z���q����x�)���oe�{�}}r�e����Tf�6�� 
^<���<��8Y�:��{�S��}|�.�,|Z��ʙ��� }@  @ 4 70@����|������M��t���y��A��ۋv���#;׼�c���so�r��  =�o}����Ͻ<}��Ϟ˛}�rǥ��Ϟ}��p u�����#��ϻ����콗�P       �z�M��J����4ѣL�����a��D�)U  F  `�~=U*S�L� `   B'�T�#�J2hd�Њ��3U*T � ��  B�R�41#I�=#F��jmL�F58���?��j�w�����_}������EU����(�� US��U_�
"��@�(����DU]_�/�������DU[�����������?�Z4����Na���$�ͥ�����on�2��y����׬�s�:m�K���y���j{H�LVYy��ޝ�۰$�*I���a�GfķdW��"��h�2��a�c�"kWFhA�#S�0�� �[ѹȤ���.A�q�M�7�=�Al�,4Y:n#nؑ�m4�r�(�Q��(��7Ef�5b�4�XK����$���ԝ�3hu���f��͝E�Z��ЗBP��h�&��t��By)BP�	Bu	BP��d%)Bj��7�fó��t�fF�Fh��<�Ԅ�^)���bTͩ���N��S�=g�]��j&��X)���ƢI�ЮG00LPȔm!#M]�̜MZ�-�0�jb�X��4��]��I�4�����!�hLPQ"	����i	��Ƴ�h�s䉆3b�B��4��$Ѭ���bˀ�
D%$U"��D"-��V�\xc�Zm(��l� ��\z�[������sx5�	���E��u�ƈ��thgI�tv5��h�LѨ�dΌ�!5�Ĥ���Gs�lﾃ}`u�Q�s�[�pkF���rp'�>N�螴��j���7mc�q=5#@��Em7��Qje��)\�־������ߎ�O�F�N��%	mp�Ȋ��];�Ge69�]��z�iOiQv]�e o6M)�\1�ՍA�`Y!����j�"H�ypk��Es$1o�8\�B��䫨�~�ƺ��r>!�*H5��$Uk��ˑͭ������7�ox�Q�H��2	1}u�9p·��V$�&:���[[̃�[ֲ�
�5M)��|]+��N��-��ј�K�$]���WC:j�~ͦ��J-	1)4��"]X������'�g]��)�L�Pw&A��]�Z���]�yb�Ek����CSx#Ơ���J5>1�Lxa��H�*F8�&��1��Iۙ�9N$��o�	�F�֐��[.������E�&��u
,�a��L�w�"O6��i�MES5V9���|ERִ���;�	��֌�������Mp�(�)v2�Ũ���BQ]-��}�N��O��;U3i��J`�]��U�D����r��$��;6>ˎ�
�2���7ּ;z��k�}�4;���[������u	N.X��fw�;F�*��ܠ�Mj�:�Z0:=�2��rt��v�f�#�׮�/#7��ѣ��n݄��ԨbkJ߱���Zw)��Y������J�-.mu�p1�{���ޝH�ȏ�i�{���v?�����.6������Zz����Ƨ�.�h���[Bj�jpV������-m50�5t' ǃ�H޸p��݃��T�əT3����w��y�o�m��߆&�)��	A�`�^Xhr:�5�5!���&�'a����iC�ֳK{��^�n3A:�(3���A�0-É���F����i��֗n���ε�o��0H��yK�y���M���e�p�J٩f���x�6G�AH�ԜKH�cy�5Q���2D���}&Z�gI7^j(��1邃z�Ʒ��u�ޚ��d� �)������-�,�b7˽30bi�7'�[�V��+t��N+����v&�]}��G����HzܻF�a�M4�V�H�h�����h�-��L�h�*$�tI�L����"rC3f2M�C�!8�Ȍ�P%E��*ziʐ��*��&	�ɂcѡJ�(�LԚ1�IjǤj	پ`��\[J�1����U-	���p�ER��.d̜�#V����m���c���	~�	5TX�f)�sJb	>�J��D.�>�5�mw�Ҏ�.$o�C���BP�%�A���1���f��^�ב��0)���Ԩ��Ѩ�BlS�f<�T�ϑKQ������n�j�(a4c-F,4đ��FNkV&��
����°��SZ�4'�'��o{��k�3�j
�}i|bc_}��Wj	9���(�QCB@��.�!�]���z�N[έ^{��<z�)�c��Z�hK� Px*o[3�������k~�A��j_`�ޡ(��lIT�r�-	���QǊM*�Bk;��5����CY��:�j��X�QER�ȪT�cbx̹m'r��pTڥFl{�}�ĺXl�,hѠ�L�ыfe�� �A�,�ELy����9�h�3ZYiL�5(cQ<�ƣ�cRر䄿-q.��PO0܊�mk&��B�$�SZ�'V�Nםo_/�K~���ޖW�DzZШ�Ћ�	k>"����5�	�L�(���b�AlTj�����)���U�A&F���� ܆1��4a�NZ���6�(J0�߻�^M���:�ѱ��a�Q��V�&����gn��r��T�9a��5ԘK�d�.� ��02l��ۡ�i����q��l�tkA�.�A���Kz�n�#�;g�֫�DL�����mL���b���j�a�4�������g�ڰy�\$B�<�Qd�2��Cl����O�f�B��PJ�I��]C��sQ���H0���N��*����w��iA|��$oKLw��;-�Z�#%�`��Ll�bh�HI�whc��r|����w(�B�Z��c�.�@��i��m�^'8��h��Cڪ'S���M&g���;�j}�7��ɨ��	�N:&(�
�KI�I�	h�`���I�c���#���&�$QQ�U�/�ސ�����YML�����̼[؜�ȋZNF�y�����OcQ%��k��!�,�<�1Ωbu��4�sm7E��`�ī����A4��Τ`b1A5��mo9>�V�ʄ�1��A�E�9𑶶���uH�cFkF��[Ȣ��iW�w�I�U�����.�[��Ͷ�����\���𓸜�M�'�Q-Cq��J|ce�SB��b�6�=okBsSB��wXH����|�F���&�Kf#KCF&�]�5��ff	v8���1&�`��LciA��hH�H;�e#an�����<�n2q0Js�:�3i��TN�V%1Abi���pH2(������Cz�֦
]
6���F$��L�.G�2d1<L}4����XŊ��l��P�np��o>Y��']�:f�|��n��A��x�)BWݥZ��3A�L�RJ"H*Ln��i�	����M^��>�C'}�:\��(v�a��h��Y�~�8-Xޱ�Q݁&I���ٙ��X�Z�,Z���F��Y���`�ve��ڇS��4k3�5�G�|���Տ[�gli�����2��~�$���>o&c��ޙ;��hƑ� '
�f2�4F�!�'a$���!��&�KԄyw������,���� �rq5j\s#�N����1,�=o�kg�H��'$U.�%�C�F�wX�&��ŵ4��ULBzH؜e���4-*��D4��	1��(�\X;tp��+��*�-�|�g�.�ժ{��{�1�,����F�!"c��Ťo(� 4i���!�2�<��<2�*ޝJ�c�̖��������K�3�zE"2!ŵ�9�qQ1-E��9�\I�hI9{�}����1�a9�]�%����wJ��w����ƷV�U���k!ie�u��r�5�Xy��,<��A:z�q�ѱ�=�����a�.��c��u��jO��$)$�����t�5	Bm6��k�_a�"�(b�bآ���-W]�f��Nw8h�7���������T�(f5�%�3f3QH����1�ٵɃN%��Pk�H@�1<��2
�`j7���y�fl�����|C�j��+�u�7f�oOpuh��zH��C]X��0�ա�V1i�o���c�d��|f���؊ګX��/��F�K�ncq��4��a3�;H�z϶��^&&�2N��.��Co|g{�ޅ�	���{|Z�c\�,Z�B�FH�/���a��Sfq}��Tl���I��Ȩ����4T%2U�0�Ħ�[҉Ԍ�IoKy�A(��Q�f�4�(bj5HE"A�%�Ϸ�&� ����Vޜ7��w1���]�4���lk���
�����5��6�GV�u��*z��:0�lJ��(J�Jr�&BP�%���/3�g`A����:��`2�\���=��@oR�BS���������)q�Q�2�!��4�KB��y�ǥ�$��N2&r���BP�0GG��y���p���i%��,LDZT��Q���J��ӆr�Q<U(�I�=`sJ�M9��8�[��I�UК�HO&A�k\삜]v�ͤ���
p��dh�=V6j�$,��9Z�ۑ5n$�3�/����Z�$��_-.��*�qT�L�H������铆h�ݢ\�b�j('�����$���kN��&��̓��3&waLZ2�f����A�E�p��[y�v3jLL���
�����f5��G~}��u��Z5Bdɩ	�Fw�{�렝��������g�؝e����a��J;�՞���MJ�zB]ϴ��⃙�b�(����I���ә���=�O$:�1z��Nü�t�'WK�c01۹�A��}t��D�d�&$���7�ﵭ,Q��ֺ�	��)1Mi���Z[J�A���vy�x|z�q�P`mZ\E*x�2$	h�4�1���k9�$�}k�Ә�';�o8�5M1o�����3N.h�aa����qDК}r`��-)t���+ͤ҄I�2�Z�ǆij�������%�����}���nj��d���K����[I�ߢP�����5j>0�I�C1�1�α04�ҚDi�tI0X�udN�$⢦D#����,5�Ϗ3�D���#��ܬl�kA�u������A�GO����t#W_-��D��xswԠ!hh]�ǏpS'�|���W�����[Mc�iAqER��պ������i�i ����� �Gl����A)�#4gs;�T����b�`h�,�q��{: ��_@�$�n5�����;�i���_�~{��h  6��` �         �`
P  $� }g@h� �[q�� 6� r���Jm ��m� )@@ݤ�          )@    � � $pm�J     ��`�p�V�m��M�j��� �6�1��V��*0�f��\�T�ҭ p�m�.���B�'VV�U�jV��IB���mm�mtm�  /N�m\9^V��lԚ�J���\ i	���N�n UJ�N�YU���i6  6�9�V��� �j�f�T���,Vp+z�F�
�j�W�UvZ
^�8�*��m��s[U@R������� 	�x�@J��U[��v���9#�s;X)�1�=EZ)g2�jۗ&��#m�P-���\�\C�m%��%���^^vZ�����{B�6Z���$ M����V���jC��ck]���� t��	�jZl$$�� �Mn� �z%Û�`��[i0f�jۀ�]������2팰6r��� -6H-� 8Zi0-�Ͷ��M�ڒA$��	6Fx���m��KS����5� �5�6�[��+�m���� -6   ��pr�[u����������L��띹W�s T��]J����ζ��*BCe�҆�;j��6T{WW�@��{FŌӲ�쪵UQ��P��[g(�ow��GGh*�.�)YV�b�8kH�lH��8v�d�H�i�ؐ�nk�8�mmm��ŷk�n���#K�	�gf�V���  [[l   �����@�&ٶ�p$��媮�"�<m̶�嚩_K�qc����&�����l��ݺ�l HK)�[�J�� ֵ�pYɒt�$�q:pp$�I�[R ��m�`jZb�6�L,RB�ڀd�m���f�m�i� Hfֱ��||�TT��նͶ ���v8m�3�	���mSJ��k��I�is,06�A#���u��,Wm�e� m�ڐ� 8  6ٶ�mn�KCm&)�i-�����6ғ.̫�9� *�I)�I�1uUR��mJ��J��V��Wg���h殬��-6 �]2�'n� 7&����J��q�����k�V�' 9F譸����WM�d&˴���|vm��-	J-6��g�K�O����Ź%���@��"m�����[�k���zt�<�|��9 V�J�.����4��t.�L��n�����t��Hr�(hV��P͆���ͫL�evgg��&�nf���J�vI�����Ib�Ö���!W�GqsB�-�Թb�AmpQ*�U��1Z���'O'NY��{t���6	V��;m�'����F�j�sˮ%Z���T��gB��K�ʪgaզj�"'hfC�-���:�&�#[4���v��%�� m(\�P���j�V�G��v�i�$��ce��p�R�T�JJ�#����*��6.�I0/^���&m�;l�6�bG �R��UPF3��U�y�nBBj�в�q�UP�(Q��UmJ.�8���@U�(�VV��n6ٷ�zw�$�� q��ٶ�I�L86ݤX�` ��  �-��5s�qJJ�I�v���鴂G;m�B@e��  
������3M�-�� �<kj��԰e˽!�^Z�a�b]�U�;U�R��J�����K̽e��wH�^j���3 ��f� H  �'gF7m��l�n�sm�6��m�s��H����� ԫ�\a�j�%�*wU[*�g���X��e��kqgj($4[Ivem�j��dm#.�۶e� ��)Uv����]] �P\�b�v�I����$/Cv�%]zڶ�u ��P�.�^ڭ�S���Y}���}omH^*�ۢPo����8��a˰�}�R�[@8���-�m��4�ۓ��=)s��q�+]UUr�\�*q1��ezL�e.�R��U*��R�Y�����>��S[v�Z4��ʹݷ	����8��!UBٖODWe:�X�x�s�-x�V�J��*�'���`�˝�rU�Ʈ�iL�9�A��nl��'B��[[*��M��]�k�z5�B+�š�/e�����I�pTE���ݴ��&�&I�,i8 -�^�r�5�U[P
��@2��@@Uu*�j��#�pԨ�6��=K;[R:괲�Ups�[�U���eܙ�~= 	km��jGU��[J���(i*��ٗfM���V�U�@J�*Ʋ�c���I���[J�R� ���5P �L�	 M�)\��`�;r���*�����m�>��n �������;]�;[*��6�vI�y�V�t0���D��kj�b5��2��5\q.���FvUy������.+n�p���v  ���U��P����4u��7hV��h:�#����p\�H��	��d�@�[%	9�lZ�b�mHM@hH�R�$�m ��$���m@T�ʪ�T�P!�sd<�IZt��A $CZ��m�Æٖ�5�n3�/G�VVw/�T�p6�ݶҝ���d�m�l-�!"� ζ*�P˘�B����D��m�$ l8��:��i�˭��b�f�Wf�j�U��H�%�T�h�撐:E�@۶��5�J�mR�����cGU���ā� t�Yj��[`�?���6�[x�cE�-�]�	�|��U�[�@V�KtRG6H� ��i�Z' ����l�ۅ���p� [Vнu�����8�nk`([v�`ai&��$;K��U6�u�A�N�v�d�Yzt�HK���P>���+�@�Z�*��YKrP�P Ԭ�;` ���n�� 6�m�L����l��Hd��ۧM�^���,HV����m�T 0m��$�C��n�Zy�p Hl,�	$ m�[RH��:i1ĳ�}=�ꪮ���66�.� ��h5�fLm!�Ŵ%�lzJ�K�u[[+��J�R�i����n�ZK�@   -����V��ڧP'WVҮ����^�'M�-�{5UJ��f������yg��-�U�R���qli &ҭ�[t�T�΄Ԣ��~g/?h�I<mU��J��zdm�t�ڳ�K��4���8� 9���ۂ�p m:�Hv�8 r�H:hͰ�I�m��R�Z)T *��1��wl��l���Ok�A���˴�'
k�����,��N�ں���]��8�nًh���  o��JZl�y]���.�	5��m� ���5�P��F�f�Q[d[���h [@p ��*U�okj�@j�j�(�U�U��X�Э��9��k����M���M�e皥y�l�(l*�9�8�<�;$�PQ\��ⲻs���-m  n�I [x$X��R ٧kp��D� �[-���kvإ��ؐn�v��n�[^U�eyvF)�Z5U��c���P^MulX�l\��wh�`��TcR���r;hb�ɖ�V�I���ir�u�    l�*�-Ғ�[_+�}ml�  6ۀ$�m< �-�cm� �m�ցm  6G;:@8�m���l�v  @[�� 8�j3��*��U�mlݤ۩y��N6ۀ�  [Cm�u�4�p�,�5��UT�*�R�m�ͷl�I�6G0�I)$��m�o![.�<��u��m�;:A���+�TxM�����k\ݰ�l�Õ6�&]{I:�8J�mn6��A��7C�Z���j5$[`v�T�p�n6�K֚:�-���[W��#��],��-��mx'@�lmZl�w�e�h �ܽd�f�H[u�   �.��Bl�W�Xb�;v�&N��6� � -����f��ɑ�ꜥP�Z��rͭ�� �ŴP�W�����uJ�UW�[ph	9�m ����}����&�C�fvL�����MJ�\T;k���u��B^��Zl����  N�!����  ��e��$�bM��  8�� mr�8��v�̱5��n�m�@
�Z���HJ��5U��$z�p�ǡ� $6�N��6ۀ $[x嵶�I/c��s�0 m��	89  6��X�F�i�-:Č�l ā{Ml�L -ɰ4u��	������V�vv־m�rB@i6�Z  	 7j^Ȧ��S^�*�V�:�$�ղ� 7;e��"�:$i�mq��:����q���<K<$C6��Y���s�/Z��͂ۑ/%�MJ�ڮ��B�N�� 6[��Ȑ�����).��/I)@GV�W紐5�[�oN�6��6���#=��Mfp��V��G��6Ͷm� �ۀ 8-�l  6��k/XhնM���  p  m �N�($�pI ��M��*�i]��V��5UT�:�Z��b^%�Z�K("@$ $8pm��u�t��`6�$ �`6�`����vY[- �`@	�[�l�� 9 �f�`�ym� �����m��kjFH��YN�GX��(�WB�3t������"�����1QU|�}�����O�����{����H����q%?ء��ҽ*�����Ԅ��`x���W�Gi����`#�t����� �
�ӳz ��M���]vȢ�i��: M!�ҝ��>�ҥ	3��}���EO��E:7���Щ���U�P0��~}� ��
�">�����5���? �x���i@��A1�`h���$�x�H$�Q0��)#"H��K��$t�C4
��y�| ��	��DN�|_ ��W�P�+iО�I���=��J�U>G�U��UC��C���G�i�G�6�>"?���l@>@�H_�К	^�P�N��rb�P��]x�
�'�.�� ���=��|"�����ۢJD$�(C��R�E��%	)JT��E��IAe�T<T�T�N�G�� �@�"$ J%"� ���B��!(&����A< � ��S�RIR�%!�� U{@��T�H
� v��=a�'Jk�����DEU�#�O�g�?���f�(�ǵ��YQ�"�Fm�V"HCP��RL�?��7��qoy�����0a���o��]&��hZ��  /Y5�� p���Z��G[7,h�Bev�%�29˹ͶV�{bd���6tm�C�.$ΐ ��=��`��6ez�����t��f����"�xc�t'A-�T�Wؤ	��\�� K� NM��nm]tl���;E'[��k��������v&ij��Q-we�U� �&t�j�W1��Pm��#��yP+�Ƿ^��h�����jZB�=7S=�'�Y��xJ���t\í�O<:N;�r�gV3��v�
��۩;f�C���.��[�ݝ[f8�=���D�n��}�^��"c��&v���NÎ;��:x�sɍ��݉�.S� �A2\X.r[S��g�7H�ᑀ(�Tvzs�Svlhn�����T�1�(fɯA��b�Íb.����BX�K̃�v�-�}�S����u��'1��T��"Ћ���Z��6�q��V4V��h����+p	t�8\�0 ��c;]ղ� �/d�1��m�hm�D��V�r]E�e0'�q��w�.5�ZIn��M�ll�Gc��l��v�I!��pj`C���܇F ж�]c��1��H�[Η9�n 6��e�+waH1p�E��Ԉ�<R�(���t�'�F�iU��s�Af��m�[UR�§(���y�� �9�[ɴ$	AY�Ga�^�� �Q� *���v�8�nV+�1nʦ�2�Q�m�i2�ئ�����(�erޓ�R��ui6��KXب^){/+�t�-u�NT9�(�\��)���{eX!�%�{c��]m\u��y7�Я1ɝN��ō�uf_m�A�Ʌ6j��E�Y���x�Hgv��2�Q!]+��0<ԽNwm7O�^�a�J����gd:��p'b؂���8� ��f7Im��\n�9evݶ����k���:f�v�k�l6ư����FE1��ݱ��/&�z쬭r�����gB��9v����u��ۭ�a��xh٭�ֵ��TO�T�V���$S�'�lQ�� :�D�C�&���*A~��� �a~����~J��咲�����x���,	[D�fꥊ����L7X�e���vöMpk˵˭�.,���M<aљ�[ �u�Lv�86��Y6�&ذf�����*n��pY��d�7t����js�n�����Q��N�nmu�{�����m���� ��805�v���D�j���V�[��$J9;�P����G:t�y��"Z0�KmQ%��Y�.b�+ԘӐc�j	�<pd�0R06ܻ����E@9�<s�@�n˔7�v��rPs�_٘�m���,\���K�QTUU%`��o��d<��{�ŀo�����p��SE(�D�I+ ��V�z��3w��f�+{���*
���L��=�����7�Xn�;�+�ڬ���V�9�;t����������-�3ӝ����dC�qs-���sQ��=��ٱز܋#e y@�1�D-$��ir���\�`�}t����uŀo���F&�UH�J����[�����f,Smqbi.,IqDG�yw�,�ܬ�ޫ ö*jxUA
j�J���uŀg����\�9�s�� �z��+쬮;*�{�X;�V�o+��q`=�TWE�������ӻ�`��;�ִϹ۠=�fg}zz��M�`�Y9����p#\���uq��t���L*<+:{S�$�W�����6���;�uŀo���ӻ�`wwUr���H�!I+��q`��`t��Xv�ױbI��s��ڬ�YU%�Z �~�����~�T�	��P��H4��z*�կ�����>���7�;�촹
�dl�[���n�3������`t��U*IR��B�J�3������`���>󠕄���B��nR�Nv$��Yy��s�a�{�ݸ����b�Ȗ�ՈST�U%`g��,wyX���;�����*��쬮;*�9�� {���3����z{�
��U4M%`����c���������t��#����� �~�}Uߞ���W�����l )(	0Im5�付�q}���@}��܏Q�� ��b�"�3���7w��g������<�b_t�jF�W�ad��-��.�"�u��σl��X@�烍]���u�5Z�VF�����n�;���s�@���3����o\J�	}B�*��U%`��`���3���7w��a�s�GX�-�W-���� o���wyX����ة��P$��D�J���ϵ�`�Հ{���3������F�H�쬭�m�9���̝�k <�V��ViA D�}0*L�$�S$TB1DY.0=�fiW���Ӈ����pıh���{�j�V�����?�t}N젴v�����(�<w+RVKwm+��F�AЄB��Llc����FҺ�mښ1���r�k��D�zfb �t��Y�r⪫q��.�T
�������[��yZ
¼Y�%�]�cI����eݖ���Ů�[l�O=�	�tx�ͦ�!�����7n��SC�sx0��A��}�~}ҝ�s�.H�뎚<:�&�[��c�f�����:��Ny�����/;#s��;8k�m��Հgw+ �w+ ��V{��&hS2(�Dʔ��gw+ �w+ �޺ ��v��rA��hIn�3���7���=��`������)B��T�����}����V���=ܬ�Q<��E J��ET��}���7�V�nՀ{�mX�����o|�E�RQI-T�VѬ��&r��[���� �0�������#ƭ�B�K <�� �w+ �o'Dd���X;����T��D���g���g�)��(C�;O�;���R�`���3���ݽeLR�2�IS5I+ �o+ ����go+ �����}�F�U� �bQ���5`|Հg���o������±��E�u�t��@y?��]�w�����n�8|��E�lC�1���\������Z\��KA[�"�a�h����$m��[���� s�uX{yXv�:cz9*P��(E"��V��V��o5`|Հg����;We��J�8Y-���n�7�v�%1Ē��I��u��s���]'$�T�(D%J�V���=��}��=���ة(�@�!MR�I+ �o+ �o+ �o+'���7�Ӳ؈7"��$r�:�h'�l�k�yX�6/1I��e�,V晲[[��T�3UIX�yX{yX=�V�޺ �Ϫ
7:�X����s�^rz_:�o5`��n"&G��)�Q0��MMJI+��Հ{w��n�+ �9۠;�u����@h�� o�~�U^���꫿=�}Wrp��q$�on��\��v��jʩ�۠����`���3w�����50tbf�a�5u����瓪����v��Kn۶����lS��OMi�m�(�k�����`��`���ݣ���F2�+eU�t��^I6s�� ��X{yXf�I�%I)MU(�������`��`�����%�Z�7ednIn�9�v�s��7���g���g��*���
����RV��V�����V���,�άY���m��Z(�r֠�n�br�eêU��HL����Ҍ���gq۲<�l@�n��	r[Q`qg���v�n����8ٮ52��w�w:�-��Ϝ��n�xxi�Ț����f�t���m�VԱ��қ�ӗvm��!���K����RWg�7g�Ӣc����;�s[S��=��s��&�I-�e�ŝ9н��dMΡ7V�	���qʚ���eĪY���$���Q�-a���7��cu�w�.�D�2g��\8u�R�nU�SUEN8����n�>��� ��V�w+��5TIrI)$IX�ܬ{yX{�X��:c��$P�Q*�V�����V~�铟5`��6�䔪��USBI+ ����oo+ ����oo+v��I*�$P�J�	+�{y|��y�}�\���t�|w�؝-n�P�e��e�ɴ���]l��`�n��::�]�G��2����j�NIT����s��w������333y�w�;���X��vV�Qˬ�{��b�`X����Н�_y������<�u(�:�X����w�{��{۝��wY���9�9�Z��QES�:��s�����wY���;���.�rA���@U�%����o�ݧ���m�weӳ�����hh�H�ū��5�;�WO.�ۛv�Ҙ�qn9�C�P��\qA8�vЄ-�"nۼ�������;���-�I�N�,���}Ͻ���R��j����wgv|��l�L���Uv�t��3����pĿ�b�g��&�"�1��A�'���Mm%	���-�;2r�����vt��]lO@t�kD�5Qx�gK�p����ݨ�P�@��0iG�o�Z<3RU��)�F���oѐXi�2�� �12���D�2BC�s�)�=҆��z`8�]��uRQ�Oy�0�(;X�ȭa��H0�d$��/g)
��C�vP�.�X[޴�c9�%#4�:0p7XC��5ܴF�a�(/w�� ΄:�N�0���1��C�N��!,�2H�-G�#��Az���]j7�C�ʑ	8��&���Bfí:g��e���;@1A<���!׽1�8�qz]h5'C`ٹ0�������ǨB ��:}�}P=E�0W��GR�� �
�U:D�A�]�>�M��6�|d���~�JR��{���l�A��ί2"2O3��m�ĥ(y��Cܥ)}�s})JRs�~�Cܥ��9�����)C�?p��l#U��Z�C�ZY�1b;�z�1b���·�JR����R����fb��,Y�ߚӂ�O��%r�KHa��t�ۙ�z{LdDخnP���u�z�S�Q��snUB�H�-�y�3b�����l�D��9���)C�=�:�)K�s��Pf ��w�Bq�QES��t�fb%/��o�?!9)C�߿~�{��.~��})JRs�~�Cܟ�a�O�r��֬�ȷ��dZ��Ҕ������R���9���)9�s��R���9��b\�z:[B�B-M]kK6f*R����R����·�JR����R���=��@� A ��a ��BXJ!����J�����<�·�Pf.�v7"Nxd��۬��1{��·�JB O��l�{�t��}ss|}�v�"���;j)[m��&�9�/i����F4�
;rŁ��C�����j�5V������������9���)C�=�:�)O��uд�'=��t=ʃ1�^dDM�䝒�m��A��<���=�R�s��)JN{���{��w���b�9�y?P�MWej��k���R����])JRs�~�Cܥ)}�s})JRs�y�Cܥ)�������l��A�����K6f R����R����|��JS�s�t�f ��w�D Ȣ��$M�t�fb/��o�)JN{�7�{��>�9�JR������)Jq�a9�9��޵���T�gc��\�H-ج�:(�ٷS��]�Z�5�^,ԓ�줂�KӾk�����5d��$�h�.3�:��(ݴJxsm	�݈�94���ђ�G��&�P]= /7\\/*�R���jyɎwT���N�p����m��!��k��q���b[F�g>�vmc.Խ�z�/tsʶ�Z1�^f�j��r��,���@�M5a\��\��$�b_��oZ�o�N[<�v5�)�']Z�v
�0d��،�O���p5����y5��n�ȵ���)JN����Cܥ)}Ϲ���)=��s��R�����JR��}�ގ�R�ADݺгfb�w���aJR{Ͼ�Cܥ)�s�k�)JO�篅�3f.�.��I�,���f�'���t=�R�g>�R����s|��JR��s})JR}�9���z5�*���ݺY�1b��}5��1.��o��)J_s�o�)JOy���{���/��Ȉ���;%��k1b]���!�R�����JR������)�����b���ԡ�婃���p�ӧ�<��hL��qcp�G*���K^����]ps��ʞ�*i��V�гfb�w���R����}·�JS����A�*�)I�~��{��=3�ά���oV��k-�{�JR��}�:��MѰ�Pv��䦳�s])JR}�9�Cܥ)}Ϲ���
��������A�ENI�ۥ�3f/?��:R����s|��²�d�������)>��~�{��9��3Y���-�Y����(�I����r���>��R����}·�J����JS�1}��v�FKiv�B͙�3�}���)I�>��r���>��R����s|��JS��o������owk%��hm�Wv�k��3��ձ<[�``vN��f\�J/p�Uڪ���e)>��~�{��/��7Ҕ�'�s��=�R�����JR��y��o{ѭ�Em��t�fb�w���b����yr���>��R����}·�JT}��@�qy'e�-�Y�3b����=�R�����Jv+�H��U��*" �R�a�!FD(Q�	W�^�B)�:��s��=�R�g9�t�)C��g6U4�l�F�гfb�w���b�I�=��r���Ϲ���)>�o���A��O�PL�P,D���u��1���|���u<�m݁݁�{��Cܥ)}Ϲ���)?������3��;Z+���3�'b������ۂ����鱷mZ%8��r��\Yk����=p���;�ĥ)�����JR��9��r���>��R����y·�JS�}s5�2�"��5�k[�JR��y�o��)J_s�o�)JOy���{��>�}�t�(��z;\�%����u�f�����s})JR{Ͼ�Cܥ)}Ϲ���A��{��͙�3}dr$灖I{��Ҕ�'���t=�R�����JR��9���(8��$��!"���* B�(]�w���);���f���[TV��K6f �]|���f �߽��{��/y�7Ҕ�'���t=�R��39?~��9sp����5EGN�n l���vT��u��s�,���ў��s�Wl�b���޿��3f#��JR���߹��)J}���JR���Gꊚh�V�MhY�1b9��})JR{�~�Cܥ)�{�k�)JW~�o��3f/��'�#p��)JOy���{��>�y�t�)I���|��JR����R���߾��TUU9"v],٘�1u�ޚ�A��>�o��)J^��JP��,���s��l�A��w��b�u��,�b�)>�o��)J^��JR���߹��)J}�s��JR��x�C!�K �q�\q0=������2V79a��Rm7ue�u���Jv�nu��qͱ�g��������w�>x����g�g:�6�iLc�#�v�p�g��G/�=�[z#�己N��K�L��C��;Z死[�' �g#q1C���û.��.Wcj�g;k�レ�,c�v���+�&3��q���<;���W ��<x[@U&���<���VG�gV�t��Q��&�m)��W7qъ�<=t8�L�؆ɝ����vf�H+�	-��X�Teu��,�ț��t�D���~�JR���߹��)J}�s��Pf �߽��f������9s��5�V���)JOy���{����s��t�)I�s��R���9�������?;l�L�I,v],٘�0�>�5Ҕ�'�s���)K�s��JR��{�:�)Kߎe��Y���޷��{�JR�Y2N{���r����߷Ҕ�'���t=�R�g��R���:?UShE��6WMf�����9�)JP	�=��r����9������'��l�A����)&�py-C���O�mn=T/f�Ѐ1���L��1�gz��n�M%U�PR=(��+mz�A�����t=�R�g��R����u�`�*��Oy�1b_w�^��"���ɣ3{�{��>Ϲ�t���b{,�&�Bڂc�ܥ'}}�{�ܥ)�5�gJR������)Js��� -1WZ�r�f �A��v{�{��=���J$I��s�Cܤf/?~�5��1/���Ζ����u�X=�R��9�t�)I�~��r����9���)9���0{��=揵��'<�+��f �A���}��3�Vy�~����)?{�~��ܥ)���5��1.w��
TE�'kr[�G�;[�����2��WkIc�å}D�M6����Dʔ����͙�3_}��
Rsϵ�`�)J{��5Ҕ�'���if����W� ���L��v�f R��>�9��~ FC%>�߿k�)JOs���)O��s])JP��fsa@h�W���٘�1q�ޚ�A�I�>��r�~W����9���])JRw�5��=�R�k�����
[f�f ����if��
}�s��JR��>�9�ܥ)���3�A���痬���(�rDݺY�1���R���ϵ�`�)J{���JR��}�:�)K���Z�4sV�e_"���s�;8ծQ6-eK�lj���p���c��܀�u��,�b�}���0{��=�\�t�)I�>��s�3=���1}�~t���Xd3]u�Z�)O}�9�)JR{�y·�JS���k�)JO��}���JR����9s�Ie�
�^�f �����Cܥ)�{�5Ҕ�'��>懹JS�Oy�1b]^����2�$�Kn��JS���k�)JN��\�r����Δ�1��3�t@�H&i"BT�(
 00I�	H�0	Ȓ��� 1|!N{'}��=�R��]d#C��:팖�f �A�}��0{��?������)JR{�s�Cܤf.>w�Y�3b���lD����e�s�v�O7�e)�-��-��)1ۀ�V4qu�(�r��Wi��t�l�A����3�)JO>��t=�R��s]�IrR��s_�`�)JpϿ�5��oFf�-oyҔ�'�}�:�)Os߹���);��s�=�R�{�s:R���<�e����7n�l�A����Mf�'}�s�JS�u�gJR��}��K6f �Gy�7$b�Uւ4[f�)F����9�ܥ)��3�)JO>��t=�P~`�}���JR���~��R[aJ˭6f �_r{�Y����(���s��%)O��~�JR����!�R���U�a���(4���ba���_vݚ��]	�'�!�%h�`�zh��!Ԧ�q�H H#��%o����ù������t�d�@������hz�4��Gӣ���h �`��2a$6�,6��EWn�i���kV`��THm�k�B����U#�%��<�형b�������d0#Lh,$���y놔Ȇ��<� �L� �l���"e��C�p��d����ic��FXDFf� ��$��{	]"=��&B��Zt��l�JD+�abS0��	�cC' ������u�~Lw��5�1K�$���uL�B	5C�R'�f��:"�fz������_���   [[k{-�L�����  ��Ԡ��Si.�t�s�㥝j���d�g*���ҭcS*��$v���Ā}֐�a#�N��`���lh̪�7W�� ;�$jn��h�f�)ZѠ�'\� W�ַj�6��%�d-�	�\X$L�yܬ�R|�b�9!dvνlm��4�����%u0�f���
,u[�B��q��;;YIr�<e���c�6ǜ�-��ݹ��Jݪe���>���\�����9,�&ж��y刋���۱�s��Q4�[9�ӏsqciv�3�����������*��D݋�)��[Q���f����!ۄep_��X���4;@&Q�c��2OJ������ޜ�l���N��[(v2Q�6]�L���n�Evơ@�3�)y�ö�Q��k{+�����M�/Q\p��4mP�t�s��T�j��+bG�˱��+izVx��p3�Rݸ"��..��3p�U�hnNz�m�[x������E��K<جu�IK�G^Iڻ�7�C����9MX�2���������l��kW��8���@�� u��av�m���Rp�o��b1����@<�'.F��@����fv�5�S�=n��+���ݝ�쬾e�H�=��J�ժ�����]t�P �6]��<��WiM��(:�����uPF�c���X� ��bSwQ���v��Vm�,�zjv͖�[���@�\N1흞�p��^\��R�7[Y��rh��}���pp}u�6�36�ny��˝�Eo:�c�5��h��L{V���&��K	���M���*t3����%��S&�h�H���|�i��������m&L�R�l�0���[�qN���8���Hv�ݛ��svl�@�f�Y`&�Z�9�۫`�-u�vHܐ��ɞȮ��(	��`��O-<����/�.1'�@gr��4m���j�71�=�=��ͪ:����o{�A^��_��t��)(O�M@O�=@W�Q;TǨ!� s;�^ot��F���p�Yq
%�SD]�Jg�/Kֱ�]U�'�C
�����J:y˩Q�<A�'jƳx�!)'�w@&ě�e�m���О���l��%:��KN����d�na�u�S��Z���1����&�^P4�+.��s]�ըܑ� ����A>3�]��5�M��V�vMĖ�gv����t��ld��KIA�Q���ĒQf~�~�]z���K.	����lu�!��b$RФ@��\GE�v^�S��p���̌o7��JR��s���)Os߹���)9�9�Cܥ)��3�)JOy�}m�L�9l�[��3f.>w�I/�NJRy�~��{��>�_�gJR��w���l�A���y��/$�B[5�JRw���!�R���s�Ҕ�	��s���)O��ߵҔ�����7@M���I�6f I.r{�Y�1)=��s��R��=�5Ҕ�I����,٘�1\� �<�X����k1������)H��{�k�)JO��7�{��=�y�t�)I�>��,�i���vmZ�`M�k��I����C�2&ѐ�<�0�z<����ݮz~#���岷���JS����JR��y�o�u{���'i,a������~nH�X��h��U���\�҂����������������lj�l�����M�y{���YIm�(G.�l���4��|:�X���n��"i�R�SB�J�}�0�n��v�����/u���L�9l�[����:�;��0�n�}�0���R�Z/k�&�D����'��џ34]��\tu�gZ=�\bW5�w'a�j�S����	Z0G���ug33}���`Ԡ��&��H���0G��v�uf��S`o�Z0wfX�i�yM!R����w�����4uwi$cĒȅ����
yݳ ��u`oCt�@R��ffh���fhvww}��ou�y�ޚ#K}�}� {�<�U���&���3�ZX����}�6�uf��zh����M9aS���Kyd�a�us�9;uшL��p�����g5~w���0��R"�T!JWf��Ձ��� �������v��7R����iR��JU`k�y��ηVy�f��zi`.:�,s*R[#��`q�ޫ�ݳ�n���0�DT�2&j���"�l9��;������`-��w�~wÀ� `ea�%��aS�E��?u��������o,�`�Jh�
�� ������� 7[Z�{��9�\&zYZ��9U��8�=��M�)2<=��N�^���<��.�qٹ"JQ@�&h"�*�5�<��Ձ�nـl�u`oC�M(J*��
�f {�U�D˯�c{���n���sSRB������;��ηV�[� �mX��ڤ(E$�B
���g[�ۭ� n��{�� �:K�R��R��JU`{u��9���w��{���=Jl
�waٙ�X%�#I{�]��(�5Q?�kU�Ud)aȭ��sn�^���`'��a��]��F��iHxf�f3g;42���� V��&��M�(s��p�Ӈ O �s�>;A��pZ�4(�#cR"PV��A �mʸG�ي�&�/5��=��VSOhf��n����g�mf����A9�+/AT������P��<<�d�1���sU�؄�0��~Y����-g�|�Uc�!Q��X�|�;K�m���pu��F4��X�W7\.J�U��*RZ��?����t�%h�=JY��ـ	1��2s4UUKLUU���Z3�� ���7w�0u�`��5
I���)�d*��g[�w[� �mX�v� �5�P�(������"�o0u�`{��0��ݦ��އ���)BTUMQU��%V3�;C;�{����lot��=��wʇ��KTQD���v䷕c����O&�B<]<la�Z�������{�֍8�b���������`l�u`n�y��Gр��v:T�E-���ލ���zk��bF!Y�{8�� u�9ם�U�����g3�<;���@q�=5OEASR�4ET��ݘ�%V���ǽ䱰>{�@mw���ؤʔ��-���19�%V�䱰G��qٝ٣����y�d�䝶��@s����9Ḿ�6� 7[VN�E%C�
Iq�Eol���\��j���E�ȁ;G��C�MWc�if$�n�j(�[+�u�t�9<����y������ �瑀��!���%�@o�{���X�b��w���]��z<�ۻ;8���TH�*���2�`�j����0���"PV!	=G��� ��{�j�m�� ��jjHRB�0 �V�����vwW��9����s��_�sw���\qECMLH4��6��S`����|��ޔ�����6 �;��=�.�9��cXm�e56[q�%�Ou,	/!\�9iهI����O4�J�y���76DD}`:�X���U_(����%��76*-^��9��^�溫�9�w���Pp=�~�FH~J�m���{�~��|n�#�>3ͼ�7i�����T$AT���3J� �>��u��3ͼ�7i�:��:�S�P� �^wιwU�k�$��Q5PERU`{u��7i��>�U� �y)�9ٖٝ�R4�CS�c�
���avݸ5�lَ[κk�����uh�=�Ot��{����훩W�}��=�`}��F��Sn��y,��q�*�]h#U���s�� ���}� ��(�vfa�k.8������bBb�,�67�l��Y�3<F���7{��0�Ӥ�B�R�Q4�J�>=�o0�nl{]� �����}=.�+�T�RIf�M̀{��0�n�{[�s��B��	J����/g��)�y���B90;%�E�gll5%�خ�t8�isbBsr�WX�A؍�9�ɵ��Lf{��s��8��e,�c����:wY�uۻ<J�mu�z�SsFM�vv��f:C�1e8Ԉ�ׇF����l��etո�{�
�c���6.�zV.ܒ/7:�:z�b�Gv|��l�9pZ�n���:��-�U�v�m�|��޷���U-�Ք.:{�1��0=Ia�sI]�u��Uq�a:��݁����
�������k�8��K�����7i���uKJ%|AJ��2Wf�������w&X��f�8������P��h�罽��ɖ��ـz[u`{�ç
�)BUUQH%,�>�����l�=-���,�,|�~��?w��ȣu���F۪�{]� ���۫��� ��u`~_�~�4"~\V�'GG�r'6�є�i��l3�c�q�6�$Ӣ��Oi�u��<LHLU}g�z;�l��Y�ln��f�k�`�:��P�$�J�i�X��w�@��  �0>A�	F#i����I��_|����6ںр}	)�wp<�caQSS4�T���`�l{vч33����-��>��� �aHș��j����7{��m76ko0���sV ��(��*SD�M]��nl�ݛ<�� [��{�h�7�x�j�Ǉ�j��)4�^�m�hef|S���eq�7m�c{gD&�T��KbN�Z#iǥB1�(���>�wf -�V��~;�����������穀�j������� [��{�h��"�ϒY�����͉����#���`��������ճfʺ1�� 4�$�H�p���s_�5�"B�� ��`0�1�i��]��=#�@�y1��'4�F
�Sj�H�ӫ�P� ��4�dvF�H֘sft!�M�!��(S�AH�,@L� kҔ�=F�b�	!��S�3����n�uz���4K�t����a�{���t�x�P��U���tX'���&���`��vx+�؜؛;UO��Q�o�t�$S�4"�*;E�E_ ��G|�c;|���NΝݜ�=�� �U`y-J%H�UUIR�Y�}Ze���� }�X������r�!I)R�*��X���>sV�u� z�,ؒ��{�
Xۊ��I,b���Ɛ�p�.�z��Kc��S��6�M����;��H�1U535 r]V��h��#� >��� �c���"[���jZ���ou� z�,��`�j�1�:SE8��DU[`l�y%�s;���U���c`�H�����SLM%6ko0{��7{�FDDD�nlt7N%LIK�j���Y��Ձ�{V6��Q`g�,�9��ƇL����"�cIu�3�z�Fp6\	�\3�.�����Zw�օ�:�M��6;����=�����`�5`k|5(�")TIU%JK# �Ss`f�� 7��w��`�OS��
IJ�IJ�)�3[y��Ձ���0u76���c"�y��.��$�}��]�����)E��$� 7XR�ɚj&��j����V��o*�۽ـ^��7�]�O��)�$X�(4�2�I�Ҡ��1
1&�!�MbI���ڟ��(���֚��&9e���c6�/��?4��6��Pl�f9j�&�L��s��p[Yem.�׃�f�Vfp �[\��1��1m6�՝����X�P�瞶�2N�Sk��V3�i뗶7Z[`�%�i�{^lp���q��]��M�
���<�/c���+$�0�Kq{�q�[E�f����d�8��|���ZrWe���ؖf~Ř��Ė/�6�i�ɲ��A��1�w+�ۘ*p�W���K/��T�˸#��+:��_}|鸽�5�LJWf�_��6�[� ��v�f q{��ӏʄc�'-z�����H�j��k�`�nn ��ĩ�)|�MTR�K0{��=��}����ݭ� =c���aMLHJJ����0u76�[�>�����Ԍ�Ibd��Ѱ>����1,���� 7����l�7\;�������[Z'�cd}Y�.���m���d�u�m�(�N��بxV��کX픊X�z�s���=����yZ���R�7�訩�Z�9k�K��s���U,K���bZ�*I"���҂p�Q�E;Qـ�޾0l��� 7X�$A!
�¤��ۮـ{������<����j�1�e*W�$I3"Wwuኈ��s7W���ﺯ~�[�U�}�t�˽�F�<�6XE%�@}�7���X�����=�TD(r��kD�#�d6�-�oH�G��;�y�82G�c����ݦ~�;z�y���۪���� �e(�wwv�� ��T*!Q2��;u�0�R��� =����݀�$�fZ*R���E5Yf�������>�&!LISS`��8�wf�fw�T����F򖍕OT�
�������� 7���Ss�|�_v{�@y|uwԶ��-vIw��j�>�;v���Ḿ�� ��闵��Ӳ`.F+�9�;n�]���f��K�����mE���bLWiN=wZc�%`v�npu76����#� j]V�j�)��*��"
���>�No���0{��1�npa��(�� �IU���� 7���|����Ձ�]8�A%/�����4� wc۪�[IF�jSa�vv�gb������7�W��t�&� �#��Ձ��� 7��ݰ��	�놲����=�e�:�I�-� �룎�-��0l2w����5�U@L�� ��u`ww<��j���s�y�OP��PJ�*�BJ�����ݙ����5.���0�R�wg`=㣥�U)>�Ji$� 7��v���Ձ��� ;�qEHMC�D�=MUX;3��Z� �5)�3wV`���5`�:HQ_LT�E1Uj� ��S`s�337�.��K�����w;@@8� 	$�,2���O�U��#G8����ڀ�z��k���ja�Z�v\�iN�n�؅�k��^rb�'ޖ���ݎ�aܖqv;v�� D
���l7eם\ۍ��7P`���ͭ���WoJv�a�ͧ�ڗ�j�sV�igqh@l�gq���R㶹�ɝI?�b�������T�.;W�L-�� F_h]ɶ��%D���]i:�[ôjFơ坤���0ݞ++��~��{�����;��3���6�E�sۉ��(��5�s�8#wC�Ta,�I�?����LL�����m�y��Ձ�˜��}�7�X��J�\$QW.���W����R��=�l�՘ ���xJ�\h#m��o|�Ͼ����0{��=�UN�A)���+.� �5)�3wV`�*��fwvh�;� ������A*P�)	*�=���ڰ3u78�7Vs�p)J��v�O<2�#�v�s��y��\��:�6�r�nͨ4�:�n'f7������=�U���%�R�ggg�y.� ^G����+$�e�@o�����!@ͮ������dD���V`�*�6��_J�x�v��5t�}�>���wgvh�WuXn�t`�$I4˄�*����y�ͫ7Ss�q�ޚq�?0d���Ee��=�U�����G�l.�>�uf �P*��z�՞����v���X�W�]v.8�x��Gm^rlݧ���P'�ۡ;d�R�3u78�7V��� 7�V�S ��351 ��p�n�{�� o6��M���z���A*P�*����V`�*��۾v���Wtl�~�48qu�'\er�Kn���Dj����ѩM�G��}�	1��q~I�.Im��/��}�3��0y�`d����s*EP��ۜ�wY8Q9-�\��W��պ���W����5&�&5]��jM]=���zh��<��Ձ����C�4I1R�A(�������a�ͫ=O�`<��<A��M1�QQ$�KEMf j�=]ΰ��g��7y� =c��
�UƂ0r��7��}6}�7�}����XA�I�0�pǋ<�f/b]�=u��>�W��#e����AYus�z5)�9��ٛ��������w:�n�U*IJUI	��d�Z]��G@O'ݥ��y
����va��4�/� �(U��X���ڰ7��}X����4zqu�'Yr�	���jU|;334ޞ]8���s���cg��~�"����Ym�zyt��Jlٙ��{V`�*�2=��=!�L�)�u6�f'��ߦ��uv`�*�ggvc>��8�(Q1.����J����ڰ3��s]��}�k����^|lW% CҀ#�L$�CA	�)�5v6��� �@!���0@&غ48y�˭��)0�]�@v3vw�i	���pZ`�IәX�
T��vH�m�d�4�y��h�i�ڏJ1)�:�J'@�gj�jT2���h��%�P��)���2S��AuF�LP; ҃���&)J� }o�w����{  ���ͭMG��\Ѯ  ޽��Հ�Ium.�L��6��[;l�L��m��.���q*�c��B;��,q����n���T9���W8��SĥBW�ҡ���z��d�͝F�WX6�Kh���Y6�(�
�@�+t'a�Zf�Ozu��@)�AV�55�7)=SnEs�˕hAtUVW��Pی��t�+*ӳV�]�(kcZ�	�]e&Wk�D6�����n���I�N;9̂;N3��s[1b��2�J��%�F�����糪A�/I��p�l�&���q���\�˺6,��^��XBq�$IR�	���Jvvz=�[��ve-R�Ur�K�kL�>�:5ɜƛ��xn�9�n��Aq�k�-�u;v8�LW.GSjѹ�	��WSz8��v�w<a�k�rK(LZ��qNu�v7bv{C���W� c�<':wO7�R��K�qr��8��ֻ���¶54�;:����	��@��R�K'@U�ub�W9�,�f,n�Zu����LD��cLx��Ռ���.A$�ģ<d6�v;�q���TE�P���@��m�]%����"�n	�m�6���t���]r1e#8�[����
�d�]��;Yz�.m<�.��g�Jϳ��j�3�4�ppሪV8v�l݌����6�9X�Cۋ:v�էh���x
�ŷ�*ٶw^�<��:��j�I9i�J�y��mn�M�Q�Y�Sİe��h������O
l�ˮY�Õ&q��yZ��%��8�l��L��g7, ��[1;�h�St���9R����n90���1���c��D��e\�suS�7S��^V��ަ��k:N�XM������퍭ّ*n�G5\�FŜ��J�v{m/n�q�4��t��vM��5��r\k��wc9�ֹK����]b�W7dwSv8;nb��j�ڴ�n�{vy�RZ�6'T��JF������6◞)�v��9xz:��j]X����)�\B�>U^�v+��t���{� ��Q�E=��� ��K�K1'�Y��yjt��Gmj�S-ve�����i��7n����s�p��.�-�d�>cIk�E����N��K��:�cY��ٽ�0�������Fe44\��z^`����CE�ax�6�,�]qY�U������W;�Y�=�t��]s.��tN���6:��z܀��v3��\��˥�I<�Tز�͡�#C�\�9�L٨���<�����w{�}����S�5�՛'F�pz�Zϲi�n^�mjI�q�<���~�,Mפ��d���E���}tz��`<�_�D@��0��R���T��Vz��`<�X�����Ib����l���2�WS �����o<��Ձ��ΰ��n��"	R�QHIU�}�y� o6��>u�l�u`w4�T�>�JJIf o6��>u�l�u`o��`~��P�)k���Jʛ(�v��U��5%vW�ݍS�r�siѻ}���o�����|U%`g����V�y�����wU��%=3�$�UCA3-75s�l$��h��g�vg�g�_f`�*�7��}7�$�qu�q�������f��.��IU�;1�/j�a%6oW����Ic�{ٍ����@q���`-�������� =c���T@���&�+����">��mՁ�����޺�8�hD�Gr��:�Ooa��vyܤ+\��O�Շ��v�!��]+j�L����1U��:[u`w���iWc�34��u`
at�=P�TQR�EUM��y,�ff���`z;WV -�]fb��9�ҷr�I.�_�M��/j�-����w�33U�Ձ��}���yP"=+I�S�A�fK�k 9�V{[���v���UV![FI�����������{[B�6н���.:�rZ%��Z��1�����l��ɹ��ϔv0���J�nJ��0GhE]q���Y��l��~����:�=/y����u`gl�K��&�H�����Y�9|�������X �5`o�����bM�;��W`�49f��-]X ����٣�ـtr�7펪�TȊ�3%b����Vv�������U�@����=D�c��`��n��"	R�QQ5IX��`
��>�����U��������O%J�>v��s�C[7N�'OVLۉ�6�U�=T������o.���:9t�F�U`Z����Y�l	��Q��d�7+�>���,O~��`|��0�TX���7R�TAUR]R���Vv��} v��Okk =.jfb����eL���;u���Ձ�z��#�_5`{�zD�AS1$�Y����gOou|������]�ϴ�D)UQ%5MLUcs��
O2^�hfܘ�)hij$'$Qu��L�'iN۝�L;s��]\�����5��^�+�u���;t8݊Kq�5&��1n�smgv�g\ 2��D�v{P[��Q��aY@.y�9�����4�n�)(ʼ�����%Su�;�V��1�Ã{�2;�lu��ru"�o��C�q��S�ڂ�	+i��Ϣ��*�ZU��f)�`�E�9F� ���ݱ��Q8��F0.�/Ol��h8��Յ�%�r�+��A�@|����B�6�䳜vv�.���"8�h蘨�$�*n� �Z�������� \���{U`�����j�����*b��U`w���|՞���5`t�s@}ӝP1�sZ33��@9{�`/�X�o0���PTK)TB�PU%`z^�X}�G�/�X�o0�ﮀ����lB�Iji�Q�����6�a�Q�il�[��@O9��Ve�~_}/�.�$EMIuJ���Ձ��� 9�_�X��,�a����v����ڏ�+#n�-�@w�{���,ϳ����V�}�]���V����vggaݚ尛���&�
��&�� ]�Vн�������{{ �:y�E��67-�~wfa���ں��6�� 5%V�qU,��SR�d�LUv���X�o0�j����oC����%J��Z���8��0��^n�y�b;0���㙴������<ݲܴC��(�,������ڰ=/y���Ձ�;�Ц��̕S33Y�$���ٝ� �n��B]6}��9�� ��4�-1R�U4��U��n��cuM�gf~a�ٝ�;5��}���� ;�5`w��UiEIH�����k ��u`g��`�j�������f��%)MR�=�� <�VN�5�t�:�;�TDQ\s�{\�s�YڔP���w�vG� ���=s����-��6�+i�іG�n���VN�5�t�:�3��0��](����Aܷ@m����1����4�K� >IU�A��ĝ1TLTCD���`[�V{�� y����� G��%��B��*�=����o���}�7�y؜_Q�w�<�Tn�
jh���UUIf y������������`렗J�B��Lb�lhpm�q��v9&k]����^�f-��D��"�ݢUڜ���s����Ձ��y�m��O��J
�IUT�`=ά�7��ڰ<�����Ƙg�G#k�(�e�K4�]ـ$��fg��n�� IuX��132�"��*	��m�ӻΰwUXs�;4}��� $�:i���a"����N�5�A��X��`��7�_
|�B
B��Ī2$���
��ʒ�g�_�V�ꚇ׃ekt�ҫ[\�䮎���+�7O[��$$�����ԛt�@iܶ��mjx��\�3�b���.vȏ`B�9�jHs�ܮ#v�uE�]q�2v�vxz�'$۳�ŋ[�����d��4��ں!�d��x�ly���gs��*t����L@f�!�nӤ�5e�dm����uMu���0�knv{Z$�@p�if��Pl��vZES+��%sb^X[���N�a�ƵЏ9�u۶y�F� �ƌ*�8��e����I�ەGHv���d�Jր>mXu��6��w[� _s�ԩV!�lM;-��=���c4@{������ ��V�f�bHP�H�QUK0͵`9�m`w5`=�� ��EA#�|�(���;����Հ�[��͵`k��U�$�Uv���V�o0͵`9�m`�T�3#�P�(�I%�E�;���(V��eD��;��RnN��{��u5S1r"T�R%5J���`�j�s���:{�X�O1LĒ�"��+Vk}�U�9���� b"`+����;63��Հl{T��%���.��H��&i+ {�� ��ua�D��`�j�����:��MJ�����Ww�t�:����6Շ���x��R�RA*R���IX��`������ ��׀����(I���Z{h�p�'���68��sطc�g�Kv���ud��Y�|<�=OQuӜ�L���� �R� ^���n���ov`g�~Ȣ�S+�7-����[���`w��0�J�)Z�f�A����fȚ��n���K0���g��v�P����z�C��:�v�ѤR�J6�p���!�|¶�`=�S���2��I�Y4���ÚKm�z�f�n`�m��Hԅb��CC����8��E��b��&����	u���kXY�I��ytv��d��X�`�fafj�� ��x��TX5Izٽ뤶uН.3(�MTC�YH���\Y�:�R���t��M�uc��b�kڪ��>;P҇h	�	���"�(�
�H=��
(6$�X�����w���>]�$my֝cLQ3Sa���3G{{� ;�U�/{U�_:�3�=JD����&�`Z���wwhwn�]�˦�_y,�;���q��,c��N���R�kx.�6+�X�iٺx��/�pۤY�{Efk��d�
��J��;�|Հ���Gр�}t�sѩ�Z���on�k[ ժ�� �ov`��`��x3���3Q$R�TL*���o0�5`w��>j��o
jh�"!QJ�f� wcV���j�V�,%ӻ�(�)���R �"v��T�=�|�u{��QPH�)J*i+ {�� �ɖ���Ϛ���8Q*R�%%*Uֺ)���yA���ՖQA@�wUָ��B�������UV��!$H��*��ϓ,�o0�5`w���]S0�LJ�*E���X��a s����_���Ϲ���m1�2�BK��.]V ��W�8j�E���Y�t�IAS*�
��J��;�9�e����AϚ�3��hu2)��3EEM����`s3;7{{��r��~�]���!~�a�ba�b��ȱD,X��fz�M[b���Gm| �ݔ��ڀوz9�5����t]Rn�l@��kg�m$�I��79��n;\[�W{8 W��;r�h�U� ��l)ڕ�g��<[�3�B���8��^4�{���m�D9�a�f+���t�\��������n�x�-��&����i�ƨ��z� 9�т�]*A<��ִ�ʜ���ͯp�d5�5��/PO�P;Q6 uֵ����Y`�{&[���<8{��r���7��ݩ���$ϱ��%�N������]<J���y��� {�� �ɖ�7��5U����K0�5`w��ԭ�����fv�wv��Ls�Ku�M15V۫� ��mg;�3�G{{� 9���t���URL$�M\�+�菣y���[� �mX��x����g�i�U�*�����Ib7�V �y���ŀ�㚪��&��LM��<q��6��u<kO���"&3 m���N�%b����J�c�eR9!%��9�z�{گ ��m��ϐ��� [�S5�5Qh�0�� {�ﵷ��ŉ/� �� ��E��}�tuW���� �mX�s42�T�J���2U]���ŀ�����@ͫ {�� y�7�C���ڴ�I%��;��� ��V ��W�3;�R��>�����f^���I����jU`s3�n�����m`/��`	Nz�*b��I*&*K���m��ݰAZ�v��:�n*��Zm0����
R��J��;�7�������0y�`9{ʚ�E*DԪ�һ�7�������Հ=�w��ˏ���1�W,�@}�{��W�s���(�2�H(kW���뺾�������
�;FU#q�.�a��� ��� �n����� ;[UJ~�-LD�L�U�o���ϫ� �ov`�*�;x��0��1L�T�%>��xQH��G;$�v�f_Q�M�l��WL��f��T�JUIL*���s������� 7�Vۭ� Go9�(��&�B��I(�<��� �mXn�x�w�l�|Oʹ"�tN���{ �~� �y+��=��/%��XO-,4$D)�4��v�w�l�u`y�y��4��2��qH ��b�LP$�� %�D������_���g���YG��r�[����/��� ��V��W�s;���?¦~���-���OE��㊅�n���W��7����Ӊ�(�q�m�ڭ�g�w����{ ��V����gwf�awM��(\0�"�����Y�ͫ ��w�l�S`b�Y����"	bZ �� ��w��H�wf o6��sU�S)U%0d�Wx�7V=o0y�aۼ� #���"f	�P�&��X����Հv�;�6y��&>��b���;�UnP����i��vZ+	N���`Q��ak���m�t�h��kbó��s�ݩ}hˉ6+�<dYN=�w��ky����W�Z��iv���P-�W-�����)\:��-T�b�<�!�� v�UZ�m�q[@���3�'��:wX:5���lȩ,��#p�z�q���Du�ݰ�%$�wۗ{-�DBp�13�;9v%�p9�\�1�GP���{����}����JO��)����;TH�9tj�5���(|��z�����ڮ���%EHJW�ͫ ��w�l�u`c�� rt(*t�!M(����y���Ձ�[� �m\��ʘ�T�*D*�i]�<�X��Ù�]�`uu��y2��%�*d!�"j�Ý�f��{� 5wU�o���>��@}�_|V��*���{ �mXn�g�����Bz��o�-+��w	]7Z�8���xqp��tkA�v�gx���c���vpe��v�;�6y��1�y�ͫ�n8z7E�Zѷeֶ}驙ĳ�#茈���a�� 7[Vۼ� #���Q0MJ�P��X����՜���]x��5�ZSTL54SLUf3;�C�j� ��׀z5)�3�����
�)�SJ*i+ ��U��;l��>[ݘ�J�����ܜ�Pn����t�iw���#��2v�ax����C�4,˯����s�A�O�t���n��7��ڰ2wy� ��wQ��ܶh���{1 7�VN�5�l�u`{�-�f$����ܗ{ �}�6�����_=��f��D�(A��͎!�D�fgk�?�٬���`f���3P�"�q�In��bğӽ��:�������ڰ=�uS�Q)U%0F)��ѩM�������{W_����9�w��w��q���U����V:@�/!�kp��C�׈��N���e3u!�'>�d]��ԨU
�)U��m� o6�wy�}���}�7�ީ�YZ�tuF7n`�*�f��]x��>Ifs�����?(Ҵ��G-�;�~��������>3��`�j�;���*&��3)U�һ�6y��3��`�{�C�ܬ���	��(��HA$�)��=����zEC�]��:��o9�}5*�&J�X�o0w��n���,��DQQ1N� �tMG��t�۴�G+���p�g�Ls�ݫ+Bm�V��*��ܗ{ �;�n���."">=����:J~*�A5L�T��{w��֙`g����﮳1 >����F裶KZ7dWx��X�o0w��n� ���I �%V+�������l���{w����֙`c��B�?$!QRL����X�y��i�{�����_�}?�F_����X�
�����)X��ZH�$ �'bk�u������6z�W� &R��ؽ*�t�L$��0� M4�f,y�*`k�٠v3����I� &�s	H�-c��%�*�
h!̱q&p�O�j�T���0b	�ë���Hi#N斉��ҳ�`�'ghvL�!L�d�������!�F%Ϡ3��T�A!�baO�m�G�}��,��46!]�tĔMDZ��*eXYa`T�%%;s�����:�j'����V�I���33{�ڸ�m��m �vӱ�^�p(�����  v��+ R"麝l���δӤ�5�蝬��L֍��J��]�U��ۦ!��s�	����6	�%����6݃X�R+�dd�m�@,�.P��``ЗEN���m��vvˡ6�AL`��iݱ���.uQ��)D�g@�"�	s��6�3�����g���� ���%�A�C���s�� �d�6�a�u�<g7l���G���xa�m�C@k*�6+��#��O`�v����=%�Ѭ�[^TU�D�I���L�/�u�s]�w���3��s�t͡��0��8��{e˻>����	#B�]1'��;%Ѷ!�N�C(UW.۵�����	������.�r�U!.4�v�ʠ�yE��F]��C��P�N�ۑ8{ٞ�9{�z66y�8���{�(vڻ����x2�݂��Y�ٻk�u�7F��rF{U�hm'd�[$pݓk�� �]�t�k�b��eVsT��L�&��m�F����rX� :�K�>�$òR\sTݮ4����g�!����Km��G�A� �Ӎ�xч������4�%#�H�q���<ղv1����n�N9��V �y�,Gj�g%$��4�(���	i�� C�a8!��-ri�i
U++m��Z�{�6�5��Y���y�6�ٕ�	ۖc
G�쎹��F7V��R�3�`z�q�0(f)l�ټd�Vዜf�c�.���L,.r��6�ln�M��z\p���v���'jc-���'h���L���e�w���Mkx��WO��˵��3��ʉ�xP2l싵�ש����vn9mr�;��;�SrJ1B�s��ɹ�XU+���v'�U��W@/0t�Z�Yԩ���/[Q���d���\�Za<&y6�vѵ����-M�sZ�bюMtva���w��@rON�nn��=�x����ݕ6;j�X㗤rX�hF�Q�[���޽����> �&�E�=��v��g�ɡ�E]	�b�!֔��_$���]��嶕�l�e,��*���WYh ��8�4j8f/1T���,ui9u�ٷ��"�=�����g�2�ѵ/+�MٻZ�b��:C=�x�c;����'����{\.@C���Ol����I��-ok��ܥA�y��8z���i[璶�����s��l�F����:Y��)��u@�g.�B��]��w,\VG����<P��D틙�$�,�,CԲ"��GdC�X4=� ���.t�V2�1�̽v�t��׳&�*�� ��W*�[� ��ﵰ>�,�7�}��X{z�Ȩ�HS1SJ�������=�� w6�ۼ��@��$MEJ�	�*��=�� w6�ۼ� �Ḿ�9�jd�*�)�b&"f���	wU�{uu�R��|g���7Z�IL5

AD�T��{w��鹰3��`sj���8ߨN�<=p����^�}����l�A���L�I�n�)Gc�����"�H[���ߕ3Wx��}�f n�\��W^�=�����U��\�@o����ؐG�zAW{���꫿��:�y�9����R�R����&R� �mX�y����=�� �p�*A��T����n�]76{�� �mX{z��35))��������R�>Գ 7R� ���x;�:��o�=�ۆ6����s=�P�l��2��^H��zN��I�?3��}�0�K�h�����ـ�U�/{U�R�X{=��%"ESTL�� �mX��x�nl�o0�7Z�� ��PR6In�=�w�������F�$�d��¦�XI� ����y�� �mX����"�*��UJ��;���oWtX��� �J�9�ǃ�W�ls����rUb��+������ڰ���t��ޖĩT�z��^LGg�<�V]�Fy��g�Kv���ɒ9��iH]�VVW�����.���U�/{U�R�s�;d{{� �9��TVJ�����}��ĳ3?yW{{� ��p|�QU1EDQ4��һ�re���� =mX��x�9��5*�%
��`?ky��U�/{U�{�wgwye;h�=��a�3"�2(���f�`�Հ=�w�>���[�ͨ��&I�TM@Ap�kZ�3=��n-v�KGn'b�6Pe�=n[�m��J��⨰#m�n�=�w���S,�o>���=��sS2�	D�A��]��2�~�� {M̀=����,�x�s����rUb�[)�>�wf �)E�������,M��8T��**IT� {M̀n�;�5�e�|g�y�9t�3#��D��X��W�s;33o+� ��ݘy=�'䶒i�w��ꭤtV�kPu�ݬ�����1�
�� hh rAR���v @ K[R���87*�Ʋd��V����<މ��@Ƶ=nx _Z�`�Cul[�ڱ���;<t��`Nw5n1a�cu@%�u�Y��m,�ǚ�3�����m�z3�gs���=��}Mn+�;�� ;P�9���r�cn9v�k�ae�Ik��*�	Ӌ1f$��ij�"4�',��Ïvz�	�ΰ��̊�-��]<ݙ:�<��*��U4���3I]*Wl��X��`���D n�;�A�����UA(�T�<�� �mX���&X{���m�Vʤr1˽�{�����"�&X��`�P�*"J�AS35IX���&X��`[Vy�MTʨ�S4Pb�WxݤX�����7}���ggvn�o��)��⊻k�۬(O�<�����n��9;q6�X����s:W�gOf��m��Z�j����ـ�U�n�U��`y2��NTү����� zڱ�]���ٞ!��	�j�{i%�6Y�uEg����r[������L����1�y�[V�wU5$�)*eL��U+��&X�<��u`�;�l�����q7d�ՠ6������y)��j�n�k|����80�<�Ekư/� �$�P�{He��۷g��^
]�]-�� i�\�D�,��u`�����,o�`s�z�)T���h��}��;��V�%�0Jl�d��&�"�	�2�j� [���ĵf�3��	 @�ȱ�a"� ��B/��(�(�
^s<���{�����V+%��%����� �[� ��w�>�q`8��r��|��EH��`u����x ���1�y�v�K��JUJQ"*S9eM���ٱ�Bt@[Wa��^�j�s�oa�����ؓ�(�c�R��h��}��>�o�`u��{�i�&�IS*"��*j� Q���ffwh�]����@�;u�gx���q����̲[�;�v`�U`�j�F���kz&�X��nK���31,O�~���s�]����k���}x�0ъ��Go��>�j���R��m�-�;�W�(�S`f�Y��U���4:f8?|δ���t��
��e�U����N�2��Ӧ���ԣ4n���{����|YBqy������lի0y*�v�V�� o%��1MR�2MT��V`�j�7����j��"" ΍��*iW��"�Y�y� ��w���9���a�S3$�DP�"����gv�ի� ;WU���f ���|�+ ��4:52)�Jҥw��Ձ��� y��{y����5����TqJ�piv�۞R{5���^��+��gڋ���������<[�F8�hͷ;)=�u���s÷m�'̏c#�x��W��P�ݔn��z9�iΌ�ggw/[v��.�sn�iV����+��=��g��Hz�D[ŝ�<�,g�g��z��vܛ���j9�[�$����k�[���`vͩѤ�t�f骂E%HBe+%Q�,�cx%�X�?���e'���K�>gtc�5m:W>3:��D-x$/m�(��46��Y�ç�����~w�`�*�o�_���fvo�P�M�u�~��V�8A�w���] oo;�:{�XϞ`�P�*��UT$D��X�گ ��SgC;;4|�v`���M�U4�T�E�!�SWxOs���ڰ��x|�̌C��K!m�~�}���$bē�wU�%�� ��S`b���1-ST����n9��j)VsE���$�n4�곐(�4�-�Z�]Q�˽�}�z�{y������|� �tT�1.�]��n�9�w��^X��A�	fp��=t*	�+��s�5�]�Ϲ��>��u�����{�5����d��nj� P�M���f������V���������M��b��h1,F��y�m� ��w�t�:�=�=�bE R��(����ڰ��xOs�}�}��s�}�'�$*�-n:�����[�@X=4�a��ç�]ڴp�ZzC��-Ydy*�6�nIn�9�w��}���|� <�V8�Ҋ)T��'�)R��:{�XϞ`�j�7���3 _{��db$uJYl�����s��ó9��4����=�dPs��t�ν<��V�-a�ZG;(�����W�HD�Rx������M'i�:{1�u �+֗�f!�C٘-i�Y>��v�}�jk̠�j)�tb�b���QJh�v�>� �'jJ��POPT���� �W���u�t�:�3���SIB(�"�Y�$��=�����6���jK0��p�I��}HJf�+ ��w�t�:�3RY�$���u�GMT��4�Q��{6%���s��r��<Ǎ29m�ꔹ�t8xe��ZZ�5�J�cvW��u�����M��� �%\���� jK� �nj��
���"I����5%����^��l���@s�}^��V�8A�w�$��=���fvp��S`f�� ���,���Kq�$�A�1c}���[B]6jK09���]�`}̻��I��"�$ɪ��)J,gff�wv]�������� �2eq0��U$��[=�K�Uz:E�i�G�ۈ��N�l�)��]��bnX�F"GT�����s���������۸�1�E4���"Q4�D�`	JQ|����3��@tr]Xwu������i���h�h�&f��P�U`	%mg3�Gv�f�=�`|��<�q��-�����b���E�޷�t��_sX�q)��b��&���k/%�3;��uwF�?s���\�9��]��AC0�|,M�!%���֟g�c�K�� ��#b�����Z�u)�s���u#<\�� ��m����IG�W6���{�n��v�w#�I��F�sU������l�n��<���-��v�Z�m�mdҼ�������7�
��D2s�Y���˒�f0���0:8Ǝ�z��En̖��W\ V�ݎ���x�v �����r�̬cUŀ�krn�-ؗ��lL���וaPZ[-�eK1f{�Q
"'4�c�O�m��6�=�/6օ�j^�F��ћ�D��V�7U��V�8G$���?zl/����.>������b��(QIL�L��)���۸��� n��69����12�~�+V�����Y���%)E��n���j���fi���j��?�;�����~��m���,{�M)������`�s`1�� �w��{{�z�W�!Q����Ҝ���;��[�V-�ʼl�N�b�$�:ٺLA4<QTL�E��$� IR,���wwo�;��,|���=�LADL�]�u���9�]i�u.	�IB.pM��XBX� JuE��-U�/2h�S�SDQMU4X	-Y�%)E�����˫ ������k"X���
������ghf��:;�V ��X	-Y�=�p�������MR��|� �L�|� n������&bR�ۖNm"�#���i���h��MG݊U� 3���:����?�}~m�_��"�Kuf �����ܺ���:%� ��j��&��%�3��� ��:;�V ��[��Ҧ�j^��"�aK0鹰��a��#�$�XX��`'8U$�H���$X[��L�|� �i���u9)ML���M�V��L��|� �*E��-U�s�Jǒ#�\���i��{=jxAs��܉ڃ����xrRw+a#&���ƛj�j�V���)-���~�������|��Ḿ�g���U@��������p�����X�Y�r]mU$�4�DD�UMQ`tw.���X�y�ki�z9�5UJ����br���:������ـy*GU����К� ��޹���S/l)��fj�j�fh�If���|`��Հn�E��䘙��*%�ܾכY���y�8�㮺z84�iI���9��)��D�MR�r��$����,-�XsL�m��89©&J�H�%)"�r�k ��q`6��ͦX�s��@��T�T��+X�kjK0�wwa��wWB��s�#�RE(�D�H����o0��X
5%X�	.ưl&�X��`*f"`����;3�33𻺾��������9����=%|�%?!��������պ���5���n,�l�ul��@#[��<>�Î]*t=�ԝ9�`C��)���u�n�]�l<Y@��G9��ݻ�c�(�l�n�8YԀs����4n{(p�
]Qus��jt��S�C��ز�Y�^�岂k�_��/�����} <����˜�l]F@cH�9`��c�������ݷZ:�=���g���]bv2��ܷZ���H��Ł9�-n�=c��tgnҴ�!6j�eç����+���Z���� �STh����uR,�Y���������hq{��Ym���nn[��9�T_;����ـj���Q�*�^�u_L�UI
����o0sL��m`�2�Ǯ)В����QR�K0֙`9m��n󸰈���0���*�d��RJ�,-�X�;���0kL�;ڦb������N�\���vn�ɹ���YtKe�#ݸ���W����kMMH�u��9+֥���}��|� ���� -�X�.P��ML��IE����_G�Fz.�ƙ`d�m`��X�zPJ�T
�f�����L���a�wo�`���UX:��6[i���?��~�yu�����g��|Xy�G5U0�)�����V�|�,���;Ze��jU�s�;v�3u1QR-58��q�#tM��ʶ�	�b�g���釴��wSE\\K�35UA5T�r��|��ͮ�Hw5}�N��_!M���`����ܰ�wm�����9¨��E)R���m�}�::�>
`���$IA0eC )�� �D!@�AC��y�}����.�����RʅU3)�SwJ���ŀ�o0yR,9��؎����51�qQ0���52��%m��7Ze��������uz��c�"��e����]�n�i$�i{;;#��cm۳�؞�u��0�I�
(����,�;Ze�����,�y�w77	@� �BU2$�`8I*���U���K0�_;�A�2��f�H���br�����k$�`�2�r�k #���}2U$(R%T�$���T�BIV3��֗^Ł��E4���
Q**QIf��,<�X�w��`��B
��=,vp�a��q��g��GDki�4�k��<v��uM��Uc%�v�-4�}�]��%m`-Ig;3���ŀjLt�qP��`SR��լu���o0֙`�w�oA��51P��ML��IE����u�X@o6� �n��}���A)Q@�STUR�u�X��x�w���y��J
��$� �|� �n���|� �n����BD\9�I@�}��SE �T�J��S-R��P!H�i��D燝�t�T�4��cO�b'A9 ��� 4N�#���RN;$fѢd��ںM��D� ���J��1u��(n�˷��Ӏ��PSC@PRP�t�$�t�@u����JB�F�J
nCJj'Pa�&zyئ��"��"�Jj$�D���%C�J)�15F�X����)��V��T0{��>�9�w�N����~O�����  ���v'(춪���]` ��k��`9U>WTդsF9�q/�)�goK$��Q�U�T$��F1����s��zٱY�q�m<G5�ۂ��`��'�.���V���n��nԹJ�Юt �a�V�ܯ#�+����p܄��[^ya�
r�:�t�ېɫs�%t���ﾥ{CR��-%�kY�Jr��X�J��(5m��۠�a��m��%>���y`6Vk( �{!���_}�n�o��z8��9�m͉�0E��n������Lm���Ӷ�O�v�]�D��wA;K�ɲvlc�.�v諣9w�
�ڍ���۞��1gn�h�8�6Xf��m��q�Ó)��/T�Y���Pg(�s��8����q=4��-�v���jZ7f�1'gp\Ԍ�8���gF�[��-<�X�&�郧IU�'e��W�PLA�R�m�5k�u#�G�Ҷ�9<CY�j�[�)A1S�Rr��*�Pz\�˭M��1�P�q�"����7	���":�(���n�	��f�*@7;��&�����6�ƛl�����V��Ju�vÝ�:v[���5��Nz
�r��<��Ų�g��@"M8���@q���n6���灗��Z��^2Oenm�7p$e���l��.S��u�8!m9[N�:2��mn����ltIٍ�x{slb�N�A�T�6X�"L�1�/l�t���Ib3��<r ��- d���-��Kś�ӵU��&�g��w6Mm�ۧ'7E��G��6���h,�d����m#9��bH�E��n�&���;�y=�}�Ӕ��S��\^^�Vp5�c=��ccpځ�C���'��]����n�c[�cx$�Ѯ5u���`�As�ضN�+�&:5´�A��[�F�[(�ZXv��
� �:6���2g�Ʊ�ސ�I�c�tі�d���=�C�V�V=�%zcX�����e��ܪtOl��kcn{tS�[���u��=t���mݎ��Ie�)j�ZJ٩��\Iw䷕$�`��?'�$�,Gh��(|�����Hz2�������*y�Yp���8ҥs�W��(-΄��\����q�n�h9��c���	�[xu;����p<�`ʞ�N��ܖ��;�����s�u�c6����)�-��;�X�ݫF�)b0v�MJ����3��lg�ūp�:s��\���n�ӥy4��̗���vOOh����럎b��e&�5�n���m٧n6����������۲������)���6�:�����3�n|rʪ�v:���VS�#PW]�t�SF�i�Xx����T����Ł�|� �i��[� ��u5�HT��H�Q`s�y�n�� �6� �n���3{�����
QRLQ3Y�{ʑ`�J��;33�n�[X��ـt���T�% ���RI�m���Ł����F�L��I*%�f!��*�n��y+k���w�� ߒW�}���*Za�����9ǫu��5ƺ@���g�u�/1t��v1�v�m�UWl�5Q��K)�;������y2�;ͻ�7Ze����u ���#Y�Zַ�u{�7˯b��d(
$RZ:N�Ϸ���}��uW��}��X�$��~?j��T*��6[i`�~�u�X��0֙`{�y��)b+i�=�n����%����@o%ـ{ʑ`�J��ڦe��	�HP�J�`k�y�n�� �6� ���7�������RZ&�S���ɪ;�H�m��S�N��8Sx���ҷlLx�P��ER�u�Xy�x�L�|����f �@��`�&�h������7��;�3D�\X�v`�X���ʩ��%P�ZWx�L���w��� }D�	�E��h�D?B�����������ߺ�zhSS
*TЩJ����L�ϝ�u��;�z�JTP$LL�3Y�-�E�Ѿ]���6�[���c��uB�Xݶ�R`ՔA�<G;z��G!�^��wj��:_S�nV��ۮ�J�D�,}�� �[���� ��,�:���EP"�p�Wx�no�� ��ـrUŀg�+���55��T�(UI*�=��0ܙ`���u��3��SE%��UL�if3���%|Xڻ� �Qa.��ޟGs���9�*d�J�*�H��������0֙`>}.�TL7���é	�d���r���;�C��͸����*W8�zzF��GivGt���lzs�{����,9�xѳ�)!ES��Y�@s�﷿�$����� }��x�����b������fk0�XjJ��fff�ޕ�`jK� �ݡIP�T�jdI"�3�w�k�s`ow<�;Ze��GR�U�@(�)+�]s�{����,=��[�+�y��o��Un*����pe�P1 ]a�g>D�Iݫir��:�Q�8�/��y�d����/n�S�8\�N�F���+�����ֵ�5��d�6��c�ub�$`�\�n��A^9�1��;lu��g���;��$۸�)�CO-e8]k�o]�2%:��b���m��u�G��	:dtf��[k<vw�����<3;H��Z3d몷Y�=���N�|'Rk����Ş���Oh��n#q;p�t��@��eq%��H�c��S����������=|hs�]s���U4R_!JT�&�`�2�1�;�5�9�;��3��6�i����**j�� ��u�U�l��kL��4�D�T�5%\\��崋}�� �*E�;�:I��{��l˾�[��*����%4os���X>n�u�l|�	w<���m�G��S�:8�a��K��<�p�g���8���c�u��m��ʬ�;Ze�c�� �\����y�s~�+��*��6[i������ım|����G�R,Ԗ`�H��e0�U�@(�+�]s������f�[�ŀ}˺��ڦj�����j�Q4����0֙`���5�9�7�yI<��J�dn�]���ƀ�����.���]�uf�T��bje��9��[K�#��C�.+e�7=�[���t�֝ؓ\�o��N�����~~�+�<�TX�՜��@-���5ktL~�REL
�U��������0�n�7xѼ��$EB�T��5Q`o�V`JlL������34<zݛ�u��t�������Hzb&�TUAUK0�n�7x��6os��v�5�"��%%V���]s����ӭՀ��US<0������:{��-���,t]��Ț�=��xÖ��"),VE,(�ǲ�]��W9�7_<�:u��o��F�g�**je*QQ4����`:�X7���V���⩢��
P��Q4� �����o���V����`='8�*A*aT����1�VmoM����}נ?$x��� |����|� �㦢X�!L
�U�ݬ�s��Z� Q��1-��ݛ�Y��UO���sź����n���t�B���:;��Hpu�1�B�Ж������r����� s�Հc|��ޛ���B�iH
�����`u��o���[�`n�y�7�ХB��EP��IIU�c|��ޛu��ηV�l6��%R�A8%k }\���|� s�փ�$�$�߿z�w�~��8;Ye#))�7s�ηV��;kzl����o�����-AR2�y����$������(ˋl3��79cY�KD�=pqV�۪RV^do����5���krln�W��.R���6�\��E�3v�u���W���XQ��8��=V�j��v��&8��C5���W����ϭ� ���1u�S��c]Q��6�+�ɘ2�(�nӁN�flh�Cn<s��T��m�r���"��m7Mȓ�����F
�����%�.)^��!YeQK�(tul�{u�{`L�뛓HJ݅����\��[��⠯!JT�&�`�7V��;kzl��0�'8�*E4J�U)*�o��۫�u��ηV��j%���0MR����>��u��ηV�{�@_>�$�UN��q�M�13�n���� Ķ�:<��`w�/�TI@+�DI.�_=��ݺݫ�u��a�Ʀ�&&aR&`
R��^����Y���Nث���k�����v�Z�$U8W�l���o��|���wU���'��(J��{���}�ϵ�3�"��@�
�|�q���o������1�V힤�����T����|�� �[� ǭX;�V��])�
P��Q4� s�Հc֬�ޫ|�� h��H�T)�J�JJ��`t��X��0:�X=��������TQU��kqn4Fț��@�R���n)��nC\�o�ʠ�T*�5J�լ }�X��0>{��%�߻������K�T�V�����y�t�u`�� �o+�O?�UR���
�Y�t�u`����Ѕ���YF�	0�4��tkX��fz��y:$C҈5"����2C�,�� ��"j�(�C�5h�$*�0���F�C,31"��2#0"d��$�4�s=L�l���X��1қ ���맶���h�m�Pa����K������h"�Đ���ó�J:�}�:b!a�ԝ(`��hՔDPzjq�-�'��:������f#&4JV�3v�	���Bw�����A�j�0n촩�J��&�H�c��c6m' ��ݷ��^bi�NS�4��Ȓ7u�`h��A���w��U6F��$��`�86_EUY�U��3�!S7��Y�Sv��=쇰<}N�}�����t��o��b��+� '�)�C��D:{6�
l =;pLG�LШ'z߀m���������b����Y�j�mUT(��܌v٠����] s��������ffff�;�67��T�EIRQ13��X��V����[� ǭX��Y;SRZ�s&Ei"Rtt7TBgzd�m�ً=^�c���5�:Ԫi���$4�T��j�c�M�b�wwvv�~呂�~�Bܥt�7G.�^�V�Z�=ڸ�7Ϟg����DԪ�P�a*U)*�~����j���~�N�V��:��P�	�WV�`[H�=�՘ǒ���ffga��HX�I��M�� �AJ噗]��t��G�%�A�Z��S@o�s��[� ǭX�\X�9���e����
'X���,jƳK�ء�ˍ���g��v��OKX��o=��mN^ܭ�ǒ� ��V��ӝ�ݛ 7ܻ0~��+-r8U!\lv٠�����;��gTX�]��%7�����7jn��"���b#
��zWE��:u��zՁ�:O*TLЕD��S`o�<�:u��zՁ�[�`{[&Z�B�*��M,��u`����u���^�Ϲ�uh^�F�%�9�����LW8�6�®���uu;1����OX�pq�p��fT�n.��8����Z��9�)Z�{1d{,�5�q�<�٠P�u�xTt�Cs�u��6���d]աI���d�M�����E��z�t���������]�;K�Z�ٮ�`�Mʘt���k/\��ճ�Bv�mtn}E�l/&��vjyΣK[<�X�kP��B�%�����$���,{�r,ݛ�y%�z]u�u/��kN�j�6����S��W��P�n�tT�RU�ϕ��[�`o�s�ηV�}�s
) �*�իX��6�j�G�� ��W������a4�<�SP�5��f ��M����ݽt=;�?p�"��D)%������1�V�����>y�s�h��R��SS$���1�V�����>��_=�9Á� ߔ��U�RM{#M���d�U :�.ʳ�A�V�x�H�MN�乩JUI)I3��X��6����=�����Dp����[�:��9�;�� ��8�*�`']s2��Z�=ս6��e�B�*��M,�:u��zՁ��Ł�|� 4�9�T�E
f�R�� ǭX�\X��0�n�<�C�Q)	R�J���,��N�V�简���������}b ܑEc�O5���Qj�ZX�^xK����涘���}�|�B\u��dr�������|���1�V����z�(*��
%EQT� ����1�V�����>y�s�h�!UR��ML�I+ ǭX��~|�ww3ó33]�r���uX	{ZeU)��R(�gv��w��� �mX=j��TW*QRP�T̪Q`{�0vg�wu`ݽV��>�W�g�v;$�T�R�(�N�f�D�����{e-������l�-F�ǈ���D�� �mX=j��޸�7Ϟ`�'8��H�L�T�I+ ǭX����� �mXy�)��(
�]%k ��q`o�<�6Հc֬��u�%A*����(�7Ϟ`W��7�W|���Op�Li�"U"�E��_xuW>��V�P4SL�35��J�vfh��� ��m`{�՘3�3G�����9�Z�0Q՟LA�mc;f�;��e����Ywj��U�ڗ\��J["�F�m�߻��s�q`o�s� �mX�EUSRL��S13��Xw;�|�� y����$�i��G��*���dm�V��9v`�*�� ������m`}�Bi�j�������&���=��`v�X��Ł���0N��UH�H�J$��X��uc`�]��J�3�{��?]�*sk���!-%Ԇ���3g�\��9����3�l�͜��3����)�����PX�҇��*��A���c&�Fƺ(�mЋ����E����6ض�@�v�q�Q]8t�+�v�������Z���S\�D���D��`���്�Y�g>�����U�����=	��m)�.Z��qg��� `�<kFv@�u!�k��e�g�8;���ؒK"X�����rX���D�Pa
���;�����Un襝G��-��vu\m亸r�PB��uj��ߝŁ�|� <�V�Z���tT��PJ�0(�J,���ڰzՁ�޸���
�q �QTEU,�sj�1�?L���m`o�v`R�"J���i�TL���zՁ�޸�7Ϟ`��`7�M$$�0N
�`��,���mX=j�;z�511)Q���Zy��r;�:#��j7����h;3hx���,��vsMɝN��M�m����՘��V�ʹ�۪�����5D�W#tr�`w޺�1�HY�K ���1M!� �w]�����\X��0Ó�UH�J�!$�RJ�1�V����� �mXy�
�j�T��]Z��o4�|�� o6��`���Q��JAP�,���ڰzՁ��Ł��?Oa��xߨ�D'T�ó���d�J���ێMd��z2�:��7���g������ڰzՁ�o<��h�)UD��D�I+ ��V����}�� 7�Vv�U4�T��L1U�`ԭ��՘���;�F$�1dOGu�� s����.�:�RJ(��e(�o<��Հgo+��q`{[U$W�)�UL�if o6�>ݫ�n�X�՘7.��"�{v���K���؁�6�ŵ�뇘�u�v*Ռ(��(�n4�VѺE��uE_�	!�mX����y��VK}�,UTL��������3D��0��~� ����~|��:�eed�ŀ�y� kmX{�X���=1)�)�i�	��wx������W���GU�t _�ZG  � U(�$���	�+��'���%UD��D�I+ ��V�uŀ�y� kmX�ULL�C�c�za�rf홞yرv�b2�8��k��IQ]x���DݡZ˭]����X��`�Հgo+�Q�ҔUT�M2�X��`�Հgo+��t��16s����-.B�Y+�{ �� ��Ձ�n�X}�0�6QU�*~I!RJ�3����o<��Հs}4�@�@���V�jV��-]� .��ޫ�?�_�uf�����W�?��3�qD�]�]u��"�*���f (�'r���y~�r���_����������������������W�����ᪿ����������o���;������2'������?�
"����?�EQ���Ӭ>�?������������W�l�"���i���_ɿ�����l~����H�?������O鿔������} (�(�*$��@�
L�
���J��B� 
$�( �B�  ��J�(��
$�J� ʉ2�% ���@�B
$�J,�!)�H��"��
���!!"�,*�2HP"�B�!(�!"H@ 0��*�!�! � H�	�����J @H*�H�2��!*��H��B��H�	0 JHBHL�@!% Ą2���+!**�$�!(HH*@HB�� DH0�K2��!	 H�H0�+(�� �$(�
� J ��"� @�! BB@����B��"H�(H�*�JI# J!*�� H(H�HB�(B�� H��!( �(���!,� BHD!�$�
HJ����� B�H� @�!(H���BB���2 C KD� BB��# BB2������! ¤� �����) J0��HH�1P�0����B4�B4� �!$�!$#J�*� �!"�ʩ B�##�BB1(�����ģB1 D#$�,�0��H2	(�	��(�0��� 
H0�$��(� H0(@�H2B2 B2�(�$� �
�0�B0�J2� ʤ#��($ H#
�00,� �ҁ0�� �@�(�����$ HH1(ҁB1#H�I�J����l�w������򈊫��������X�������QW_�ֵ�~���u��}<�������w�^��
"����������k��a��EU�DEU�#�����DU_��<���b�*���掿����ٙ��͜s޳;���|�߇��*���������DU_���ᑿ�g�������QW�}���*������gfQ���������g��W_������<��~��aןϰQW���������f���>�_��~�����EU��?��C}�y�(�������[�����A�7�����e5�{ ����� �s2}p��Q��9-�P *�  �#G� נ� h       �U� � hA@�4 �@ h�%�ҀHt:Ҁ�;��*�J(�JE$*���M�Ԩ)x   wB�Pt����(��`>��A����w0r��<�
� �}��`M����U�wwx>�m����� �r�9ڕV����k{�Uy�E[���e}�үm�`9�ϷM�۾;�|��>���`}x  �>�� U[ �(�u�x��6���o�M4��r����gJz���(�^�����iJ9��.`tS��4 w4�)�xP�� ��ҁ�{�z ��g�
}�� s�[�s��S���r��J^`iѥ��zP��Vm�����J-� .YOM ހ �@�P ��
��������`rg`=����}�.m:>��s�������[>���N j�}��q�>�{j]�yA������y{���
U}�;�����!���eЮ  �ϐ}@� 7n��=���|�>�݇#�`}Y�+�x����fh��;����{�B����3�ظ 1�6��}����}>	�@�������l��`-�>�^{ٴ >�}����m��
��.�o��Ϡ���<�y��}WU�s���o@�}u���������
[��;�8  '��<���G�f��>��c�\A˹�O�����A��tw0:o{�<    ��SmJJ�2�D�*��4�� dh ��O*�*i���C@�Oi��oJ�@  S�j�3MUSM�ɐ�"B�*TMD2��������l�_���f��pΏs��u�UQW�w�Ut"�
��U�*�*��*��?�TUS���S���a���?��a�t��y6JD���n��U$�_�g�0�������,�G,����~ʵ��q	u9��^i��Ke��4��P�R]���j�k����4K�a%�w5	u�l�6HB�Bu�	$�1K�q��v�C�/^�	t B�LY�ZB���X��RF�-!,+��ןo?h��P���J[w����|#�r�g�� �-��"����ǜ�B�,%w�y��$�KK�(@�Ņ&�`^��$y��e	r7`H��PfV|�(��PQ�ϴ6u�(��pԯ���f�:}�uZ��sx+���Qҙ\I"~�?ѥ۠��c�vn�ju���"�ke
�\H$�~B���cLb�#d����?a��:H0dOѧp���a�%� GT��!N�Ln{�Y����BX@��,ЗB��YҒ'%�8\8ؖp/\&�����Ѕ�Tɭ��#~��f��t�ޭ5��TR��Tp��\�Aǃ浇�8k��w�5܅?\�1a!�u��$�O O�ᰄ)�&���2��6���B�# �e�@��E�9�\A$��� R���������(d!�P�!ό���۸�6�;z���%�O�M#C4��p�rhI�i���_��c?Z�ܛ!d�M��1�"BHٜ�������j���w�f?p�I�f�oF���cȲh�Lt<���
F����J!,)�(B�.�H2V�ЀF�+̙�%ɨ��"�RHbH��j��e��˄.CXę�!a[�A�:6p5�~����3�����9�{c�.$�K�hŃ��ԕ�40!X��a�s6�p�5�aYI�|g���aX�#HHHIY��s؁��;��˸�^c�h���]&��
JZD��J2Bh@ -���8�9,�Lt�uʜ�����ad�,$�����0%aU�B`�r��Ͼ!p���p��HƘB��ς6)HY��H��5�C2$��I@!Й?��1#OߍB�XđbJo�`k{ֵ�/��$8YO����/T�� $���oa����IO��2J����'��m�K D�
�a0!W
?f���&�hu�n�;���K�U#B	I��f~9�����\\
��\����#G,]�B�0�&��j:]�a�fA4��ͤX���H������h��� ��nBq$8K���%��#�Y�x0�,�����\i�#T�Z0��\!�7�P�R	i�$��	�UH5

A��k�Y`��"bR	\4݄�l�/gXK4�9Ì,�Y�Iq%эH1bI V	@��c^b�#ӓ�_�yf���O�.�&��~��߹�����;&	(�	�A�	��B�&�}��\+�����_ŷ���Mj�F�R��+��*@� FI�Xy�xh�A��,�P-@� 1���2��a?�����]NfH[�s��O�8#H�r0ֶ0��	��$!C�t�\��T�!Lq�%d���K�������f�����r�B���,6C5e$�:h6Y�%���7����:9tl�����#p)���K�ټ���������!�u�iI�S����Yw���0�d.�u�Q�xB��6�d�JJlu�I�a?�.���FFXW2h�$��CR�)�%�y�g�~k>R,r������u���2��)GB�J`�i�`Ƙ��kZ0�)�`Mh�B�F⛅Ѷo5
�U @ȑ!p"R5$$�4ˁ���y��dbNh�\4ī��4m���¸�J�����
V��3Z�IL�aMF�h�!�0�4���,
��m��G�p�c���M�,�$$	a
KBR�.$�%�.�M��
��h m��v���9#!�+%�vv<9$8K4g�'d�k�F��bcZ�i�L5�d*c�6l�
�!
�&�k�) �E����U��1-�2޹���2Vz��6��	���	%e#�!H\��CMwXVw.f�謴�K8�;i�Bp���%�q���$>h�@'�	C��#�X�^i�7�0!3[ω�RO��-!M��	!ZP����ܒ�	fb3.�X�FI0XZi�BC]]�C�ߪ��U��cV��s�u�
�_>����6p���h%4Xi1�85�6XF��R��� ��aHS
B����XC]g���s�C���3��{ۜ���"I�.�`R8nGl��D��q�_�f�~��ۄ��0�H�S�!~kH�S�J��
�+��M�;�r^o�*F�!�8�S4���.i�h&�L*~�~	��4�X�!�M�g74D ���8s[N�1e��\�6@�o\va�|2��#� �����f�@��7,`C4C�~4B�Oߨ�	!BA��`Ҙ��$$�E�.&���y�ܗ�8~$��l�Ffa'pi�F+U�a$��%Ym���!FA�1����I��A��af?�Ce�JL�#��8^m$�at���ŀMl���z?�of����L�c$1���[�%�C��]n�R~˪s��P�&%�W	���%2r�~i����7)1 Y�R�)�����7n���)
C!xsi*�h��I\���>=���fl1!�����h��B%R�cL���\�S	p�-�����9��P��<#�h~0������S�B�RIM2�A�
ŕ50p�?���0����hM[��!��ai���l�����~ԇ�.2����)�[�m�$���O	F)0H�ML�a
1��S ]f����З�d�-��.Ja��$�����Y�gn�o)%��Hqӟ��2�xx��X��y<�MỾ]��y�Y1.�F�Gz!�� �#{2h-&��dSF D�F�["�i�H�:ă���K�*�`V�Ζ���+C��
D�i�\5���C5XH��$&hY�������tm�i(`ʒ� 3E�hHbH\e!f�q�`�LF�$&�P�4?M}��~0��^��Ԅ�I �3F�7KM�8��8ĩ�.70�	�K�	�8殦d��tp��@(B!%���B:d`q�!~��$p#dH��i$�F�LP�G�%�KĄ����IȔėB�w�~�d-�9SGvN���	bCR�	�!�n�*JbA#�
D�C2���� B���,��x�Mc%�4�$	���ā9��W!� Xi�B��R�s�'!w�K#]�����-+�Mi�H�dCBc��!�	
�o�C,֫���`~Ic Ʉ
E�F�sN����Z,���������:9�$�(�:`��j R��o��(ư��d�<��l�~	r�9��Y���_����o�����y!�P�����S��$i�7RV\nl���K��̰տ"����q2��?B���P�Q��!.HB����)$�2a�@�LѶ"�ٲq!�
�
�bP�6�@�Xԉ�"ԅcCk�'!L!fas7�~Rk�Jo&������ߍ�~z�c �>���6`���,jW��g5�0�#ڐ1�	e�H��KeR�m!R����������$t:t�
�(B��X	!�@���4K��7�s�>�8�\nHLq%�����M�oE�����"SS%� j!��F\arB4�M��c.�1n0�[�B��#m����1$���%����&~��I�[�R`C���Ӕ����P� 81.�4ˌb��,[#�ٌ.!�
��X¬?h����xF�i��aIo�d��~���>8Jd�����"נ|�B�
��$IcBjğ�T�ܹ��g��p!R$8�'�l޲����2�X~�|�.�_ׇ�����	����0"����8[0�B����*¤(�
0H`��4�5�C	�&f�ɣWSDM� q!L�"H��`h�Ǒ(d�$P�D��I.&���6~�� V�2H���LѶ]�]g��5	;�Sg������c��6�`B�)�+�*��X���A�w! F��H$
�B,�I�Ib�CD"~���/V�~ѳ�m��\e��62jB5� Is|�$��C��]0$@���������㌸i7�A�4��h���5�g6JWE�ų`iRP��󅄎h�2�		mdRX���a�H��+B�� �K��1�`29� D�4��LL�*�q�aG^Ja!r������Û����@�r��8h�����M��ށ�~��p�M C�~�#dc�	���hI��>6�
;��l�?a�p�,1�!�8p�\��y���eiR�B^�:s�9��}ꪪ��UUUUjU�����W*�UUUU�
�UT*��������U������*������U�Ub����������UUTֻV�YUe���B�UVت��m2��P6����˶�j��+�^�
�T�tUQ^�ćl5U@AD�u���F�h貏9�hk�;1�\��]�n�p����h9��^v�m'�.�a&]��@���K����m81[@T�	�RTlR�uN�A�6���d�@��1n��9�-�X��b5��)�V�:w�0p�[*ٵڝt��k3W�������
�mU]���r�*�m�ڪ��V�U�瓸�-U���,��5R�UA�JDK�<�A۫�UUU�s�TY�L�qJ��K:����y�J�FB�����49j��(v�uWR�UR�WUV7 ؖ��pRlp��jMЭU�Zv�`�$��K� W)�R@�Um*�J�/m++.����F�-����rnzU�ʤ.�n�Vj�jV��*���l說�*����U���
�*�	z��ѻuM����؉Y`h�C������lTUU��Yn��f҆�5n�	�G\.Ħ����P���f�V��v�n���j���,�U-e@�ڨ
�tU@N�S�6��*��u�PPv��������gjZۨ�6�Ņe���l:C5*n�R�sUuUyV�b���-i.
�kRUUJ�@z�a�n�eVHU �tVX��ăd .�UUPUmV�U*�We�ꫪB`*^Zny�����*�Q
�Sb��*��īUZ ��PVݹiv%���@n�
ڮVIU����V���V]�d��Uҁ��2��V�B�Z�gFy�-�^�i��W��� *���jH��Ԭ�M����.%x8��ڶ�U�� Z�����꭪���R���e���+U�iG�3Jˌ2��� ��n%R̚�
(
��U��#���7lenvz:��MU�%*�[��5v6��J�[V�ik�q����UQ^6��^eN@��*�U�^]���U�U6�`-"���Uj� *�j��;L�$4�j��W���UnX
�-t|��'7��d�-u ���tUUUR�j���W2廞d�'f��EZ����P��ؖ^Z�C毭��Bj�r�UV�c�;5d�5UU �R��N�E61K'8�tdht�@@.�j�O-�;k���ۦ��U]��1��p�[�m�5�*�T�X�]�����1�� >�g��m� �J���[����j����� 6�n��⺮����l���%�jU���(
����X�]����D���<�	ȖH��m5�J�������V�������T�j��+g$b(��Tfj�ꪫ/+*�dUZ�����V�en8�U����S��vS�p�q�UUUUV<c-b���V�Z��UUj
�
������U�Z����-��C��UUUPUUU�5UUUUUUUUUUUUUU1�8�*�T�f���ej�'�A!5P��]��s�������t������+UWT�U:����A�U�*�*ڪ��U� h�m�-��h�V��*�� �ʴ��T�U]*�MmV� �/2�,m�EO;-+�[��"�AV���UڭHY{s��:��kV�@Y2�X
��U��\bU�+jBj������
��x�ٶ��U�uUR�J�l��.Ij�U�-UT�����(
���T
��4�J�HMR�ڶ��s[UP
��+]J���ras��ܥRԯ5UQV4����UuKUTiUvZ�jk��Q��K۹��W5�PIR�R��KJx1��Z���5Ut�
6M���UR�Q+Z�wR��/-�
�[j���d�6%Z�����ݪ�U���-UUUJ�[PgUJ� � {FҭRjT��wu. ��"���}UUUUR�UT�V��^�*��
Z���j��v�6�Rej�GC/\0UUU�PV��54�V^Ͱ�='�u*���UwU��7�)��U:�^Xm㪪U[O�6*���s���wn��������9�X;i �iV���ZhW\�UH,a@�r���+-�� vE	Yz��۟*f���Nr�zB1U+.��KqY�zLvL��9^8�mTe,aCu؁�t�OwƙE�]�y�
]��{���\�q]���ԕ�����|�[Q�n�-�
�pI\p�mT�kUzͪ��������T=�Ů4�f�j�V����������*����\�R��]���QT����r�r�l����UUU*�UUT�9Z3m���&��U� �(�Pᗥj�V�]��T
�eP����/5=��R�U���)t�UAUS9�.ט]��\�^���,�!m��UUV�oCA�������s0 	Uj�+j��ꪪ�̶�b WkP����|<|�̪�s+UUU*�UUU�T�UWE�t�*������UV��(�UuTR�e���US������j�NM��O=�
�� �u֫-�V��K���9@������V�][UuUC�nYI ���ST��UV7p[@r��W[ j�j 
���]V���n�&���V���UT�)�+L��Z��j��1̮m 'F۩Z��j�ګ�����
��P��Q�6����V�UU��ljZ�M��V�HMmQE[PT�0ʵS�֮.BU���I�U��Z�}�۔�Ѷ�UUUt8�U�V���UAYQ��5UUR�UT�uU�V�pu�*]b�8�嶬k���T����*D�98a�ۮ��d���B��Z�n����꺪몥e�f��U]�a�ң��ڒ 6jX�b���z�u�KVL,$�����z����S��]nln�ݏQ�ATtswP9J��4�H�A�2��U,x::�(6Ⴊ���	������z��6��(X���]u�aC�O-)�
��-8N����ٮUP�V��ȪQۣ��4d�_!j��5-]��	vL���2Ҭ�q��uUUUT�W �N%YA�j
�TQ�C-�]UU� e����rk��䖪��V���lU �J�Ur�l��KZ���)M�T���G-
���uU*@[U[UR�x���EA������■��]]�悪���UU.�+�ʪ��/��UUQ�Uj��Z�����J��h���2�1�MWJ�Y���檪�U��5UU��Q�
��-������V����(*��������j�^�A	��e[U怪��⪕j6
��U��T
������@������UV�lm�Y)��� ÙZ�`*�U�j�@��������MUT7�.�T����UA@A]RSʶ�j�i\�Q���k�x(��*U�v�'�檪��U*�UA����W�˻HMU	k�� ��ym���c�s�!j	YZ֪�iAj��nV��M]*��9���+�UV5-Z�,�UīV�d���g�U��z�$MU*�WmW\q�UV*j��*�YZ��8#��9	�O�|?}���B-t�WV��Z�Av��ܣJ�@WU�U�	�`�8�ku/h#WW �a5�5�'�`�v���e�:h��'YW�s��ӡ�
��
9I��9�����誫6-�������P��v�@,lU���M�[Lp]*�j��-�ER�UQ�X%yj��V�QH�a�'ո��F�URUU,*�
�ܙ��Զ���ij�el��b�.5Ke*��`���J��LQAX�A'U��E���|�w��?=C�]�*�b�V��B�����o+�8e�jU��Z�UT�UUUh�T�UJw���[6m+�UUJ�+O#UUUT�U:�N��2����*�W������J3�ɤj�j��-u]PT�UR�@U[) l+J�P*�U*��Z�����)�60�T��UT�ٹ��UWK����u�4'DF� ݠ�J��\�������6�$�p]UU+h�X�m�������r�]P 9j��P��l� ��*�U�����j
���۞7J��uUUm��ڀ�ڪ���� G���]��Utl�\��5V�h�mST�D�T9������&y4�Ԥ�A�U{j���������d%���Uj��UU*�V��j�^4U�O�{ J3ۥ��ڪ��6P��R��� *��Xj��:����ꪮ�Z��B�Ci�t;,�h�@�*5�n�erb�����}�����Um:q�/mV��
���qM���_t	���p���V�e�Uyj����+UPEF^ej�W��*l���*��������#�U�`8K�[�����h�ܪ�U[j���Ѵ��:8��r�G=�^O�*TZ��g���s�g;���h���4�P U]U@���UT�ڃ��e:Q�UΌ��U,�@ȴ���:��J�Q��c�S*ʖZ���By�T�ɮGY��j��8���V���.)��UAV�,t���"��X�V�e���UUU���kj�̪�j�Wl��UUUU[���*���e����ګhS5c�UXĴ��꾪�]B�UUQ���(�9v�jt[p�Z������A֪�GW0UUh5Z��^j��-�`�$Z�`%X
�/QGl��uh*UUW��������A����n�j�V���jq@UUUUUUl�UJ�ò�UUյUR��UUU�*˰��kj��^i^ݔ&����wn�kUȵIR�Y\��6��
���������Z�jX��<���v`�@5j'7欖�"�R[s_�UR��$8��-"��?ʘ�x*"Pگ��|��Q���ҊuU1Pۤ��A؈\A_�0���T�|��C`qz$?
�A?�E��X&�t(@ʆ��
���� @�@b�T0�~��E����J�G���*�x��^uU�blTW��@B(�.h?����5�w�~N��\Pb��(� ��A �E?# Ab?  ��G��	� �@�/ƃ� �)\ ?!�����*#�qP�� ��h�D٭؇�P8�pQOȡD&��6
=���PE:'ȉ�F(���:"����|!8િ�T�)� �EW}��u�D���+�G�B�R1v�� ���?*��G�0Qh�}�C�C�@��z�BA ��|��آ&;F�P�B���@:�ѱP٥ �q 8 N(�����DT�EX@X�EbC�4EH� 邥@���?|
�*��|7��H|����������Љ��Q
"X��P��H���{֘۲	R�U,Uv�,Ye���Ԛ��(���f�s�������.7f����@�Z�<��G���v78������r�k�%(ɴ��/7���*Gcs�5�t%�q1��ԗ*��5�0	����얞D��3��8�.R퓋�� ���V�F�F�n���4�n��;)Cm��4���.�	�R�1PL;j����E��0-�h�후ʜl;Ѷ`�/:����$:e���1�9K��L�N\m�<��,����l�ŏ.� F�3���"�1Z�1ZH��f���l m<���&@5�biV��ڂzv	��t�m�̔iک곡A.sv�R��u�T�����&J��vm���Wh&�cë&�ѲE��5$rlM�	U���ns���Ldզ�ev�i��V.�#�/fD:ɒK�i]�8C<;���d�lv��8KXڑ�愳=\�٢*Z���YXY��;+WBl��(���k"��^�ܚ�N�d�8�4��k��@�-�-Ô�8��ݻ1�����������Ԫ{.J�c���Yԩ��bt>���P�2mtG*5V��f�7��pt��u�x�n��6�����+�M�a���NȬr�%�^ʠ��v�-�,�<��
f��.�K� �ݐ5�V�XmV��J,�@v�p���4�c�\�͊�j�������bm�UV���@���qj1P�cg��5�Q��%
ι KM��=�{yD��cU���H��s<q��hM�0<���t�Yty��]Z�:{���l�ĩ-�V;R6ָ7lp^{b#��|��_Q��9:度(@�(z6�h����M��F�T�����B���*Q��E��T�n�]r:U�vs��8�N�aF�O<�!�Н��#�nb�v���axn��aQs����ٔ�#sw)�kp��e���2�d^u�s��$`�y��(ql]�j'4�KZ}��`�8��F�s�a9�s�q��E�Mf=����T��FX�I!��EM���8�E:	��
�.����H����o.�����N*r��;JF��M�I�^ж�m���u�nѷ+- j4VUj�40�-c$m�ڧF!:E�,kG���q�:79df�vo3�F����ԧN�6}d䶷X�c<��x�3����oE������������y�J���*$�B�j��!�����N�vƧ7S��ll����6#�#�ݒd�R�-��gݔE]��y��N.�<���v^�)�.��h�i���~�zۜ��|��~��;��1�)�c�����+=�Uq"lO��~�����:Q����n���v� ��p�;ۑ`����L��$��*M[�Wm�ـw�"�����X�S��W@�T�MӶ������X�����qtԥ^��J�B�N�Y���8:����We�5�c� ��Ԏ�y|<�6�+n�o�7}����w�"��c�5l����hwc�`���������(��b @�f�`� ���}�r�I9�c�;�2��͵R�ڤ����l�;ۑ`۱��R[��V��M�Qb���nʷt�nǀw�e`����B!��ce&��;o �d��;�N{r, �v<�9$����v��輷&�h;��t�g.�X6���T�tgx����R�ud��,u>6��7n�t���܋ >�ǀw�e`�J ���ҫ��ـw�"�����Xݭp�Us�����+I4��;m� ��<��+��)�hU�/�Eb��HP+��3�5ٹ'����?^l�QP�tR���M���+ ���{r, ���e��E�v���`�{r, ���ɕ�w�c�a�S:��7�p١�[�v5G&:�6�l�UlP5kt>��<�N��[Sum6`�Ȱ����L����;6�$����N��k ;��ɕ�w��X{r,����e��lt���w�e`���R[��, �<�up�q���!ۦ����a'�����'��'���"�"����E����'���OKI�]c�Wm���;ۑ`wc�;�2���q��rrH}��}�<6�-������.�em�]Z2�e^�;w1b��	m���v:M4�_ l�x{&V��`�ȰJ촥���i[v�x{&V�u�X{r, ��x�S��.��&0v� ����� wv<��+ ;��U,n�m���6�`{�����'��ɕ�}�r�ٵ��|vRwN�X���UUn��W�n����X����QH�E?#��	�B� �qp! b��0!;�:eђ�槣�9x���f���^H��lu+��8{<]+qq��+�l."����LEC�M�<;t���\�;8�=�
�Z�z�y�\,�D�[�Z��F���d��n5[�aj�Ӣ�Z.��l�]{/�l�9��ok����ݪP��XU��V�u�Gy5�2��b�u��}���Nwv�Q5d���ꤷ������-<���Q��w�l��;��g�|!=�s�΁���p�ʚ�C���t甙�'�["E�|e��ut�o@�{�X�\k �nE��ǀ��l�L��!7M�XۮZ����, ݞx{&V t	(�T6��uv�m��� w��ɕ�ouư�	q��N�I��k ;ݏ �d��>�r��܋ 4��J]n�V��n��;�2��\��w�"��ǀz��UWw�E�W^{�LѼtN����n�h�,�γ�%�<3e�3d�Jn�#�x��M�@n����X�����|�w���6r6_�t#�giUo@��y���!��D7�U�Q �hX�p�>"	�I��zܓ��훒~�����vmA,n�]��I�;m`wc�;�2��\k �nE�w�I4�q����ӻo�\�-�{��7c�X{r, ��x:�i8�ۤ&�� �uưr�_�� �<��L�R$.�΄��(YK ����Yq�'��^�b�[��/.{O �ez��n��MӚX{r, ��x{&V��`��i�4���M6� wv<�9�$n��X�~k �nE�Waj*��&��o �d��>�k�\�UJ�eUd������\����T��6�v� ����� wv<��+ ���D�n�v趭&ݬ�� wv<��+ ���v22Ս��N��<.� �:ٳ���ϧ��Y�xYg��p��=j�	�t]��I�;m`wc�;�2���Z�;ۑ`�M(��v��ݷ�w�eg���$n����� wv<�UW8�{W{��M�Bn�n�����܋ ;��ɕ�IDIRm;t�����w�"��ǀw��7%O� N*�";����]�>�]K����v:M4�X����L����;ۑ`J��wjXƑc�܇l=�H%k�s���ܖ[)qq��%U-R5���l4J���]��>y�g@�nJX{r, ��x�.�O��݉�C�X�rR�U$j�����od��;'��n�v�n�۷K �/ ;���+ �nJXf���+j�RwJۼ ��x�L��)`Se��T9e2�N�]'m��2���K �/ 7v<�S�9U �� ���$5%�j:��4a�e�&9�}��C��ۺ@����z'�7rl����ksv�Q�s����Kfα��(��Z��+e0hK��rUЃ�1����yT%�Z�#+-�EbL��G� .a�n����V����G�����/ʧZ�t�Z�Ip�C��z�r�O3��tq/��N՘�y���4e�M-�hJ���RBQ�#E��\%M��(�pU�l�ɭ[5�&�.ji-�KT)/e�5!�7r�~[�~-�8\9��u�un����*Ee*�Y���}��|�}�twc�7�e`����6��N�V�`Se��ǀod��>�%,��Hջv�'m	��w����+ �\�����\�)QV­��V��7�e`K���6^ n�x[���]��J�> ��a�%�U���$��y��I�)�I/�:v^��\��m]1�,%H��]p��OH��F����<���t�On(i��K�Kn�]�I%����I�)���r�����t����6�و:vݶ���w\�`��mDx.��rc1$�c�K�KU�W�$��$��b769�_} ?����^���ߺo ���}���+�u�[��^���ߺo ���}� ��|o��l�gi(���>�$�^�x�In�|�K�c1$���W���*�ǵ��/�C,4]j9���v�w8���+��H��.��,ݮu�bt���6��g8��*�� ;�������� z�������x ~���g`�%�L�������s�m�����7~7������6���[�0�Wj(�:� |��=����x���b^���4F���?!�Mʬ��)F�H�Q���B�K��v���7ͱ.[~N����-�|@g�؝�}M~5�����Vq�!����'�I�HX�P��D��t3���&#?(���q"�!�c$8��f���lN�o!�d��P�?�"�-Bns���UƑ��́�
,�(J�w�T�� ���~t��UOȱV>Lں�@�Κ ��b>`Py����&���N�*D���j���Q1���.���?��^
�U���(:UuN�? �(/�D�@]�)��pO���� =@���R�`�D��߷�s��{� ߻���2�g0�䒊�+ĒKwc�䒗�,ė������{�۳�Cŗf�@i�� ����%/fY�$��`��$����$�ӓ���}t�fk�k�KhK������.�ˎ�4l�t��(��v�@���l��[��_���~�_ z��=����}'� w�����I���.�X�]| =����߶����� ;����w����rrI��l���!�ڊ/�I/+�W�$�����%/fY�$��{O} ���g8�D�*�� ?}�u�[os��&������"� �H	bh��U0�4��E1G������뛶��~/}m����4Zv��䒗�,Ē]�ʮV���Iy\�I$�ݼĒ�n�'J����S�7監k�9 ��cY3�G������|q]��)]���K������@:m��$�����$���1$�vaR�wL�[�;+O} �t� �ߺ��ofY�$��`��$��@Wx���줘��x�In�y�IE�*�$����$�v�ݼ��������6+�����f$��=��䒊�+ĒKd��H��=�+ R���O} ��z��I)�y��IKٖbI)WϸQ�%��_�u@�����a�L�M� sd����n�Nq��1�Ku����w�w1oYƋ�t�Wi^�d�تr�-��]���刅٬-�`%%Ł���ET�rFxCj�WN�s�f�ј2�u�t/.`¨&��E�6�@���#6�����f6�K�����c�7e,�S1((v�Y[��ǋ���k23���]�2�p[p�1���,�|���y.~߂c�����kl���R�a��Ph��m�:��ttc�sk��v3]A�8;utԝ؛�I-W<�I-�?�I){2� ?u�a��~�D�f(��x�IM���IKٖbI)�J_|�Q^�x ~���z �W�����w~�ĒS\���$����$��#��[^�l�Wj�ξ ������b�I$����$���1$�۸T�]�,
;9���tߺo ����@;{2�I%5�K�K�J)��n�-y7����9)��f�}��l�f�˹�,<Ur����f��fێ�e7������2�I%5�K�*��w����x�Kt<���H�f�W�@;�w�|�����QW�14�9)}�IE{�I%6G���s�l|v��1Ⲃ�.� u��{�M���>�96�����@>���| �l��v���`�L��@:o�7��Sd|�R�e��Jk���$���#x�b"QSx �޾����k�I)�J_|�Q^�x�In�+�N����3v�B�������\�t�EC��m˞�<�Bi�7��W�����w���$��)}�IE{�I%6G��%�׮�2�ڹ�d� �������^$�Sd|�S\�bI/�y>�7L�\�eO} �t� w������0���F4����r�s����1�Jvdk�J^�w�6�u��d� w���w�|/����S�@:n�� �^����H�QӶ��$��b1$��]���w�$z��� ��_} �xU��5�e#�-@nT�2��a�,�u&�`�[��2�/[�27+(��K��y����ާ�$���$��b1$���DIRh�S)��� ����@;׾������~�D�f%hݴ�$��#�䒑�F$��nF��$�wz> �?���+�"��W�@$s�$�����I(�Ex��9\ڮr��#ͦ�Y.��뜠n�tt3)]���O-������;r, �#�&�ŀ{��rl��w�+%˼t���r�8p(��q֍��5l0M��^Q��p��\�ʞ�~���dx�ذ����w]����X6G�M�� �k�`�"�>�e�16�Wm�m�X�5� �� ov<HS�V�����6��k�;r, ��x�U/G<�@�(��N�'n��`�"�=UJl��K�X�5�uQ�!!^�D�[�$�B ب�`H�!I$$���䄖�|���*�AE��tg�^M-�k��g9V��{Csec[�gH�!��^0�s�&
:^���N��kb%6C�c�6�<�ݐ�$ka��]��dn+��kٌn�4f��[��y�8=%f�f^صۑ�n#&�)�x�����HU�ͨSU�4�4��Dq���eYiYqeF��j�P� �pE�	s�<�\�ûY1�$GF��;R6�~����O_OAՉ,�e��(G�5��2�T�ź�KO�D��0]nlmڶ�i�hc�m`�y�ob�>���Ȱ�JR$�V�Um]�M�m�Y��\�$v���~���ǟ�^�^2��v;e�����~0	ۑa�$M�x�<��
j1�	�W"G)��r{�o|�ހ~���@&�x�9T��k ��J��]��I�+��l� �Ur�����?5�O�ޞ[}���st6Je�ĥ��i�3Z���q!��a8F�-BgVʄ dw�'9�<�|��銬v���o�I�}5ư	ۑz�_ ==�{�(~�T��Bm��Zܓ��]����1M�<`���@�!� o�M�o>�w$;���	�{�H4JA�&ӷI�j�X���dx~��I�w���*V�����X6G��ǀ}5ư�r, Һ��i5m�V�ݤ���c�=\�9�L�_ݹ�dx�@���Sj�ջ
cI"�+Uq��]�\i�t�:s<a�n�Y�3��ԛ��Ze[��l�]��}5ư�{ M������
j1�
�i�c���ob�W*������<�����ڔ+Qիj�b�� M��߾�<mX�D��]_��oWrO��y`v$�Ve�)�n�m�~K�<��?5�}�ذl� �JV�������������/�==�>y��>�|�6��CE��%��!����`�](h��o'��G��k<���\Rm;t�����w��`� }����:��F�[CcC�� M��ݑ�Mq���� 4��Kwm�V�ݤ���#�>��X{{ M��vr4�l�ݎ��V��>��X{{ M��NUU󚫕O�s�	H�	��ZR0"D	�d��V!�!T# # �$4���#Iʥ��Nr�U+�]�<d)�[ev�v�;m���� &���d��'�����[�����!�b���2sѧ�ۧ�0�5����^;g�����k��YI�+m`��엀}5ư��,wRIEyt�e;m�M����5�w�"�	�<�G���j�|m��ճ ��X{r, �#�;��u����M�n��ն�?-��, ����r,Us�^��ߚ�<��=�3F����o@<��@�s�������w���v�Xr������\ڪBݩB0��$��CC�K��,#N O�8��W"qI��~��JbYt��X�QM(~A�&��hh5��S���>`�H(w�����␦3?�@�mCPX+f���yK��D����..�_���F1p����b�1����$�Fa��`P��"�`F2��ߎ� @ce��"l�v��5-���aޯtJ2!��l!!��)A5��o0�SaL3��ц�1��ˢ����0b�@�ZH!���~�E�l����+)
��(�͑�B1�����H<Fp�1�a"@�(ht����! �"~m8~c� E#	�R�~:�p�����INp�w~�����U@WUKjkkv�Pgh�F���ک�tT���ٱ6W�u�X��-];��'RC���&��;��m�/`���Pd�U�\i��#��`�ݓ$n�zۓ�i�v7�S���ǅ�-��ng����ja�A�-Km1͇��Ci�r�޻[I�:ͬ�e9ݱ߽=����׮7ו�p��h;ZӠ�:�k�1���CX���+fz�t�sh����Nʙ6J�u��c����	V��#p�CD��׳Xe�M&�ќ !�������@��iȷTeQ-IY��lE��;ԑ��Q�P�N�m�Z�&S��RnQo�-�U���v�O�gf��a{t���Y��C�vO�\4JȜ�%����lҦm��+�R�eX���O+�n�Dvdg�h��@�Þ�Z8��Ge����x����F�ХqO[v6�ٵj��'�8���s�Wt�J�SěOP�AU۴Ƚ0�Z� �\M��d�l]7�홶&OG<���2M�{</" �W&��D$�hku�u�b�h�hƞMgN2��c��MN�\�s=����-�F��q�ӆ��i�P��7R�q��[eMv�eI8�
9��n��1��upq��ں�f����4��p:Ix	0�����iι;g(<�n�k�`@r��ѫ8�XE@ۖ��X��&�V���+��K<t-�xD3��������J��谛�,x�����EYQس��))b!BeJ�n-��Y\���s��q�5[�Μ7�W�7G �wu�b��F��[��UJu`k۶��ν�rVh����C���v�q�*s�.�
�IÉ�k���]���������s����`yٰvי�����f&)
hP�
-2bijY�.88��U5�Ms�o�� ��d�.�2��P� :�'G*��y����t"�YA�#n�eSKe0��i��ڠ�&��ܧ=tX.P�0�ږ��(?(0�h)�:�$���U(�/��Fl�_��2٫�Y�]kJb���V�7:u���d{ �
7���v�x��6Bv�J�Un49+�7'�(�A�K�tE����s�Z���N�wm��͗��n0
�n�B�����rq�,�q���n{Z�@A���nݸ�dĢ��y���&���J�CU�@`:svD뱙����y`Җ�����-�.�\ZF�	 u�k����Od�G�Nu�����A�Uq5��C���E9J.]2�0J=g���R��~b3�}e�v�Um]�M����ߖ���7nE����< ��<Ӳ��ݎ�����>��Y��~�=���`�~��ˑg�;���Vڢ���c��%�� &���U�~������o�?�`�R�F:Wl�I�+��=\K��x���}5�yoӒ��ǖ߿t
O��i�r���"�=U��w�<��I~��	�<��y&먹��#�١�p%9Cs��i�Τ$��*��:�nS�����-��6�v����~k ݹ�_�r�K������2%�bw�_��i��/!y��~9��Q��S��bX�'{�z�9(aH�1,H$��T�PH�&�X�]����Kı>����Kı?{���ӑ?���2%��=����h�ֹ��'��NJrS����^��Kı>����K�,O������Kı;�{�iȖ%�bS��~�Pv��M�+�'�����������iȖ%�b~�w�]�"X�%���޻ND�,�9?�����"X�%�~����<n�G��'��NJrS�绿j�9ı,�׽v��bX�%�{�m9ı,O��z�9ı,g߭i���Mn����fa�WbO9p�U�����U�<!vw'vGt}������
��T���^B���~����^Kľ�}��"X�%����]��#�"X�'���]�"X�%������h�Cd���^B������r(X�%����]�"X�%����j�9ı,N�^��r'�2&D�'�~�Ow��qō��O㒜��;�����Kı>�w�]�"X�<��*�`*H����v��bX�%�{�m9ı,O{��=�ֲkZ5s5n���"X� �r'���]�"X�%��k���9ı,K����r%�`D  X�{��n!"����K�(�S)��r[���z�ybH�N��u��Kı>��ͧ"X�%����j�9ı,Oǻ��/�A6�V�{=�b����J݉N�g6�OZ�f��]��p}�]�9�ղD�����ı,K����r%�bX�{��ӑ,K���ߵv��bX�'{�z�9^B�������ô�2;_9=�,K����6��bX�'������Kı;�{�iȖ%�b_w��ӑ��/!yﾺ�k��.c�/���B%�b}��ڻND�,K�׽v��bX�%�{�m9ı,O��siȔ�%9>��t��G
�G+{��p�,� ��=��]�"X�%����m9ı,O��siȖ%��O�B ��] �O�?�O}�j�9ı,Og��_k.��5����j�9ı,K����r%�bX?{^��r%�bX�{���ӑ,K��u�]�"X�%������W�MHY,�O;7p�;V;�爦01��s���ƞ`خH�X�,L�r{y�^B�~�����Kı>�w�]�"X�%���޻ND�,K������bX�'�zl��.���O9=���/!y?}�>nӐ�"dL�b{����ND�,K�{���r%�bX�{^��r%�bX�������xl�S�Oo!y�^N�^��r%�bX��ﵴ�Kı>����Kı>�w�]�"X�%��;��u�R�m�9<������x{;�fӑ,K�����ӑ,K���ߵv��bX�'{�z�9ı,�'o��0�5i�3�������O��z�9ı,?����?�v��X�%��k���9ı,Og{��r%�bX�E�?>=��Zֵd�ӗ�w�ڱ����-�l[�,�T�(�N��V��e�X��QI�X���z[��O�Q��t�].B�/5F�<��]��,C@�N�
����T_e���6��Em)f欈���bZjUK�����f��6iS���W)�Z��Hu[�u�a�ӊ�z�5�2r��E��{hY�n-�;9.�:��	�&_�M���7y�љd�jL�b�%��c�]��i&"��!��
��5��SO��ݰx�;���O㒜��'������Kı;�{�iȖ%�b_�ﵰ�_�2%�bw�_��iȖ%�NO�~�}�$x�쮚�;��rS���'{�z�9�P�DȖ%�}���"X�%���]�"X�%�߽�jm9�^B�w~�Jo�f�:���<����bX��w��r%�bX�{^��r%�X�'~�����Kı;�{�i��/!y���J}�5�b�e�,K�>����Kı;���M�"X�%���޻ND�,D�/~�9=���/!y>�}|>����nӑ,K����56��bX��Q����v��X�%�}�kiȖ%�b}�{�iȖ%�b|{]�e�\��2s��:ڙ򵺮{�4<j�@��}�|�k�v�`�({�Ns��s�x �[�ry��%�bX����v��bX�%�{�m9ı,O�׽v���bX�'~����Oo!y�^N��̖߰��n֮ӑ,KĽ�}��!��d�|����%�bo��ӑ,K��{���r%�bX����O�
@\��,J};��.]fd�CR��ֳiȖ%�b}�����Kı=����ND�@��u�]�"X�%�~�}��"X�%�~��L�\�̗Yu����ND�,D�{y��Kı;�w�iȖ%�b_��kiȖ%��ES"}�����Kı?����.D#���j�����%9)��뾻ND�,K���[ND�,K���M�"X�%��wy��Kı�0C���0LPt�E­ò\N���џGG���>j�&x�����~z�?:�{Y�.kWiȖ%�b_��kiȖ%�b~����Kı=��=v*r%�bX����Kı;�Y,��5.CY�Z-�kiȖ%�b~����?�"X����fӑ,K������Kı/�����ı=��}����7�Oo!y�^O��g�iȖ%�bw��ӑ,q�@"@bE��`L��;���iȖ%�b}���iȖ%�b~�����Pj����w���B��s�,N�]��r%�bX���ٴ�Kı?{���r%�`@r'��������%9?o���q�
EZ��r%�bX���ٴ�Kİ_���6��bX�'{�g�iȖ%�c;׿r{y�^B��v��mP�n3*�� t];2��X=Z�]�6l��B��9٧��U!�αr����{��7����]�"X�%������r%�bX���9ı,N�}��r%���/!�﮻�bj�Gq��'��ı,N�^�fӑElK��u�]�"X�%��｛ND�,K���M�"��,Oy���iӚ���k	�f�iȖ%�b{����r%�bX���ٴ�K���o�iȖ%�bw��{6��bX�'s�Ź=�30�B��jm9İF��w�ͧ"X�%���ߦӑ,K��u��m9İ>��"l��ߦӑ,K��ݲYw���f�kY35�ND�,K���]�"X�%������r%�bX��w��Kı;���iȖ%�b �����䟍i�e��h����[��Fś<F�f���^8[���k��k�y'�O�TV%ɜ���rS�������?�iȖ%�bw�ߦӑ,K��w�͡Ȗ%�b~����Kı?e�N��(5V�gg;�Oo!y�^N����r	bX�'s��m9ı,O���6��bX�'{�g�iȟ�Tȅ�?}��vj��	�����/!xX��fӑ,K���o�iȖ?��"dO{_���ND�,K����ӑ-�/!y	�w}���n��w���K��?{���r%�bX�ͧ"X�%���~�ND�,K��{6��/!y�~��ͱ5v�����ږ%�bw��{6��bX�'{�z�9ı,N�}��r%�bX�{���p�%9)��ϟ����Gd�U`����nVpp��GD�\�L���4u�88/un��`x�0��oα�}�rVb��gi�39���꣥�tc��t�RöA���n��6�G�p�3͞J$h��.�e͸$�{���At<v�fOv�}Mk�ި���wn;Tm�D�sҋu���3@Qƭ.������j�1�c��`��t/�$��yi���`+Lr���%�ڷ�]�Y1�O q�m��Zv(�gXk�:�Y��e�V�s��xrS��������w���,K��{6��bX�'��~�ND�,K�׳ٴ�Kı;����f�]e�֦ӑ,K��w�ͧ"X�%���ߦӑ,K��u��m9ı,O���m9ı,N��K.��֍k&f�iȖ%�b~���Kı;�{=�ND�,K��~�ND�,K��{6��bX�'|vM���������^B���~�o9=�bX�'���6��bX�'s��m9İ?��̉����6��bX�'�yg�ݡj*����w���%9)��{�M�"X�%��｛ND�,K�}�M�"X�%������r%�bX�g'����ዡ.͙�ʳW�AnKU�Ê��Z�%ٝ��D��1k�5���mI�
FPʟܟJrS����}��'��N%���ߦӑ,K����{6Ȗ%�b}���iȖ%�b_���칗Wk)�u�浴�Kı?w���rLHP�?�	T���	��(1��+`�R*F�a�+��bX��[��m9ı,N����ND�,K������%�c�~��_�Zj���7�Oo!y
�'�׳ٴ�Kı>�w��K�`�dL�������Kı>�������/!y����71�e2�*�x��bX�'���6��bX�%���m9ı,O�׽v��bX 6'�׳ٴ�Kı;����f�]e�֦ӑ,K��{�ͧ"X�%��~���Kı>���ͧ"X�%��{�M�"X�%����&jap�Ff��w��8��*Z@ʓj:�uc���T���;99�+�۴��e�6wy?�%�b~���Kı>���ͧ"X�%��{�M��*@T�"X���{ﻼ��%9)�NO�����j��]k.�v��bX�'�׽��r%�bX�w���Kı=��iȖ%�b~���O��dL�b}����٥��l����^B���}�{<�Ȗ%�b{=�fӑ,`H��$iB�M���iH�S!z�j�.Gg�������"�m�C����2
�+9(^!�� !�l�*JK��x���DbJ47��ކ
S@~������*�RXȑ�0��HF,�mJKFXR��?ي��)�ViB*@&��I,`F�F��p6�4�m��G�i$`S�1>	��~c�
`J��
&�®�i��(h�*~��G�Abm:�`�t/Q D��E���S����?D�7�o��Kħ*G<�9_�r��G)n�J�[��M,��Ѵ�K�,Og���r%�bX���z�9ı,O��{Y��Kı>�}�iȖ%�b_��sٙ�W55�j]L���r%�bX���z�9ı,N���]�"X�%��{�ND�,K���6��bX�'�{���s.�:a���U�.�X:N��4<��GN�l<7&�+�;Va7D��Xu!-eux��X�%��o�.ӑ,K�����"X�%�}����"X�%������Oo!y�^N��y�Ս�S*��kWiȖ%�b}���ӑ,KĽ���ӑ,K���{�iȖ%�b~�}̛ND�,K���.Ofa���Y�Ѵ�Kı/�w��r%�bX���z�9��@XdL����̛ND�,K����"X�%��ݲۻ욆�Z0�Z�ӑ,K���{�iȖ%�b~�}̛ND�,K���6��bX�L�&}��[ND�,K�:M�L
جh�S�Oo!y�^O���t�r%�bX�}�p�r%�bX���m9ı,O�k޻ND�,K�z'�ݽ��IU�0!,6\
�1�;7f<�����>�8� �v�h��%�t*n�Y�d�~�bX�'{��ND�,K��}��"X�%���{�iȖ%�b~�}̛ND�,K��s=p�CD֡�2K�Ѵ�Kı/�w��r%�bX��׽v��bX�'���ɴ�Kı>����ı/����M\��ɩu�3Z�r%�bX��׽v��bX�'���ɴ�Kı>����Kı/�ﵴ�Kı=����˩rkYm��]k5v��bY�"Dȟw�߲m9ı,N���6��bX�%���[ND�,K����ӑ,K���=�F�.�sY�BfkSiȖ%�b}�}�iȖ%�a�,s������Kı>�ӑ,K���jm9ı,O�I�B�*'��"CA�b�4!�V��P�ÓK�m�{�|R0�,��UQ�$��Hޙ\O�!�8w�W���\�\���4&�%�;��ۯ����ʗ3�1���٫I�+�6I�:�����G�Ӱ���݋�lLd,a�!��[���m�P�a�-َ�,QW	�]����h C��J�/q�/Z�qQ��Y�sJ���J\��XQ�Y�<��c�`��V�br�)-�����h-�Ns�'$�O5��h�-�!�R l�n�d��綟[���SB�n�g�g�^���0�B�.�h�~�bX�%����"X�%���{�iȖ%�bw��56��bX�'{�p�r%�bX���[w�˨k!u�u�m9ı,O�׽v��X�%��{���r%�bX��}�iȖ%�b_}�ki�%�bX���oٔL��*���Oo!y�^N��޷�OjX�%����6��b�b_}�kiȖ%�b~����Kı?d���Y,�ˍ�kZ�jm9ı,N����Kı/��kiȖ%�b~����K�lO��sSiȖ%�b_��g�����3Tٞr{y�^B�}ߟ�,K�{^��r%�bX�{��ӑ,K��{�ND�,K�CW�]�RfWh�q(��`�]�
���E��.�yu�Y��S�۝�ȺXYsZ�r%�bX���z�9ı,O��sSiȖ%�bw���"X�%�{��[ND�,K���֮��Z�-�eֳWiȖ%�b}�{��NB��S�$"@'��F�iA�mK�,O{���"X�%�}��m9ı,O�k޻ND�,K�u��H]j�Z���m9ı,O��m9ı,K߽�m9�[������Kı;�{9��Kı;�����k!u�W4m9ĲD�{�M�$��צĐI���n	  �w���Ky�^N���}�ٱ�4|���,K�}�M�"X�%����ͧ"X�%��{�ND�,K��{[ND�%9)��C���XِH����f��*���썕�C�8w�&��9PJSp!ڒr���{��|@t�ѹ�
�'y>��%9?~���ӑ,K�����ӑ,KĽ����9ı,O�{~�ND�,K�O��e%��q��f�5��Kı>����Kı/~����Kı?}��m9ı,N���m9ı�w�|h��35���'�����b^���ӑ,K������K.���[U�%6��lD$K������Kı?}�p�r%�bY�~��߱�L�Ѧ���'�����"~����r%�bX�w��ӑ,K�����ӑ,K [������b[�^O��M���k�P�o���B�X�'������KİE����ӑ,KĽ�}��"X�%���o�iȅ�/!y>�}/�q�6�Fk���B���0�wwYi�����UdL���\$;����jB�W5��&f�6��bX�'�w�6��bX�%��m9ı,O�k޻���L�bX����56��bX�'�������k!n��4m9ı,K�w��r(%�b~�^��r%�bX�w��ӑ,K�����ӑ,B����->�nlu��/���B�X�'��]�"X�%��}�jm9�ı>����Kı/}�kiȔ�%9>�����8�x�����9,K[�����r%�bX�}�p�r%�bX��ﵴ�K���p��2 -�K����Kı>���~Ġ�ns�����/!y���}�iȖ%�b����ӑ,K������Kı>��M�"X�%�����>��[0�B�i��Kl(׍q<�V��mY�L�-�[��0<}��{�e�zwh��3FIu�6��bX�%��m9ı,O�k޻ND�,K�����r%�bX�}�p�r%�bX��}{칓WY�0Թ�浴�Kı?g��m9�@���L�bw�����r%�bX�￸m9ı,K�w��r'�DNI�LrS��_e����i�u]�ND�,K����ӑ,K�����"X�%�{��[ND�,K�}�f��rS�������w_�!*��!��ND�,DB�����ӑ,KĽ�}��"X�%��>��iȖ%� X�w��ӑ,K��|x�/�����WY�6��bX�%��m9ı,?�Ec�����O�,K�￿����Kı?w���Kı>U�~A�TjEZ�U��K���:�4�[٬��|K�ۦ@��Od�#��}>3�]��P�����C+p�M���!n���ֲ�[��g�U�6W����	�޲���ݞY�D����5�p���)�ZFq��&ȼ��U�zۚ84�:��b�l�]&��NODڸ�Al�ףwv��ΠVsZ3��:.P�CRE�ĸ��q-��d��8醂��O�s�s���;'c.��3�2S��=����R�!G8�0�vè0����rn{\�I$��B���#�Vi\���rX�%���w��9ı,O��sSiȖ%�b~��iȖ%�b^���ӑ��/!y;�����]c�+��r{xX�%��}�jm9�	\��,O����iȖ%�b_{�[ND�,K��}�NE[ı?d��}��Xe��5��jm9ı,O��m9ı,K�w��r%�bX�����9ı,O��sSiȖ%�b_ݽ�f3Vjꙣ%�f��"X� X��ﵴ�Kı?g{��r%�bX�w��ӑ,K���{���Kı/a�g�6��4ڙ|���������|����bX�'������Kı?w���Kı/}�kiȖ%�bw��g�f�f��m��t3k�r�V	5Ư3�
$��f�p��!a}}����)ݹ�v���ND�,K�����r%�bX���p�r%�bX��ﵰ�P���,K�k��iȖ%�bw�����f�.j�Z��֦ӑ,K�����Ӑ�p"�_ �Tf�ı.��kiȖ%�b}����Kı>��M��8^B�����;�������"X�%�{��[ND�,K���]�"X�(�ș����ӑ,K��}��iȖ%�bw�Ym��MCY�]f���K��?{]��r%�bX�w��ӑ,K�����"X��{��[ND�,K���L����:ֲ�ӑ,K����56��bX���}���~�bX�%������Kı?{]��r%�bX����%�5	�3]��:�OU.�6;�hx����sk�{�``�5���ԝ��|L�o�ߛ�oq������"X�%�{��[ND�,K���]�"X�%��}�jm9ķ����N��&y�fy���/!Ľ�}��"X�%����ӑ,K����56��bX�'~�m9�/!y���|`G3h�je���^%����ӑ,K����56��c�������d�ȟ����"X�%�{���r%�bX�g��f��ɭal�u���r%�`؟{��ӑ,K�����"X�%�}��[ND�,������9ı,N�y��3J�ɜ�m�����/!y����ٴ�Kİo��kiȖ%�b~����Kı>�}�M�"X�%�{�,:]�Yc�CHH5��]#�kO\�;Y�$^8|��WO\*H�g�w��]4=�t�6��bX�%�{�m9ı,O��}v��bX�'�﹩��Kı;�}�iȖ%�b{��-�_��Z0��kiȖ%�b~����?�dL�bw�����r%�bX�￸m9ı,K����r%�bX��Hn�Φ��:ֲ�ӑ,K����56��bX�'~�m9�ľ�}��"X�%����ӑ,K���v�Y.��fkW5���K�lN��p�r%�bX��ﵴ�Kı?{]��r%�`o�J��E��!U@��8������������K�/!���V�$�3��9=���/%�}��[ND�,K� �����v��X�%���o�WiȖ%�bw����=���/!y���@K�1�lͼ+�X�1/Db\��kuk��5�
�b�P���;V�&V��je���^B���羻ND�,K�w~��r%�bX����ت�%�bX��ﵴ�Kĳ���t�#n��\�.O9=���/!�w~��r�"dK����ӑ,KĿ������bX�'�k��NF{9�&9)�翧OL�yss�͕���Kı=�o�m9ı,K����r%��ؖ'�k��ND�,K�w'���B�����>���ڹn ��jm9ĳ� dL������Kı>�׿�ӑ,K���ߵv��bX*��߻�M�"X�%��d�~�]CY�]f���Kı?g���r%�bX�{���ӑ,K���ߦӑ,Kľ�}��"X�%���G��@�3ZQ}Zh0�P6:D�R	��A�l�	�y&���H�@�GQBO��$R!��@>#F4��ʆ�!��?F�Aċ�6&CFBJ��C_ M!�����<^(-�b
�*
�+T-۩g-�J�	nxk1j��n{�Y;X�H�0
]�f/v���C�S���sZH���t烗h�Jd��ҍ�L�]���\����h{r�H�Nي�<:5�p�qF����$ܾaywf��N�(��L�M����nT���y;=��qD<h�� M�@��B�QS�Zd'���p�9�kuR9y�2��&Ҧ���� %f�bG�JÔƀ��u��e͒�+�ӌ-ŉ�Ӌ�5����*��jݶV{��蛢3�ٓ=NT���A�#[���l�Ի�h�� �&ΐ�9Tm�8��x�؝���3�9��Y���mĎۨ�g�d�̻��7;f���[��b6��
�J��D�1%��ݝ�a;eb`e܌k��7��y��RݘRY�qF����-H�a��@���I�۰`�<�.p�]�]���q�uݳ�@�m����i k�rI�;R�s�7QS�q=f��ڗ[�V�x��= ��@r�Mۇ���u��͞{���]�Uaݫ���Ydʕ��Q�N���T��<�i��5�S#۵�V+����=a��%����XŸm�����d�+t]@��M�t���o\>������)��#�뚫���.%�:�L�\899�-d� �Ϛ+WNC��@;\��A�-��nU��ć��06��0���A� �c;��፛�q�;Dg�$���#���ٮrv	��C]e$${u�$u\a\]l ���MqӶ��ro����V�]/5�W4�U�P������7	���ͩ]vڋ0�qk �Ґ\[Q�HH���v��m.�l�q�,�v��� ݨV��`�ɜhNݝ�]=�����El�q�m�N� aJ
ݙ,��`v;sZ�8f��ClW a�[O�ul��u�`�M� �{�k��HO{Z6���96x�� uhCО뙩��ˮE^A�G���j6�mElA`��'$�����$���)�S��t@z�B�E8(�mPJ�UOӜ��䜟ӾswT���y�(��L�DvX%�ڌL��v���$Z�JZ[�K���*��	)zI��S�٩������i7�iyCN��f�ڷ.��n���^��F��2���-���8�ᛣ��Mnu����7(��dc0mwf0�V,���^��ka�������\)��.��Sҽ�A4u&���"ؓ%�6,�Yn&?���w�u��6�Bڸ�I/��� �͓uץ3\�
�q�.���2�ua�9$�y,Hy#����Z���m9ı,O{���ӑ,K���ߦӑ,Kľ�}���?DȖ%��{�6��bX�'�'����Dk�;(��'�����/'wϮӑ,Kľ�}��"X�%��=�fӑ,K���ߵv��ؖ%�w�>��n+s��o���B�����ﵴ�Kı?g���r%�bX�{���ӑ,K���ߦӑ,KĽ�C�����9.���O㒜��)��{�ͧ"X�%����j�9ı,N���m9İ������bX�'���}���t��.���^B��������Kı>����r%�bX��ﵴ�Kı?g���r%�bY����M��]�3�r�h%��<"�zōi����5g5����`�w�z]����{5�5t�kZ�ND�,K�w~�ND�,K������bX�'���ͧ"X�%����j�9ı,O�=-�Y�L����jm9ı,K����r>@��>�ڇ"X�&�^�m9ı,Ow���ӑ,K�����l�����������z厱��9|�Ȗ%�b~�wٴ�Kı>�w�]�"X�X�'~��6��bX�%�{�m9ı,Ow�f�Mi�iֵ35�ND�,�RD�������Kı=�o�m9ı,K����r%�`�X����m9ı,O�'a�e��j�4�3Z�֮ӑ,K���ߦӑ,K�s��y�W�� ���;K�R���F5�hgǡ�Gg��Z�s��n�Q�,�uvF眈���2Cy���m;#�>]���ƿr�r��]���� /���n؝���>]���ư�\0vG��+�I�G������U��n���~k ���q�U�UV.Ur�W+�N��nǀl��hv������6���9�qM�� =����ǀl�5�oj$���\I��0vG�z��qw���'������'����в�]3��D�L�ػ�Ni����ssXÓZ�����vE*����իo >��8���Ur�@{}�z@�q����t���6G�UU$M�� {}�M�?Us�I��Qy!�n�v�6�6?;#��_�UWf���{���� �u]*���i�|��f�q/o���y�#�a4B"$��`U�~^"=D����=7$�N�{�Y��N��m� �v<dq�{�;#�?s��{Z�v]ש�]�����I�2=-�z��1���7=4�Q�0��{��4;{F�.���g/�?{��zߟ_ ����c�&�KT�J�j��I�����UU��\��~��< �����ư�A)E�v�k�1�f N�����q)�?5�M��&���7J�v��շ�M� �k ��s��K��<ހ/q����wm�#�`����g��=��������w����F�tv��V�Ɗ�`+^������$��Oe�j��t�Q����j�����;+;O\���kR�Xr�ѹbM�4NÓ��	4��P�n�:%d5Ŷ;UoPp�d[Z����+$gZ���)��g��Ƌ�vD�t���U�ۢy��]�*N N�'
k�G���� t�rI�.��u�s��m\����6g��6���x��@y?��N{�'&��>m�7-%Q�G���u.Y
��ɗ*�t���.q��sb�-�qBUi�!���.ݦ���~0vG�I�UW�UUW;a�ߟ���V�;E����m�;#�ܪ���x����7�៫��W)"-(^^V���v��� w�� �k�n�� 6�[J�Z���Wv��U\�)I2Z�7|�`� >����7j۱�X�`�s���� w���$�Z�"�d���n��B���	0ݻM���>������.:0�s�s�Ξ�WE��vr�l�	� }$x�>k�����9>`���Ӡ{��p[�՗P�h�.k[�Nw��`�& +IG-`���<�U��?Us��'�����x��z����@�����	� }6<����h�v�ڱ���~��W��r���~0�����c�$�R���V���M[��f M��W*�w���=�׀ou� �U�!�|�av���hPŴ�(wv�t�'�r�<ͫ)���݌�6���9m��c�$�R��z�@zO<�7��l�]3�s��o���d����D��`���>Se窹ʯ�Wg��z���o��۶"�;�=�?� M���*% ��hW����f��}{��w�,���V��Лf����xT�� ��K�;��N�J���2���;w�|�K�7n)xw\0RK���;/��4Ն"�b�9�#iǛ<-}���w����QQ"v�C�R�u��E�W��ح��I~^����%�-���V�@�7n�Ս�� ��r��Ĉ��^��z�ۊ^z�
�~�l���n�j�0��^�^�qK�7u� �t������V� �I/ �uİ�p�+�]��Ur��I��s�᾿|zߛ�k�t�]-3�v����7u� 7v< �H�	���z��
c`���դr�s�a�t��'4��r鰧����!�O�ӆ����i���p�ݏ >�<{&��)e�mڵ�v��0�c��G�od��;�ឪ���z���n�)۫�v� v{� �Ɂ���� �O<a�S�o�����{&�� ���{��W����G�OZ1�uv��0�`��y�����$�ﻻ7$�ʤO��T ����ٳ1�,���,n�V�ݺ������1�5��;=ùK�Dن���[s͑�*cN5poaSezB��8����ms�{,�d�R�� 	vu���ES��q��L0+�3D2Mp�hQ���J̖��	��B3%i�##�׌XC��=nFݬ�sp��5�t������t�	n!��,dշ��l��S0��J���R��
l�M
�XݝZh{9�rs�q���JOda�R�1��@�=u��Z���8[Qe�Wi�
@\y�c=�]��l��~0���1w\0](Z�`ҶZb�V� �dy�q#�=��6G� ���#e��^�t�n�R���o ��b0�`u� >���Z)Wv�ӻ�l�����p��� �و�7�,��m���]&ـM� �H�	ݘ�w\0�m�7h�U�Âc�F��Ey�����u<܋�\.�~�_s��~�.Z�����}�<wf# ��7\0�h�T�|v��;��	ݙf�W�V�,zDz�������=����ǀ|���ARN�;V�m�`�ᇪ�#���6{����n�]��vն`��I�و��_��W�{���
������1]
ـI���W&�|���?f�`����:�T��r��la�X�\ʬ
�&�@�#��6{8�Bl�rs��-�p������O~�`��vk��W���x�Y���6��sN����þ�'%�������xݎZ�7�,��ݖ��vـn� }6<7��V�ݪ�U\��"kb@�6ҔdD�q'�S]�$�0D�@��'�t�@�tmQ����
o�5Px��^!�������T��f���{ q`�b�c�1�7�SP���N��(f@+p�JJB��3��e�!��LO�:u� BHO���@��H�*%������7bb���1
�q�L�Wi�&�LCF�T� �k�~6l?(S�GL]7��U�	�P:&��B@#"� ���
�C��D��"��y��Ȉ`�t��:E���o.��χ@���.����y��;'C�$��J�r�{��6~�`��n���[��sŎ��?�x��@���$��s�^���t{��I�m��,gcf�d���g�M�����%�'�_U�Z�9�G*�b.�-Q�n��}��G� �u� >�?�\�W�;�~0�%ߛ�Cc�ݵm�{���H;�y��?�g�W8����Z��j�Э���׀}��M���v�	�V7hJݶ����]�g���u�'��k�r	��,X��	HDV6` �+�b�/ ݫ%���wV�e�`��w��Eݗ�}��uMTR�\�Ivv�9��:�9��Z�1G��v�'Q�-ݦ)W����·��G���?@n�� ��/ ��� ��������WƝ]��`we窹I������3�r���Py,�be;|m�����;�~��%'�� ��X}�C�-�����g$��&x�$��I�s�[��, ��v�Эc�ݵm��p�?W*������'��z�I��k�rN �)� ~#���U��~)��nj��hx���ll�e�,n(̷��a��u��
6FF˭�tn]x�n��F	���]�����S�2$��Z�l��۬����Z7F�R�É���kf8t����yb:!A�:������9�*�έf$�q��t�:u�����Sr)u\�9�S�ۅG�iKF�B���s\C�h���<<pXh�g��,��«�E���\ն躦�a�[n{sh��ND5�.Pѭ��뮍�\*(uI�g�$��gv�\�[t�'��}��ˑ`��n�v�
��Ս��wn��;.E�n��0�<�＜��Iɱ��_a��tβ���y�0���r�T��{� �_���AK�����;.�l����qI�����ˑ`��ob�+���.Z��˶`�G�{���o���H�`�� �6R�t����E&]��� �����)�絼���{��w��K�^�i����wm��"�7u� ݎ�������DP�ؕ6��e۷md���f��#�O�U
P$
"G`���������N����{ W۷j4����wm[f�������R[�X���:���ݛ�n���{��N[����@�\��7u��9\�7�� ��BG��V�I+n��xe�Xꪩ&x�	�~0�#�7u��#VZnݮ%wV�v{��V]��ر� u�8�5 �y��V$g#�'V�][�I�`��oc� }$�Uϐo��M��icE�whM� �� �H��p�7u�=U�H�ްWuyl\�um�l���xf�p@! E����ٹ'߻���>�iN1���:t����r��g�H�`��I�Ul�%M�n�v�6`��oc� }$xf�`�f�|���4�.��
��qJ^��8I.��X�XQ�}7��k��׻r�? �Lt��M��z~� �H��p�7u� �-�WcWmZwv��`�G��$o��I�{3�r�I_�%��U��Un�ݷ�o��n����?�{� �j�(�Wn�ں�hu�ou� ����7��N���KBY��� tD��'��?N����>��or]�kVe�v��0��~��{��7���7u���O�y��4�h�7P��R�{����
��$J����cx��^*�v�^f˖����>������n뇹\����0~��Ӡ~��#}�]�<b�;�|��n����Iy�竗f�
��Һ�ZWL	#�woF-ݼ��� s��KIX�;�v�0�p�>RK�;5���$���'�����ۻ�`)%���n���UUs���>)];�&�v�n�j��S�v�$�Z-��;r��v�wA�]݊N��xM�[7jq������8�:��(XPA]�<e�e�)&_X��Ɣ�b�l1�3���+۬����Cl,��[f���./�;��B��k��[]�y�݃FcbM�;Z����j��e��mY�S"�V�n�nM���#8�C�ַ�8�u����������0(�ќ�S�O��s�qX#v(At�[%�+R�f���E*�4���fN�M�[�n��	���7u� �� �H���\��V�][�I�`��oc��^ٮ�H�����-2���0	�~0�����%���$~0͔	Yyl\�um�l��+�/_�߯ ����`��l6�S���V����ٮ�`��I�GjYq��Co�-�1��RY�2u�	�]��u{//8�����V�ɉq1B(��-������C{0�#�;5� 9��!h���YsY�jnI����1�� �ǹT�'�� �G� ��-H$�eZi7i��`�G�vk���II�o��v�$�l`��ݻo�\�U~����~0{��oc� }$xe�jQn�5t��M� ���+�+��ߎ�o�ߞٮ�o���2ӣDa�G�:�SK���-cў����f��	��RjWC6����u�V�m������ ��w\0͔$�Yt�.����ꤍ�~0	#�oc���jYLl�c�Wv�����rO��]��؂�H���j�@�<_Ur�y� vO<�A��BT�v���M���U�RL�}�|���vk� Wۨ�aWCc����f ov<�\����k����7��� �����Jhvd�5H��Lj KqflǠ����d��L���F�tPe�>@ٙܐRR	��|���>��ou�ܮW+��y�/�/[WE[�nջw�vk��� �����y���U$o�)��&���I�`c����Uĺ�=x�?�����ui���l�� �I/ ���.VQE�I� !�(*F �HH� F# F*�	DD�$! ���D��T<
��znI��Ė��T�.[x�Ixf�`��M� �����n���)�8[���l���d�*>$��y��k�TL�r'nU�b7Ze;;.����`��M��W9��o���o-��~'�b�Q��[���M� �I/ ��z��U$�^�-P��V'm� ;��I��w\0	�� �Yn�m�v�m�W*���M������$��巽�J|��Jvr�m��������#�3�9W��p�O�F[���,�DY  �Gq�
O�6;P޷���#���/	��K.
����G����k�ő�L�����B��"�R,�,!"�N�`�z��@08$ ������R!�iq`Y�:%0�[�]����
�'��!J�#B�?#� ?-B)�!17�� @�LU:�	�0�D�**�IϘĄ��@����$�iE�D�diG4�ӴbI �M ��&U�[\FՉ"�Ѹ 3CS��rmV�d$�B1�#(��I�Ѩ���D��	�$^��-aX��>�T�mT"��j���eAۭ%���[d�oh)���nכ�m�u�</$��e��D�� ��pa�1`�(.n�w��y{����RCV^����4m��u�Ɨ4h���
�99�<��U�,��C1��G��,a퓜­t��٧��Y7%���N�w�`�}���s��&�. "#�N�`���ֹ@j]�#x���� \dn�,s�p�������l� ������LQV��r�GD��@A����u��p��Us&Z��'�Ԩ�[vAڏ]�@�v1�*�҈Ul8��*]�JV�#UN!��
荞q/Dtmйؐ{UU�ꆮx5@,��k��VZZ�� �dͰ��j���I��i���1��Iښ�Ǳ��3È�s��M��d����LVP�qr"����vWn^��6&����)��ǁ9�6�����S&���U���g�Q����#�:<"���J��Ӂ8w3S��O;�1dNt�n�=T���� Q1k��^ױs��"ᱳ�]�'8�)�S����g�r�*�/<һ`ePv;��m���k�dZ��8΋��z0��lX���L�`�2mv���,�l�u7\z��5��qsxZٟ6����jG60���� O-3n�<�� �m�&�r�ns��ن�p��*����,-pl(O9������ZB,֊��=�7r������q��z�]2r�:�GQù�F.��Q*���!t��m �n\��G$�c2�͓Z9�[h�PĴj]w\e����0'u��cE�����AAll�d8��b�Yde0�rc[����;�ح�����6�
nb7)=������W���i�ꥰ����D%��xD�7K��GE6l;mf�5��9 9�0*����r�z�D'���뻰��6�g��J_:�=����ث�؜��ʄn���t�3��5iM�Z��;oi��ge��[vBz���4�.f���,K�$�SkK�^���؝]�����H � �W�Qs�l(�?�����,��֫�\�!J���&!0���-T]�ٹ3j3p�"RO&jֽG���;K�%�{dXe룲6(�Q���v%�#v���c=n�Ѹ9:��2�5ƏX����aq	�F�iT�c��u��;��76�S�:yzi#���*�35&uNꬭ�뛳�еS1�
4�ۅ��6+���!j����6S.J�C�kkMP�99ɤ�q�a��X�;��OV.4iuc.1!%�J!��nj@	T� \H�&ـw�� >� }$�s��l=<��~_�,ch�v��l��ǀ|���ou� ���s��x���k�m�}�<{��`�c�6�Ll�c�Wv��Sfx�$�� }6<��K�����*��	Si��m6`��M� >�<{��ۅ�QuwJ��]*N�]n�-�D�)����ͮY,�j�0-�n����K���bv�> ��� >�<��ܪ����=�����;ֳZ�5�krI����Q��4����`�� >�~�$I~�z��X�BV�۶�	���7u� >� }$x�J�J��v���&ـn� }6< �H�=Jl����e�۲�ںM� >� }$x�\0�p�?Us���Q�2�wn�`�]�+��u��uȮGi��3s]�g�heG=9ܕ�w�۾�T��+��	������7��n�����'���q��v��;���`��M� >�<�I��z�"�N��ճ �?���$�%b���)�d��T�� Nw������7$�>�""���bv�0?r��Ļ������`{��~���ߌ����~v"ݎ۶���>Se��p�7�ᅷ�������Ĭ�m@��ӧ�X��nA�l���6{Npb����n�ؗv4�&���7��ou� >��r��^��eˢ�����][,M� ��z���RA�O<��׀ou�?$M�	/VYM�-;.��`}<����p�7��vHT��+��	��M� ���fV�W+�nrrs��e���>~?A��$s�[x�\0�2���͏ �M>��	-��3K���-�Z8	����ó;���Ŷ+c���F^�n$����kZn5nճ�'�����͏�W�&�� +�#�ҵCc�X�۬ ��< ٱ��`$���Ur�UU�����z��9��h��?_}�t�>�=��r���� ��� �v��-݅�4
�v���`I��vG���s�9�}�t߿:m�p2��S�y�v`���r�w���z��\0r��R���;~���]EkU�����I�vL�,��4c�	.�
6�:p!�nO)�'�绠��:�b����Aݱ�97�P�\$�q鑲�p.���y��'S`j�*�X%�����V_����+<��F`�$��3��6CR;Og�d�mѲ��]�P,�4;m�Dv�w:Alu[���btkT��ꅵd�4Щ��,-��A++��]t����e�S�B��v��Z�<��:vݫq�9�q[�2i�K�����N�Ӡ�� Oo�j�^���9_ ������R�Ƹ���;o �$���f̬ ��<��RG|{�����v���ۼv?͙X~��G}<��=x��J�� m;t�nճ ٳ+ >� l��=\R9���B�Cc�X�۬ �H�fǀn�ŀo~���?�P�����%�4�2��I׍RNӐ�.]Ŵ�H��v�˱un�)����ݻv��i[o�	��n�ŀI�+�+� ;�y���B������[˚ַ$����wcV�@�5q�;>�X�dx&ǀwuڲ����Z-�m��I�+ >�<=�U${�� �����e���i+n��#�"�/ ݽ� �fV�eH�Ƹ���+o �l���r�s��=�� �H��%+1�tЭ��N�tR %s�=;�e�v܋,�:Þ��Swu��������Ʈ����`��Iv^�u���N�!���N�{��U$���-��v�, ��TV
���b��f }$x]���ʛ6�H�l�`��� ��?.� VW+�\.��,��GmYi�n�wv�x�W+�׳׀Is� �fV }$x�/h�j�4
�v����`I��I��	#vKP��w"Q���9�n^Z5��X�\v%:�)tT�Or��ZYD��NIw\N�eu�ȍ�������#�"�^�{��!De�؝4��n��#�^�W*�v���%�,w]?��$l�@�1�Lwunһo ���^�{$�X�����I��v���ۼW� {���ܓ����f䓝�u�>��H��Tf
�y��srN}�m3:$6��C�+k �fV }$xSe��"�?Um^�/;V����[�H�섀ۆ.9��ӭ�*R:+s�vU�+�6�3��]�w9	V�ং�n�*π}�{��)���\?W*�A�Oe`z�E��4�m4컷xSe���X�2�O��y�s���/��.>qn���.�7ny`l��>]�����>��]"Rt��E���X�2��d�)��=U�UR�s� �^)/Y�Sbt�wCn��d�)����,M�^[��כ���A�k�Dw��ګ�-#�wA���2i�a��v3]���9���$�P3���-X�]p�RV:`N�ƅ�Q1S�;��͜{#'�Wg+=9T�S���0���nk8͋�g��y��1���>�n�հ��.u<��uk�ͭy�-�]��?�W�b���Mi� L�zƽ	�7���lm"(�D�ژ�y���$��I��������شC�/a�X�Q�ڃʹe�b��-�9�;u���-v�EŹ�ջwm�����;�ذ	$���r���N|���ﻠy����&H�7g`��X�e`.�xRK�;ۭJ�4$�v�؛X�e`ݑ���Uq//{׀n���
�uK�t66+;n����I/ �nE�I&V�Q�M�i��n�ն����~���r�f~���߿e`{��-@�.���]1j4�P�+)���:��� �4RVmmc���
��O�>�Ȱ	6e`{��M��wuڴ@N�;�LcM��2�V��*��@��G�m���O{��l�{׀}�៫��9ĉ�T����v��]������"�/Ur��K��ޞ��$���Zul�wV�;��?s��/_�� ��� �fV }ݏ ���E��[)��l�w�}�p�$ٕ�wc�"�/ �#j]�˶�i��I��l��sr;=p�Xn�ZؼƘ��Mb��2��I�c�iU�BM�m�6π������xSe�w\0�۸�
�66��M�X�v<)�����2�ܓ��z},�ȓj���e|��}߳rN~�]����'5�����h��ZE;@�°у�����N�i6��������$>i���N�~�``�F~��X�"�#	%�?l - q�##��L�B�)�Ɩ��bZ�c���8�)-!G��IZ�vp8|�P4r���H+
J���%%h���+�dc�c�џ���:j�ʻA4���h�B���q�WB�Ȉ��1 >QI�G����>���'߻�nI����6�&4�]��m�v�,M�X�v<s��U%�O<}׭�[��Z.�M�X�2���x;#�>����g'��6��v�s
��lֆ�����4 �N� m�Շ����&t�^0�YN�t˻��_ wg� N���{��'$����߽����5���uv��	���ŀMٕ�vG�}ZJ�2鉔��j��;�ذ	�2��W9\H��� =��v�u�Tn�m;he��X���/z{�������~�Y$�9���O-���wΔ�DS`�۬ ��<ܪ�W�W9_��~��%���$ٕ�}
�j���U��ӫ8��x���3���{]Z9�ő��]J�y��Vl�m�n���)����,M�X�dx{{Eڸƕ�:Wm]�x{{~�s����+�v~���X���E6^~H��unբ�ݵ�{��X�dxz��%����7ny`7�J��GZ���Y���I-����~��~���� �fV$��ӫ�;��i�o �l��s��V�_��e`ݑ�I� �m��`�"�J��s�M�瓜��|݆��l&b]�^����d�=��ӓv��M�j�4��\��/n���v�ƨ�����-�f�6L�cnΫcgF�μP�u�*{p��N�nv{��D�,�k�f`��s����9:��V^2,g�f�\�H7z�Cs\�Wv?.}_r��G���{�xA�vI;1/60�����.��0��sC٫�ge�K��rNs�A�������[R�V��&a��̛?a��k�i3����ԎX�;WLl�o�����v\��&ɕ�����W�<��x��y*�hM���[f6L� �dx[%��p�	�r�`�4�WE�� >��x{��%6?����l���V���v+o������z�	���&ɕ�M� �oKm$�i��j��7��~�秽�|�O<-��	���rR�^��ؓ3��(͹QćM@�d6l���m��vvə�g7$.z���M�+ >������	���'�#�%�N�ue�Zn���U:��U*���pCS޼H�`d��$�����N��m��E�^��~��8��������擑,�b��l�w��W+�����}��?{�� �H��K�7�Z�Jn�e�C-�M��2��#�"�/ ������(�\痯F�l�4A�����
\��N��3�7m�u%Qo��˥1Q�Y���E$�w\?s���=�{+ �U��ٚ���_-�;��>���{޾0{�����=�������۱+`�ڶ����� �L�.��ʺ$xSe�H��[�M]�M��`~��{�V w���"�^��{P�YtS��Ym�i���� ��z��_�I�I2�ܮW;^��g��:uV��v..v�.�mۗ�8{a�$t�ul�\���<qj�4k���2Gi�U_�?_?~���p�&ɕ�I��T+�_-_eۼw\3�RG��������K�7�Z�Jn�e�C-�M��2��#�"�/ �� NԸ���V�n�<�}<�)�^����,D7?�C�"Y���rN�c޺M[7i��V��x�\0	�e`�c�	%\i'@��LSۯHG`�1˶y9�m���Ga�Y;u�ү�s�>��vؕ�0Wm]�6?�2���l��}#�[�-զ�˦�M��2������{P%,�)�N��ai���ǀdx~���9IM������	6k-:�S���m��$x�\0�e`�c�'4�8��W��o ����W�~������� 6H�	U�(��h1 �XDpb��4�Fwgb�9Hԃˌ:��� �J%=v�����v���F�㫊�&`��d�z�4�V�l/ab#`1���{m��	\&f��nWqq����\N�UFθx4�������W-q�iѸXC7��,�
ַg�.s��k�.z����&V-{P�e�싼������1D��d�e�� �=I�S��,\`���%�S\�Ԗí���p\��[�a���� <m0J���#gW������V��."�wM*lt�m�Cl����+ >� l��s��+� �s� =�/̰M5nˤ�u�M�=��q ���6��L�e]i��:n�Iح� �#�7u� �&V }$x���.��V4�]����5n��6I��I l��H���ui���i��6I��I l����`�iP��ڌK��n\<n�� z�E�n�x�s����8��jx�b��YV�ÙAk >�<T���ذ�e`vj��&U��N�m�����"H��6I��Iz�=�z�뢙|.�݊��G� �&V }$x�%�ۭJ�:v˶�[��`$��>Se���ٞ0m�y�	����t�n���x�G�n��L���Np���j$xC:]lҰxʦ��îϋMm��I�V{"��d�_�u��!�7i�e�w�~�����l�+��$����i[�-�R���m�������"�^ l��#�����v�V%n�	�{+ �I/�UUR���*i�W��P���xWv^��*#)Qn���t�n����d� ջ/�s����_��ߓ�{���k;�Rm�X���x��e�$���� ���Vb-'tm\�㉋: ��F�ղ��;�Q�wr�O8�H]e�<7'h�,YZ��۲��e`)%�����m�M6`$��U$M�y`����p���"�,CM[��&�`o�X�G�w�� �&V���'c7i�j���~�J{�xd�X��J��߽x��U۠�
jյM���8`$��;ۑ`�<z�~�v�ȋ6��%s2}wI���8��{���^�T�C��*�ч�m��E�i��d�X{r, �#�~�w�z�t<���{e5��-Y�>v�X�G�w�� �&V&�-V[�ʻ�i��X�G�w��s�O{�X��� ��I8�!�����0�8`$��:�%�#���*2�
Ɔ[��0�e`�%����䟻��7$᯴E81x�19MJJ$�~�r :L0!��eN*9H� �!	@BO�%�@`"4���;a+��ă�i68�Q%�0b|���@]�_�Ȏ:�8E�����l� ���0��� b#�N
`�
�L�МEu���AV��� E�6��~O���kU��."p��! �0��>VS������x�궶���@�U uuPqWPq�Є�.������`eV-��T�x1ڷ�0k��ÞgX�P��ض};���>��PJ�B�%�qY`���Ղ�pp�s��km6�VCn��2�	�jS�����.Z6�]�z��<3X7���t�Y.�c��Hg�^��\F�ܔK����:�������e�E�� �,XE�b�Hᶖ��")�'��8y�g{ U�L��Z�h�ÜI�����Ez�W2�ڸ�r��ɜ�]�p��n�+k/ah�r���|�#�5���0�0� Q��F��
3�c魘&Ij
����w;��-d6���W��,Y��H�;2�mtmIf��^��$�V�Ol�s�`��l.'o3k�#�8waݝȩ��T�N1O�Jhy���8�c[FQVPϳĆ�سp�[).���G��J)��k��¸7h;H+wz�����jQ���zZٖ��!�7`�/"T�r����ć�6|�(�$�8�S�'�w�ٲ���ͺ�6ͦ��<'!���v}RV�U/Ih�Zq�C�0�(����u%q�4���ݞ�g�h�].���C�ɵ��\��SR�]��k�e�֨�[lL,�WK��D&��Z�6�Ov;��v@A.�V��2kiڌ����MN�;q�+�8x�kv�E�C�T�ږ؃��N��zV�W8����V��[q����,�܍%�����S��Zu�B����U���v�)�h�LDjE+�1�`�a������*.H�m�R6��<Y��Ϛ�����Ɵ<i��k��tT�5rqu][���8�3g(��7c�v���,&7Y�]X�h�g�;�B�۵ʭ^�Ԏ��ᕃ���69��iA�.c�r]�S�fp-:{��#����g���B�t� �v�:5׏9��a�{Q�&ďdx=K�&:ٞ���cMv��t�QR]@p���+*�d�>5���i���2��p�s��.{�йP�Su!k����*����>:�yE�E�� ��������t~ OȘ?
�i�I���m�S�t�a�D�B�i��ٺ��{���.��;,{�r�����$���ݣ[��/����8�:ڰ<t��:�e֥�Lc��xC�bu��]�np�����[�d+{�7�Xڍ�1W�.��'\'Js�v��u0�~���%�aa�A� 1!��&V�΍G�l]<7=��a,),b]��f͹慉(0�F�W ���������Ns\O�Lqsdy�\qb�W��ٹ��ɞ�����{�ݎ��R�ks6�Vx��<T���`$��;��Pnڶ6�n���x�%��`$���#���vT^B�@��շm��$�~X�2��\��$w}�E�z�	�L��-ڴ]6�l�6I��vG�j�^��ŀw�
���Z��Гu�vG�{���z�v��L�[}���n4Z�Y��&����ë��v^!�;�c0�BN�v.6��[!�.-�wM:v���<��� �&V }�+H�rˡ���]�xWv^Dt,!�@y�f��lܒw����G��ʪ�RGT*/RMؕ��[�v� �������<�v^��T�hM5n��M����g�����ջ/ �L��Juv�cm;v�]��H���x�e`�#�>}���]<D�\�SL7FY�J��G�6�fы�X�%�L�5�BX��ñ�ڶ�����,I2����U~�����~OE�)�u4Z�:�I�����Iw�x�{� ��y#v�G���iۡ&� ;=�H���W�h(@b�� �J#JCZ�]ﵹ�'�{�7$�~�Ĩ��e't�Ӷ� I#�;�p�$�+ >� ��I9e���펕�xw\0{����g��I���ٺՌ�6A�І�dф��v3ɮS���n�V�L��t4k8�qFƈ�hl�$�+ >� I#�;��oo�v5�536��g���������}�<d~0	$��7jS��۶�7i�V���:���wu� ݓ+ >� |WV�J`�v�Э�W9\�R�3��=��l��r�\�S���ŀN�Bݔ�nբ�6��ٕ�l� �^��wi�u��S��P�g�M�@nJ�uBI������� ��p�ˢMF���\�՝ ���@�^��vL�n��:L�v��:����H��O{+ >�ǀJ�$���c�v�
��w\0�2��9ʮRGvy���^�J�R�i��v���&Vݹ�$��d����m5n��ջu�wnE�uI/ ��/ ݓ+ ޛ8���)�L����;��^�u�ƽݝ�# T���ϵGL��g;m�K*v�t��/V^��\f(7lc���s���O\A�G�fPMc˴%4Cr������U�/]��+�]e-՘�����en����-�l����u�nćj n��s<]wbsy�8���BF{*(z{&+�X�Vu��D�&�����#��C���*S��'4ӷ�4/S��A@��sĂ���M,�n��Z����X�Z���E�Ą��˳DT�������o��/ ݓ+ ݹ |Wv�R�X!�ݴ���:����"O{+ ���uI/ ��Bݔ�nբ麷n��2�ۑ`RK�:���N֕��;v[�tZn�ۑ`RK�>�Ȱ=\�+������x�H��e't���Ixݽ� ݓ+ ���`ͭ��mq�vB�ɮ��i�Z嗃r������|p0Pg��nv�pz��ֽ���?�o�<��2��{�$�V�i)#
5��\ށ��vv�I'�NNM��n,�Ixݽ� �D�Aҡ�պ��V���ob�:����q.��,O{+ ݩN�j�[t�Ӧ��XT���{�&V�ob����)@����V��v�,��s�{�W�wny`RK�$�J#-P�ҥO���u+��V:�E�\��U+���=(�Is:� ��-��)�ݫE�h���&V��ŀuI/�U_ �߼�mB������t�7X{{�$��܋ ݓ+ �'2ӫe't�[XT���r,�U2_-?�j���ٹ'߳���JЈ�e������>�Ȱ�2���,�IxZTPT��&��v��&V��ŀuI/ ��"������;���6ġf�[�dsu7��ŤJ�O%Ҥk��#�AE�n�J�f]իun���,�Ixݹ�A'��X��u�պ��ݧM���%�v�,vT��>��X�]Z�(����n��{ݕ2��{ղ^�O���Z.�E��=Kg�pܓ���]�?_��ܟ�u��X5ʬ�ϧVݭ*"��6[m��7Xݽ� ��/ ���`�1���O�����>�e��b���
 �^��p.��!F��n��ជ�tg���%͸���������v�,�&# ���`]"Je�]1�Э��ob�;�b0�{��/=IB��I�i��wm`=�F�ob�>[%�v�,�"�J�cV����F�ob�>[%�v�,s�UJO{�`W�׬V�ۧv�46��>RK�>��X옌��ŀv�+�*�Q^�{/���qV�C��ôP�%L�Y� ��3L���@�;2^S]��B������!sJ�d8ċV.S�P��p<��#/Z�ŷl���voC�[�:�mƠ������!l�v;.�V�Y��<J�'��e{#ˬrS�#e��]���;Ufr9�q��f��s޵�d��RYp�K����)��]���NؗT#�df[3E��DG$�'Y�MSiiF2���0HV!�A1h�7-��N��;=
��`�4�`��V�FݝU��y�~�`�b0�{�^;vSe��˦�m�vLF�ob�>Se�v�, ���E���&�M� ���`)���{���M���u�%trۛ���I/���۠|���z�LF��u�,է�^�e��m	��>��X�LF�ob�>Se�}��4/���dvb�g	]B��X�f�m��5~��������^bm�J��s��	����`�ϯ����`g��X�l �SLi�Tջh�>��X�È���S��,�߻��}��n�7�b0ڔ��շN�:hm��|���>��X�LF�ob�:��m)@�Ҷ�v� ���`�1ݽ� �M��N�R�)�������>�1{{�ݗ�}ۑ`��Iw��25�x�y�s����(��J��M+j�Eh�JW�\��F���U�*� �ob�>[���r,��M���iղ��4ƭ��/ ��"�>�1{{��$���L|.�&� ��"�>�1w�qp����8�?k$$��ȹ2�k�I0���~t�A�d�	��a�;���7�!i�|���$5�C�'1So��GG8R�$w��*��l�:F١Ӱ�!�2�d����!���$`Ya+��>�)L)�&�W��&�2`� ��0 !��Rc��S�$$�--�Hm4§&+�`SRKp>��PJ
���HB`H����/�f���"BX�����!#
IeI?p��
�Rvࡤ^ �@�� ��QnI��,c$ �abX�K!���֏��T�V! F@�ZB,�ab@��IR�M"a��?6�kKH�#: gH��X~!���HRRXĉ4�D���P� P. �LN"���I�TJ���:��:PX/��Q�@�����d�e¥;t�+v;�����UU�^�/}X��,�v^��Ns����-��{��Q���ʙ���ŀun��>�Ȱ	ئV v%��J����+2���j8�W�5p��f_ug�����Eԛ�g+y-)tEK �ݗ�}ۑ`�L�UW9ʮ|�v���G�z�X!��c�xݹ;��;�ذ��x�2�aM��v;�� ���w��`-�xݎSkJ�-�ۤۦZm�{{۹'/�w7$���ry���E��%	 IRc 1Hȑ#��H	 �H��)a 0`�	A$)P*E�������nI��ęrӫe;�i�[X�l�����$ٌ�>��X�t��gȵv�c�E�Kt�n�`��s��G4��6�n�r�W-=r�ZJ��*c嫦Э��wg��	�1�ݽ���r�A�'� ���N�t�&�'nݺ�'d�g�UUĎ��,�O^[}���'�NNI���{��!�����fճ׀|�e�wfV;&3 �����RLwi�m�� �n��>�̬M���ݗ�us���@��v�v� ��2�	6c0�v^�/PA��K ) 3���񙎪��<��k�}mz#���ּ�z�nې�����Z8]���V�sIØ74�͓8���y����CŻm����u&Þɬv�UD۶�TWvN�;��Q�4t��D*�����9�ɇ�B��޸���ag��6:v���i�u�;�^�a�a��rk��4�sm	��ە�����۵��]v���Cc�R�R}$�$�{�m������[�v[�M[��uu\<��rl�E�6XGW��-Hj��L�Ga�
��{��z�˻/ �M��}ݙXSkJ��v&�0�ـ|�����x�ٕ�I�����G�ޠ���[)�ջ�v�����>�̬<��=��;�<�	]"H)�1r��hV� ��2�	6c0�{�/ �dU):ӡ���n�`l�`v�,�6^�ve`H�:n�M���t��;R�ģ�˫7Y�yp�NyNl(�����.�6\��f�ob�>[����+ ���}R��Wr��M4&�v��ݗ����A^�����͛�w�{�M�9�>��:��R��V�Wm�n���+ ���}�ذ�� ��­աݎ�n�	�1�ݽ� �n��>�̬ ����v&�*�l�>��X�v^�ve`�c0s��W���1�c3*��A�`��n�Z;)�y�9g첒p;Fظ�kW��d��/3���Rz���+ ���}�ذ��$��j�+w�}ݙX����� �n��$�*�զ��m��nٹ'w��ܓ����sG�c��Pi�z���V�"BCT�n���wn��{�ݗ�}ݙX�E��}��~�"%�[}?~�����9�wg����啀}�ذ�Z�wj��vb�v�r��$燵������6%�8�.jjj��;;�..�v��g��ٕ�}$YXݽ� �n����,*�Z��&� �d2��{�ݗ�}ݙX6��-4Ӥ�e��Xݽ� �n��>�̬�"��'d����]1�ջ�v��ݗ�}ݙX;�ݛ�H�$�$�< �	@C���w$��v�j�u1ˆ�En���+ �H���{�ݗ�}����_��_�Fg]3Y-ئ�����狜h�M���/2�2%�Y�2t\��M�;mۯ��啀}�ذ��W>Aݞ��5��&1�uwWm�u�}�ذ������>�,��UURGk�u��;i�4Ӷ��=x�ٕ�}$YXݽ� ꮊX���һm;w��W)wg�����V�ob�>[��]���C���`�^V�ob�>[����+ ��s������\5�pU.��'6�ڗ
��]�=�*6Al�V���K�)YH�ax�	�� &�kFZ`�u���[�^r�2D����i���B2�=��p�Y;����ٸwcWb�Tر�e��֜�� ��;nڎ� iJ�̤j݈ծ�
]���V�6��A���{.[T��c��,�`����9�h�\F��K�]Ki3-ˬ2ڂ���E�>����E���Iθ��rl�6���N�7N�{�����9v����zK&tU���-۬{s� �M��}ݙX�/+ ������ݪ�t���>Se�wfV;%�`v�,k�I4�q����B�x�ٕ�N�yXݽ� �n��6YD��vq�'nݺ�'u8`m�XWv^�ve`A��*T�j�*�m&��܋ ����;ݙX���)]
S*�N�k��tmk��i;89�v���(�ݦŢ��ù�7`��T�vЭ4�XWv^����'u8~�|��~��"����XRi[lv�rO߾���P~94-��XGQ �
�� 1	 2N�۬0�"�:���vTB���wLu�N�p�>�Ȱ���ٕ�kmB�cM�7vƓf�nE�uwe��̬wS���Xݫ�v��Ӷ��ݗ�wve`��0��<��~���E�֪�%�%p��Ԙ���������7����A�Ks����޶c^��WM�[���=��N�p�>ۑ`]�x�������[�۬wS��܋ ����;�2����V�U�i6`mȰ��,;�9ʣ��AB��f����rO�v�rN|e�����i���;�ذݙX��r,W6ZR��aJҷv�wfV;�� �\� �ob�?w杗��;$��Y�q�+rb:P�<����y�N9�E=6�@����WFk�K��I��lO�����ŀn���	���h����cI� �\�<��s� �{+ ���}� �7j�ݪ�t�w��`�2�	�N��X��"q���[X�*�����lO���:�\G
�*�Ɗ���D��PGz�]���*"un�t5l��'u8`)%���X�̬������tƛW���F��%��=�������sZ��F{6��F����M��m��{���ݗ�n���9�lO��W^J�ĩ��M�w�uwe�"I�����������9߰J��3�;�Oe`��0�Ȱ��VʈO��C��I7X��r, ���ɕ����]��vݱ�ـw�"�3���g�@�Θ���"���������������UEZ*�*��*����������������E��!B AP�B,�T"AP�U,�B��0T"�AP�0T EP�	 dQDXAP�AP�BBT �T B(�T "�P��B ,*�T  �P��B�T"	B T"�AP�)B)B*�B(�P��AP��B
 �P��T"�T"T AP�E�����AP�!P�)B !B�B(�B*T �T#AP�	 cB$B,EB"�T ���B"0T"��P���T �B ,��P��EB �T �B
T"#P��B
,EB(B"!P�AP��P�P��#P��P�P�T!P�	BE@@T$BAP�EB@T"0T"��T"
�P��@T"���B(U�@T"�T!B,BP�"@T" AP�,`*��UE_�QUE_�EU|*�*�UQW�*���誢������*��*���(����"����UE_��PVI��[�1@�sV` �����^���� �     P(    ����     � Х /��� } � �
   �� i@GZ  � ���  k����ڀR�  �4h[PrA�    =��@h�hQ��6�8:���ft�8����{����Gۧ�"}����; �_^��{�����` 7{�����-�>�>>�}÷�y��Ϯ��P��P>�OMz9t^�w�5�n��kͺ{h  ���A�+CZ�2��T6���l����-U��O}�lN@o�������ϡ�'UOs:)��
}8۾0=��� E�p�9��=������a����`���FO ��A�aѺ���� wP � �W{��-�}��@}g�Q��4����n�gJ
g`t�;4ow=4�73�:���.�g� ���F�h�ܦ�  �@iwp:P��`
�� �l�)����P飝����>�{���wpt4�u�N���� r��h5������aKۼ���y�f �ﺏO}�(9�7�����y������m����� {� !��,�;�P�M7�����/Kͼ�;�z^���q��p��> $�>�  x�]����|��w����`t݀gݵ�epm6�=2W�E5U�vg�d0  ���M�օ�(�n۸�7�����0�B�s�l��t9�N@0  ��SmJJ�1 �تT��j�  Lʤ��UT�@h2d0�?i����P   ���%* �"B�*T$F��G��'�����X�����������{���;�� ��5��� 
��PT�dW�� 
����*�O�}����D���l�&�Y�?�5
D����DJ1M���E�7!K�XO����}����R�t��s�����eI����NH�L(KH�H��������}^@���˚�a,Bp�HhX��N�'�!��ge�ݩe�	d���3�$�)%��J�����O��D�(�9��5���@��3I�v�Hj	L�"I��p�>��p���5�
B��?����(±�
@�E�0����S�	e12s�BK�%LM~��'8�c3[�.%��T%�e��k5��Z��y���ЂD8	��5�57����.m`\5R�L�%p��L�u�>�!f
���a����^�(H$F�gs���J�E����f�0��.�ӷD�dd"@�rw{##8�HK5rd��g�lČB�bJ��.h%�������� B�#t}�����'�\G��Ր�s�,�=�˩u:�K�~^����0!d]gߞs�ye�+�d�,���SI$c$��K�֥֘XR\�7ŭ�@�_�$�) ~~d(`I#.�y�nh���L9L�WF��Z$�D�h����bV\H�!,p���^w1��D�3���I,�D�E��0�L'��pp�GK
`�h�$�����9���ۀ�Zd�B���g��a��(JZ���0������2�@���:v���	A�h��4CIc�i&�'H|a@��@��, ŲH�$���˧l)�H:7�T T���$��et����L�l��!l���܃�ֶ!�5p���1�Z���t���T�J�P>ńx�D��IO�)�.2@�v���Ĕ�BX�0�!R��.��5	��B�X�aB�2X]5s�٨A�`�ZF���d$�ܒ&�ӽ�Z�JCP��Ck!D�w�@�#%�D�eR%����L�&�ȚV#�\`�3{�+��5�e��߾JG22Y�5s��	M˒�~�/��֊�Җ�!@��$�h�:����?^ɺ�eR�)���H�&$X�i�j�]oi��f� �@ŉ$x@��0Ѻ22;�gz��G1�����h�1�B���:v�>��r�X���K����?>��l`�%#�bHF�FI�Ѭ�vG������k�Ѯs��K��g�B���� ��8,j=]p?��|��ILʓ
��M�ۄ�io�.a��1%�4R�߫�n�����,��Y�%��Y�HB�?���z/>�����0�JR��c�JƘD��/Ü�Fl�kp�S���G�4�F���"HKB8�p!���̬�d a�k\�rY^s_�~%/ �!	anz��7���Y�h�Ȼ
Q�TX��!p�n%�"ЁV]�.jM��JB�! �XF��s&����f��2��	M[�Ü�%�����±�-"�,2tP�q����8l�aP#`Px@H$O��$���X��@���b��?J�6O�)$,���$$�q86��k��>��#���!L�T�csf�V��HD"D��B���B$!e��N`�g�>]~�t��v1�B�-��	HV%yu�o �R%��#L6�NB��s4:w	5�L!|}�W	98b|p�0�B�`t4���2�K�w���&���d!>���8�3L.kpև��H�e�	�6JƤ�/!ax3JX^B�`�-�����2���O���9��*�F�%��g/��/$��̙�jD�X������-�h¶!J�U��_ȏ2r�/GO��0!$k
iep��lgXq���������o��fO���a���!.1����%bA��6˛99�٘�5��
~�u�%�bL.(bC��,5�5�)�2%H������4%HHX%Rj��j�,�B���+(H�$er!.L	cL$�u���Ǖ��������1��,�D�����Q�:�G�0 �! ���R���$�F��  �
@��C4���?	7��Ѣ�Ϟӡ+kω_��e	��!$BH@���
B0%!2̈́(I��1!�h��d$f�KsR�E�A�$XsL�K��o���dB<��!�6'7�_�40ѳL���f�p�����F�\aM�}��m�r�4m��:��K�8;�*��,j�˾2��&o_]�T��ԅ9�!7����Q�H4ל�z~�G���S�\�Z>�7������O��}>�A�$e!n�%�%ĈQ0b0>����f��� 7F�&� �eѴ�
�
@���Y�N��>�+f�͜��U&�4�I�ӌ0�l>�)R�i�K��M?����k�� ~H�����o|�o[�8�Z����E�/�ｬ}[V���);;]��k�������V4�ʐ�� �K�[�]WYn��f�
�������~��Y�5�P��
c
0�5��&�a� @���F��4هѕ�XYyg��@l�decX�Y!-,�-�1�C���_4�>�$�Lnm�\4f�!3-55�LW����7����߷/	���F%��B��6{���%�g�<�~��CwrtϮ��YsS�1�J����Y����aHXg�.��@�N���}$�,,)���2Y	
����#!w��f�G�$���>�Z�'�P}|��.|g���3���1$\!L��B��!� �BF�K)���,-r�4���?���#c���R��$h���$'��0�������~�M�?2�%��T��D�/�(f��%q%0)�����5��\��2?~�r\�% Y!�[8KǄI���+��@�C[7��lptn%X���8o&�b����;�\R$���&�8�,RU�o`\0�����8C>��8P�
������� �F-nm$X�bӥO�0#@�OYn�!'	`�q��
�^��H��!��ҝ�� CL���a! D
8J�2�����fٚ޳0#H�D�ٲ24�W�Y��Y4Ͳ��Cy��B�61�B�R<'N0c�i���	�kC�8~m�$��y��a����߿	��@��@b�B"E`

X��K�6�0��T�tB�#A�4	�@�H�c�~	��q��m�°�y.�F�m�\6��~�|j B���V!���ąRRUđ��O���5�w+���h�1F.k�
�$�Hd���D$B�g#��4n�H�PIX\�I!�w���**J��H@�	�v۟/���X�����9y��\�4S��vq���M�����.���5�JJH�ۅ٣��>�9�e�B�,aL��,-��k��B'"E�4�Ĭi�al�f��5e֩	ė\�??c�n�ܱ>8_��R�q���0�4�C���-P!p����3H@!���4��J#he�SA�~%�h��!B�h!C0�ko'���kb0(c��"Rh���&�HÂAX�-��)��j�"Xd������ٛf����&�bDMs�$����Iy�X�F����Z�q�4�	II�O��a�B�`Jm��4�0���$		�F4$#Ю�ܠB5�&乨F.���5��P�0X�ɦk4�rXA�IY	d�4f�nO�h��,��B�Jf��g�c�����wӅ�r��٦����I�H�cHd��R�����м7��8h�ߎS\�d&����Z�WO��ܫ��-t����]|��N�ݗ@�3�[~�~��j�[��y��]}�>xL2�z1��_��_�+N?2렝�$(���ŉ4F�jK�t8F�+�#����(`��Iɤٰ�������!W�(l��h��011(B��j���M0�*Y �����7��3�c�޿O�?<�W4r��s��wwk��H���!!u�Y߇������a���>�XK]č�����7Li�e�r�xs9�]�[�9�;�|�,��%�#
BFD��+����\�l~]�p��0���n�l����2��\�����9�p�v��HK&bi��^�˷�?h��R��i�59�W��`Y�$&�^LHH�����~������5,����bS)��!u��|jN}�����Ņ���y���e6�4�@��0	 � H�$�����aM�$$	m��FR����ile� %�$��5���k_Li�s_}���@���4��5_��Mg�atp��P��H�HP����e��!.%�S��\�I,�i�,ļ�h��G�e ���^B|�y��UVڪ�UUUUUUUUUUUUJ�UUUUUUU[UUUUUUUUUUUUUUUUUJ��UUUUUUUU*�������������UUUUUAUTUUZ����ڪ�%��V�����pΈVkj��W���6�j���x��h��ت�@����U+��bւ��UX�\B`���b%7SU�v���j�������C�6��4UR��R��ST�[�T��U[J�O0UU`�j���0P;*�S��S�'b�UU^�U��[M��uF��mmJD��$�]kjݔ�+:%C��se�d���*�+���Ug�G�ت�O#b�`��V^Z�jv�aؐ+���c��b�Jk����ej�H�%UuRe�����έ7U�j�j�k��ۀ[A������s�-� �����c�� ���V��vUy���,��V�*��������P���+1@-��k �m��ʧ���j �VX �C`�s�e��k�eZt�qU*�]�Z��0LJ�U��U�KA]l ��C�5R�er�]UP$���V���VUZ�����v�Y���7r��Z���
�Bhp�u�2s��.�ݵ�j�� :�l��^�cj�2Q�Jǎx88S���)�HL�V�T�*�2ԫR��+�uv�uI�n*�h���~��QD򺳩j��
�`*BP8�:����ڪ�ʵUJ�*�Tjutҡ�%���m<*�UU]U*�ʪ���`$:�ڤ,ҫU�U:s4�f�m�SﶪU���(Q��GM���ykm��݉ݑ[v�Tb�Tf��SI���+xj�٤&�*���Vێ�E[]Ums�j[R��[���F6��
�j�`M�UPlT>v��e�G:-��*�m.֩�`�2��(��>�꺪��C���
�K��>²�l��+̪
�U�]��rа[	�\��Ş{L� ���MV�VʻU*�[  [U[*ښ�q����]�J�UN��ڎ�"ĔLJ�l��WUU��lQEʅe����V�%��KUU����}PC���P��Ky��������|��UUr�=O' ��xe�����^kj�Mk�U-WUT�zö�[
�UBE�7J�UU[.�uUYM�*�m@b����aT�@��t�\f%�v�1��)��71=�	ګv�3�PAt��I^@W������V���^v抪����v3P�,�d��T�Ut����vibɾO��ݝ���ޛ5X��9�RS�"��<6_/�ڵM��A7;�yB���{u�r98怌��R�j�f {[�R�[��p>�6k�5Un����ꪷm��,0�lV�U�����wZ����bZ�U�<��r�M%�6+���>���ڬ㦪�eP �:"K���`�����,d�F���5%,Yj�U�b���7�疸tN���]������[�%��S�К�j��8�t�R���Z��n������Y��T��)�UUuWTl���0f�ݰt�v�j����*e%G;l�V��6�UJ[uŞ�����UU, i��`@�UP*����#���v�6�*�h��y����v�4��TRJ�54�)����U[uʳeQ�Ht ���(��5��%�N��^�&t  �@*�V��NW$�����ݵR�J�S�@�-Q<ހ��s��m�V����hė^Q5������[6���7"��d4�zUwd#3&"���m{U@�3e�����(���8�U]c��m�<3�岶\�;=���tD����Z
������UUUT-UUWUJ�	����q�!=�_w�_T�9d���ڪ�����Z(�t_��*�9!U��kj��k�������;e$��U*�Έ
�@P��V���CV��NK������p�T�uWUU\�T�]P�'�kyR�l�l�T�U�e�� ��U]���Ҭ�k��VQ�� �.�������j@P�OIj��h6ET   0%Ų�ѽi.V����\PP�Uң�i��Pnˬ5ŵuN�'�_}��\�X�UYUʬU���팓j�eM��Z�@R�,UB�3�U�:8+�F���A�C5T�UR�HMUmUUUmUUQG[Hq�ή��@�ݸ��Y%mW�5�T�t�Uj�
Z�5*�UUWUU��J�R�Ur��Bj��!N
մҭUuuN�!V2�4VԵT�[�UU)-H�i���*�����SUUUUC�j���tmUUUU�Ì5m�u@UUUP�r�E�U���U[N�B�+[��*��j������v�^ؗ�U�u���Rٕ�uR� ѫ��
�R�
V���`�.�����V�ʪ���;ނ��j
��Vժ��^Mhk��V
;$e%ePt>u
�AK�U�9���M�m�F�V��W6��UT�m
�pM!6�UTjj����t���j��eZU�6�nҭUW@��R^��UPT�WT��KJ�Ҩqn��
����Pr�T��j8SMM�ZC�-����
����@N�HJ�J���UUUV�KU@�5@U ��U�eZ���1���jڬbڛnMUV�UX��l��`)mMU[J�����f�*�ȪCW�^��+r6결���h����J�$M�W�mYE^�趄.YZ��
ڤ'�eZ���  '����������
���J�UUWU@+;*��U++T��	핥k������LJd�%�m���UUUUV�*\@;��#�G!��x6M�i�]!p2(����E���FSP�X�9�Y��Wv7��Cy�t�b7;�mTl�	���v�,jܵ�$�F��媯+�[ ��u��:u�"�2�7U��rx�\k�UV*�b��!nX���sԃ��f�1qm1��mp�p��.��#n�k�U�SmT�V�ʇ򀮵l�j��
��4�T���Sb�^S"��J��UUUU(�j��"��UT�V�Y�j�����^Z��U[�W!0U*�NZZ��붡6�H��u[�[G^Ld1��(;k��pܹ��6uF��T۷��R�(Z��T�a檠 *�`���uQ�4΢��T�y��U�	Cm�Z��j����L��UPR��e�VV�-m5Ȳ5T*��XŌ&��K�UUUѶ��h��0o6e�n�,m�(�L��
����WL [m��`�U@UsUW+�RY5մ-[UT���UU�
� UA��au�ři��J�ꨀx�&>�o��C����$Q����u�WL�j+ZUUPpV����+dm��U.ͺڕYvj�O*�[*�*���̀�E���R�	[V���UWUU��D�hVUڞ]��+h
�����5YEV��@���UU=�ea�T����ת���m�Z��eAP��V����TT�ګj��:Z�U��AV����t` � :�U��8*S+��:OWc�H!�T�Ş%vj���;]�j�����d*�{fVڪ�ݥy����m �UUS˳UPb�WUP
�;r�@U[Z���T��h�"�Bb�P)V�V��x�*�R�0ҭ[UUU*�F�U����骁8j�����m�����m�UZ����v��������gst�c9]���,�ڢ�۩U`���N�ȏ4l
3���h����Ҩ5u@����K��PpYw�MZ����
�Q �S��U�����PmTRW!@�m�TUՖ����aV������UUUmUUUUU������j������
�j�I ��j�����#`j�j��U
�j��N ��
������
����yN+���(8�,1z�ꪪ�b�����	��ȁջuUUuT9�V��Z���P��X��-U�U��\K��Q��`�P(�sR��mMڡ˵Sjݩj�[��`p.]W8E��[UUS����R��UU*�k�B�W5UUT�PCm�b

�Pt\�Ͱ�jݪ��lUK�����U���	��XŵJ�*�:㊪�SmUL ��[mʀ�v��}��qU�6٠��U��
����ڪ�j�
��હ^v����������Z��*�H5Ul���+TpV�P�kt�̖Y���j������
�hjmUUTfj����UUU*�WUg� 1EUR	�ګ��T��j��'����`���T��4�;T�KC������j�h�f畢��iɖ��6�*�V��+JgF[t�J�T
�a��m�
����6*��P*���U`-���J��V
^U������UPUUO$�lUUT�Pl�5Ϊ����V6�%�j���ŋ��
�UUU[R���~��,�����9V���X���M�WR�-R��Y��їg�s��Z�3%
���b�q�Vj�	U��V���qU[a�v�SUPm�W �Vy�b��r�a^��Z�e�:����.CUc6`9"�D4X�ڨ;�V+
(���UUUm������!�oTʵT��*�@Vʪ�j�����R�TƝUUW*�UU]K�L8j���
�*���/&nݝ�४��PZ��j�������
P *���-UR���ہ�<U����nKE���������UUZ��������k`*U��U�����SUUQ�e�j���ꭕj�j�th��U�^��(j����I@�!$�UUm�kj��
���9ڥZ�V[U�	��ڱPT*�%��n!����\�uU��UJ�۾�^_�[j��V�c6ኪ�*��������Z��8��I��������U�`]��u�L��N�O����>E���?�T�
o�&���(�����B�!�J�T@�@،4��^N�������`iZ.��j<G��Ё�D&�������8)��1H�H��4���P�'Ab�O��	Ph���HpD8�~E��Yt��4*mQM���U_����"<�Ȃ|��T �P\:�:���c��U"�808���@��*JWH��ʸu ~A���!�� ���`@�~?=  � M��6���c	R��x+�G�C�@6 	�t�Q~L�!�Sh� iF� �q��_������@6Q?$)�tUM%D��X�A�p��P�D;������pD�TS��M$b#?���X2!A��S_�A8!���/SiD�!��G�A�A�@1�@(B+)��$$(�"� |��P��P�BF�n"|$ $Qb��(�����?"���s?(�80A$dVE���BE(�� �T� S�"�A#�E>
����5T4�/ �ç�!b�𑀧�P@\Q���"Pj'����U�%J�Q��pIН$���t�����m�⪭��UUJ��U[��/-Uir[�g��(lF��x����i�.vq�9�Sk�v����6z[�s#�.%R��"pر����I"eq \d�c��m�<M#�P	���X��8S	�Y�`�t�F[bڌX�;jbЛX�0�kO`��a�I5.�;p�5�(����d�8��F��g�jܩ�"gn��S�6x3]c:x��F�7D;w'#��"�-��s�;�����) ӷi]�Br8� ���w')�d:x�-�8�u�)�)6��rt/!Y�����&e6���ޮ��ta�deyvP�>�Gii�C�Qr��seD33+�*��S��vW@��; n�Z��%ؙa&�IfJ�KoT*��U��둋�x�]l�iL�mL�*��s�\�����Ru��Zqb��Ѵ�m����l�Q�^��c#M�v�� �u�2�9C�˴��dN����ەٰ�qjCQUcB�6X�-%p�[tm�*y`����^1�����
� kD����S=I�MiU����PmDc*�#@��:M�VSZ^<V]�6h�����T�&5F�9k��
��x�#ma���X4ҴP�L@l� tN��4J�\�б��ڨ:vE^����V����=ab��jV��h�9��mk��FH@��i���BE�K��eX�,��%B�m�r�n1cqm��������k�T؍�vfr���t=�aFUM���61tm�m�hjT�!H6h%��9�N�Uڞ�C�-�!�1k�l��y�qmcc(�Un���n{��w�'^��SS�W:^}��WM\B�Ԕ�xln�(���Q�p�̮���S		Нlq�e;�᪞^�h頂ƺR���jgC�(����Ί�[pvģY"��J]Vh�ZFP��`Qb��,r�ٲ�#ClXɫ�����\v�*B���[m϶Ud�NFe���[�Hͭ����d�4�j�WS��۫'O��'Ft��{;��]�bQ< ? ����.: A�!�U�����u����(��F*�F'��k��MHe�D��H�`Gk��\Ѭ"�)��i-��E���uA��qm��v�M۷!�5���ǡ-��Mv.ws��н�O�ѳ��l*�9��I�Nn�k��3�3�֤��\�a��)��%ٗaX	����l�c�:�'��ƍ�:�k
�],v
:̊`6h�庹�Hj1h�o�Ǧ� *�M�-�T]Bٚ��'�%Q����%�3)ai�.>y��v� w`�����&Lc�'a�e7G���ɺ�}�z0>��_�U���~0 �#�ul.�[|Wl�;*�,�r�T�����|�`�� ݫ�v�;m]���Wm`RK�7�� ݎe^ŀҶ��.��j�������p�;*�,�IxԻEm�*�Ҵ;I6`�� �ذ�%���/vߧROܟ}<��&�)�e���$�������ʑ�7�����)���-ص�91�S�Jƨ��π�U�,�Ix�8`�� ޕ|�Ւ�]�j���ַ$�{���%Gj&)D��BUs���c��;5� ;+c�;.�e�bt�I���ۼ{0�ᇫ�I�x�{׀j��v���tӥl�m��p�����%�5� �7R%][�V��0elxT����n��\�W9���<�'F8�\�]���h��5��.���ȡ�ݲu�g%c�T�"�j������^�\0��+c��[J�Mڵm��V� ٮ�p����RK�r��H�5Z��`�5C�]jnI��^��O�}�nua�,j@"KX#�`�""�y����nI��]��ޖ�(��:��j��l����RK�6k� n���斬�]�;Uv�xT�����< �[���-��i^V�5��0ᘹ^%=�Ne|��@nt��j�J�� 1�"��ؚj�ݻ�6k� n��elxT��R�.�Uv��t��vـ�<�G����5{޼Mp�"ԉWWN��[tҷx��<�/W���uI��;*�X�j�ݫ�m�-�x��|�e�{�ں��x�)W bX�q]	�&[����|Vҵ�nիlV��x��|�e�������U\�Hx��v	t��5�� <�fݻ��0kc4���gzg��JL���	�����e������׀j�c�>[��|�ޏ�+l�y1*uiX��w�j�c�>[��	5� �n��;�/��d*��ګ-���ݗ�I����Qlx��mU�bt�I���ۼr�Kޙ� $�x��<�$�T��]���+b�l�ݏ �%�O?����x�ᄘ?�tHČC���@>i�cT] 4X��	$�4&���X�+�
8H�DH��e�5�Mӻc��]08j�FZ,�stOf��x�<J;d.���+l�Y.�؋�hg�k-�<����X��z6���q&
��a
�н@l���m�cm�v�����["t��1Q�%vpB�E!efe�V+�/�;���f@���(`�PN���?��}���]�iH�bŝdy�u��Ѳ����.��]A��2��[3�����9$d�@�z�5�&������\�z�4ҙ��a��%�+ֹ���laCL�Sf���n����������	5� 7v<���T�v�n�ڶ�����)#ޏ� I<�Qlx�V�R��ڵm�hV� �\0{�������#��b�,���;��0=U\Jl��"�x���	5� �횔LJ�ZV5Ci��j�c��ǀI����W9\�wh	��Wj�9%��a��U��	HFCD��󆆶�4��2R��LV�"hPE�m�������ݏ�U\��E��<����<�t2�MSN��7u�7����q���P(�HT:�DC�/��_Y��e`-ۏ >�{��@�^Uwv4��vـI=��j���#�7u� !���N�:��|��`{��*�����}�<w\0ݙXe\#m]�M�j� �H�UT�<|��X�ˏ ����v&�"�<�S���SX��*P��9N9v�Xw�8&&�ge#ua��\��ܽ�<}:�y2�]� }$xȕ�bD���pwI6`�2�ܪ���������p�6�f��V��:�V� ��q��G�)�U]�s���6�\0ݙX{E_!j�"�ӵĝ��I���̬Weǀ}.��]Gi��M5Mݷ�n���+ ��q��G�}�{�2�:)�\eQY�t�n�l=e�=<a��ݰz0��=�l���H�li��J� �ٕ�j���#�7u� !���N�:���n�`�.<�r���x���7veg��I���I�5wcm������x�`ݙX�ˏ &�)(�n�v�ĭ�w\0�̬Weǁ*�����!�HT7s��$�gO���&�^�&���+ �K�_�����7u��o�<�9TD��%�J�*YyPa�9�e֕�K�ɩ]����V��E��ZV�Z�_�������wve`�|�� �WN�v� }�<�\�H�?��Weǀ}���N���M5Mݷ�n��ٕ�j����]�]�EV��N��Wm�wfV�����G�n� B�D�RuuwV����`�.< �dx�`ݙX�\��Q\�UU�v��T<[�jp�6�љ`Xݲ���f��m����k���od�뮂��;lq�`c���^Yl�&j��*�n���;,s�;�94�bՕͲ�Ysm%H�H�qU)z���BMy6%p��4�ע���Ìd�b��ݹ瀹��]]�gO�!l�$2������ĳZ�*k.��Ь�]/F��`;�=�d0�6�3W35����\����Esw�1�b�#X�i���������`��g���[)2�8�uW2�T\Eh�U���p�7u� ����5v\x4�IbNۻv�V��`��wve`�.<�{d�v����q��ـwve`�.<��`]�R��S�J+V� ��q�lp�7u� ����;�*�VA���$����I3��l���5vo^�x{g�{�6� kf�)�u��ڳ���t#;��#v��x��STv:^��ᔚj�&�w\0�̬We�ꮧ]Os��ݷ��t��6�!���?}�vo��(���dp0���q�9�W�Ϲ������Mp�;����&���un��b�X������wfV�Q��ؓ��ݦ���}#���v8`��x:P��'mݻm�V��w\0��j���� �9�UT�R��5�ݶ�M�ZWի3HU���=���Ҋn5�^$m8nt�5X�@ӻBt�V�'���j���� ���횔LJ���`�����G��UU$o��`#�nɕ��W7h��VxE��k�&����wu����Q9L�kEv�A�pǊ��� �M_�@�fؤ�'{@�.�xJ���Г>@�~��C5����X��0W1�d6�RĤtf���w���p�pӁ"' ���
B"J��bR�f��1�ā,nu��--��t���a�����;"��8u�`���ńjB w@�������@�!�D6�E���,��K�MsZ`FU����6?������^��[�%�1��4pU����hM�֐�4 --SZ5�In��J�u�������z=A? �5 )ĀD����+����ClU�#��~�V�ձ�۩wQӻt2�MU�� ���&V��G��r���� �g�z���i��J� ݓ+ ��#�;#���ܮW)x5K�	%���uR������v-�	wJ0�EbYX��*��5��F�,�31Q6g�=Z��vG����I=��z�qz���N�t�M+o �G���̬WT�=U\�B��X���ݶիV�d~0ݙX����b�����MU���)=�$��_{[�~�uٹ4pJā`� �D�0��X�?�?�@!��PP�W�o���rO�ɝ��R�M5B��X��+��r����{��wu� ��շkR­����'\�TU����'f�."���V��[F�؊�}���x��5�ז�~���}���&V��G�wn����t2�MU�ـwu� �ɕ�j����j��]Ժ�v�uvһl�;�e`��ݎ�� �wbi�un��e۬Wv��;�� ���wd��%)�ciݧv:m��fݎ�wfx���V���gj�Er��!$!�|/w�h����Y�%�`�A��p�lѱ��K��N��k���+G*�z�lT4B���J�bb�q�(gRq�rsm\���b�X�y�\�ag���f��1l������Rmdm&1۷e��7X��J��X<�^�&bԁvv��{#�:�%'(�T�&6n���[15Ph��ӹCH;R���Ķ���(�+�K�b]m$�E6���۲�/e�nfY�n��$q��˺^�nv]B�qx	�w����j֍���Zc��m�h�d���wd��7��0��vF*Wi"XҦ��f�&V���wc��u� ކ�Q1*O��T]ݺ�7u8`��}��wd��;�*�VA���ZV��8`v8`�e`��0�KLt�t2�e$�0�0ܩ=��$���;�� ;��I��ry|ܔ#��ûN��wr,��g�y�gl@��Z��f.��Y�1ͻ)�>�｝wS��=Uʪ����l�����칥eQH���<��}��>I�rq�0&��| ��3�צ�}�znI��~�<��N�:�?���b��n=��0�0��Uq-��V$O� oJ%˱1��m�h�f;��Xf��8`��Wuh%��*h-� ݓ+ �bp�;#�����N}�~�>U�Sa��8�4	[@��FLv�h�U��-���	�tGm�ص�^)����5E�ۯ���~0��ou� ݓ+ �����dj�5�jـvG{��X{��c�n��-��M��l�7��nɕ��r�9C"�@X�DB	��D�|�M�	�D33��rnI�����:�Z]�EV��;hVـn���;؜0����`7Uڍ��t�)�� �bp�=U]�{��c�n�ݛ�y_���-ԅ���f[�Y0*K��t8nŊ���.2��%�6qظ��u�ʩZ�Zwc��-6|W���7��n���>�N�P��&7v�]�X�\3�$l����S�wnE��Uq#}�*Uv��v�4ـl����ӆ��R[/�X��`�k����5E�۬s�]���l�y`ݙ[���j�"A`�Q�"tx�#�����=��e��r�2C6� {��x�S��y7��w�9�m�ޛܛ���/�Os�%�u�5q��o1�{�lι���K��\Ю�%�&̴n�Z1Όnel�9?~ �ϻ���]�>��I.�Y��$��E��%ۺ���&9�%6f� ��y��Ϻ����I%�����%�fU�I%��+v8b�u��� ?s���� �ל<�����ϻ���s�'� Y��c��òUf�m� �ל<���w7`�}�� �u�]o~�y彀9e|����Pwm}�Ijٕx�Kܮl��w�%��f+m���o9m�Qt�EҔ�A���aV"`%�H*���v���uBųD��yEjĤ褑�K��r�W����\�1z�f�W���.��q�m��܇`)P�{c���ug/2qi]��u$�+���h�)�֍דcS�YuCY�9I�89��+�9�y��6�`-F�۷d�@���0tX����an���^Ý���6a��j]����2��Z�V��î1O>h�Iչ��nJ�jK�-f����t�I)�!\�i��y]�����a�Dtg���}��G��ҽ-�t8�v�<;J�`���$��~����%�3I}�E��%�fU�I.�7)Dĩ>+C�n��$�&`g�s������[�����������s��N����ǧ]~�����m� ���x��;���I6��＞x�������w9��`��煿��*�����7m������[o�����|�$��w�Ǟ {��ƿ�%6f� ��9�����{���� ���xճ*�$��r����ڷwf�6(,z�Al0�&�V��
��l1�k�+��f�7nva���;3����v��޼���y޿I<�y��O< '7'�4�*�췰��8y�I��՟�����e�i� D��H�"5Q
!�_/����������{�9�m��x��:��YC�.�ud��Kn{,Ē]ݟW�/ܯ�m����I%��x��CkosJ�WZ�^��m�9����~N�=y�� �o^}潀�o;�΁�3c3� ޼N��ʪ����庒R��,ĒSd���$� �܎}[���v�dp���k��@��#E��ᩭف(��`�os,�˔�&_$��~������1$��>�s����?'`��}�+���W'� ~ϻ���Q�kV�{���9m�������ל<��ԛc���]���]vJl�ݶ�w���[m�����q_�#"����M��	3������-�����ݶ����c�e��.�s<�������q��� ��� s�s��=��5J����&�ĒS\��Iwf3IM����^'`5���u]F,��/'	�	�ru�v%ݻLs��.�j�r�E4�E� �hl��ud����������]�ĒS\��KjF*WevT�ڦK��y�'� �x���� ~��e� ����ÃB:͂7l�< ?z�; 9��x6����� }Ͼ�y�=�n�u��[e; &��$�u�F$��O��W]��9��
`�p���+$
��"@`E!!	�$ !'�D(#�$�14��U�ֿwWv�~�|�0l�9<���w�`�O��Ilq�I%�Ⱦ�$�t{��Ka+	�`��3� z���<>��m���rt�Qi���g}y�,(�� �����$�8�$���_���u���e� ^66�G-nZ�3� x�7���{�{ל���{z����{��L���j���T� ���< =�;oa��N������>~N������v�戗 ;�ͷ�ߺwr����7m�����9�m�w]�ݷ�W�ֿ����y����i���*R�;-� �9�'9m�ʡ�����_������y�m�w��ݶݝI�a1�)6���02*D���턁*f͊m ���1	�R�&<˹�h7����(�L�5l�`@�78o�������M��%4�a�A#�	JR4���a# q>���K�S�5�H���C���#)�|f��I�� �AtC��	0��M�B ���c�"@8g8r�h���i��o���D� �daHl�j�
.��p�8Aa�a�����&��|+ �(@��(�F�	�h� Jf��.`B�5"�sD��:p5�������! �Z��p�h!L	p �i0	�Ą%ܛ b�"C�ZcE`0�B�P�xp��A
���o�|�w6ǂJJ��� �������p h"��#x�rKd�g<��ު��)UU@���mX�d *��x�<D:�ӂ���m��^ּz���l��1vǥ��gl�jޮ��l��λN�$Y�"�mJ�v��8\�m�1V�x�Ә�wl�3�"���[������m�Qg�l��������f*�9�M;\���=�U���O$�ag��GGY����i�p��f��@cl� F��.eql�.ح1e�:{[]A�&I���O3�m�Cc��t����툰ӵa!ݺT�=n3Q�Z���)^Z��[�]�=���d�B���4�]��$���0ȅK�˚�춸J�{�Gn^3Eg�d�\se]"��|�Q9���#��$�P⣚�JU����)RW:4$�=�;�d��ہ�-���j�+�m���{.��'m��h�9��s[Z!��ц� 'f0/m��Q��fۍ>Rn�7Y7#�ayvNSkq��e	ó`AE �EP)v����%���n�.L�±����H�dlT�	B%����r�+�����0Z��ۉ���t!��AT����<�K�WGd�rf
�; �ux)u��mf�X�
b���Vح���\��L��	ٸw���e��Z��X�fo#aP�����Z�T���}��~�b<>�S�q�l'<g��F�BlA�q�K����Z�/��mn�cNQz�-����^7A�xp���f$E�PL2Ѻ�J6��F�8j��.�2VX&�����x�&�fsׅ��0�;%t'���`C��q�L�v�N7\o9��!��kB���	�z�B��Ԯ��,�]F��1�[�=oE]�.�T�4A�QF8B��0*��k� W���6����9	T���|�F-�03��m��C����܎��v�v�L�xYF;AK*�V"�л��di���^3,E�{A�a�i��0%�d�2�+g={�!��Cl+���r �c�KZ�M��eǮm$�3�㷒���UT�.L��Iӧp5��$0E?qTj�]��H����6�-6��~EC����sz�Ϧ��Ւ�X�q��7&�Y3v�v�ص�|��ң׍�iF"z�u[=���1�7c{�GMr�D��t�7)�^q�pv]�ۓ�s9XN4Wm ���魍��ٖ���1���Vn��I�a���Sf��&�R�]�9n¸�^0��k
Vu��g�����^ +�lF)�G�u����@�ͥ9�aU����r���g��\�h�L�u�"�U�v�.\Ն���E��Xf9�B��>�����f������`ܓ��@DP�&�n�<F�g�v�~��kIlr/�I%�c1$��>��I.�Y�uה]�[e; =��y�u$��i{��f$���߾��I%�Ƴ�ʫ�K��w>jу`����>��� l������ʯ�ʪm�~�Ē^��~_|�[����^E(;[���Ӥ�������?'`�y�� �u�]mϾ�/�l�Z��3� x�; �TC�߽~���{z����{��Ӹ{��1�b�5�@�R�hJ1�h&P�*[e�I���[�2�(��;�xO3�s\�+`�k�]��|�Kd�bI.�ϫ�W�u�]O}@>�?�� >���	�7+��k59�m�w���6�HP�$��C�!������r�o��j��o>��9� fa���%��޲�+����yϼ�x	-�5�{����{<}�I)�c1$����V���fy�I6����������$�Lf$�W��7=��_|�S�_����r'N2��{��|������I-��W�$����$%�UEjZ]t�r(c�l�F��v�#&9z3�Cs�w7j|�����ٿ��;�3*J��S���<��+ $��W9_�\턞���{��b�牴Tٴ�zϾ����s������=��ly������v{�j��;lcm;-�u��{��;ݙXmo*�¢��M�{^�$����rN�'�eR�F#.S�t��'N�}�����{��>�X^�s���9��&����L�݊�n�{���ʮW���|^������7e'*�N���R̵��u; ^�[���hF!�^�`\�k*PaR-��UY�X��`e�4!1;o�;��XSe����U|�����Q^h�ĩ>]�LWn����r�6y��zy��2��7��**v�5n��p�	6<<��{+ ������[���M�f�W)/zy��{+ ��������1��J�h�*0@�>S��k����7$��i�i�wVڻim��e`����y��	6< �um��v۫��v��Bs��׋p��k;=i0�S�^�WgAHkqͣ(�n˷i�&���xv8`�ݓ+ ��U�i�+�|�t&� ���ʤ�ޞx�{+ �l� ޔ��Hi�[n�;�`�����"�/ ��� ٵZ,��B���fV�x{0M� �@��I>]�Nһu�E6^�V��ē�ﵹ'������M�iD	��S�9ʹ��(��)-d�i���'tAu�jv�⊺2��^�\�[��g�v1��6��ݞwl�V�C��#B��!��n�ݖ8�0Kn��Qø4��(�1��8�����8�ؑyȽf��ݶn9�e����	Q�it��م�Ù)��{r򤅎�&�r��ƻ���e���eӃ�ϱ��9���Cc{m�J�`�d!�[���I�t���q"|�5���Hi��I�ɵQ�X!69�v.�ew\������ts�m5�ջ�{��lx{&Wꯐyzz���ŵCbt�I��l�	6<�9č�{+ ����Kذۭ����wVڻim�ݙXSe��Iw�<�ޞxV���r��v��-]���W��׀w�<�M�ܮR�=�`��W�n�J�]�w�}/b�?s��W��9W���>����XSe�[qJ��P�,�m �k�!V�m)�.L!�b��|p�j�������Ľ��ɕ�*m|�O<{�+ �l�r��W>A�\��=�^�b.�V�ݷ�ovec
HD1P�*rz�~�}~��	6<���U~�W*�vo���T���S���`��~��{�9�U${�� �=��vQ�vYQS�m5�ջ��*��]�X�O<{�+�~��?߿�@����ˠ�eIT�sz&ǀove`M��}/b�;��ݼAH\m�(��� ��k�>⭂5M9���=�j��ǻ��~���/4,"��=��E6^�����9_ =��j��]�2ӫ���Z�u�E6^yU�~�w�rI�w�ܓ��wf� ��{��7cE�
�t&� �y`���,T]���6��u�}��j�׀�2Ճ�[l�Bma<���}��;�}�rN���nO��E��{��?T��"��cV]�j��7�2�W9U�z�޿��y`ݏ �ʮ�������JU-6� v���i����tl�F-x3�9i�Bz��[kdh�[���n��}��>��`ݏ�s��W�&�e`��i++ʮݴp�n���Y�qB�=��[�w��f䝿�����"9�������:L��Bv� ~��<{�+W9ļ�޼���vI���M+�h�i���*��� ��z���X�� _�*; _7�{��$��tEڵ�N�һbWn��%�Kذnǀove`�ʪڃSʄ>$]Z�JlM��R]�.��*`˰���A��%��i�fۨ���cwb��M��������fǀovez��o�x�G��Ut����	�y"l�V���{����I��6?�����;t���\��߲��%������w��ߖ ~��<����6�X�ٝ��G�߾��z� M���̬�7�
�EWn�8[�x��, ���n̬.�x�w��8�}����h4j�5ءh�`bݭ��%y�;6��imB��9ŕj�Z�8L烊��:���z. ��h.Ϋ;�����q�ͬ�D���5�#]j��ڿ/��A6�I$t�eX��hzغ���<[���v����+�9����*�q����C�Q}Pͷ5�8��c@�.bc��1�8I�qm����3��VF�ƭ�0���u��htn4�Ν�%������Қ$���] હ��:O,�y�lt���+����:L��Bv�@&���>ݙX]����Xd�LLt�m��i��>�2��H��z�	�<�nǀuCij�ҺWl۬.�x��,=I�� 鱗�	R�U�n��
v�n�=Jk�X����+���s�*�9�����~��Ut۫��t&����w��W�yo�x��,m�Gv5vM�x1���nxT5j��5��^��=�>�|X���Ph5A��,�%�qp�	�����e`vK�7��~�r�A�'� �Q~̻fV�8�3�{~������$@��	$��D)�А�*#bCO1�+M���00�/���%Q)� ��_۟���`��� �veg�UUI��hW�V��p�n�˞X[����s��U\����e`�����:�m��:L��Bv���ٕ�E�/�\�r�c�X��2��2��E�T���>ݙX���UW�}��˞X[���{S��6�s�@�'G:�{]�d׀�yr�`�L<Rk1JFc�:����5���2\l	Du�[�^��ŀE�/�W9��\�s����?���]����J�;c�xeȰ�e��� ��^~�s���UʻD����n��X&��{߯ ݎ�>��� \x`��^��4�P����:�ޛ�Aq��9��Qp�42�M(h̀D��x��t�N�, �m���$?'!�������^�A�WI�!�Јf�Nմ#!��7� �h�L��ԡ��A�R��mX~��g��N�<~+��M��tZѵ��ȡ���x�	@���N���A�v#�T��*��P`�S�����|�R"����mD](���~Pv�@l�\��[�� ���J�D��+�Lj�m	���9�'��`S޼��X[%�($i-һlC
BM��x�����$���rO��vnI����	�r89+J��84�BdqXlTr�3�==%m���.E��~�uǄ��Y(���߿^�l�_��v��?~x��_�ۡ�t�I���w�E�^6L� �#��y#d�S.�ӵm�]�IۼO{+ 'dx~�W?U�=���?}���}=���q�1���fwoӠ�}�=�E�/j����R}X��r��B�aN�o ;�<ܯ\�����e`� �ʪ��=w�42���x�=��Ju��6�1�����d�'`�E���G��w�2ٲ�Z��������X�c�s��y��#ܺ�t��ZM�[��&V l���#�5M���$6����]�i0�$�`����UU%�� ��e`��s����%d.W�N�������ߟ ���׀wd���ٮn�ݺL��M+o �6^���?s�����@=���nI9�{��>f��q�E P�?�!&� �cUB�� :SZLt{}�YK�]&�P@i�st�Tb�ɦ5f�9HL��g`ݪ�m��Vzo98�����d� t͖Z���;{^S�l�n2데��ȯ�g��[�&�8u-F$(�[Mĥ�1qM9.�CQ2�=v��3vSr`ݤ�^�S��vBD�Pb�g�2έ�ulA�8q��Ba�J�SY�]��P�4J]4k<=\ڵ�E�O+�n٩p�B���f�����"/�Gj��vϜ1^h��xib,�ˊ��(��n<=����0�4;�Qi��wg����4��T������V l�������5i����V��N�ݺ��z�\H;=�E���;�2���$z�tK�.������y���������\���� ��~x��D��˺m���Se�ݙX�c��*��v{� ����+�Lj�m
��ݙX���qOO?�;=�j�/ �%�n�ۥ�	[�h�kif%@�ϸ��k���C������)��r˩DT�1�	J�| ��x���Se���W9���X���u��&�1U��=��I$�}T��P�JAVI�@\D?� u�~���f�{��7$�w��p7��4�ۤ�V�m����;�2��W+��$OO< ���6:�*�Nշav�'n�;^�9U\��懲OO< �v�J�s��[se��DUڿX�E�N�ݺ�� }�<T�xwgg@'�o�ޗ^5�a�U�b��.-cf�U-��[e�H4�Ҍқ,�(���:Y�/��]�&�N�m��;=�j�/ ����9UU�zy��z�+b�hi;o �6^�ٕ�6< �dy�W9I�#ܺ�t��ZM�[�d�V o~�6�D(�(1�BW*�W9�Uz�T��g��'� 'P�F�v����� }�<T�x��-��V��q�U��ӱ�X�x���Ur_���6Oe`͏ >4�1�[��سt�j��ڸ6y��#;�D7;.�7j_cv\iWD6�]E`�n�m����;�2�f���U��U]�7߿<��?�[�]���N��ݙY�s��OO< ����l�V���W,v"էv� 6lx����*�.����?��W�v'n�t�oܪ�K��xe�� ��_QUU¸.� �T��+e�6�wv� �nE�{�U[�> �<�]��	����k���aD�n�b�an4�]����GJ/ӸB-:�[���!_8�cZ�7wvπ�G� ;���_�vy��	�^U��v��f wv<�+�������?~�}��0�p�����r�����q�U�|��&��?~��f�`wc�6l�m:hWJ�M�j��z�\����o�� ��x��*�������~u�ҫt˷l�hk �+ ���W)l�%�� �nE�mUWtP���P��
I�N��I����R
�j�)@�0��[=��VGR	� �5������K��p��*:�cm4�uI�HQH���g���7i<dٱf���Y�L+֭#v�^��S�h�g��c�v.�D���nv6�ۮ-�C�y
U��;X0����`i�n��h�1�������!���֋s�QŶ�k��\�ژ����ِ��K@"�m�&s����G�Ӥ�:N�I����o.2кX��Ҝbt��c�v݁��eZ�p�|=[&��X���ݞ���yc�ZVҵn� ��ߞ�r,�d�X�ѵqںN��L�M��n܋?�U��ʻ7ߟ� ��~���Ǟ�$JF�Ը�i�t�+wv���� �+ ;��r,k��V�����f��}�}X�y��"��U�r��U^��ߌ �B���b�lC
BM� wv<v�X�0	�et��=���L2���\۱Sf�ܫB�ha
�$������CMe�㾻>��u�v:�o�=/�X�0	�e~�Us���{ߞ�߿e[N�Ҳ�gm`���ބ�RUS�j���f����r,�$zu�J�LWN؛l�7��V wv<?s�\�R_���?Zj*N�i[Jպ��Il�x��,��%���%�*��]&�n��M��n܋ �]�� o��|�נ|�oo��y�����2�8x���lk�-��I�R�ֻ��@f�0o������t�+v����� ;$x�����mwP�V����wwv� �窒�� ������m/*�b�lC
V����� ݎ~�.�S���X&��5�}���'��u�Q�v(��Ӷ�X�x�?r����`����<�J\�������M
�U����0�p�?r���?�$�x���t�o=vJڳVb��w36�\3Ҩ��ػ��y���ô/-��]��R��=����Ӷ&��> ����$p�>�� �E]ҵ):V����x����~������o���I0ۣj�.�t��eӶ�$p�>��߹˿߿?� {����씸��.�WN��qw����� 7v<����bo�n�30�!/QN �G�\���H�8t�J˷i+k �8`����ʮU���Ϡ~���0	/b�>���;�0�h��J��.��u��:���l �D3y���5��mc�갵�m�Jـlx�� ��/Ur��A�y��7�N;�>Zv�i6�	#�~�~���.�߯ߖ�ߟ� $���'��i�%t���HM��s� �0�UU�${�� ���n�Դ�t�t퉺wm`~�9���x�zy�#��r������/����i��	6<�%�Xv�, �r.7T���	R��IE��G*�7q�@(��(P��C�f f���@Sx��t� �
�`�!���������"T �@V����Q$ 
��!G�
�����q@����tI�HBU���"kD@#��"%���K#�S� �Z)�å��z�~⪭�)���UU��t�*�/f�<aA�jH0���"��([Ex�5�V�e�I�7U�n��^ƌ6�nx cI�NԼ�W)�6SUU$�8���T�ݛ�eu9�iY��b��r�1���[��z��=����a�PI99M�Z���n�=��z�6^�8An#8�\�=�(��J{�8Ӎ��S�g!8n��d�wNe�awl�J<���j�iuۻ+.�nƱ^�ɰ��ݓ�T��e�N{-�T�2�=k��`&�O�d�ì筧qnr �n��$��XͶ�k��ع4Gh�*
�rc��Eh�n�v7mm91u�s.L4��E^�E	��������m��Ƿr��&xa��6a�Y`8vAc{J��S��ڗ����A����4��k\{Bk�k�����)q�Amn�q��#(o PЗr5��*��khn� b�Ƞ��T��Nl*�*�����dQ�n��]��v��4'P�;#�Tݵ��m��0�c�xe��蹆����۳.ه�� �`JꭷGl\sR�۩	4srN��*�G�	���Mf�iJ١q@��
4*�ᶙ����Aֆ*:c���(q  C��[RW[��dㆌ+rO6A�a=fI�Z�� l8n��'�
_5M�*b�+��mE�OO���l��Ƴ��#�6�Ìk2�����T[I�`��h;"X11]�ʙb�l-[ͪh 9K`H�i�ؙ���cm���;�6eV ƻ(�n�2J [.�l+�V�"Y��#����n�t�Z쏂l��q�,ݪ��ׅm���� +��.�:ŕ8�gp�u^hҐ�����ƞD�OT��ؒ�U�"�=�J�+�C�n0�P���O��ŝA.��q�A%�25���-�݊)���z'�:x�8�����X	�h�4�3b�ۃ3P�v▔�d���]kXD,1c�e�Ժ����xu�5nX���&7�I9ȁ�)O�+�(8+��G��N��|"t�7���D: ~M�,�Pt
�� ^���f)��Ls93v�g.z{vi��g�g� wbw685"�WT�L��<;:֧X�le�d[B��1��^"�ڻ"�N��E��L#�J�4A'k�/]&��wY6"�6R��HV���*Y�]f�s���-���`]7J�z�Fp�`qS�(��8�ܣC��v��x�Zg�+��8v�8�;N�A�j��W^�)�*t[z2�d߮�q��㱯qB؅��T�b]��J�0F.ml�cv�nM���T#�rmٴ\������%�Xv�/Us��<��o�K��2n���$�� ��ŀE6^�܋?W��]��y%��˦���v���	���E6^�܋ ��, Ӵ��6'm���[kܪKޞxe�� ��,W)ls� �Q8�^wEZv�i6���X��`�ذO=z�p���V�2`��ѪK�U�9.��[�|���z)Ik�:�i��h��p��U�������׀wob�	6?ܮ|����H]O+�X���7Iۼ�v�_�!��� �'��krO��z�M��E����r��i��"�/ �nE����R^^��e�,K�j�J�N��L�v���\]��X��� ��Ł����%�O<����R��]ձ[������=��*�c�Y���!,K������bX�'��޻ND���5����z�q�m���ɦ+CnSK̐����a�X`���n�祳-��i5��s5�\�m9ı,O����9ı,K�w��r%�bX���z�?� ��ı?���ٴ�Kı/�K�a��r��������NJrS����ki�"�ș������ND�,K�?���ND�,K�뾻NE ,K���뼗/�2�4Xe�ֶ��bX�'��޻ND�,K��}v��c60�A'��7Q3��ӑ,KĿ�ﵴ�Kı=���5��[�2]j3Y���K�F����]�"X�%��u�]�"X�%�}��[ND�,K�u�]�"X�%����fdѩ�5��Z5����Kı>�w��KıP��}��"X�%�����ӑ,K����]�"X�%���C^�ݙ�v쎐l��Z2���2j�`tf%�5��ن�u��\���s�vs�I�A��x�Kı/��kiȖ%�b~���Kı=�w�j��bX�'���<���צ�5�﬿aM=�cH��9ı,O�׽v��%�b{��ӑ,K���ߦӑ,Kľ�}��""�L�b}�����ɫ��f��ff�ӑ,K���׿�ӑ,K���ߦӑ,��Dȗ�����r%�bX�{_��iȖ%�bx���s0�a�t�zk�_�K!z}�ߟ��9ı,K����m9ı,O�׽v��bX�?���0���4�_��� t"�Q�O��{��9ı�俽�����r��PT�'Ò��K������bX�'��޻ND�,K��}v��bX�'���6��bY�^���O��~��J�y�80��#�g 7!�B�-f�޸H`�����d׽��}�.�\�F�{���%9)��������Kı=�w�iȖ%�b}���iȖ%�b{=�fӑ,K����2k.��
d�j�Y���Kı=��i��2&D�;�o�m9ı,O����m9ı,O�׽v��bX�t�����n[2'�>^��צ��{�M�"X�%���}�ND�D�,O�׽v��bX�'���m9ĳ������7����w���NJ%���}�ND�,K�u�]�"X�%����ͧ"X�*��{�M�"Y�NJr~����̨�2��|9(�%�����ӑ,K��#���]��%�bw����r%�bX��ﵴ�Kı ���H�}ffng3/�+e�M�=���lY�������<'d�[љ��D{`�<�X�-�F�'�{!@
�m�Q�$'�����Ƣ#�ѳ��RX�Qi���m8�HuG�)����j"��\\��@01CF�n�����aMv���Q�Օ!	�Q�Ж�ܹ�<�r��gm[Zl���2� ,��Mi(���A�ب�%���k2ۙ ��_�_η~�e�ն�z����ȝk�=�{Lrў���Ϫ �7#s9IT�5jm2\��OJrS���{��r%�bX�w]��r%�bX��ﵰ�V ��ı>����ӑ5�Mz~�}�~���0�Ο/Mı>���?�c�2%����m9ı,O�����Kı=��ͧ����;�/B�צ�����܌P�ɚ��r%�bX���fӑ,K���{�iȖ4X�'�����H�����I�;��/fe�2\�n	 �蟻�z�9ı,O}�siȖ%�b}�w�iȖ%�b{;�fӑ,Kzk�����*f�I�Q�Q�t�zk�D�=��ͧ"X�%�w]��r%�bX���ٴ�Kı?w^��r%�NJr_�z{g���lC�RTY��Ĵ.V����@�y�X�q>ܣS�hG\��5�m9ı,O����9ı,Og{��r%�bX���z�?�c�&D�,O��siȖ%�bg��Ɍ��2�ul�j�9ı,Og{��r@ ��m�"n%����]�"X�%����ͧ"X�%��u�]�"/wN7B�ק�Y}�?���)��bX�'�����r%�bX����m9ı,O����9ı,O���m�^�z���~��ք�0n�7#���K��D����ND�,K�׿�ӑ,K��;�fӑ,K���{�iȖ%�bx�I|Y��\�kY�\ֶ��bX�'��}v��bX�'��{6��bX�'��޻ND�,K��{[ND�,K����4Y�2I�X$S�33\���4���Pa\@fK�Tq�m�gdiI�mFdT4֋�t��5�'s��ٴ�Kı?w^��r%�bX�����r%�bX�w]��r%�bX�zC��\��kY�!5sY��Kı?w^��r�@�DȖ%￿���Kı;�{��9ı,O���m>^��wCt/Mz~���´uԚ��]�"X�%�{���m9ı,O����9�ʿ� ������O������y�ND�,K�����^�z����k�Ƥ�i��h
�9ı,O����9ı,N�}��r%�bX���z�9İ?��3�߿>t�zk�^���{}ԧS�Xms��Y��Kı;���iȖ%�b~���Kı/�����Kı>��ٴ�Kı)���/�����1֮�̫��Mn�Ć���-�@�]N-����6����J�V�p'�>^��צ�?����r%�bX��{��r%�bX�g{��r%�bX���ٴ�Kı/���a�mf����rS����{��Ӑ��DȖ's��ͧ"X�%�����m9ı,O�׽v��bX���}�n���(L�O���5�b}��iȖ%�b{;�fӑ,K���{�iȖ%�b_w��ӑ,K����P?f\��U���rS��,Og}��r%�bX���z�9ı,K����r%�`i�T<H��u"w����r%�bX��̗'���h�M\�m9ı,O�׽v��bX����ki�%�bX��{�6��bX�'���m9ı,K������K�%4ĎRk��`�F��g����/i_cvWB6�Y��c��ӑ,Kľｭ�"X�%��w�ͧ"X�%��｛ND�,K�u�^�|9)�NJr{����\16rU)W[ND�,K��}�ND�,K��{6��bX�'��޻ND�,K����O�%9)�NO���cp�E��mnsiȖ%�b{;�fӑ,K���{�iȖ?���/������Kı:{��Ο/Mzk�^��e�
zJ�V�nf�iȖ%�b~���Kı/��kiȖ%�b}��iȖ%�� �ȟ����m9ı,K��Iip�53��]f�ӑ,Kľｭ�"X�%��w�ͧ"X�%��｛ND�,K�u�]�"X�%��_ �E�,F�F �o=�O7Q�͵�96.����^[G0%���F06"i�r�8{p��\�	�
�*����ͨ����a��\�%�]�`K���Jd@�Y��h�/�Ę��(]� Xb(B�MF��[�@ �KkU�g�>��PAѫ�Gb�!iMp,�
�Z,jڤ�)��� S�K�;����e�ʎ[GRR��Y���X4��YL���Y0շ_ xJ��k</�Дe��k5��6�\0\�,�s*u����'	 ��r-��\:z$�x�־O�,K��=�fӑ,K��w�ͧ"X�%�����ӑ,Kľ���W�)�r��ۄ���J�m���m9ı,Og}��r�G"dK�k���9ı,K����m9ı,O���m9ı,OzC��[���k4d&�k6��bX�'��޻ND�,K������bX�'���6��bX�%�}�m9ı,O}�p�k5dː�f�73WiȖ%�b_w��ӑ,K��;�fӑ,Kľｭ�"X�%�����ӑ,K������rh���j]jYu�m9ı,O���m9ı,K����r%�bX���z�9ı,K����r%�bX�gm�e��u���b��ane��<Z���%*:����æ��8�#Ln�����w���NKľｭ�"X�%�����ӑ,Kľｭ�"X�%��{�M�"X��ק�Y~������O���,K�u�]�!�) B"���  O�}q,K���m9ı,O���6��bX�%�}�m9���%�=��-��e�n��'Òı,K����r%�bX�w���r%�ؖ%�}�m9ı,O�׽v��צ�5��}�n���L�O���bX�w���r%�bX������Kı?w^��r%�b-�}�{[NNJrS���i��~�eʮ�*w��Kı/��kiȖ%�a��$~������Kı/������Kı>�w��Kı?�><�ֳ$2�d̪�N��H����0p[!tRm�R�TưfX����;�qlc�QX�/�?�%�b}���M�"X�%�}�{[ND�,K��~��'�ı/������/Mzk�^�����[i�ɦ�v��bX�%�}�m9 ı>�w��Kı/��kiȖ%�b~���'Ò���'�����g%R�Z�ӑ,K���ߦӑ,K��w�ͧ"X�{�	'�.�|�HH�A�~+.�!!&��'�
P)H'�Ҫn�A|����i���hL!Fd�)��~5�G�!��͑hO���s��x�A���X�� ����J�i�qwFY{�8�D8h8'�0qu��Ɉ�a$]�%�%��GI]�פ@� a� ЯU�� ɉȼ��Mi�s��x@�, �
$�j�7���+�a��G��к���09$�BA�$^R,,*B�K��RE���%%�([+���$U�pCb�|6	#J	�W��T"�EOʅQ�v $>A6qʆ�S��P0bT���&s���r%�bX��w��r%�bX���ٓ=���.��Z�ND�,�P���^��ͧ"X�%�����6��bX�%�}�m9ı,O���m9ı,O����&��Z�ֵ�s5�ND�,K�}�M�"X�%��)3�����~�bX�'}��M�"X�%�}�{[ND�,K��z�t��ko�#e�e���	Q���φ��]�ӝ�ʖ��l�������:|�4Kľｭ�"X�%��w~�ND�,K���� r%�bX����ӑ,K����|�3�2k.��3Z�r%�bX��w��?��DȖ%�������bX�'���]�"X�%�}�y�'�s����'�y?O���ʵ�jm9ı,K����r%�bX����WiȖ%�b_w��ӑ,K�ｿM�"X�%��=7�[���k4d5nk[ND�,V���o=v��bX�%�}�m9ı,N����r%�`EG�(@H�A��G�hU��� &�A�Q9�^����bX�z����c)�ɦ��:|�5�X������Kı;���iȖ%�b{=�fӑ,K���o=v��bk�^����7;,��T%8feb��Rg�Z���rFs�i�-�4�0uԳ��I��3Y�u�eֵ��Kı;���iȖ%�b{=�fӑ,K���o=v��bX�%���m9ı,O���d�{S.����u���Kı=���i��bX����ӑ,Kľ����"X�%��w~�ND�ʙ����?�Q���<���צ�5�������r%�bX������KlK���6��bX�'���m9ı,O|�}v�FV��;����צ�5��{[ND�,K���6��bX�'���m9ı �?w���ӑ,K����|�3�2k.��3Z�r%�bX�����Kİ�c������~�bX�'�����ӑ,Kľ����"X�%�E7	���@V+�,bTh&
�)o����Jen���[1ڮ�H�%�c�q���<��r�y�)<���8A�U�5#7W<��=�!p�-9Y��O�ې��qX��6�2��6��1�Z�CNv��q@����ٚ8�W�Xv2A�)�s�nx8j��m)��	[v	����r�,����g�D7�x��.������8q��F�ҫ+^9���D��,c��&�0����UP��&S�WN��L��q�:��E��7m�]�' ��#W��5�*�O9�q�w���ٕ3AY��Kı=��iȖ%�b~��]�"X�%�}�{[ND�,K���6��bX�'���Y.OK��Ѩj�k[ND�,K�}�j�9ı,K�{��r%�bX�����Kı/��kiȟʄș�����2jh�2�.�k)nkWiȖ%�b_����m9ı,N����r%��ș�kiȖ%�b}���j�9ı,O����1�sQD�����NJI�Jr{�o�iȖ%�b_{��ӑ,K���oڻND�,K������bX�'����c<k&���Yu���Kı/��kiȖ%�b"���]�"X�%�}�{[ND�,K���6��bX��9��>1`]�m�i�| �l�-`�ܶ�u�"z�s��������i@#��(��Q5��35��"X�%���ߵv��bX�%�}�m9ı,O{��� ��L�bX������r%�bX�����n&�f�fj��]�"X�%�}�{[NB���)	ѩ�ب��,Os���r%�bX��w��r%�bX����ӑ,K����|�3�2jf���m9ı,O{���r%�bX������Kı?{��]�"X�%��{~�ND�,�'����m*�eL�*w���NJ*"g�������bX�'������Kı=�o�iȖ%�!b{�ߦӑ,K�����%��f��2Y�ͧ"X�%����z�9ı,?��s�m?D�,K�����ND�,K��{6��bX�'�I��Rfa&���tv�u8%ju��p��=��y)^�C�ƍ��cg�1+�Yj�y>��%��{~�ND�,K���6��bX�'���l�Kı?{��ӑ,JrS����.cnj)�y>��bX�����Kı=���iȖ%�b~���M�"X�%��{~�NAZrS���w�����8f-Ij���rX�%�����ND�,K�����K��+� �F�������Kı=����Kı>�|{܅Q�X����Mgv�?�����Kı=�o�iȖ%�b{�ߦӑ,Kľ����"X�%�ߵ=�b2�Q�[�O���5�O}��M�"X�%��G���M��%�b_����m9ı,O��ߦӑ,K�~��a�n�0�`V�`�=qW+�gFL<�}�W��U7����������'2�Y��356��X�%������ӑ,Kľ����"X�%��޾��Kı=���iȖ%�bw�Ox��kZ�kZ��MkSiȖ%�b_w��ӑı?{��6��bX�'���m9ı,O{���r%�bX���yd�=,ֳFCW3Z�r%�bX����ND�,K�{�6��`6%��w~�ND�,K��{[ND�,K����&�I�!u�YKn�m9ı,Ow���Kı=���iȖ%�b_}�kiȖ%��
:?�?����ʁ��$r��f!:E� _�SJ���=����"X�%������1ssQIngy>��%�ﹴ�KİOg��m9ı,O����"X�%����6��bX����Oށ;�� g�!�(���݊ѓq�w�=\T�Ԛ�˭���4t�����2��渟�X�%�����ͧ"X�%������Kı=�����D`���,K����ӑ,K��	����0��\U���rS����������'�,K��{�ND�,K�ﹴ�Kı=�{ٴ�H,�=��e��%̳%���A=��fĐI���&��'�{>��iȖ%�b~ﯸy���Mzk����ݷ�h!�8ʳiȖ%�bw��6��bX�'��{6��bX�'����ӑ,K�=�����JrS������Ci��*f���"X�%����ͧ"X�%������Kı=���ӑ,K���m9ı,LM ���^�I�I��D\�a�Y����[�����)�qѵ�`��x�\��]�32��[�s���llڶaA@�[kmn3���m��r�m��8u��T�0��m��P�غ���ml�mB�dN����1�#��;`�0�5�W����/�V�qN;msB���lQ&�3�C��#�m�N���H'rL��2I;��5�����e-�Ӻ|�Xy� ��Ri�B����gE�ܚ�Eag�-1�\$@��g������P��Qs1��'�%9(�'{��ND�,K��m9ı,N����r%�bX�Ͻ��r%�NJr}����h�1+��mY�O�%8X�'��p�r%�bX��w��Kı=�{ٴ�Kı?w��6��S���������6梒���|9,K�﻿M�"X�%����ͧ"X�ș�_�ND�,K�����rS�����z{Ln��bԥS���bY��0r'�����ND�,K�_�ND�,K��m9ı,I�3���G)�r�tJ���,t��K�fӑ,K���_p�r%�bX��}�iȖ%�bw�ߦӑ,K��}�fӑ,K���[O{0��4[�bU����5��:���x;�=K��3r73�$�c��]&�uKVw���NJ%����6��bX�'}��m9ı,Og��m9ı,O����"X��ק��_�zXh!�8ʳΟ/MzX�'{�p�rQ���B *��S�9��Ϯӑ,K��{}�iȖ%�bw���"X�%�ߵ}�P��
��e�t�zk�^�����]�"X�%�����ӑ,�!�2'����iȖ%�b{���6��bX�'���Y.OK5�ѐˬ��r%�g�)Ȟ����m9ı,O{��ӑ,K��}�ND�,K��}v���%9)�����Ҙ�����|ı,N����Kİ�D�>����i�%�bX��׿�ӑ,K��}}�iȖ%�b gН����ˬ�pZa�hF��j�*Y�2ʺsz���m�-���=�\*B�m6�9�f�>t��5�X������Kı;��iȖ%�b}�_p�r%�bX��}�iȖ%�b}���&3Ʋh�n���6��bX�%��m9,K������Kı;���ӑ,K���ND�%9)��C�����b�,\���rX�%��}}�iȖ%�bw���"X��`
6�PB!"��!RAj�*�*)�8��P�7=��m9ı,O���6��bk�^��g��v#+Aq���:|�5���@����m9ı,O{���ӑ,K���]�"X�%�����Ο/Mzk�^�K����)����+�iȖ%�bw���"X�%��! S�����~�bX�'���m9ı,N����Kı>�_Oe�4�-�6X$SteR�8�l��GR%��{i�NU+²�0�
ث���'Òı,N���r%�bX�ﯸm9ı,N���A9ı,N����Kı=�����f��2��fӑ,K������?��L�b{���6��bX�'����m9ı,N���r'�TȖ'}���&��,�]kU�u�iȖ%�b{���6��bX�'}�p�r%�X�'s��m9ı,O���ND�,K�Oo��fhչ���B�Ѵ�Kı;�{�ӑ,K��{�ͧ"X�%��}}�iȖ%��
�SPl(E Ad$a��԰E)�\�BP�PJ�e����D�N����r%�NJr{�=�7��5�6�w���NK���]�"X�%��N��iȖ%�bw���"X�%��w~�ND�5�M?��=��[��$���Q���3q�L,�x��ڰ�2'��c��:�kSSZ֮j�9ı,N�w~�ND�,K��m9ı,O{��� �%�bX�����Kı<g�{V�jL��j�՚֦ӑ,K���ND�,K���6��bX�'}���9ı,N�w~�ND�,K�>���AM�U�t�zk�^���߾�6��bX�'����9ı,N�w~�ND�,K���ND�,K����.�[uB՝��rS���Na;����9ı,OOo�m9ı,O���m9ıD�=���ӑ,K���Jg����a�Y���Kı;���m9ı,O���m9ı,O{���Kı>���Kı8��X�<-#>8F14h���Uq1���HQ WL$d>0�?�$f�,�H;� ��4��,b l5�>�7���C��L�϶��$���5%I��6Ec�P��>"O��$?]�6�x�T�� �`���Rl���$��<��zu����f�0���T"���.i��2�(�v�i5�Ȗ������c	$�# ���,b��T
�R0c�E	|��O��l�~Q�M�~.�2#%	Wh�¤��R�7�� �-U��:�R̓?�Umn�Pb��������Y��m���$�w'��`�û&j�j�k�WQyb��2�6�5ذ\[��`�U.9�=�+=�;�'�4�;��Q����]h-�D�Ջ��4���-�t�ń��]�Pܚw ��Ӭl�f�j98  ��'TU��J1�vu��l����b����W�aX���k�фSuNr����r�l���I�@�M"�+������v� v2��ѷov�����;�q)3�����b�����cd���<�n�=���IEm��,Ɓ}m�	Yfy��`T�
g���r%�˲����h�!����As����s�8���5�6w0��$x7l%-gh�D�Pq����:�;jmmL��r�v��Q�I�ʠ1���5	��ڀ崚D��6h��vh�R���B�5�����ѵ � éݻ]R��[�-TmJd0i��j�U��M�<)��"n�θ��N��ӄg�l�)6b�%P����	8���\�q�@��2 ���X)�=v+�-�u�=�n�6\-3��K��"*M-h݅ta��\f���lC�A-����m�6-�ND3�Q�sݭ�P;Rl�]�F#*�:��x+ֺ����tS˵�� h���N9��"7��=o;W�U�:C[C�!(��#`\x�	�s��e��[���<k&Ʃ�d�;�f���2q�x�@��R8.`��ב)`� �\8;`�ʎ�6��̈́��h�%��wcr&�p����azک���t��]�rInSuX�vq�46�Dz��(jj�KMU������C���\�у��]6u�y�:2-Kl��%涸0�g!gm3��Oő��L����+�Ρq�=X1���&e�5����Z4�)L�t�	�R1��Z�u�V��*�m/e��a��PVĠ+1Y4N���� ��#/kg�uk G�I�+�]'p!�܁���U�Y�Z��5��1����C@�����
E�4� �  iS�?'�&��DS�~;��YKL���.kV�3M��İ���\q@�e�3�0ݙ^��]�ڝ�.ѷ 몏YE��h2�jb��kx��e�tΖ�\$�Ѥ��WXR��W	a�� M��M�g�jHj�	�'A!j�zZ*w</[rk��'eݶϤz3��e�
�s<&��yz�.��0�D�b��Q9�u2����l)�pNt��z���-s�Oz͇��]d\ٶ<��䛜���l�^�&�%�҄rJb���[fb�f���=	����N�E�V3d��ew�O��^���=�{�ӑ,K����ND�,K�뾻�~��,K�����NDצ�5�����o��h&r[p�:|�,K����ND�,K�뾻ND�,K��ߦӑ,K���{�ӐKı;���&3Ʋh�n�e�ND�,K�뾻ND�,K��ߦӑ,K���{�ӑ,K����N��%9>�y=�k����7��"X�"2'����6��bX�'�����Kı=���ӑ,K���>;�yz���^�����f�E0�Z��r%�bX�����Kı=���iȖ%�b}�w�iȖ%�b}���m9ı,O�x��m�&&h)�.ӳV�wkŮ5;��їq�;��Mع���V�SDq�g�>^��צ�=�{�ND�,K�k��ND�,K�N��a���"X�'����iȖ%�oO޷�����L�r�:|�5�K�k��NC�(���8�&�X�z~ߦӑ,K����ND�,K�{�6��bX�'��]�i��j�a����r%�bX�zw~�ND�,K�{�6��bX�'���m9ı,O����9ı,O�����nB�Z�j�ӑ,K�����"X�%����6��bX�'���6��bX%��v��iȖ%�b}��zeѩ�����K�6��bX�'��p�r%�bX+�o��i�%�bX������r%�bX�����Kı?�?��M��ett	�Z�X��-H�vS^vD�m)�υ�g��q���/�g>�Ӯ@�.�6��X�%�����m9ı,O��ߦӑ,K��������2%�bw��iȖ%�b}����n��ѭjjkZ��]�"X�%��ݻ��r%�bX�����Kı=����Kı>����Kı<}����je���˫��M�"X�%�߽�ND�,K�{~�ND���}�O� Z�Y@�00�T #F"$���SH���O�;�o�iȖ%�b~��~�ND�,K�=�'��Lֲ��\��h�r%�g��02'���6��bX�'����K{�^������ݬ��=����lT�v�� �{���Nɕ�N�����4ˤ!��6��i-�n��Ad!X��R	v1�k��gV�>����n¦����������7�e`���W+� ����;#���f	���&ov�s�����'A~�?��<g��Α�Ӧ]�M;(V� �߼��K�>�{6L�WIJ������wV;k ;$y$��v�I������@��4(/�z�=ՀuQ��ɥc���cm�`�e`v�XeȰ�n(U�Av�m�����l	�꓎��[�"�bS��w۬JJ��1sN)�j�Tsz�{�g@��"�;.E��kny`�U���ڧmZV�`v�,�6^�v�,Ͼ{����9���~��m\�u@�z��~X��ذ�\��RSg����,o7��*����)�m����X�fV�ob��+�9W��ߖ���N�:�����5m`ݙX��*��s��;�X��ذ�TW�ʿL<�պm_�3��t����q:�䬰��tڻ=�с�.n�1�m��u�@� t�j}��+�;8�vWk�q���8mv�6��8
�N���xۣ0@��8��f� M�=7��鹀^��^�C���Sh�VȺ�V�ؽ��G;9w���}θ����pBM� �����v�qm��$g|a�Obm>\��0 �Cf�^-4ږ.���$��~�M���s��=��69u�z�z��N`<�6I�S:�M�!<��.�;f�ZӦ]�M;*պ�'��X����^��\���-=J��ɫN�'uc��wc�>�{;�+ ��"��H�������c-�m��۞X�̬?W9Ļ�<���x��ԁ�����:n��&ɕ�}�ذwc��W9G��ώ���k������wm���X]�x��ذ	ݙX��9�T���R
�a�.��F]���-�hQv�2�`M���[��Q%g(V�i,��-�����X�̯�U\��wny`��wIY�]"�i��>��ş���Ă �~Sc���w|�Xv�X]�xۮ�S�N�*�63�[X�̬��Ň��\K�g� �m�,�#�KI��M;*պ�>��X;��Wob�'ve`t��_#��t���m`�ǀ{��r�Z��{g���{ݭ(�|I]�Pr��%�z+����م�[�]ή`R�:�Mn�l� �\顙��Dɕz��y�����΁�ob�"���%w��Q�����:n��'veg��W9I۞X�x��ذ��)eZ�wj�v�m��ob��������U9t8�j�m�B*��"�����.�7d��;�eԲ��m�`[k��W+�y�,��<��2��{7�N�+ ���LN��>��ŀI�+ ���`����q�݅:�����k]�T�4z��`����p8F�5]� pB��eɶߤ���{7c3�n*�$.o�>���g@���`�c�>��ŀ}�t�Zt�[I�e��`v�,����s�vz����}����$E�R�|��۫b���y�t�� ��2��r,*?��O���r+����t���O�{�nI�}��rN~ϻw'@��B~H�NvI'z����=�y����.ڱr���+ ���`������`]�sQ�c0����i�#6��".��(�J�AƷc�����5b(��A���wO<��_f��v�[u�6_�, ���v�/�s��v{+ ݌���`+l���X�v<`wfV�nE�����D���g�5t�����wK�X�ٕ�}ۑ`����]\�c�%bm�e
��>�̬��ŀwc��+�����;����b�i�e��`v�X�v<`wfV�W;r�;]SmZ8'�#Xw^���HGO�O.i0�]�%����x�����/�ݪ�Xګ�'{��a=s;�=(�!�@f9�y�7lq����9B�׮�t�Is��`�4���!�)�ڙ�-;{q�w�,Սs��n�US��1�Z�X�+�!-��m�
P�	e+-����q�٣��h���X+\�ΰټnq����;��ݭ
�$zF{;�wf��`1�j�L�ۆ��ZhʆuZ�x���u�r[�.8��t��븻e)jQ�����t�� ��2��U�U��l6_�� ����o�;�\����q绠~�xݹ }�~�W=[˗�\l,n��m[� ݞxݹ�����]�?~x�^�xQ�R�RmҴ�v����܋ >� ���^ w���]K���-��� }���s���^�} �ߞ�nE�M*Tʻ��I[Tvݩ^�:fvwg��{3f�]e����@0Ӷ:�ˀ�n4��*h$�U����{������r, ��<��W)��I\�֩�Y���'?}�o��$d���1�&ƿ�DM>T>�g��X��<��e��$w��t�l�;��ݿy`wc���Uq-�'� ;=�j�)Z�Gj�Չ1����r�-�� ݲz���v�X��ڻ�v�i�-���7c�>��}��`wc�?r��J���(٘J��5K��0/2��N�y7bwg�@��y��t����Y�w���C��*�@����t��, ��x�ݏ �!RX�����v�ݳ �ob��ǀ|����8g��ĉ��^�I'e
�&���d��>F�x]]i\%�|�s����Gr� �����&��2� D!F@�F0� X{�9��%�JY�w�v�I��1zl?~?�X�6~V6�` ��jh~��}�(��P�֞'�GZ�g�b]j6�F�D+"cu0G�1�&������6�[5���6q�xzU0�|�u�? �?";>Ez����!�Qh��H �PC���^*�Z��}o��� ��X�Z5t+ ���T1�������ܮr��<���~�c��C��E�x�0��, ��x�ݏ �ʥ
5yx���u����7�l�Sr�s��F��ۈ�s>U���2�L�C12\��>������ǀ|������W;a����R���;��HI�v� wv<�ʪH�$��;=����tm]ʻM���o ���l�X~�*���� l�x���b�acwmڱ6�?r�UK�g��?��x�U�u�z�3{�<W�bn��Mګ�f���s��~�*������5��}��E���:�m�E�˫L��C�u�ߏU��[���i�'IÛ�uN\�P'v�Ŷ|�<�	�$�� ��v�j�VA]&�cm��Iy��s����r�Uvo�ߖ��� �v<�\�RGd|�S�4"���Ս��s� ��{��$vO<�g�x��"�2ح��N���\�r�zL��� ��K�>[��P�]���v�Ę�ـuwe���W9^�{��[�^��	�Э"$z+jŌ (.�	�w2q4�d̒}��U�Ǜ�5�Zz�r� �ٺ��uɴ<�ֱU;$��@���a[&���av��S��gE��[��R��Ɖ������ۇBtvPiK��K�h�ѫv�I��L� ͮ�fm���	P-�2��)
��m�KY�rNű�Ћ��k6�ɴ4��.�K���n@�H�qEdŭV�-�:7�,\Ph�]�/<��z(���N�q�Ӻ}��o
|��-u�h0Z=�l��C�h h6y���3�{^�!'���l+6+\�9ށ����/d������W�5l��[W/Ը�j��n�e��>]���8`]�x{d��DB��4��i&�U�k �c���Ň�ʮ%�g�xv��vk.v�vP��j�6`Uqn��n��^�����h;�wPCWI�m�{d��~��s����7|�`�N�|g�_Iy�Τ6�,M`�DQ����1�4��.8�N,�c�6W�6֯7N.MZcj�� �k���{��\�U|�v�z�	���n�lV�e���'���f�" ��l���뇻�e`�{׀vk����TMZubL�6`l�X{d���W)-���7���"�m��:�Ӷ;�u��UU~�r��0���	<�f�`vL�k�{r�-Swmج�x{�e�Xݓ+ ��%��)9WB|.�_���m0�2���0�wi�N]�4�A7b�[�]�I�Ա�"��)��m�zO,�ɕ�ol��Us� ݏ��������[����}�2�ܮq"m������:���s�9\��=^�w_�5t����X���^���Q�
�og)}�O�xwfV�ɜn���J����n��8`��`�X��/ ݸ ��L�+h��l�;/b�=Uʪ������g�x{0��r��E�0�D2s-t���T\��{^v8rY4C�9��#e���!��2��d��n����V��K�;��v^ŀK<�����+�:�q﻿�I-7|�`�X{&V~H��r���-Sj�B����~0�ذ�L�{�}��zO=�h����m����N_���nI�����>����ɤZ�H��D�|(9�w������م�4d�n�T[f�ɕ�~��z�w������>y=�v�4ָF�MeY�n� 
5�D���e�[k*l���f�y�Iǐ�7򡫤�V��&��^���\0�L��8�:��ҧVյcw�w�� �/ �d��7�Ix��E�e�[E��f�{�ɕ��Ur�W*���߯ ���`J��Qn�$�N��;�2��^����,*7h���ն��;�X��/ �\��U'�~�~X{&V W+�syJ�Dͦ���#D$I���y�i�1��9:`y���m��*�q�;J�Z���7��l�NQk��.��K@�'��a7�`�z�۠����a^{=5�cOP �yU� �+���Y7:�کI՘	-j�Ӎ�"wfN�L�;��u'���Έ��Q�n,��@��mjv$�[�;#!:�D�O��u5;�:}N+�A�V���-k�D��&��\�\O�M�zKYm
m,�� �`b*i��	�-�AG�bP!Y+cLmզ!�]�	��[�R�;�=�e�X{&W�W9\��&��^�x�궮��ݫ�`Se竜�)#w���&��^���Yp�V�.�&�����+ ��%��p�;5� �ւb��!�MpB�X��/ �c�����+ ��g�V촩յm[wx{0ۑ`�X{��n���\�]��3B�]f�7�ma�c%dGrO�B3�CZpR�6�fh[�(�,`Ķ+h��l�7c��ɕ�w�%����P�]��e��Bl�;�2�k��6k����c��r,*7h���ն��;�X{r]��p��)/�Xｕ�v�W���-Sj�Wn� �c��r,��+�)n�z� �<T�[��ݫ�`�"�;�2����;��z�U[!�_;M	RƁ]�)���]�V��ؖ�t�"�V[O��ta�U(��\W�6`�9<������;ے� �c�k��L�h&+�R��+u�w��0>�^�eȰ�L��ɜn�[�Hum[V�����f�_��܀�	���T����� �0�L�Wy\�_*�5μ��.���*�2ح�Ui6`�K��G�w�%��\�*����^".�^Bl��)�w�� �n�z��7|�`�K���{e�Su��5��(�̥(�G�3��.��#6fi̈́м� ��(J�-`�]]���$��;��j�/ �d��;]��]���v�Zn� �c��r,��+ �U��H�<T�[��ݫ�`_���L��IW�w�� �u,-�M�I�M�{&V�nGx{0=UU��*���_�` 	�w�զ�![��܎��8`�� �d��$�S����ƪ�̰ne�S.ck	V=�5���˷iC`��� �9��gkH��9]�>����y���;�2�ʯ�wo�w�l<��U�e�[V��l�7c��ɕ�}ۑ����U�E�*'v�$�Bl�;�2��r;�;��n�*7h���t�M�N���nGx{0�� �d��6�W���-Sj�+�� �c��Ix{&V;��}_]:8QUC$�u @��\�hJ���D���B�$�bA)�"'G%T0�>`�Q\ȝϔ?3�:;C�k5L]"��  T"b;h�ҥ�F��i��FD�Ѣ�f �	G!� IT����@�!�4�	����?�������Fh�H��� �0!۟�`�;����ĪB5�7HD`П����3�$�7�󾪪�*��UUB�*�����
���L֊�6��)]�&ˋ<F,ٛ��3h���st�ۗs���H��j��,�lv'��v�݇n�\X�@Z�F�[5�ɭc1�`�2�F0cq�EW�̃^�;f�aC�䱉¬ۃ�&7aW���<Q[J]�`�H�f.9$66���#�l��.�;[Uʋ�n)Y���;��$�ct�n,����\Թ�m�7R	߇�_&���r\L��vԬYeؕy�<��D�y����ۢ�,j8Be�u�Z+�#��@�0m����(�v!�����;�Jp��Kn�4v�[9Ҵ�m��5c����AU�GqrnkKgg���\t=�m�۲^[m
�ol��,���UN>>~����,�]�������ݑN$+�\Pe+
��J�m2gR	;O�V�;�k/&��0�m�xG�X�f�j�l:�:89w;�^T���v�A=�P �%6��u�Wcb��n�B�ۢ�+�LMC!�e�c[{\L��:D�0�uќ&q���po�����8*�X2] ,��{d)L)�ˡ	4���e%@5e�3����Ig���$�����&7l��G&܄^ڣ��MsH�qf�.pd�5�1�\1�u�fsC20t�p.�����lg2��6����"��L.�Cs�ys�tT6:shU.c!������kU�i+T�3�p�GG���<�:�W���j�N�;�ӫ�y6�����$�3���w)9T-��S���7`�c����*�S��n��,�d�T�$p�gv�fm����g�����;UL���y��ې3�Q��OkhH�[si��Y����#[J �Ӭ����+d#��p;{eU�n��3���K�v��q���t�N��E[��>Yբ��;h�yv3�u�sӍUt�+��R2�ܡ]�o; S�sQ��\6�ÀWB��G]wdN��N����Ŵк�kp�X01հ��)��t�Q!����B*)T@��M
W�S�*G��B�,E�'��@�g��w�a�J�g
8��٦�Y�ff��F���P�r�7{wq���b
m^QИ2�(���l�Au�Kn{`Ո�Yh���t4��phq�R^6d2�2� ˰8a�YH�s�X%g���q��^5��w]�D'������X��cQ.sA�%�%j5�l�K�7@G!ӣvNv�f6٥C-�(��#
:f�(;T�Gb%�b[,��t�6fm�e3D`�9;>�rN�O�6'�F6;c�=����U`�G����GS �~�=��c*ha�e�nK����#�l�^�� �d��'c���8`Jeԫ�C��e�ۼ��+ ��-`�p�"�/?U$M(�W~)Zb�B�X�?Z�;�ᇪ������� �����&q�v;I�ڻM�X{0�K�;�2�	�j,�G�J�L�+j�ZM�]��sw������;��o@�q�PZL��tmr�.��`��8��x�.��5H])l�A��Yt5��j��I�����X�j,��Se�Q�Eʺ�t�M�N��I;������ mb�P�$�W-���nǀw�eg�ʪ���T���!��6��IZk ���j���;�2��� ��j���nՅ�0=U�R�z��{+ �����8`m2�R�Nʺl��ݻ�;�2��� �c���/ �ꭕn���Fu�۵"��S;;�	�UQ
ź��F����c�
�0l�T�����|����;��oob�r��A��e`�>y����&ݷ��<��ԓ���|`��V�cQ`�t�ڹL��mZ2�jnI����rO߻ݛ��I��V0"x�@ �T-;�}�_�`}�~0Ү��TB�i&$�X{&V�n)x{0��X��ۢS��ul��N���n)x{0�̬��+ ���$RvЕ4����^�&8pKz�U�KR��»�R�,�WIw]V�6Z��J�;�;��ove`�Xݸ���R���amڰ�f�ٕ��RF����;����7c�&�.�+��.�(�j�`�e`v◀n�{�+ ޕ��wPCE����u��W9T���׀I�� �ve`}K�r(UIx�Q?w��nIϾ��ɬ�ڥV�ڶ���� �ve`�e`v�K��QEL,M4�e!r�L}ٮ����t�k�χY�e�vt��G
��u ƃJڵV�f�ٕ�vI��}ۊ^�0Ү��TB�hM%v� �+=\�$w|ז'��{�+ ��[tJL�ulWt$�`v5�0�UW8���}�e`�d�4����mRV��7c��ٕ�vI��}ۊ^ҵJM&閛J���fV�&V�n)x�p�UNY�]`�x$�Y�JNv�*���uat���ZG'Gn�4f��6J�2��@��Xؽ�VĤ\�b��J��e��җ&���xS��ʭ6c@9G9�W��! a{'����g陸D�sCa���[a�Rі�BN��ɴ$q����<AJй�BP�M�e��,�Y�.{<��$e��쵎xY�R��`����J���������{���<�R"&XEK��l<+e�7����>K��ʻН�PC\��C��)�.�y�1�������>}�K�7c��ٕ�oJ�һ�!��\I]��>��/ ݎ۳+ �+?��7Ϟt�i��WI���k �������;$��>�����Vժ��0�fV�&V�u��=ʮs�Og�iV�h�!7`�۬�L���Q`�� �ve`���uJ�H� ��4x`YD�n��l���\ϩ��6`��	���Ş��{%v�u����}�2��2��D��r[1se���y篧Y�NI�g*��a����'ve`wZ� �颕m&閛J��۳+ �+UR]�ז'��{d�W`�X:���u�vI��}�j,v8`n̬M(�+�4�)�	]��>��W9\����;'���2���۵���vq���˛,�G�zSY,\���МYN�2g6W�h�ۚ��1�[�Zށ瞾��ٕ�vI��|����%*��W��Vժ��0�fV�&V�u����v�n�]��I�	�]��;$��>��Up��Z}�9M�n,�ٕ�w�Kn�I�N��wE�� ���XeȰ�fV�����x�3΁��&�
�XeȰ�fV�&V�u���D9J�|J��m�ڎ�uL��2�ue0�v����p^Rx6.E���t��n�i�����ٕ�nɕ�}�j/r�A��y`l�z����e4��n��2���ז��y`n̬�@�]�M��Wn� ���vL��|�Z��ue�5cn���qo����?d�X�W8̅!L�dj�������IK:u��4��T��N��&Vٮ��7nE�z���-��]�X���H������-�+\�%ʽ���"\����܏\��D��vX�)���M%m������w�r,�{t��j�յwue�Xw]ŀn܋ �k��&V��N>4ؕ16����7nE�}5� �w]ŀu4�v�n���WWv����8`�w�\�$�z��z�1�~�i^h�i����wu�Xv�X�\0��s��ߴ��~b�p�f�S8���m̩��m b2#u���u�-�]>�`�	�1��-kL�r�c4����Z��j]ų��]c��v�eMZ��ꗭ�����+�;�]Rˈ%�;F�	h����	� ���k�-<�⸃c���vL��x\"ݼ!�D�y����Dqf�T�j4�:��zv�֠��i�t,43l�	vc.)��w���O����ҼH�3�؅�l�F�f"Ys�ʗ�D��ٽqf6���$(�e���;���Ȱ��`��}/��V�.��&�m�Xv�X�`��vk��	J�D���4��\k ���0�wݹ�P�V�*$�@��`~�r�T�{<`#�,�r,/l�����z��ulWt�l�;5�X�Ȱ	�p�;#������Ik�maɃ�	��=Ul��C�y�����ݳ>\�hG�m�E���6�V&Е�_�D�ߺ��;����XQ����2�i]�m`�ᾨ`�`��@����+���0 ��v�R���Ut�@�ـwc�ٮ��;�� �k�6��(WƝ��)]�f��q`��}5� ���W�E�JW|iX��Xv8`Mp�;�� �븰�r�ۡ]�n���v��i�nF.]g�%į�|���l�X:9.,�չ�7wM+j�X�0��`��wu�^��?�X�*�v�@�J�0�p�;-l��0	��N�)tJL�un��-[0�[/ ����Wy2�Nk�Q&�U�:�
�r4��Q���xN� h �h"�Dݬ�]]�HE�E����,�#Q*�Z��؃�N��ÇS2^~Gi�cBD��Cf�c�NQN�ߴ&�'��b2�I��ѻCtti�f����$P��!ϣ$�������I?~>���򿘜9�_�66���u�b��u�#�� ��>�H%#H"�IFY�Mg�H]pX0$ @�+j�h��Q�D�D-�`��Jp2 �D���䅌�BH �����R����sRϏ��~eM�ؤfB�H,D��4��c�6G�h�+�C\Z1x~�E�b,!��1`	���SJ�/QQ�/D0?<	V&�:Q�|@:�&� b"Q:�׊�Z�}��r��`GB��-�ƪ���w��r�Kg�����wc����ݿ޻淪�寧a�e�]�a��8`��wml��0�J�h�������[�n�U�I�V�fg:0���n���Ki�/�H��Gm=���0�[/ ��W*�ϐw�~0	��Q�|I�M��ݶ`�[/ ��p�7c����QjҥJq�V6���8`�� ݎe���v�¬����2�j�&����}�uٹ'���ܞ_����i`��s���nI���e̘z�m��6�v8`�[/ ��8`+J%�
�k����%Lskث:�sx�mӞ
��l4�0�1�	��%ӫm�|�l�;��^�0�p��I<-�>~��y��?6��QJc;�;��=U��q#���l��wml<��N���Y����ئ���~0�p�;��^�0��ڻ���j��[f�����S׀wc��zZ[J6RN�m�� ���xv8`H�wc�u\N�[$�^�ސ����R]L N��v�I�ےR�;�u��Bv�ӓ���q�S�m��<��C�@�qۧ�6�==��)�Ů�H��rk�͹���ǔ�h�N]:��gmӳ(a�'Z���,�gE�C�q&�g{�����a3���\�ɝ�d�c!1�fh6�ps)?W�L|�j��ӵ��Ɛ��ϻF7�*���sn��y��	��ܳ��nٞ��̺���$���A��7jG./)a�h�f���Z+�[m䬦�\v�iDN���T�Uci������0�p�;��^ڗ
��Swt�i��6`H�wc�ݵ���p���RD^�hEz��մ&ـl��woc�=UĶy��7���'n��;EӦ���ـwoc��0�p�;�� �Tq��hWm�ݎf�`��woc�V�ʴ�!�n��,��8����2�HF��$������{�;�������[	F�an1�������|����{���u[Wa,���pv	� ����TJ��.R��\���s����U|�w����p�;5� �KKTtĝ�m�� ���xv8`��wc����J�R�8ҫm�ݎf�`��woc���q]Je�e��X�0�p�;�� ���xv8`���s|S<� �XƠ^G-�A���ԅ��.�)^-�.�6���re!�)�.iU>翟v�;�;�� ��v�K.X[����0��w�wc�7\0�p�$*8�ƛJ�m�]�x~�7$��k�r��E�)� [�/��~0�s����ڻ�[ݫlV�[0	��wc��{���u[WbS�M5��	� ��ܪ��w�<�`u� ��[-�m��0���ݣJ�*�K��*�[LHNۮt;<0��v8��]@E�R�a�[ݷ�7�o ��n�`��}�|�i\wV��j�m�xv8`u� ����;�;R�˺��L�i��6`u� ����;�;�� �ܩE݈�V�7m$�0�p�&�˼����/c��b�Q�	��'����s��}_�@�a��b��av�m��=͞����ݎ[}���=�}���;��a��k��JG/��h�N1t<��#�WmXZ�6e��wI����w�<�`u� ��m��>�+j�lwv��Z�l�&�ݎ��w�wc�{��W8����Z�t�e�6`<�`���%������--Q�v!�R���UW+���]�<�`��wc�����F�.����wxv8`u� ��m��6�;ʡQ�K$�{���I�-��f���%�յ��.^��6�:+#�1���2Cs��\��M��]7>��&H���8Ggq�^yw=+�|�r�ã�c,�umF< �3�3�T�pN5�Im��'zl;���.A��on�=ۋ9n����Ɇ#$��V n��2@�M��@v��[��xJ��1�f�]�ha��@#F�]����m*0�,-,vV6���%����w��ચU99r�3!2k5�Mu�ú��C��a�hur�p]�xv�7mO��a�jwI�Sj�4LU<�?����X`oe�ݎ�V�wqU��7CbVـwc�6�]���vk�T�K�Wuv�.����;�� ���0�\%:��b�m�wm<�0�p�;�� 7v'�}�V��j���[b�jـvk�ݎ��<�0�\��^��|]�ۊz��d�F� �j��w�~���냧*�8eAu�R:.���h<Ѧ �}�~� �؞ݎ�� �G� �(��tĝ�m�� 7v'�T�r��t����@sk���+�/��p�W9��>p�7u� ���W�E�#�˧j�ݶ�ݎf�`����;#�Q��*�j��ـvk�ݎ��<�0���X�ݺvЭ� �� �؞ݎf�`�jn�cIIY�62	M(ٖ)f�p�����SѺ"�¾�L�*8�!��y�N�y�נ}��vk�ݎ®�X�iS�i���ݎf�`�����m��\E��ڶ�jճ �G$��uٹ�b~P 	�CJ$��<{0��ZD�ӥj�`�0�p�����p�>�� �KZK�%N�+���0v�<�0�p�;�� ��Ի^J��e�yw#����Զ��<�TXy���8���dF�Z�l�u�%�0h��<�����o���p�7j�,��V]F;L�i��N��>�� ݎ�^ŀv\� �+B�EV+�V�[f�0ڽ� ��A[��ul.�]���0=\�r�����y`H�7%ã � |ªA	B
R�F*|��_�7$�L�v�q�j퍴*�k ���p�7j�,��C��'Į� cj���#C�c(���k��r�/<�.A�f��ѭ����[b�+k �Gv8`�{������ �-���]:V�i&�v8g�����X���oc�z������z�S�Jƨ���}W<�ˑ`��n�zU�KVKAwM�����ˑ`��n���b�;.�e�c�ʶ����{0�2�W�{� �ܪ�UW9���U�� U�A Uj��" 
���*����*��(��"�TX
�X
�@`*@��A*
�F���Eb*V�
�
�Qb�E@��DP��D���B( �� ��@
�"*D�"�
�V"�`*��"�"�� *�b��F�
� X�,Q�F�(�H
�A��D ����
�X",H��H
�",
�b�� *�"�"*",�"��B�",DH���@��@D�"�T��@T�"�B(� *"�",H
���0EO���*�� U�DU��P@^ 
����*��" ������ 
����*��DU�" ����d�Mf(�����f�A@��̟\���64�k(  �@�n��U@��H4��@ � 
I��(�   <�T��
���UD@TQQEP �HD�T�*� HHED�D�EB�UAE� ��$�   ��( 
   �c`_}�f�n3��}�O�����x }7�y��=��zy:|�H/ d}�  7�Ň' =� �K�,\��w9by� �Y<�q�������� �      Hf ϫ鹝����zk�Z��p��!ێ�h�{p��y`u����S[:�['�u�bi� �����W�� <���oN�.���ǳ��;qO|� ӽ)2�lN]=��v^�绍[��    @P����;���o��.���^�� V��1��8�ݗ'��u=}��)��듽�����9� ���O��y���������םo>����|[�JO�P4��9�)���q�c�����=@�    
)�w =�Su��y�ڜM����8t�AAe�AL@)�� Y�)�� t@=(��:P\��*�h�AB�8 ;��*\���f4�� �Jh(w �gE)L����(�� �#JP (  �  �� Δ�b�����@�e(��#G� >���rݾ���h�;�Wܠ��r�9:� ��p��x���(z>�y�.�{{ͩ8}�=:FN���  zBM��@ 4 i�4���M�#@�=U*'�$` �'�T�Oe   �����R�i�42DHSeJSP� ��M�����?��?�C����Tw>�K���$�DB�j��@EUР����U� "�������S�O���h�B~)R$��6˰��rXl�?���|l$����fBM��JB�!��D)-�� �S ]��\�%X��4	�#�%��h�&2 IJ!	 UkQ��La.	" mH�� �X	�&��d@�"4&�'�	�i��PJ%A�Ҧ��c.�����)r$(�:��Ԥ.o�g5i�9��J��\�� �(F: R]��M	Ӹڴ�V�s�I�ml!$,�N�Xp1Ӣ8��B.�@�U����?0ֿ���<�Ë��p�%&h�.(
��,�k|xXU�A)���l)���J�����AB;��IV�M!R��̦�~Ĕ�}$�.��3x�t��E!p$~��G_�0���^&M&�uj)�Z�*�yH�ŕ��.�uF�/m��!"9M&�4�p%�K"A�$5�o��X�`Z�XP#A����Zk	x�����[�2�滿B�^�d	"�2��DJbp"�T~C!�4���X���D�E]�~
��%TU8�;gra��2�)_��$�h��k����̦k��B�].����\��4��6�~W�g���Ԑ�y�_�ύ47ȑ�>�dsM	��5*lֺ��F���*�	A�!LP���D���a0�m����d�RIp%0!)h��H����c�� �!ωqԬ	��If�#B,$ka�O�0�v0�*�$d�F`�B~��~�~!�$c�ɰ͡kD����@aa�!	4\��vGZ��đ�L�d"Fn����˸�VF��O���B���C&�ƣ���A!4�	k-�F�
A��hٰ܇��J�� ��1���É"Jc$d.�nMJ�B�����G�)
HC�5��~捲�!Y���Q��I8� ��!��a:b�0"E��5�2n_Ą*B�� &$Y.Jo�B�5\�C���J�������!�mw	$��!8�W{˅K���0�#l�����{�g H�^���S4ƎH˰��ς���g8�v��}�����$H�d,Xᡅ�%ȕ�SD4F���Ԍp�"	V!L X�HS ����0�3|�r�$H˚���D1�]7�F*�sP����a������wm]�}��/<�z����J&�C�M	�@�GY��ۉ��2D�#(O��Ø�ɨ��[�*Q6��%�p68HH��`Y�2�\��n��sz�F��y.��2�+&��D�&��AJ��݋��*�y�쐔�$�لa�t�ĭ���ƌcF�X2m�L�f�qM[��;�4�HD'pME;T�jӝ��@ܹ��L4D��������HH�`�4ӹ$���eH���i��3�)��r�P�&:#\$tr\�.kr�a
�#�,D�)��W50bAk�����Ă���E��hl�H�ϓGӱ��d�>H�>�X��BŁ��Ԣ��7���9�M�y��L��4!��vfCuÏ濝�,Ja{�A*��zp��O�����
aT:��ڡ-��q������&��;�{�UD�'iK���J �P�Ӹ�	MB��(�Jj�ma��IT�uUt�X�Y��2�K�F$ C��"t>�� S �X�B��T0#B#4?���sy6~�p#p���H<6�F��0$�#$?;��~	q�����3sm��mq W\B1!\#C�����Q�HŁ�ed���I~!a!H�D̒�l��9�a��#aLi�0%7�ѥ.l�2n���.��֍s?y2��q�p������U�L o�!�a*I�׍]�(�2eP�P�H��"!�|@�0!2N�Q���i�$hi&}������}��9��Ą
H�i��I$		��� %0؁D�HRSh��$w��V���/W~e{�9%�jRr����J}u괝��T������L��4�$#��Xcm
�H��5�1�=�@�$���s��oZ։�Fe�l칧b&���[PҏȔL�T���R�v}��<	L5ǖLѵ�۩���dk�����]&�o�o��C���W	sI+�U!u���yMH��*E�
"A		T�&i����D��^e[X�(BD" #E,JL�&k�CSP�2�e0&g5��w��)T�^���e�b���t�
-q�p!L51!�h���T���U�k��F�$
ƍ�^$k�
��k �����ߵ2���R!\ �)��!��~&i4dj4�.~�Lփ��4e>����?2���G$Qk4��5I����� l�I��B@��@�B���!���v�Se��"�CYX�P�� ���4���-
m
�w����y���Ep�6��@��XGE�E
g�%LB���եexs��Y#1XF: �5��ߺ�:w��oa*F�jB�#L���T��0�Ԑ�l��a	@���! UB-<� ��h�Û$8�����IZ�)N�B���h�� \l��u�*�s���5���Hw�R,�P�1�)Y����G���?$�I�량e�� B���R�Y	� �H�d,���~�`)�l!LNh��o�q� �6�ߴR[d�f`Is0�W0@����]�5��\��(�����q�5`�6��bB�>0��qx���9�eO�6)!Ma�N�h���Gg�$�K���B0! �"�{���ݙا7O����l�m	$��*3^�6u���ۓ���e��6hJ3��!q�L&o��|?}�{�!HXP	���F�l��w�(dX�J�����vB�)��bF��e��4BY4K���xD�%�3P���$�/a"OǱ��%L�!MU�e�&�]���@D�<ՍaW�u���*};o�������D!	�KD!
h%*�J�i	K/r�BF�w!!6�0�\4�Bσe1IB�H�B�"�'�'^*��*$�� �]������1�����d! ��E�ZR&K�1i�	&��/xf!X]HV�	`E�0!I�mx�:��� �M��rB�l�/p� �I��B\%V3��դ
c���E#ni�����`d��F� ���8�R��°hr%�X4cSA�Jf�W0������P����5�6Ϻ\~�bP��ņ���C�i$i��0�sf�q�,5*nnd�LG�P+�I!1u��9�h�σ�+��ǒ��"R eW�r�ς	0R�1i!!!	ˣ�Ґ����!��Da"D�4����~�4��y�R0!FA�E����L.e���Y��4~�>�i�g߹�`�����F~����X@���%?~�@��m$c-'��}\4N6��d�@���^I3N����,p Q�H�1�4B� b�)
�d
@����ä5���ad5�bD�
 �n�a�Z6�q6�i�z��X�R��)�SI�L��ϭ��~��' �\��.m7u�����Ml�p���4;�,�J4�$'�M�7�V��*��`��jS!^鋥���e	S�%r�$c3D��l��iZ� &�	j�p�W^#ȝM�(ߴ�C��rF:K�.rV��p/�3|��~�8p��C��j����6�")y4bX��d	 �N�Z�Z��ӢƉ��%T�"@Q*,t�HX0��%	I�d!t]O�O��K;�$Ɯ%1�p�I�JS@9ej���H%�44KF$�|>���ljJbƉ��&�WY-�Y��*B$YB��jB�c! �.�@C�����;���Y�&�3W����'"�D�D!$%L� A���l��c�Ѻ���HEM;PJ"S@��ژ���"_���A^���ymJ^���T��E������@��;�W!B\��5d3�4�Lc5�g��Z���۵�*�&��S	L�\���a�~��%�<!p�
bJ�� F1ĕ���Dh`�@(�f�f��8CY�$��!$d�0 A�@�$j�1���Ԍ'�T�?|BJ`B1�#��K��d�n��-�h�a���!u	+ �A�F?�p�~�?���!"�P@��(���m��d   ��� -��m�     l�`�    m�  �     m�                                                             �� �             m��� p                  �a�       հ           �  �[�m                            �|      U��׵K,�N��2���V6��m[ 4��H�R��&Ī�ҭnٶ��[@|��o�i"��U���cm�;m�(.u,�
�i�q�ڙ0���YR轍+kj�*t ��v�]Ya��pk�52���6��lv�u��ʌ�[F�+ۯ�>�]��0wgX4Ѳì&�U�A��Y����	��z��qs=��%R��KvV�	VSRuR�t����QJKj��9�t�����[t�G�uU �� ��궀��f�����B�*ؠ�c-�2�usTl��Q��ꭕ��v˷*���U��v����}���۶�:�m��`8��VW�*�HMU��W+�EWA��[���fYUy@��6���m۷km���4�:�  z�����7�Mڂ��#֜�V���n(��}c|0q]nq-Kv8��R�X�'mC*=�yq;f+pr�Z�^kQF��-!1�M�N���Z��"�XÌ�j�U8:�vh�ll����ДN��66�mͰ��n�V�֒YCZ��BD���+��͠ږ�*m��Ywj�M����ٶ$u�8�4ur�jۛf����@*�@���pGj�a�Um@l V�*��D�ڨb��T
�r�i#n�q��M�[F<9Ғ�Ҽq�M��g��-��v�d�h ���u�����АJ6�[V�F����Ҫ��TC��j�H�kA���V�PpK�,i�y@z�@E��6I �[�E����P6ͮP&�pm�h�lͺM�.�l �fv8}7��;f��8pݤ�.�*���2��Pp�@Ti�v��pSWMv���@�n�*���T
�չ����#]��v �k���@8  I�k��`"���V�ܸ[m�m�Ž%�ؠ
��X%@jٲ�j�0�$��D.���f�j���V��d����}���!r�_�hWݞνQ�1z�oݲi1��ċiӥ��k�[m�|>��G � ��n�N���m���e:zv�FM�)`�
�^��Wj�lnBq�8Σif���7e��Yv�U˳s���r�*һM��ʛPBm�եt�'CA��YR����@�`
����Qm �W.�۰�E��v�8�v�b��-UR�E��ƀ���c��PⲎw��ge�
�k����5A�F�j��.�mU [,�̼Z�8�j�RZr�J��*��̗C��m!5z� �bc m��_^��j҇,T��R��$Ar��ko �&��[p	�G9���r�sb�H�l2�cZpl�n��KJm�f6�M���mYV"�v54�1��UUUU����3 J5T��gM��v�W�vR"�� ��m��һb�xu5�@UR��n�}�}SHt��޲j��JqmM�t�m����4����1� p�k���Vi���R��P$l �UW[���&0�W*��2�)�*�	D���Ɣ� 5�a�6 �����W4���J��g�5m���'�V¶�*	�=J��hUj��XN���&b[n�d�x5Kcb֍���pcWm�q�u��o�XO�&��ֶ�@`�řH�X�-��� ��\�I7h ��mG�+I�7�,��E����鶬l���>��j�cB�NN�i6n݁��''��$ӥ�"`���|�,M�ت�i`���qm6̓��ln7gYk5��N�
L��Qg����X1���R�M��p�+uK��U�S�Uj�j�[�4�� ٬a�U����ꪮ%*8*��6I�#P�ճ�L�,�c#��86ٴ�p�E��Ӭ�k�!!�#h���Kukי�Č�mٰgk����V@6�m� R��ƅiYZu��ضZ�9��mm� q l��]�jF��i�Zf�  e�e�*�5;<�u�*w\��	}J�l�*۵K�ݺG�4JT��T������[y5����m�٩l�n�KU�Q��}}��&"Wd)�յR�R��M�R�J[,����Z�)�E!�b֤�H+ee�gER�K]�t���p ZvλmrN�H[S��\-�8������[s��Z 
�s6ݲ�sc�J[l�puR���q�Iy �.� �u�����2�F��Yvh�wmP^�bM�鵲-�h��@(Sm��-U'b*��@6��֮�BC���>ļ�)��q��Z8����THv�u]Ut���+�'>�-j�WV���z�٩ɕI٪۩V�(.���f��m� ���:��UyN'��[V��$�� ��6U]��8*��)	��	��m5�����vn3��,���]a���m��נtr˲�F��sdSFԛ���P YsE����*�[\�:�t+0O;<�UM�yZ�U���79���Rt��	  �� �6ż5n�0^����� Z�[4^ͷv�6�(U�!L'l�xZ����m� ���2��W*lU*�
�mݲ��mm ���Ƴ\ �amq���_}ڜ�V�H�S�(��V���d06���r��WS�f�j�����	��	�y�i^k�''��(km����  �m��m����}��߷m��m�Ŵ ��8�I��M�����t�k�/6��n[l�jWT�,���'sn@�,�:�}}�|�?-
��M�݃m� � h:��n�kkc����\d$8h��`m�Z�:ާI�x��ug�B��c��WP�`&F��ev�ЂV�U��jv�h �]26� \�j�[:��0N�Ӂ&�2�լ�ܑ  �	6�	,��wh�*�6읹Z��`*�^3�Q����6f�J��A�,�֮�i	���4��� �/j�7��P��� �b�UT�TN�Zum �ꋵI�  ޝ.� m��$��M�u �hXg��aU�j�Z��� ܫE�sSj�ڶU����N�@&��t��;Z� p^�Kz�H�!*�j�>V�ޤ�O�|$ 6�p&��i�m����5-  �h�E�!��6[�_i�n��Q*�.���[S�긵\��	���L�m��x.VZ x���YP�l�D���m�8 �3v��  ���%�p��	Vک^��@ZL��i�UU��������T���J�q�2��Qj��ݳ�K#v`e:�t�fn�@�,u�P��`T��ᬎ�[�fݷ^E�ڵ���2���H�85�]6[[���^v�� �]��Iz���yX�!W�������mh��\��P�^"]k�n�[�F���.e ه-V�K�k�]/�#;�$Ք�wG��H؃l@�8��mU�hM$�I�滧gmy��k[%@j���8� *��ݷ�����3m�UUT�7C�Ug�ieo��\
�o�ٰ �`n�� ��
�ڶ�ge���gn�j�ڭW5��n�5�E0���HUUT�U��=�V��M�.� ��[�[K��V��Js��h
�r��[A��V�nXg�"M�h��v�[I	�l-� 6ͤ�l�`��l �l����pH m.����/6�(q��� 6�T$��ծ�[B@9�� 6�mZl�Wlm��L�6d
�f�Wevgݶhp�;]5E6    ���`��$۝M� �Np$���Id�}�Ϡ6�$ ݰ6���LȽM� ې
uH6�[A`�Z�U������U*��I{)l�6�6]6����6̮k3��Ď"i�m� !���  ���m�%���ĉ $$-�V�c\l�8  C�.����@ m��7^�6�����H�kh  I6��8�m[d�`  �kd����-� �$  Hv�l��׀ � �	Ƨl�p8r@h����� �8��&�
�]�Z�Ut�fU�Z�`r��,��m�����0
���V��j��%$��v�d������W�@^�7Y�V��t7n�u�w,�p�E�HKsH��M!6�U�UC����v�����5[wkrl$ � p  I}h��^ж�]���� 8  ���5J6���6�K�ܐp�� k�ᶶ�̫�^�givy�����I�Ӷ��a�G[�`ŶOh��m&8[U][&F��v���YS��j#
��UuJ��u��תM  luܝ7[+�DĹ�6Ze���Lt�U_�����{��UO(�UO�x #EC�ت ���� h�t�y*�����< CZ`�E0`!@S�B*�����`�N*��.�8�@8��AP�,]�Uv�1�@"��*|��b�
8<h��_�(� �H1 (u>CJ�mU5���¥U�%8�`��W� *� �="�� �7C�<��z"T؋�4��x &��("'@�?��E
�"�0@��� �N��@�
p���Cj�U�M*H ��� �(~F ��>P��l� �� ��D~��P*� �� `���X�|`@��j'PP���P�!�O�	��V�)��H*ƛ>b�Y 1@�D$C�pj�����`q "AX�b�ʫ�jhGI��q6 ����B,�`��b�TW�R$z@� �A�~D8(�T:(��w��� >���Q����V@�T
�*� �Z#�E*�XDQ¡F")Ȉ4 ��b�P�Ou�{���6o�-hl��($�6�           � ��   6�   l     l�lۯ9ۮ�8��n��cm�ɶ�ݕws�N(-tc.�ケ�ֵ�lB�Q�M�ΊEt�Yz�W�w ٮ1�Kdu$�,\u��oC�F�V;dT]���HX�bg��cu���@��39�m����nƵ��X��kl��68�\�ڳ��t����� k�K��ڸ�f%W�r, oi���� Qe�y-�=�I��L�q�m�5�V��[��i��[b}!eܙu͵Tр�W��rm�%'�>-vUp+����i��;x]]I��:]3�u�Ps���n۶ME<�e�,�c��֪�1˚�9����Z�N�Q��,����q��["��z:��-t,9r�mw-����V������ƥ@StȜ��P�k`�%�U1
ͥ���d���99�Hva�[Z������&���ر�����8����Vu\���7�q*�:�;/k�mݸ-c�5��� Snq6 
ᇶ�7"��ۯL��z��xC��T� �W�Ԑ��� 3��,�V�Ps[!����M�h�A��&�X�Yvm 2�҆E��k�N�;�e�88ZIA�m[�Ԏ1U�U�y�9��YBvz�f��TR��v�nqp�5��C�G5a�u՞Ӹ��j�S`;O*�����.�ɞP�srm���:V;]X}��<�S�;v­�מH���v��qmuͲn��Y9n���p\8�R��t�u�aij'��Q�N�{Me�JW���m�:4"Q��+�h;	�,��m]Y�̜���x^��[�hKV\�W2��EC/ZuAή�K�e��Ӷ��Z9P�<�b0s��N�RDʧaO&4k��F��Ť6ێ����b�	����uk]@5@vx�泉c	��Rއv�
�5���p�g/Pkc����Ǎ�H0����/��Wh*�
�D4(h!^�����r�k35�k@ ��lxi5����OV�k9\v�-."��P��h'V���Y&o.�Oo`�"� �q�k������+��+N�v�B����I-�t{�f���ƙcbѫ���v��D6��4a�i�,m�Β��uÑ����n�Mi|�f�����tp���t�Ż[1�Z*G8gN']u;���؆�s[�a&L��f����`Z��96�7gv�����4�Ř�<C1��~��!��)�{����ݟ��;�ZX��R��m�To1�@�v��33>V��~��YM��1�Ɓ�6�pR-����)�~���=]�@��$0�W���;�����S@�v����v�P��#��h�uwM�ӻ�`n����"";�n���.��8Oh�P8���rc�ᣔ���y#=��^y`�W�m0�d,u�R���- ��h�S@�K)��bCA@�Ly$�@/u��P��R@�R�B]�wn��_�ڴ^΢#Q(�M�F)&���eaf������y�6c��bd �bdMG��h�j�*�@�������ǹRH�<iGz������7�zl�|X(IB������7@��Weǎ\u,ث%��Gs^^���N�r�.�� WY^�B`�L��"��ߞ���Z���:��@��81�����7���Z�+�=�`gr�TD$��X�Ƶ#u.���T���?�z���$�*#��(̅E� B��Eģq�`�;�7>�;��>���;�M�:4��AAHh_U��f���Zz�h^�Hh(I�O$�h�Y�u}V�޲�W�h{�ZDD�2@`�o9u����^�ZN�vKwWg��{.���dxw]��=X�(�D�)RO�_��h�)�u}V�z��s�\fH�lL��Šw���(����v�ͫ�=�`s�M=ɉH�x�4���^�O��+�-���@��[�hm�ࣛ ��v�oM��ϋ�J9R������۰3e�ANLԪ$&A�Ǡu}V�޲�W�hW��6!$���n�6��jP9�t虥2�7�F��[�K��sq��;�-���WcU�;Nۓs�Q����/}>4���<�W�u}V��bx��ѥ�

C@�����z^������bCA@�Lxۏ@�^����@�YM��������J9yIH�>���h��/uz������ˌ����8����9{��?^��ܓ�ϻw$����������)Q���7UM��m��08u� �ݻ'MU�R������//`{F���p���[}�-!�6u�z�%�9JK��G2p�:�1-<UkB�tQ���tM�J��b2�5W+��<A]\�+�tx�G:9b�]�xV�����J"����<s��]�n'b�kٔe��n6���� h��6�k��Eu�V��k�b�ܼn���K����q��{�r��jCA�3.�+�q����#�^ɣZw`��&�˲�nӆS]��ѵy�dĤm<xȜ^��= ��4��Z��Z��*�hCm�rl��U�&�����`u�2l�H��[� ��Ɯ���h��h�נ�f�����U�(�jx܋@�]�@�ֽ ��4Wj�;�O�Y�(,�X9�˭z��h�ՠ~�ՠ}����ש�G�v�u<��Mƒ3�8��!)uui�m�y�褳�<�ni�p�Wdy)�m��ڰ>��v2s������́�W�
]S�t��'L�m���7�D$�1bv�b	U�#�V�֣K��=T�"`�}'�Ͽ]�?+�= ��4�>E�c�Ȣ�h�Š~���9[^�w����h�P�J�T���r�JuN�b"'���`��@��Z�������$��Ӊ8���h]�@�_U�r�^�z��IcX�@�K&,&�$Q��qWc��]�n�ex�v8G2��l�� ���=�#�@�v���h�נr������U�Q8����ڷ�H����*���Z��<Byf4���"���נr��'��30RJ!������y�otJt �A��H�Vנz�V�u�h�נr�Zdm�7o�����Z�٠r�^�����C����v��O�c��v�5��=�O*��������\�gQW��BGiل\�����u�h�נr���ڴꌸ��	���*eS�����z�f=ݛ�|���@�4�$� M��n=����ՠm�.��\�0�S�!����|����@;ﾚ��U�%	ZI%
���3Q�>
5�7"�[f��e���*�|�Wj�=yV�863�?�rb|�˲��eCN�gt�8Ǣ��f�u�S�u�p���XBCJI�w;V�˭z��h��@�;���A����}̛؆����wf��g1�~�L���r&�"iǠz�V��mzs�h�ՠ{�.3$r2'��Z����ՠw;V���Z�Tr$)$O�q��ՠw;n䟻��ܓ��{��qj) �^������Nm� �kX����.�{f��Ȋ�f�'E'�>�"�]_�˷���4:-�����ذ����p�#��n�^1ѵuXL��vx���/[׶�c��I7�Z\x�;&�K��m:�Ѫsys��BL��#���4uTm׵���x�: �r��'�~>��*�H칭��M�wWJlKԮ���\����K<)�Bhjubq��������{����y�;�h'B��q��0U=Xfzsl��0��ҧm[�ƪ�g@lZ׀��m8ۋ@����Zyڴ�j�?/#81�#�@�!z��h�j�;��@�^���vd�26F�G�ȴ�h�է��.__���?�Z��?䚣M���q��ՠy^�@�v���z�ݔPh�d�<�@�^��fw���*�zs�h��fE�	�fA�g��K� rEgWݳ�l�rv��uˉ�ZG!�pMƛQA����Z/Z��s��.0��ٰ:�`j����)�H�9�`u��7���LP�'&L�;��Z��h���İNH�'��;��@�}V���Z/Z�w�Iv%rD M��n-��Z��h�k�;��@��� uH�#	�@�v���zs�h���>Ϻ�~�2%���#كba�x�͵�!n�Ϸm]�����s֘�{-���!��<nE�
���Z�Jh�ՠ{��I�4ډ8!����[�g���G}gƁ�?�Z/Z�#�(�ѐM�T�)��3��`gWtي�lA�%0!A�F߃Z֥X�H�e̴#@�Lҟ8�~�8\۵��h���b2Q��$
�}�6�e`R^pYf+�|q�f���苠��MF��-tXj Z4�t� hҠ��h!�]~5�.��jho�B:b�9$�hL�1�C�3�v�4B)Y@�����?��K$��'>W�����Y@^���C���)P��"p᠔vbb'�ƃS�P6s�#C%�Y��L3�C=���`l�#m�A�4�� ���a���)�i��&���M9��I E�cA@ځ�&j�\z�1 ٭��֌`�����xw�i��V �7eIX�H�hU�?*��h'����4!�� '�u	@��A�	τ:�*t@ +E~ϯ}�@���@���mA7mE�4�s���d���;J"v�]��W.}��q�)�N-��zs��d���Nc�5DB���kn[���9���Wb;m͹��O�Q1��۞Qu֎��Z%n��O[^M��P��g����O��'���s�����6r%���"(�q������?�;���@�����տff$yr(`�r<��D��;���@��^���Z���ó%0q�"�7"�9zנw;V�?^��ܘE:@� ��X%N�D�ֻw$��p�/f\ˤ�ۏ@�v��yڴWj�<�����(�Ɖ����c�!�6鶬J\g����6ƹݺxy��s6����`�u�)��ȿ���=�ڴ/Z��j�<�:�PMƙ&F9&���Z.���j��٠wc]�#dN1(�Z.���j�*��@�v����@� ��6�#�@�v��Z�Wj�*�@�1.j�Q�M��Z^���ՠU�^��]�`bQ��J$�����m��m�B@ ���f��M���Ț�m�5#Qbv���7`��'U�����w,��1��vѱh5(�lvT3�n��"��:�1Dp@;���� �^��ƌ�/n7oiN�v���Tp�=r[�Uc��.�vhwe�d�X�s�$� �ZG����6�k�	�'km��.˔�$�s��6DԛxM�g����o=0�%�����������*�O�1*�Dl\�خk[iz���{Y�/<9��B�)���nR"Da�B`��}ϾZ]���ՠ������Lq6I�r-����j��f��ֽ���'f4ډ8!���v� ��h]k�*�@;���ȤCO"��f��ֽ���s�h]��n
8�$�ڒh]k�*�@�;V�_[4ܮT�&񤉶Н���<mnókk=8�����ܛ�;fpWQ˚cY$ȞLd�L�DМz]��vs�gٕ�B��ݛ��k	�a4�U)�:u`f�t����G�M0�vNoU�ӻ�BP���L����1�s534�{�VϹ�f�$��ߞ�����?/"�ar�rh]k�*�@�;V�_[4�òVE���I�Wuz�ڬ>̫��ɰ6"5mh鹑�h=8OhηK�L�b�a�z����h�9ݺ��Fr�N؀�'����q��"�������˭z]����E2)�ȴ�٠yu�@�����Z�g_���4�2&�z�Z�'o�w7Q "�b!"���A0�,O�С�3;۹'o�w7$�᮸�7�$��)�Wuz�ڴ
�k�<�נ~���nq��¦��������{�<�7f����ٷ�?/�Ԇ��F�{r��Y:/#��uxEZݮrt!џ[/I��J�!���-�S�d�mŠ��˭z]���j�?/"�dQ��`�94.��wW�{��@/���a��(5�<#�$z]���j��f��ֽ�w;1��F7E#�=�ՠN��u�'��{���)�$`���B
N
qT�ow7$��Y�[;]j̸�h�l�<�נr�@�;V�����������q�qtJ`�s�V�����)@g�oMvǲ�&����u1W7�lN4��$�}��=�uz�ڴ��h��Vd�ܑ�)�˺���Z��4.�������!9��z�ڴ��i���K���Uo�@��`�n�#��mŠ������:wz�>I(��}6N�u��K�% �����2l������;���>̫��BP@����A��h��C��}��u�$�`  � � ��m"�����5�c\;uʾ��m��qիry���{]2p��R��u��;7v����qulE��Y]���κN��nr�}�Q���^Ka�9��Ph�6�ڍ�b��h.�� �읧���mۏol���rܷu�/jzϋ�P�ms�ۆ�n��]���e��[q��gkȡNz6qv��ZM&�qk�sv[�N��&���{����@r\s��7%q���ܦu��-�ֻa��t%�׬�v0�-Y��v�H�n$�$~��{�k��f��ֽ�y��n4cqdR=��^����"#�)��{�`c�zl}�M�P�aݿ�x��H�������@��^��o^f́ܓvl�WrL��j\�EL����Q�P��o�6�����fM������wj��R�dTI5T�f�j�U6_{�`jP�r���ۻV˭z��H�F�!���o6��u�W�G:��0T�^ӁN�;��Q�����ލ�܉$�K�q��>���l�<���f~AU�=��U���M���nI9��[~�R4��,B-���ꉰ&���ܓ���nI��Z������0BNM��U�r�@��uz��4�òPj"Ha )�˺������������<����҉cqdR=���M����v�ݜ�`c�rla#ߟ��s��Iҧg�ڧ��0lqǇ�.��b�9�7g�������K�����(��G�����U�U�^�����N��T�t�h�:�m��ޛ�DD�w��{�~z޶h��\d$���Njìgo;�F�X�$���$$��Dd(����Vl�]�ϻ�J�I
8�<qɠ~�:� �����U��@���$��F�!7z޶h��� ��4�gW��B$rq��p%쉳>z���+�n8��Χ�r��v;"ʽ>�ص�Ftf�v5�eoM�go;�F�X�s�=��eX5$0��@=z�����z٠~��Q��VLm�7JI�~�:� �[4�3�;����4�\i��R"&$z޶h���rI��w[���dH5
i�REؔ��
���G����d��U�����.�M�������v���sk�}�3f�9ܳ@�C�&�O�'��&L�hYv�����ND���נD㛲\U��Z:A�89>��gI&&�qD����4�gW�~�j�BQ����;��x	V���)���n��Q�W�(��;�Ł�]���y���đ]"`�&�c�@����?y�Z}���~�����"�(��,�	H�>��]�����4�e�a���s}Vq�^h�L��HuN�9�r�BP��ܳޟ�Ǜ�9}�ܓ�l ~�h 0�@��0`s�6�VA(� ��h �#"�E�E�C+ �LF��22�*R� �1q�`�H�Q�:�`fGD2��a�Ӎ(��3��s*���~ 4) ����0X��������c"����lF���[ ��@�Lq5F@$*\2H�0��W8J�� 1 Cn�BI�X�ه�!���"jeޛ�a�j�i q`F~X1����.�!>��`BL?��0B�F1���+��t�f���Gđ����ZB08�A�x�����?�i�B��j�D��ͦ�Zt�*�`sm�m$             7m�@  �ٶ     [@ m       ��ˮ���Ԡ�Z�Lj�ۉ��ϳ�ؔ��D;p�;O%ی&�۳i��lVR��&.z�ip!�s:�r9�6m 0�ucx��Ŷ����ws���M���捑uc������<:���\�KR���k'��"���ȩ��V��}؜|11��DN�DΦ�OalT��a̭�Ͷ4�dL��f������OH[��l����S��(BG�Y4Fm�3�[��\ꃓF� �t�a�B�>�����v ��]�ܞՁ���s����;l܆�]V4=U�6�'0mup ���BQu*�[��o(�;<)�v�S�����mk��3SvX�.��9��-�躶Ʊ�T�<��:����䰜�x����Ûѹo8�țn԰lF����[n�l��۪��ك��]�x�ʸ�0]�y�8���<�k&���k3�]���#��w[���-�Rlm�Kks��-��vG%ɵ�\8�m�;mƭ���]�hLl�aؚ)�u�r��㙪��ny�@ѫX��A2\q5�.۵���a�1��v)���K��V�;<&Γ�	�2�j��;h݆�y���vtG:�a�:�2��Ϗ7c ꎮ�J]�N����q�qۋ������ݑ.�yxNsu�eݺj�g�ui'�� Xsn�	ۡ&�B-r�uX�i�M6�6c�#'�;:�{�Z�������q��Og.}e;��?o�6���`��5Q�n�f� )FN�:]*1*�.��.Rb��͎�gv�vvt+�6nU�#�f�bj�$6�q�X�l]7*���*���]!� �:����v�[5�J�A3��ۂ�d�L��#�����
��U ckS<w��N�N���0�n1�F�[(	d g�� ��:ͯ7@#�-[�����ݩ�(�؄zRP ���R���y�{�?(xx*~8à�F"#�"lPSG� �ALU�>��o���䍶  ��p�P	z��t��K��n������*��;���s�Վ�s��e\���-���5���ݍ��1��k&V2c�H�vtl��[��c�!�km��Ƿ u�0�[N��n�Y���m5��\g�J���dfl@���}�톈��-�a����W-��l]2�N�#	��QK��q��]��5�9�A��9�lmۃ���Ӯ�lo���{�w������;�������_a������s�T�v`X�W0�:tn{n�����|��j�����?�Ͽ�@��W�~^������~���	�ٟD�J&%M�ǝɿȄ��N��M�no����w'~��+�}�QA�c�N=˯�@;�r��B��(����:����R��9T6ښmӒ�ՇСB����͓6l<�M���C�k5�܃@�j�l���f�l}&d��IB�w6x�~�/uz���RY�h1'w"pHy�N5�g�m�Ll�i^^ڴd�S�ٝ�k�������*朂m���&��|��6��ʰ>fO�y$�}!ܓޛ�Y��Բ�)�2:n�37��D(N!BB�P�1�P��4 j������`w�f̀s�ʽ�	��c�.F��[� �죺��3�#���@�w�~���d��P��S3UV�v����6�?�&��Q
gپ� ���2/KuL� U:v}�������o|��s�`{6C��`u����g<{=	.��!��䍍g��,e�ː���;��ޗ��ֵ29�'�$�ߵ��I_u��$���S�DB�D/��y��m����S��%�T�T��m����5(���ܚz��m��zs����.K��̷�A�Z����)�R�j����M=sm������5�)�GY�������{���r�~>tHe�9eT�N���#�IEV{~��6�N���}��8��j��N^�M���M>D������$��"$��J���|�gv�um���^�m��ߚ����I�|�}�a��Bu�ѽ��#lZ �9�L�ǳ��w_v~���F�ڇURq��{Y��m��ю���>��a/��\�ۏRI{�P����j��'"�m��2��"f[�r��o�6��m�����ʛ���]߰WK��? ?�/Nq��}�Sm���k5���mM���z�*����$�����q��%�+}�m��[��6���eM���D%�M(�a(K�w��{��6�OٵMQRꨉ����$��:�ߒK���O���KϾ����^]w���&�Đ�(����t8�4gY��a4�k�띺�vV$kF�ʭ�EŻԪi�t�!����6w(�V�o����o���j��ɖ�v�_8�z�)��ܕLM�2�d�V�o����=ДB���^�[m���>q�ϲ�uz�L�{��޲��R�R�c��q��+m��o�Wq�aB��;�k�m�����o���]2����5L���Q3����6�ݣ][m�����6��^��o�O��&�P��I9��$z©�$������{��ݯ[-��}]��6��G;���ӻ��~k'��~  �I   �72����;-f6�目ڞ��;8�Ѷ�5�s�u�=+Bv6ij{���hږ�r[x���s<b7kn8��v#��n�2-v�]�b�����2ְ��2�p�t+�_���;��7^�a˔�`y�J�'�������9��ՉۧX�]:��4e�T�v� rG
� K������y�-�CҜmō}�ۊG��$���˖���y�����]=�ȅ��o����wn�jlMY��݅}�Q��Z/������?���e��m����<����z��f�m�����#�1�4���$���jI+��~��^�*ޤ�W�g��6ы��/���sU474�m�����6��T�f���e����6�em��m�"��449t�!���z�D�n���m����8�}�e��z���s�����ՑL[7%S��]�k3.�7m��߻�����?�S�$������$�dU�I%޻E$Hb-�l�&�W�b��6��xr�2��ɑ�x�i�j�yۿ{����ۯ���Vv�{!S�ͷ�[l��}����m����Τ�(\P?����?�ӿ���W�CF�-�~�ݼ�VC�:��5�^oZ���m���_8�}�e�����(�	*�o�+�ۏ�nZp��� ~�����+��ǩB�3�[l��{��|�m���\��YM�2�����m�$�S?m�q��+m��o�Wq�(�$�U�\盶�U����"E�8�hp���$���jI.��~I/\���!~����$�>w �읧k���-mƲub��ऌ=89琍�N��%��{��s�����pI�_�I^����Iz�Z�K��V��_}-���N�m��ODj��j��i��)��(�US}�o��m����m���w9��S2�dKͩ��je���3C��N��8�}��m��(��x�@�?����޼���'�$�N�)� ��~����{���m��]��-��ϻsv�*J!L�o5��Zȭ"]2j���f�;m��Wq󍷰�$����<m���l�%y�ũ$��h�M�D�X��-��.�V;�e��nu�f���v����0=���أ�M�ǎF'"��$�'�=I%����o;9i�$��L�����;8�ʗ&�:�S�&���m��w+��JL�ܝ�����]��L�&oСB�BJ�����&U5U5.e�D�j����׭��o>����JfuL���m��ͮq��f)*�S���K���[oa)���q����7m�����9m�*�xxw���e����=�449t�f�8�x�z��$��Y��Iy۬ԒWӪ��$�ٞ��~��HhqF SvE.��ۍ3��\>Ӻ���oi$��%s���y��~�F(�%#~I%�w����$���jI+��}���I\n�ޤ���J�b�dH�	��q���˒�̷����6�)�ٛm����s�Iy*�xי�*�&j�����-�߲�Ϝm����ͷ脼���7���%_���Ԓ_��1+M���br.q����6f�m��6y���s.Km��N���^wcL�����8ޤ���ry��Ԕv�y'm�k5��3ܙ�m�N�N����~~~�` �� WnDlkR�\:p{&h�c����+n��bEg���j�)�=ZpθV�ǻl���28�a���@�fj����Xs��c,�u�vj۹��%����ݭ��[�Aw��g�q��Jq�[�Q�Y�h2�q�E[�ߞ�|?t�6h�g;%�W9fi��0���Bu�e�&���Jq��.L�iҎ0���R7DW�(ۻ�SS"`��N�SML�y�k;n���7*�F�i�rn]KwE�"�޿ӻ�:i2�EUT�J�����oӾ�-��}]��6�T�rga%ɖ���_8�d>�$P�A��Bq��J�u_�}���q��Ͷ��k5���d�m�̊x#"hhME�M���Iv7սI%�Ϋ���co���$��~_�$�gLE{�G�X�TͶ�g���6�em��m���>q���������_��ͺ��S���Od*�q����e���v�_�6�T��Ͷ��ޯ��+B$�����7Ja!�Q������4v:���m��=]� ���V��s�=F7&BD܈Ԓ]��~��^��oRI~���=撶}�Ԓ^�/��7�Pǚ�K���-����o�?����[�P��j<�PH��TK���$"�H��q 嘚"@�U�% �@�e�"R�)�7̯�����V�-��}]��l.T?_�U~�!�f_�����s����[-�B�IUW�����x���m���T���$�c��$�t��M��Wq��y���z���w�����?�}�2E	$�6ӈԒWӪ��$�I(����6���k�o���[m�S��v���8�x��D���s�B�^O]��ɐ����)�`��{����Go���$�f��6�Sݵ6�o����o���z�(K���o�8�x���j�f�:k	&=I%�ޯ���Q�$�Ӫ��&�O2�ߢ"!/$�������sN�T���T󍷻^�[m��]��:Y
Ӂ��a�,XI�������æ��2#�b�'�$$��B�HBM1��0^$0���h?�<�}��МT�	��d�;	R$Q>(%_����~ ������	��������iy�7����/s["����2C3X\H@c�A�J�"�^�5�$��0N��f��0�*����N!�:)�qC��@��8�	𦪡� QS� U4�P��tE6����m����8�4b�c�t����ff���:��@�+k�:�����s@��FU��dr19����zS@�{�����興Y�2�h��{�β�<���rn1� ��h[ه �/R-�Y��]<���ʠ�hmYކ�o����h�w4����p��h����P�F1����[��u}V��õh�ՠ2�r&�M��h��vӘ�Ԕ(o{;���smXvV�LX&��&��?g��@�v�3zՇBP�%S�zl.��OZn���X��@�v��빠^v��}9���P�hSmKMT����A��9�6���v��^v�:�7az^��k�Ǧ��$�i��F��Ɯ_��nh��@��v��h�)�c�d#Mɚ�j�?e�M�h�t2�)��cn4��@���4�ՠw��h��@��m��B)2A�Ð��	�V�3�ZX��vv��u\�H1�,�@�t����DnV��-�����c�!GI��T?A�)J�(Q�_Ͽ>��  08x N�[ѦL��A/Id�Ӯ��e^�ڵ��M�������Y�y��l�݈Sg���9w4�cv4�6�ɋh��Ny�q���>zv�e)�P�G3��`�(���締Y�U�-Ƀvݹ��3)�Ƒ*����ʃ�?c��r�k�'\NI�����rHki�=�t/a��IqpM����2�H����¥{ON��o�{��������F���z���SІs�'��r�"b��oe֜��9ٶ[���a�8y�Tni����mHP/Ϫ�?e�M�h��=�ë��,I��	ȴץ�@��Z�)�^v���#���F/�$n(1F�r-���h���g�_W��@��}�|K�N8�4G�4�3�XX��v3���6=��ve�_L�����e��]�`}i�� ܝ�`gݬ,}�.���DD�+Ͳ�F�g�M���n��[Uf�v`=/L���{n.ݨ���Y���o����{9��ϻ��"Gwgu�ݣ[c�T��Ђ�,�҅
�R"�@��b�	���"Q	ѹ��`f��9�k �*EȲI�"��Z�]���Zj��(o�2��3���9��	*�j�өs2敇�P�)�ޔ�ei`}���Q	)���3`��}����*$�Z�t����Z�]��ڴ�H¤��x�5����`�1��u��k����&�.�&�[�'����}���w�M���Q�7�Z��@�빠~����B�0�L�,�aZ�\ӥ-9�&ꝁٽj���=ƾ,�ޛ�DD��_���Q���7&hs�-�:Y��r(AZҠ��^?(��!/��M�;���v^&eM̺�NE�~�JhϪ�/��h}�����~4��|�Q2Rc��rW�v�K{���3r��9�k>��X9�ʻ�Gm��)��n-v�M�cz�f�[K��,e՗!][�v�]*�68ḿٽj���Ł�5�����$���O��7|�z����:�L�4��V�D6}�V�l�>�Z�>�����ME�'!�~�Jh]�O�31=��7kK��'�%K�$���3E��DCͭ�`owmX̬,�	� I@�D(QSƾ,���UP�*i̡74��2Ձ�D(��Ӏum�Wj�=�)#HȌMd�@gˏ.�nE\�=z�!�=��9�= U��Kǳ���w�U�C�.��eT�׀�.�Ɓ�ڿ������?�҆6�SsE�ŝ�/b^IB��}>�77֬�V��	B��=�=T���ꤩ uE���y���j��ea`qgk �Z"�A$�i�b�-��31^��3v��8������6�]�F�m:���t�\̹�`w2��=
"#�5�^I;�������ܓ�P�W���ץ�??E�F�  h�����- �θ���ƓsVp��i7V�ε�M��v��єc���Nsm�;�0���I�Z5ۤs�NwgГ��-h���s+���v���9���VWq�=u��s�b;#!�F�U�"�悴�&�C�u���:�xmç]EŢ�bg���R�R�#�ݺ.��)]&\�9�y�ΓWbN`㋍�б���.�WBDn��9m֮I�c=��Z�l��l]nD��಍�3�v�qƘ�kFCU��EAV�q(��t�T�Q�}�}�z�V�{�4�)�~����u��rH�]��d�;�^Q
d��x�7}^,a���6w���T�%J�Ne	'��Y�wYM�:S@�v��w�M:sQTT��,6!�m�`}�V��9���%�f�Ł�g�����P��x'�:S@�v���4�)�������1L��vpm�sW'���f��o�n5�wn�*�ڮH��b��fA�H6`)���Z�h�V��\a�2��[�5S)�S*i���6ewM��kVDB�BQv=���?R�h�տ��߳�$rEK���vf֖�v���B��}��v�w]��`�hȔPܺj�f����zX��v}9��^fޖV�&?������p�=]�@�fg���~ߧƁ�t����H� ����粻�r��Arr�k���B��g�#.UJ���96����7�F�_YM޲�q��3��n���Kp�'��YM�bG�,��;���Jo���'�m�!���N�,��'���f��Т`��I�JU1-J"%%�ͫ,�V�>���s$PMS&D���<�ޖ�+K�Қ�t��{-r")$pX(��_�o�>9�X���?���������w&óQ`�jzg-�WF��<��f�T�����^~����6ԇ�;�>4��M�e4���=�WJ:)9S5.SsM�����<��7=^,f׋��a`qdu1�܍D�(���޲��Ji�%�Y�{�ύ��e��&dX�o�h��P����`wr��9�kD*C1P�LW]�o�rO��}!ĺrSp�u5L�3��`~P�_�BQ���>�3���!�:ndn�v�y��[�W����[�����ͧ���ώk��`x <�xțxC#���4��Kr�������(����Ł���U'2E�2d@��Nc�/$�L�ͯ{kŁ�;X_�M�V��E*uUD̔�uE������;XY�Q��V��ƀ[VI$QF�jCC���/K�2��;�VJ���`}�'�8�(�D��h�Қ�e4�|X���:#.(�ȄA����"X9�E*C�����NPM �b�5C5!Q"~`�	:@��"�0	 	�!��R�i����Rw���G�{���E~��#Pf�I� to��pM@��W�_e��K+���m�-��            �t� ͳl     � ��v�    �����Y=�U�#���R�1�$�y^;{=TNnog��:�����m;���N-��N����1��OmK�"��a�y۱��j�t�����օ7�V���P��M�`�q�#���Lb�iH4���j@�|�Z��bc�9Y:��W���v;<g	J�њ�8HI�%�-����d���g�k�.�na�ܷP<V1�A����l�G-Ƶ�ms�dGNq�,��;�$��ĝv�n�++Ӷ�u�uV�g)��VCIm e��gj��'K�4� �k�
6p%�ݶ���Rg�G�m(tn�u>�ܵnpa�9�&��봘���mrY^�苳����,�xH6!	�{{i�!]6�8����&�qpF���e�-cY1�iݗ�Y\�e(	��j#eq]�g�:1�)�m��C�՞;U��p-�����u[1��q��۠�V\����+C5�g�bx�n,Ke��u��l�$6�f�[`�p��]T�u��;e���s��tf��b�.m�j9�k�ܐh�ģ<�B;t��Ujn@w�m�r�t�p�Z+����f�X7	q����Ti�8�t��(ͶQ�E��E+0���Fʽb��7e�vV͹��1��i]]�R�a���z;K�7]mfӂq��Zr�0O8�6`ay��)�9\mL�[W.\m��Q=onNN��#&��q�+���;�ا��n6��v�B��1-^:�,�:�F.��[��8�fNAn S�ez��j��A�=��Pggt�cF�9�a|�Tpm[u�;0myS��-���[���[���ʵX:�GmR�n���j#,vvôxm�����N�Ľv6��m�wn��e���V\����v�a��TX=nկU̼�	J���������ؠ���F�s:.� 0(hS���)�ꮅ>E�|(u@���ࡊ�QҊ� Uz�e�/v�o� 	 �۷Z���k�]<��c�^����	�Ph�;g��e^ٌ�i�J�m�W�i�n�e�smn)�'�'l��#nc,��l<k;n�췳N�.^�ݭ�W�]^�p��(*:�n-1�r�
�+��v�z%��bp<��b�Z�����lr�g�B<���}hN]�_C�U5�q��L�ס[VnG��,9��u����ݩ�ѻ[y2��(m=��u��˚83�a���ä��\h��{�w���o���;�,��>�f�,�||�/Hg�?��K'��o�<m7�G&�}Қ�JXõ��w�ʿ%舙:�Ư.j�'�Di�h����t��w��f�,,�AUĵ@��S4��!?����;�ڰ3���!��zXwg��&��D6`) ����Jh���?S�4/uDq�fLp�ۀ��\�`g����V#M�[r�#�L����q9�Kz%T��ͩj�UT�tQ3U�ͯ�e4��M ����mXTI#n\�����3��节)B�IDBj5(��&��,36�����Cg݂u5�4�t鲪���>�+K ��ʳ�"{ܭ,�kK�Le)�ԩ��K�f�(M���`or��>��J^���[Q����6��#�@��Ł�DBߺ�<|s����`�ߛ@!g�a���/W=n�v7d�r6$(�m��=]�r:+q��=y�U\���+,�|X]�� ��D(^����`dm/�~T	���M2�����$�gwj���i`}�V�M�wkT�sD4Sr:Ke�n��;5�cJ�"�(؄��y�`v���jމm9m��c*���(S���X�?��k�@=�f�[V9$MF�jC@�s���D,������;�_)]���Id�2kY�0�u#%xayϣ�l�<���ڶ�C'@7��ם`�5Mk�k��37��ٯ��G�3~lc��I�S-:�D���ʽ��g�gƁ���?S�4�E6,m�G�\����ϻXX��z�$�g�6�X���5�����EC��.f�$�ۗ����ZX~�U��B�%q
I�1�ux������gŁ���D첥�*��C�,�k��77��ٯ�ݯ��D.��K�l����!8L��d�����.���B�㶕����c=6��{n�;�_}�^��Ѥ-��}�����=���;�,ط�[U)�m�ܲ[vf�/�舉����`{׋ ��ʰ�ƌc�۩�u5U-��_b�şD(����}�|h��W�̂QD�#��;�,3y�����(��߯������7�q�kdx��Y�vs���s������GB�;5<0�� !��!ғ�ιӺ�qOm=���1]�g;c֍$:Ɯ�=6[Oli�O3�1�'*u8�ݷ���@�e�Ui{r��;Y6�=�;^WuC��a��qc��n�g���o)f胤ӝʎ�q�c\�@ٷm���=Oq��p�nW���M�r�D7:M�uu��&YҤt����؆�n;\�N㮮�<u4U4'C�t�Ӓ�uD,_DBIy��4'�cv1ɹ��G�f�bӳ�1�Ş����r�:���k�+����߀���X�|Xڟ�/�(�Y@no���Y^�T�P�)K�����X_�!������6�����!(����g�_R�T1:n��2�߹?� ��vlD�up��s���V�&H�U UC�DD)���`}��M���Ł����n�h�2�:)�)�`nV��BI,����gܟŀno;;��nj���\'bw`pC坕�L]�;y����l���f�p�"@ER!
���??���c��V߻��y$��C���`bȗ��Pɗ UKl�3u>/�BiD	%p�"a�y����=����D%�$�N�k�3�5*e�RT���37�`~�)�~�)�{�%4�Ufō2�f� �v���;���3~n�ŀfo;Ҳ9r�I�SJF��e���Ł���`���������-՗;����F]�#��F�8�:����sa�άZ�ݸzL�-+��On�ŀfo;�ϋ�ϋٯ�R��)�2�,3y�Т!B�3�o��������S!���6T����ܲ[vw����k�̅	 �#O�!t����ܒ}���@?��T�RH�J&ڐ�?^��=�����o>,Y<��2�Cm�e����`��������k�@�iT��б
@��lLwn�.��[�N�k%�ѷ7XSإA��ŭx�,S�,Q�ㆀw���YM��M��)�wr�6&�P��o �M�Y��(l�r��;��K ��ʽl����q@��"`������=ݒ���4�e4g�/�#l�7#�8X�����o>,%D(�	C��U��q`f��T����nGD̦� ��v���_n�Łٲ�k= t���ݷg��oItlsncu�l۴is�Ō�κj!:뤵���m
��`{y�`{��`f�|X���)RQI#MF�jC@�zS@�vJX��79�Dɫb���P�2�C�9��>4��i�bW�����@���n<mb��4��h�+����TBO����31�WL��&4��$�@�YM��MײY�$�����Z�F @"�����=����I�;���!�  �p�z��^ź�c6���486��cFΠ�m�U�֗Nri����v�G�L]l�<n-�droZ�l݆���sY,�se�H`�N�Rp#'<Q��넸Y7LX�'P��<���Yݡ6� '����gu�ţL�+n}@��XB�Tu��goX^2]"�u���Rl��%�h=I�b۷'%P&�v��ɩ$�(P����Ȝ�jS�2U����p'F��n�Ɏ��g6�@��Y���\���$ib��n�����d��w���e4g�/�T�������4^U��D6�ڰ3�ZX��>��3���0r"1%���4���?]|Xڟ�[�-�&�*��۰79�`{9�`v*� ��v��Q�4�i��4޲��;V�{�f�{�4��*J�ك�Y��ٷ'n� �٭ǅ�g�ȩ�M��K�
�ޗ�QN���r!�-���U�6����)�~���?_��(�[�Y���ܒ~��u���(B Ċ�#�J W�ɛ�7$��uٰ/�ڴw*�bnM�I�gk���s���U�6�����m�eK���e���Ł���l3l�=zS@�y��j�&����'qWt�B��'w�~~��`{9�`j��Z�ӗ-���E���H�(�5qnW�m��~�=}�Y�v����9��n^\�r"02H�o��z���������gƀ{����G"l�AI4�_����ŀfo; �[�=#n�t���T�X�|X�_tB9�:���0�A5R�> 46pb!H'�wf�D>���.ȉ�FL�C��,��F:��$
��$6U&0#�L��2���!�^��X��i
��x	�X�4*f�5��d0�����hM���)��� �[�򣸲(�<�1\؃�ء��q?��@�Ma8C�V�J�vTV�� v ��c8
=�!߀�O�C�v(D�ȪtQ��G�0���%�
w�`gs��őS��!�.D�m�$������7{�`vk���YM���B��N<mdn,n�u��D}�7��`v-|X��n��1���M��u;yzx�8�𙛭rt�=] �	��wl�� ���U�ٯ��ϋ�k��37���Y�`S��m:�R�h�9�V���z������/�S@�y��u���9&��/��4��4��?z�h�n�<i��6) �����ٹ'?w]����`$H��K"�
�Q�(��gm4�e�$�H6H����Jh�e4��M ��� �RC�8�Ӹ�a�����R���F.�B۞B;sh(ڡ�;/�X�Q5B����ϋqk��37����1dT�.3"J2
I$4�Δ�{��9���ϲ��P�g{�铣�S-T˕T� ����(����X��Ɓ��SchjM�I�~��g>,b�ŇТ&w{�`d��6�2���e��=���?$�j�����krN~ϻw$�y���P.1� �� �B��^]{Z��f` �� %���i=�[L�x+�l=vʎ��mt�X�6��g�u۩��g7��m�6*F�"C�k��[gOA��u���yݮ6U	�ۓ����=�<�vb�wiʫ�K;s9ovӦ��$	n�
�l�&i���h�s)�np�<k��jю{r��6g�:����Ì���#`���ʀf�a;1C��]��5������W[�g%�('l�A��G�N�m̲ih�ܽ���;�=�5��0=������fퟫ�����0�s�Xf�=��6����A�m��6) �����c�9�V>]�/��D�wW�:�m��ʡ�d�������|Y�$��j����׊b��rH�Mš�No��`f����eoM��=��dIFAG�Hh��)�}���O�{��h�e4���A��2<��nu꣎�۲�=sϳ�yu�xx�;u�z�<�r����T��%�U2�37���ׅ�ϲ���Օ����m����R���m��|[W
D(�I,"!R� � ���U~@�-����\����`zVƮ*]6�����h�e4�t���H�M�Y�{á�R`��NG�8h�Q	�V^���Ձ��aa���ޖq~�m��0�(��!��Y��DF}���3~��Ł���:uB���6M�������r�߯�)�����[N.Pu�Z<�t�å�5ԩG�I�ܭ,}���ߗk��{�V��}7$���R�YM��)��Y�~��߱#������Fۂ�B��\�,3y��Ij�!B�I*�[4�=�S@���`)���Q`�1�h|�u�h�ߖ���S@�gJh�E���M�I�~���?z�X�v����U��	��Sn[L(��u�nxeh��ˮ�l�qѱd�O[��Y��L������t�eN]�����o���t��{�f����@��C�k ��p�;�Қ�u��Қ�YM�:�6�́!��{����k���s���Z��j�%��9R()&�������S@�gK7'W��~_$�!U��⅔bH�\A��P�#@�E "
�U*"pH#9����x�ϜPrIi��4޲���ŀfo;ݯ��K�K�CsT��ԡ� ��5����>v<luۮ�]���2�$��i�1�	�I�^�>43y��||�!/Hf��,�9�>I�Q`�1�h��h�Jh�e4�t���䎵fb�p�_��`g�zXf�=+#T��mb��4޲�{�M ����v�Ȩί"I���<I�@�h����`vWt��|XBM(D(�PLJ��U�6������m��! �����֒8���ۺ%4V:�iۇ+�Up���A��]���mr�n��:��[g!���}�2sh�؝��'WT�D������fI�"C��'k��n2z1����M�:-��[���n�[m�v"���*��kM��a�tu&k�E�+�!��Hæ<s�9v\#�зN�g�\�b�`��M���-��AԤ�DBW	E�$��U
�)�s���Z�2Z��1Y�%�ݴ��z苶3��4�"cfB)��4�j�?z�h�Jh��T���Q�A�4�j�?z�h�Jh��o�� ������$�F�qŠ{��f�� ��vg>,ȩ�tP��ˡ��UE���f��`��3�h�e4��Zȓj,�4��4�)�~���/����i�9�n���ɹ����"k���� 3G9���5�[n8����������\����>ߟŁ��Ł۩�`������S�S�*UP���e�����$�$��	%�.;��w��`g�XX�U�ȓn�p�/vJh�ܫ<�7������ZX}�e����TS�lUE��Q��f��g�ŁϲS@��S@?vZ�Ɉj8�nrK>����K�.���=�W� ��ʰ=��ho
�3B�4����0底M�`y���͸�!�yT���usv�!����rIi��?����/���z٠_YM�����7��4�+�Ca��Ձ������,w!�%��6��H1�@=z��ڴ���ٮ�` @���Ab�
�iDj���Y�~�&䛿Z�3uu�n��ƪf�-�ТB{��vwkK>閬��U�ƾ�����%��R�杁߲��5BQ�٧�_ g��`gӘ���]:&I#yѺїdC=l��y���y�Z��F�:s�Ͱ��`�N}��{jz-�Oo�ߟ���V����B^����X�'��\�qE:���4��*��f�kK����Ϻe���a�qiT�2]M9��(���7�ZX}���Q���`�}4�ҙ\PrIi��4z�,�]j�3;��(�B�PЄ)� $L(���Rʐ
I�ʀ`y���ܓ�gu/�Ժ˙�'��/v]� ������=�.�m���i��3���k�e�\;�;n��:<���͹��\s�J�*�6-b���lD{KRmXgs�;9�`fs��K�uϷ4� ���DcI�NI�_[����Ł۫�Xv�)�%lr�}�&�6dƜ��^�|h�.�z������j�,yl�I#Ĝ4ݗs@=z�����1^�~4ꏵ7��!�H�%�f�z������>,�]j����t�I�!D�|0�?H���ґ�Hk12D��C�M�	
n �bB	B3&5S_j�f+�"�aP�M�t�$%ںK�(�1��1�"����GZ!#D3}
'�ă�c������Ͽa�(���"�!���I�iFF����'�ظ��~�;�2+W\e�A���ᒡ�Y��?���]R�08�r�$�U�EN1��7��C��$�Q��+m�M1ʙm�9�h-��            �@  �n�     5�  �l      ��6��([�j�ơ���۴6���^:����
���Ӳ�N-t���9%5ɻq�]���8�{���[ �^�� `Q���=dv�ˮɯwGb7�@�vmh��Zٸ���nܙ�(�\�`4�-=8r)�v-v,����5�I���t�v��+�`����B'����T��x6x5,�'���Y-�n���2�ٮ��"i:�s;n�Q�ca�a�.Ch��bg��+�s=��gH-��6�tDn��k�9ZN��Grsx�q��:4����d���*[��8[��`���8�l+��S9���8�rC�[ny�8g6��<=��!<B�A�7]Z�l��b1H�w*&NXѺ6�ܻ���.sk�i�lK�<�NCs��g�A�>BUҺv�ŰS�����s��u��G:ˣE����������]l�lq.]ìy*��nt� �[��2툀�x�3�a��:��(�s$N���p"�ͨ�6����{\�L��Cr]��p��/Y �,�v��!��$�ln�:��Ym��s!&:,��A =*Hf�g:N�(�s��g j��t:�l��.C���][[q�6�V���}��T{qk.x����n՛;�Y:$R\�:*�Z`Me�Gr�����p�tul���8�۷�ر��@J�ybٱ��J��u��@�<=�c�������F�-��n�9=]��k�ɋc'N�U]�=���q���1�\c]p11�6`J�79�n�೻� �pc0P��Y�MuK{gj��P+��[����j����=+��;�BL�iH�k�MKѤ(������uWl������h���w�,��j��HFC$���T����<�D��gȳ��֝5�&��Y��׈�u�,�������qm]�u�2͓5o,4kZ5l$�.f�|��T#��qG�/ ���"�z���Ax��z~�"8��BP�DDZ��rT�m��m��m��:m�&�qm�j����'�L�1Hq�+�Oi����jꍜ&뭫O ��iܘ-�����c����uXp�{w.݇Uɫ:6��0�Gܚ�.�FpSu ⳻n)`y����K�Xz��Ms���n�P}'O�l���ud���z�BS�s��[��.��ݞۚ5·1�h��J�4r��q�'n�:�]jjߕQ��I7�ur�ur�@�V�;tẍ�v������A�{FG��,g�����@��nNN�n�߲��3�Yk�_H�z�=�5�]S��Em�3@�˹�Uֽ��������pQ����Hh�.�WZ��w4�S@��	@U9��d��T�=	7�ݫ{�j���)�^컚���vdp�Ͷ�$��/���=�S@��w4�l�:��Pg���e�}���JvNM�]�F��1��9�楬z��{V�n��9w\�+7�n��`�����~�Ձ�/X��Ss"���SsE����V�%�����	BPHf�;��Ձ�ϋ��]M���BD�,s4�l�/���=�S@��w4���8$H�R&I&��۹�{�����w4�l���e��)i����e4�]j�3{����j��"S��R�fY����7^v7>k�th�程�bmRى�w#�#M��N��Ay�"��6߿��mX�̫>̵��;�ZX�bc�����l�䙠�f�}n��˹�{�u!�?�m<IɲN��vnI���sL �B))b���8�)��~�w4�[4�=�ˎ&�6dƜ����$��zX��՞L��O��W�,K�=���iȖ%�bw���ڕM̊���M��&Bd&B�ż[ND�,K��{[ND�,K�{�6��bX�'���6��bX�'�z�~~�&����-�A���#��Nw%�.�b�;��t���vU_��o�7�����l���iȖ%�b_��kiȖ%�b{�{�ӑ,K���ߦ��~��,��^�^�\!2!2�o�.�b*�n]j�ֵ��"X�%���NC�A9"X�����ӑ,K�����ND�,K�}�fӐ[ı+������j��.\Ҹ\!2!2��ٴ�Kı=ޞ��Kı?g��m9ı,O���m9ı,O�z��ʗ3CtL�p�Bd&Bd,�[�iȖ%�b~ϻ��r%�bX���p�r%�`tO�#Dx���7���6��bX�'O�[wI|\�32k0֍�"X�%��>�iȖ%�b~���iȖ%�b~����r%�bX��V�\.�	��7oJ�lT�H��.6\�͏l�t�sٍq��ֺ�����k��&f��8zM�r=�Y�����{��"~���iȖ%�b~����r%�bX��Opؼ�bX�'���ͧ"X�%���	g���)�3Z6��bX�'﻿M�!��"dK����iȖ%�b}���m9ı,O���m9�  DȖ'{����Ys!��kX[��ND�,K����iȖ%�b~ϻ��r%����>�����Kı>��6��bX�'�z�r�\�]jkV�i�6��bX�'���ͧ"X�%�����"X�%�����iȖ%���AȞ����ӑ,KĿw���)��U3.����p��L��_n���Kİ�A#�}���ı,O{���"X�%��>�iȖ%�bww��??_�D�l �)�`8u(�*���ft�$�F��L��vH��,[�r�I�Em�R�T:�D���.{+��ݡ���9�)�:4\�f�Ѷѳmmˑ 퓇���7;,]�+?�}���V!�5��S��"t�����A��t�ҹ6Ս4�4r$J���̽aĽ��S�jKm�D�)��ms8{p[�ѵ��X*�Ҳ�h�u��K�	"�ն�攩���
ffA�;l�a��؍ԝ���۞qm�ՊS];��z=RQS55M�nf�B�!2!{r��Ȗ%�bw�=�iȖ%�b~ϻ�ڼ�bX�'���m9ı,O�{���c�.�虢�p��L��[���ӑ,K���wٴ�Kı=���iȖ%�b~����O���,O�ͻ����c3&�h�r%�bX�g}��ND�,K�{�6��bؖ'��ND�,K�v{�ӑ,K���5�]TL�.Q5357�&Bd&B����"X�%�����ӑ,K��ݞ��Kű?g��m9ı,O�}�[�.��L�h˚Ѵ�Kı?}�p�r%�bX����6��bX�'���ͧ"X�%���ND�,K!yD%�x�f[t��7T"�j�T��Ad,l��*�����n�;�=�-��v�5��`M��NfERꪓuK��!2!2�Oq\.D�,K�}�fӑ,K�����"X�%�����ӑ,K�����\��њ�Y%��iȖ%�b~ϻ��r�l )'P�j�h��'�'}���r%�bX���p�r%�bX����6��bX�%���I�H*���uL�U7�&Bd&B�wx�"X�%�����ӑ,��ݞ��Kı?g��m9ı,J���=�SY��jܶ�h�r%�bX���m9ı,N���ND�,K�}�fӑ,K���{�ӑ,K���]�ؚlr���T�L��L���x�9ı,A��wٴ�Kı?{���Kı?}�p�r%�bX�3�����Gc6[t�m�ד/a��u{9vL=a����[/Hg��K��Gb�e��Fӑ,K���wٴ�Kı?{���Kı?}�p�r%�bX����6��bX�'�Hk�˖�N�̘L�fk6��bX�'�{�6���bX�'��ND�,K�v{�ӑ,K���wٴ�Kı?a�����S)���M�"X�%�����ӑ,K��}=�iȖ0��C��!�)P+�q��5U��?�bfk�ͧ"X�%��w~�ND�,K����M��[(��M�+��!1(@'���m9ı,O��}�ND�,K���6��bX�'��ND�	��1��L̲JUU,M\.�
ı?g��m9ı,O{���r%�bX���m9ı,Ow���r%�oq������i�q��ٟ�ᛜ�g��﮾)�Iȷ]���rṙڬ�&���www_W�D�UML˪d���_�	�����m9ı,O�w�6��bX�'���m9ı,O��}�ND�,K��h�i����s-˪.L��L��sxm9DB�$Ot����H'��}�BE$N���7�,K�w	�5m����mִm9ı,Ot����Kı?g}��r%�bX����Kı>�}�iȖ%�by�wI|\�2橚�ӑ,K?�9�{��6��bX�'����6��bX�'��m9İ>U=C�!�����iȖ%�b~�C^�\�Zu���ff�iȖ%�b{�ߦӑ,K�����"X�%����"X�%��=�f�p��L��^��t=�ܶ��'s��//Qzu�����=�L5��g��a6y��<Uf�j[�.��Lɩ�f���Kı=�p�r%�bX���p�r%��L���l�^Q|B�!2����p��L��[��0�����SM��p�ı,Ot��m9ı,O���6��bX�'���m9ı,N��p�r
�%�b}�g��n�M�e�4m9ı,O���6��bX�'���m9ı,O{���Kı=���\!2!2��A4K��̕L�ֳiȖ%�b{�ߦӑ,K����ND�,K�=�ND�,�6w6nL��L��q-�j�jj�˹u���Kı=���ӑ,K��O{�ӑ,K��{�ͧ"X�%�ϻ�+�����$,߾�J����m��4R@ �λ��-*�#�9aj��T����4�wbֲ{���<%�������m�.ѓu5�ڷ���Ul��<�g�S���)v�G/���#�2#�{7<�
٬`�F�1�p3����p����n�	[�`,m�ny�b�ظr�:�g����˃λ#���*�YvB:7m���{�����`ֺmW\ɢ�-�ɭ!4�!Dٛ�5��Pq�Σ��8x��1�'8/U�ɻs�^vy�]&.���:��k�f�+]�=���2X�'�=��iȖ%�b{=�fӑ,K�������B ~��,K����6��bX�'���t����fd�3Z6��bX�'���m9ı,O��m9ı,O{���Kı;��p�r%�bX�zMOz�Y�:����Y��Kı?{���Kı;���iȖ(�%�ߎ��ӑ,K���l�.�	�����j�D���@�f�m9ı,N��p�r%�bX���m9ı,O���m9ı,Wۛ�p�Bd&Bd,�fA&�s#�UN��h�r%�bX���m9ı,?���{�6��X�%�����m9ı,N��p�r%�bX���Ӛ�L�d�cu��ώu� �����-��D����q���#���<��6�7}��oq�ı>�wٴ�Kı?{���Kı;���iȖ%�bw���JB���{��N�P麡��\/�%�b~�}�i�_(17H$���R#�P��?!�� H��b{|��"X�%����ӑ,K���ߦӑ?�*dKǵ��u4���+��!2!o���m9ı,N�w�6��c�C"dN�o�m9ı,O����iȖ%!2v2�=RPɚ��sT�L��-�߻=�iȖ%�b}�o�iȖ%�b~���iȖ%�bw���"X�%�����|e�2��ɭND�,K�{~�ND�,K���ND�,K���m9ı,N���ND�!2�3B�jF�	ۥHmJ��#�K�����'pՋ�Y��!�"Kv����}���,֝a�asR�ӑ,K���{�ӑ,K��}�ND�,K�v{�ӑ,K���ߦӑ,K���=/��L�K��2�m9ı,N����Kı=�g�m9ı,O���m9ı,O}�p�rX�%�ߵfA&��I�UM7SJ�p��L��[�7�ӑ,K���ߦӑ,b��!|�LW��|�.��q	'�lBF)$�	�C���5�uL$�$B�*Y��3f��P��
D�޴6�&�<��U(�>�C�C�TJ ��	�<D>UC��G���7߽�ND�,K���m9ı,O��=y�啪
��&���	��	���z\.�K���{�ӑ,K��}�ND�,@,N���ND�,K���ª$����C�T\.�	�����\�bX�'{�p�r%�bX����6�!2!2woK��!2!{7�����`I֓���+��q�1���[q�謄�"��7W7h������b�1����%�bX�����"X�%�߻=�iȖ%�b}�o�a�T?DȦBd.���\!2!2�V�yIC����KnkFӑ,K��ݞ��Kı>����Kı?{���Kı;�{�ӑ,K���Yf�2�rj�֍�"X�%����M�"X�%�����"X
%����6��bX�'~���"X�%�ޓW��eUEJ�2��担�!3�JH]����Kı=���ND�,K�v{�ӑ,K ��@�q/������!2!}&-	�Ii�&j��"X�%����6��bX��$Q=�O����Kı;�����Kı?{���Kı=��sX[HL��ND�<��^8��Ϙ9�0v�ۜt絛b��lP/>�dϳ��u0M�{���ou�bw��p�r%�bX�{���r%�bX���p�r%�bX���iȖ)��pZ�G)�hQT��W�'ı>����?��&DȖ'����6��bX�'����iȖ%�bw��p�r%�bX����0�k5��uu���r%�bX���p�r%�bX���iȖ?��ș�����K�L�����\!2!2[��mSEM=j��Lִm9ı��}�ND�,K�v{�ӑ,K���ߦӑ,K���{�ӑ,K��λ�xɩ�����KsZ�r%�bX����6��HL��興#=�x�_�	�����iȖ%�b^���ӑ,K��;U>	���#�Qj�7Ow{��{�ױ����� 	  	 ��9n���gR]=�p�1&��8<��	���چ�uPqN�u�Z�����l����N3���w�����a��h=V��]���M�N�8��-b�2�s�ۗ;��zv�E�w��Y���:.�=�u(��)4�+��~��:�Na;6�GJx��m�=r\��ɖ�t�,�ǽ{���=�i��O������n���;x�n���j��n�=�F�nū��T�җS���K!p��L��Y�_��"X�%�ｿM�"X�%���޻9ı,O}��ND�,K�&����LuL3��56��bX�'���6��bX�'{�z�9ı,O}��ND�,K�{~�ND�,K(���&�1ʖ�*i������$.�^��r%�bX����6��`�b}�o�iȖ%�b_}�kiȖ%�HYҲ%��̒��SM�S�\!2?!$%$/f��\.�	��=��p�BbX�%������bX�'{�z�9�L��Y�ۙnX=e7T��W�+ı>����Kİ��{[ND�,K�׽v��bX�'����L��L��u����,�IH庌�p����k�����Fu�˶��ya@� G�4Jj�54�fi���&Bd&B{�ڴ�Kı;�{�iȖ%�b{��p�
��"X�'���6��bX�Bk�G��(�55NI�.��L��N'{�z�9�)HdD�~� �Mı=��p�r%�bX����m9ı,K��m9ı,N��yg����53Y-�5v��bX�'����"X�%����M�"X�"ș�=�\!2!2�{��p��L��Z���/���\��5�iȖ%�ʬQ2'���6��bX�%����[ND�,K�׽v��bX�'~;�ND�,K�$׭��LuL3���ND�,K���[ND�,K�k޻ND�,K���"X�%����ND�&Bd.�K��Sd�qTL�JT�4^�yy�>���*vG�l�9����R��o������o���T�Ԏ\ֶ��bX�'~׽v��bX�'�;�ND�,K�w�6ȳ�L�bX�����ӑ,K�����yT�r��SM�S�\!2!2�f��r¬r&D�;���ND�,K�w���r%�bX��^��r'�Er*HL��/\�r�~e7T�	�+���bX�����"X�%�}�kiȖ<_�L�8��5�?���]�"X�%��p�r%�bX����a�f�W33W5�ͧ"X�02&w���ӑ,K��u��v��bX�'���ӑ,K��=�fӑ,K���dɫ��j��Y�m9ı,N��z�9ı,��g�m9ı,O���m9ı,K������bX�%�{�zۨOvz.c�6�����9=!t�#�v��"4�hE�K"uϙ��tCjp{���D�,O�v{�ӑ,K��=�fӑ,KĿ��kiȖ%�bw�{�iȖ%�b~~�L�Yu��5rkFӑ,K��=�fӐ�R�L�b_���m9ı,Ow_��iȖ%�b~���6����2%��3_�g����0����m9ı,K�����"X�%�ߵ�]�"X�%����p�r%�bX�f����	��	����[sNU4��kiȖ%��'~׽v��bX�'�=�iȖ%�b}��iȖ%��8�p�<�A���K�o�m9ı,O}5�)뫖���Y�sZ�ND�,K�ݞ��Kİ�H�_��ͧ�%�b_���m9ı,N��z�9ı,OǴI�K��e�-�Ѭ�g�eG7H=�lE�suo�����c�ۧ��ʹ�������|h(6Ʈ���7���x�;���ͧ"X�%�w��ӑ,K�����ӑ,K���g�m9ĳ�oq���ߨ���`Z*�����7��b_�ﵴ�Kı;����Kı?}��ND�,K��}�ND�)	��+u�N�ꦜ�H���\!2�bw�{�iȖ%�b~���6��c�(�r&D�{�6��bX�%����ӑ,K��C]�<d5u�&a2���r%�bX�����"X�%��{�ͧ"X�%�w��ӑ,K���~�\!2!2c7�rpn���䧓Z6��bX�'���6��bX��s�{�[O�,K��u��v��bX�'�=�iȖ%�b~h��'�Ќ� �uVd������Ԇ�   8u�X0���Z kG��ɻV�U̓��ʑٗU���q�]�jMl�H;m�(x�i1���h�kS�T�۳����lg��Fݭ��}��;](c ��:��N�]ӝz�h�k��9P66b�Y�A�N�;T&����8i�_m4�aœ5d��m�GNaM����G	
�4Bl�Ð�$��F��m��s:m=Pg��ч����R�9�ι2!۪��ڗ��<��ŷN�,(];�Fl&I�c=�Rz<���ɭgS�,KĿ���m9ı,N��z�9ı,O�v{���P��dFBd,�o��p��L��O��Ayˢ�R�R�Z�r%�bX��^��r�	"dK��p�r%�bX���fӑ,KĿ��kiȖ%�bw�]v�2ښt�i��w�&Bd&B��o�"X�%��{�ͧ"X�%�w��ӑ,K�����ӑ,K���w2��]6U6*���	��	��;�fӑ,KĿ��kiȖ%�bw�{�iȖ%�X�����"X�%�s5l�R�SSM�UUSp�Bd&Bd'������bX�'~׽v��bX�'�=�iȖ%�b}��iȖ%�b���~���ny��q��B�/<h���s�l7Dr��}�Z�k3������8��]�3D�k[ND�,K�k޻ND�,K�ݞ��Kı>�wٰ9ı,K������bX�'z�I�!�fh�	��ӑ,K���g�m9���"X�{��ӑ,KĿw��ӑ,K�����ӑ?�S*dK����u.�%9*���	��	����m9ı,K������`�%�ߵ�]�"X�%��g���Kı;�C^��j���榳[ND�,�`dL��\!2!2�{��p��L��]���m9İ?�dN�{��ӑ,K�OW�yˢ�4���L��N'~׽v��bX�'ݞߦӑ,K����6��bX�%������bX���
fX{�2��KBniSD�Ssi{X"ݹ���b�unwD[�]ū��t=���;�K�4努�����/�L��L��z�Zr%�bX�{��ӑ,KĿ{��ÈA�I�{�M�$ޝ��nY/�6U6&UQj(A��T+!i	��K���m9ı,N��z�9ı,O�=�M�"ؖ%�{�_S
j�չ�jff���bX�%������bX�'~׽v��c�O��:"Q�"�X�q�xH��w���m9ı,O���6��bX�'p�ajjj�Z�ɚ&�Z�r%�bX��^��r%�bX�v{~�ND�,K��}�ND�,�B�3�����r%�bX��i��"�SHr"[�w�&Bd&B�~�ND�,K�=����i�%�bX������r%�bX��^��r%�bX������!�`uRv`F���p\<��b�"�^\��b��5	�:��w�I>�K356��bX�'���6��bX�%������bX�'~׽v��bX�'ݞߦӑ,K��Iz�a���	�˭fӑ,KĿ{��ӑı,N��z�9ı,O�=�M�"X���]�͛���!<^�N���h��p��L��[��;�� �,O��~�ND�,K��}�ND�,K��{[ND�,K����ԷY0ֵ�Zչ�]�"X�b|w���r%�bX�{]��r%�bX�����r%�` ��p�u������ӑ,K����2����M�M�꨸\!2 �>����Kı/�����Kı;����Kı>;��m9ĳ�ow��?x�.�oIm��{�v�`p��]����Ͷ���p���mp��(�x�:�[�kS5�]�"X�%�~ｭ�"X�%�ߵ�]�"X�%���o�a��C�L�bX���fӑ,K�����>��7U4�EMU��	��	�����D�,K�ߦӑ,K����ӑ,KĿw��ӑ,K��CW��:�C��Ӹ\!2!2Vm��Kı>����K�,K�}�m9ı,N��z�9ı,O���0t�L"s4\.�	���Y�iȖ%�b_��kiȖ%�bw�{�iȖ%�b|w���r%�bX��!�[�5\̙p�����r%�bX�����r%�bX��^��r%�bX���6��bX�'��}v��bX�'I��><�D���$!SP2 Q*�	&�b#��CS�t1 ��A�; �b�Qp�GH��""�O��iR�I�veR)��(Qv�?1�H�C��M�����8l�BAB�O��@���jX�`CG�J(s ��
�Í^�� DJ�M�L��$��J�U�$�����~�2ۑ,���h��            -�  6Ͱ    Z� �v�      !��^��?�����b \OX�s�f瞮��/�ŵg��GG[��Y%�.2�Qd��Me�EU]�m��Ȣ����W&�F�d�x��c=j��[`���j��x�A��.+b��婠b�6%��I�Zu�m�`[�m<L�����lqQd��m��.��=��m2#-�.��X�7�7���	�A�]�͆^M�t�؄��['Fuż��{=��������v+K��ݩ��cwV�s��g�}�x�F猥�5��O#��6����M>Y΍�1)e�"p���uJfVx�Wmڮ5��y�呩 BT����t�789!��N�`|0��n:��[��͇��t;���K�bղ�	�9�]0)�e�tb;$.��֦py���΅R��n�,Z�7\�91�Eζ�`�<q)�_>��j�dl�&�;�j��c���J�n{tS�l8^�{i$m�˱�s�y'�m����e[8�eM�+��WQ�WB���=s�G/�ܺ.�C��q�
��	����\NA��V��s�%�v��՗ t:A@zV{3�)A�#=[5����gH�6��%N�6��"Vx{np��"8�% �6xx0��QOh���%�_�i���D�ee,���^1��#���Vt68��5����s�k����Q�8�f�g ��厊�8��Ϯ�4Z����ySYgu�l���s5�j�9���2�0���tV\�U���(ܩ��"Eٔ�P���P ���RհdDq�S5���d
B���\����u:�]��v�Ru�W%�#tp����j��EiI4dĹ#��`)V1��^]3���À]N�U��ɞ�m��u�<co;qћb�m�h�Eۀb�=�-�ڀ�KX���l^��%Jk�wp�A:���s;�tK7Ee&�.�_�~|
�
�����U("8���|���`|(���u��  h��:���h�|6 �����^�6��dgcZ�n%g����o��_R��ɓ`3�� ������Kl�.%Շ0m2h�nLpmĎ�m{'Y'�;I��wkY]�nqr���q����ݹ<�N�oI\eNlpWe'�K	�\���t�#V�sv9�]�qv�%1�4��$���\��ie@��âb�7
�������:�h���z���;����ݝ�ݗ��ӎ�mv8Ny�3���X�o�۟�k��۱V��,K������ӑ,K������r%�bX�{]��r%�bX��{�p�Bd&Bd,²5��˕SRUSsUv��bX�'ݞߦӑ,K����ӑ,KĿ{��ӑ,K��������B�!{�na�M?2��lVkZ�ND�,K�����r%�bX��{��r%��C"dOw_��iȖ%��Y�����	��	��f�IN��T��\.kWiȖ%�b_��kiȖ%�bw�{�iȖ%�b}���m9İlO����9ı,N����h�Z�\��k5��"X�%�{����"X�%��g���Kı>����Kı/�����Kı?�=�kVf4�x�!�x�n��.�W'*��k��v{u;3��:����e.˻r5�����K������r%�bX�{]��r%�bX��{��r%�bX��{��r%�bX����^�]��l���r%�bX�{]��r�P� ^4��Ȗ%��m9ı,K�w��r%�bX�v{~�ND�@*d��[�y�M	�.BhuN�p��N%�{�����"X�%�{����"X�%��g���Kı>����K��	�26'f������L��ؗ�{��r%�bX�v{~�ND�,K�k��ND�,�FdL������!2!2�[���ʩ�*�\�U��Kı>;��m9ı,O����9ı,K�}�m9ı,K�����!2!2�ǧ*h��M2���m.�zLr:kX������z��8�`3p�g]�չ�d[p��ճZ�7Z��r%�bX�w]��r%�bX�����r%�bX��}�l?�!�&D�,N�����r%�bY	�OxR�P)*i�r��;��!2�~ｭ�!���,K������Kı;�����Kı>���K!I
H]K~G�rܒ�sE4:n�x�1,K�ｭ�"X�%��g���K�q��Е�B�(�%SD������v��bX�%��}��"R����s;�U,nZ*�"����İlO�=�M�"X�%��u�]�"X�%�~����"X�%�w��ӑ,K���}��4K��a�-���ND�,K�뾻ND�,K��{[ND�,K�ｭ�"X�%��g���Kı/{;�5mr�F�u�ep����� ��k�ձ�c�Q�wI�"K��-}��ۙ��K�\�����	��	��wv�9ı,K������bX�'ݞߦӑ,K����ӑ,KĿI�bvJ��nh��p��L��O�ݫND�,K�ߦӑ,K����ӑ,KĿw��ӑ,K��f��j�.UMIUR檮L��L��6�m9ı,O����9ı,K���m9ı,K߽�m9ı,O{��Ip���SZ��Z��r%�g�RB�^��.�	��	��\!2 �/~����K��3"}�~����%T�RT�t�9�v����f��,��������-� (9�Xز��9�h��4n��'c@�.���usp։9w/G��*]������@�S@�}V�z�4fs:�j)�fӓ@�S��- ��h�h���Lj<i�7E��g���̫5$���ݫ�mi`^�R���4��H��٠�٠{:�h��hE�����J@�I4�[4gYM��� �Z�I���{~�6���l ��> < .�n��%V�kف�[{�V�^;Xk�Uآ�V�8�y[�3��t�	�c<���4(�#Q[�����ő�-%*]�!��FN��.������6S�����{[u�{��nٻ��ڒ �t���k��V������m���b���Wɞ��yg�ڞ]�`���ط1�u���j`����ټ5�i<�-Q	4�{�yҙ���44**y��{	��cٓ�Dy�l��n�s����l�_ndo#��4���ύ��� �[4�[4y(�<x��������g��Д6�ڰ�v��r����nk֥T�RT�t�9�v�ݫ �[4gYM�����ʿ��	��M��s�1o>,�ޛ�%��nՁԞ,�2�tD!�U��S@�>�@;�������Is������c���k��+��es��<����]��--d݋]xy��lY��m���hu�@;���l�����z�1SEM2[� ��v�P�D$�n��˵�`{9�`l���r��R�h��h�e4�?��}>4߾�����"m��1�Ӓh�e4޲��l�{��-�@+�Iˡ���MQ`s�,���y������=��h�V�D�4Ly0?������cI�n���ƹݺxLІ*gdz6�Ǒ�c#�D��4�٠�֬�r��Iq�����ֵn�:�532�R��ټ�[ϋٯ� Ͷh1vu��P0�94gYM�s�����ȡ ��~��9g~��@>���;��q�� �N<I�m���k��7{��{7�����`v�:+"�7��w[4�����S@���;��RD�!H6��S�yy�X������9,�cn͓��h��R��P��Y	�MǠ��h��0�9�kP��>}͛�N@����UN�[��݁���=���=9�V��4�(s&&��A)!�{�)�zsz����,�ŀv���:�әsI�e��(����3~��Y��JP��!)IG�����oC�R�F�Ȥz����{�4{�4?��`j��rekn)�3��!�i����J4��,y%��N�}q�3�-0�,��ܝ\#%�	��o�b�f�,NoV�~��@����Aǉ5��h���=9�V��v�k���2}���"��D�yu���[4���=��<��q�ŒG�@M6��=������35�a�ZQ����m��6�M�4�,�����2���=�����J1%�}s��� �����u���&v�Bs�_Z��l�[K��-��ul������g�#�N���u�۳pJB\�Ӈ��=3�� �]�!���&%y.Y[k�ƹ��k�:vy��cl�ϵ��[㫞���v��fy�7���� ��/5������q�Q�n9֡����.k�+�ef9���sJ[*��Ş\�%'4�4O���K�٪#TDZ�A�� P'�t�u�t��Y���u�ݛ�3�0gv��Dl%t�4�L���p�Ec��|w�|h�h�l�?x���Z0��$���h�h�[4�,���t��ʆu2(�Ƣ��6��=������35�`{+�l���.�N�Ȅ9���J�+u��|h�h�l�=��š��ĚB�h���z٠��@��ڴ�봑�dM�c���0æC�k�&3��ձm�9�$��rf�<��`0�i���cc��~ � o��~��,{����:���)l&j[V���[�; �0�D"�Hq��Z��M���@���Tm�	�m�4�U�{�)�~�h�[4ԏ�Lm")��-��M���@?z٠~��4���djHD�9�ڴ�����)�~�Jh��ZD�'���h,u�q�e�ٶ�O-����q컛��2]�>�Sպ%GmD�����4ה����)�_;V�ً��҄�f)&���|X�|X�� �o;:7�)� �N<I�ӆ���)�~�է��b_�%0 D�HHL�!!�K����?=�B0!)%-��"^;�|ρ������Oٌ6Z����ɉ�'BGP�H���$ҍ�Dk(B���B�,�	��bCI�0��Y�����H�A(@O���Đ9��m��D�"`��BBA�!��h�M��&ڬ�F��q��
�l��X���D����Y�dG���@�X`��5H�묨��"��8p�L��^�ъ��/��5��C�?�M�H���S?�@�H13�@�ۄA���R%��C,�!ن���h��lH�LNj֒�sf��bD�%����k����ڢ��� ���� �Gf��� �_��UV��!	�t4l z��L(��	d����=�<�Ċꞡ��X�Ƥn�v� ��@��R��$������dj��
��U��s`��`{6_�_����ܭ�?5�����h�����ӷ=�T��v�wB[mw��0�[N�>y�T��USv�e�`{5�`nWt��BP� {��@��G��?��E �5!�~�Jh�j�{��?z�M �r��a��"'��h�j�{��?^R��YM˳���QƛQDE�����l�,g>,-B�(�!( V�h�\#A�B	$���@��H��0��	Ga+��m���1KtU:	���@�yJh�e4�j�{��߽߼�?{R6N�r�a�=lr#�{&�iݕ����C�v뗚Mv�^�^^x�X!ǉ4�p����_;V�{�g�ٙ���{�Ɓ{05�8,kԍ�@ϧ1ިI%�{�Vێ��9�V���5��s�R�*����`�l�?^R��YM�v��w��TI��R$ܚ��)�~���?Wj��@�xBciH,mHh������7w����|XDB=�߭�??$H�` 9Mké@%�8D늍���U�nF􈦍r��ީWmg �=[r�O�dۛ-�rf��m�Cq�)���؄m��KKm�;k(Q�z.=e�Vэ�9��>q�=���ͦḹ,��fu�::���@MW�T�6�����
F�S�II*�4+�p��t�65�Kv��]�u'b��wJ.��0��s�nF��cۃ��*VR�q�ǿ�wr%�e�mƴ�+�DM��/`�K����|��Ԓ7n����K�.��M�$�<���U�y������@�ܥ4��h]�DG��@�Z��4�*Z�Қ�j�;1wP�����U���cv3�����N���{���ŸA(�x�i�������yڴ��h�T��`�����Ғ8h��@;�f�{�K@�zS@;�P�,k,��d�LIvcn
7��4v5���nv�t��k�¼��2[�pE����ѨM����h�)M��M�ڴq��Q&�jH����9߮�7�'�(QKA�0��%un�����7w���ä	ى6��6�4��h��hwY�~�R��Uq���D��O#��?Wj��@�ܥ4��h]��#��Dڊ,�@;���r��9�XX��v�S����L����{K�Í���z�Ns��9��m����\�길�OR�HLiB!����Z�Ɓ}e4�ڴ���=��ŹQ8�&�4�_t���v� ��4�U��w��\pCI���hf�SQIBR�Q1���ڰ;y�`d�UrN]�SNl�y��V�{�4Wj�:��1�mƠT�������j�����Ӏwgu��l�;ܩ����9�,q�'��zLr;>��!!q��\�m�a`5q]C��Ds�p�v�`�h�Ajf��YM��h�נw�[����Ȇ����4I��h�נw�[����?/e�#��D�$ȴ]k�;֭���h�V����\iB!�I���6��|X��6�H���t��H�/D�s9�ܓaw�$��dS4[)�Z�Z.�6}��X	>�ۉiҔ�c�	��9�AP�2��:XN5n�w[	�l���Ҍ�lm'���|���V}��lq��֖3�I3�20i8�m��/�[��ՠ\��{�DCgq�-�n��2:�`ow]�2s����7wmX�#M�")���ՠZ�Z��h֭� �mcdC_�HƞI"�-v��w4�Jh�V����R��߀ 4R@ ����]]�m,��^��F��v�����y�.^L���&���֜c��V9�Zpn*ݷn6۞�Ϙ�ɾ7�pXn�aN{R�k6i9��l^�څ|�m:J�&��*��i):3������ľN[�S��z��Հ�:����f���b���݁�H-]�����.@z˲��^���&%���u�:nʹ��{���}ލI�BQ���*�ԩe.��B��N�6ڸt厯�&m�G+� \]\݆tI�C�pqțD�E�=��s@����k�h��@��|�4��F6`�4�Jh�V�k�m��=��ŹN8�&b#��k�h�U��-��V�mi`s)�y%6I2L�4)�y�Z��h�e4]�@������a&8�IŠ[e4Բ��ՠ^}V���fǉ��ɑ�1��p�6.A�u*r��[.�zs�mv+�g����0Y�!�D��lN�YM�j�/>�@��h�l�iD�%2[,���K�m$�%vu�\��S@�K)��O��""y$�@����)�~�e4]�@���Dj%��I��h�M�[)�Z�Zs�����Y$cfG�[)�Z�Zs�m��?ZG�$��O	���7>�wSs�(�����<�me��S�k&�Z���@3/3p�-v�����w4��S@�p1�Uā����Z��Z��h����k�h����!�Lӛ��Ձ����J<���B��$��W\���6j5&�U1)#���~β��ՠ{�U�w[��wR<�P�h�_�Hh����{���r��8�+b75���!95��.vN�[zJz�F˚���wn�j`��rdxy�K�C�E�]�h�S@���h�ՠU��"5�D�$�ȴ�)�${���w�y�Zfs�q�,�1�ㆁ��S@�v����)�}��)N�6榦SR2���P��������I���f��4��`E�E�P�H`(X�H��GW���ܓ���f���m8)�y�Zu��?R�h�ՠ~�J)"Mb2&�sƱ<��k���\s�kۃ���ݜ�盩r��w=�k��#��9�@qh�S@�K)�z��TDq�������*�S�D��YM�ڴϪ�;����_��y�� �4����/>�@�YM �S& �XD�I�y�Zu��?R�h�ՠr�u�G"m`�Zu��&��M��:P}ٰ<�%
""#�(W�� EU��@EU�*������ "��� "���(���
�V(��"�(���@",�"� ����B(�",�"�H�,UH",UV� "*A", ",Ub���"��, �"�B� b��� ��X�,F�b��T ��P ���"�B� b
�U�"�",P�"�X",T ��B(��*B(�`��X",U�*�(���,`�� 
��, ��H���"�"
�� �H�,�"Ȃ� �� �H� ������������� "��@EU�*�W��U_�U�@EU��W�DU_�"��@U�1AY&SYH�2��Y�hP��3'� ax� ��4 (     P � �@P���B�@��   >�T���
�)���H}��F��$�H@��k5$ H PE}h���Q ` (��J�		v�    �u�@A�t�<v����@}�{�)�G��( =��JQG͔�x�|O��|{��w��w�y�p��l�W�  �(���y�=��B�8t��**�k�R�bR���
[<t3g�w2�̓�;j��  |� }�]�� 5�s�u�iU;o�kͨ�����l*���[}�ͯ�G6�m]�U}��W U��[���}y�p >��
�6�W�� }�U�\��j���Z�6R�]:�]��w����}��W�f�!�e\��Ҹ��� ��j�P��iy`=^�Twg��{[Wf�Z�3�ޚ��ld�@͎���|���:ncJ�{�����}zÀ v<�97X}��}�[7y����s��j�5W�@-�7ū́�v�< ��� J eA��]�����ћ}鎆����Q�:�yB'�;����������-�6|�;����{������ ���z=�Bv���s���>��bN����� ��=���݀l-���{�z�:��s���r����nPR������)@�����)@͔���j����;����R���  F�3J �����ӭ�)J[�(�)���R�Q�((q���n�t�7w���P �Ҕ)��  S�6Ԥ�@4Ǫ�EOʚ D�*�*ڨhF�Oi���TP  5O�j�Om)R�  "(&)IDb�&�qO���?�g���.g����T�m�R�Nr\���� "�����\*����h�����_���TU7���俿���d1��2_lap��%�+��VH�FX�VRIXY%��*��.o_fSg�7���!�?m��LÙ����c `�e6R���&C���!��s&G�>ֱ��b����(CA��0B�ˢ@�X�EĒd����a����°Ô B���M:Ȅ	5ns�dB�t5���Ji7#
ICNS,� A���	
ƙaL1$BH�c��%2wB�2�p�ecu!.3P�C.�6��$2c�a��$ME?��q��B>�ⓅPf)p�IH5.	�.��MKn6�O/��<�k4&���&e�aL`��8R"@��HY`C�SzԐ!h��pGp��o�G�� �!	\�i���������N�V�����ӽ,�#D�8��$`B�jˣss{�$0`A�~!!�\�sQ��σ.vSZӁtЅ��A�ܻ�����!	14:��k��xnaL�B:H�2�L(��2ˌ�!�L`�))BB1!!)*p�Z�5�LW�N�thT%�)&%%r�a
|�,	
�q���$���Ia���Y� Cz>�e�Nf�1�I�_�&�˼��l(B���$�ػfa%H��	�0"�"D���3p�å�nL�jk�\���BѨC\d�3��,�:��!����*J�`o�%�iF�����_��F���Ўp���gn�cW�����.�0^3����%��7�c�ԋ�H��rhbT��B&7�h>��� X������Đ�I�i�^�;�%>c{ă�B:l���aR혟��&2�������d̸g�1�댗��J`���M�HuϦ3#�3)p�Hᅐ�F1aH��CA�i�\��LĤHJa�S J`�!dea����D�\K��y�`�hR#B�F���N.�x0��H��q��!�s���z?%�f�(a�����ki��F����$#	��Sd(�����pkd���[0��XЖ#�bIH��H�	
���p�FB�cL�4M�lԆ�Sd
�#��A��R�����'���{����S��&��ٹ�����H��P�V@��
��!p���B����(bV`��>(F�+�ԅaR,ak��{�
#07�o�Fm�w��-f1�oa	RQ"A���%̹e3���]kC��&>�\i�-��#�7?F��B&����4�J��@#�U�]g�3��8������K�feك)�A�˖��1�J21�`�;�C�60 D�Cg�����ĎB$VVX�$XH���H%�[�����$�F��$�A#��!1��d�����.F"��(� R6&0��4�Yq���B�\�@�"Ptw�z7>�rP�LC5i��>ld�!V%�
8`S	
 ˩>�'c�B��%1
��%�1
ʅ#��2@ � EIN���&�`�b%pD��;�3�P�δ��1Ѷ5R5�P�A����X��B�eSϜR$R Q�cHk7B`�U���Қcp[�'T�\M��:!f!R���N���/�Zδ��m4L�K&fd�0q>6�@�	i�	
D�(J���"@9!��0B�y	Č$#W9��:M�%є�D���0�FB$��aP�M��H8r��#�܋1��V�� S�O�!�I$d�_��ð�!33����ހ�f����
�K#�DJ�V)B4��ٻ���:���C��7���a
a#\dJ!�oN��VK��&H�JCVS�D�Z@�̘�넟_��n�J�J`�n&i'�̗�p0�|W;yHh~l.L�c�O�����Zr��� ���c�|�������gR�4wL�/
t�a��>�9��2�!E�	2�`��� �0�c@�eT�l�,�fD�IdJ���q
���� m�Ӊ�+@�C��5	D1bB�B=��@����Q�1���u�@�4A)+�$.N��L���d)LMI�%�i��)D��ZA%��tla\	erH`(B9HЅ R'��8J,bB�$BaH�Y�Eб���Bp%�~��4�9	!p�ɣ%�1��c��y�D�k��I�4ؙ3gg�P �8��a]#�a�ۮ���d�F	l��7����&^;�K`�ذ�-ލ0�η��q��詶H�;yrf?G��{����ON�?3��;�˼�M�G��Mɧr3ǚ����������R����������2$HB�K��$�k���Ą���*Hhb�"Ha�������y3����$��#&*JoX�E�"���������0k_gHܴ5�~#L!�HP���2`�t�`��2�H�Ru]b/B̻��F0k(B�$�#�d�p���9���E��e���d��!��/�d�ٸ�H�n2F.a��\gi[	��>�C��1�>���w� ��xH}�bs�`]M�q����+�Z�)��F%�aL���pJ�y�\Hٌ�y�;�3�\:�1�mؑ
LoD��4���-pHg.�o���#����.��H� $p���Mo!	��]��5�Jd�3�Is��_qouY�5�	&��N��	�t �JB��ą2B�����:�l��4|�j��`����v�
��1jA��Pß�}�&2���lM�aXq���i��8ow���Б�I�����D�����8��ы)p`ɱ�2ė�f�l��2�K!��\j�4��[>��`�	##T�-�Ա12�1�A*B�6�u�ɨY��d,Yͻ���#�Ѷk�%�J`�I�b�HF6�1$A��i��o3z��R,~���|D��� #FJ�J���t�d��5s,nIro�5�3Q������q���9��k5� X@�����
�G$i'L}.pn}��
`�`���-��R%,T�T+�Ӌu^�؂r�`����X�d�cB D3	$dK!.{7a21��Bˊ<f�J�H20��i�$
�����:�0+!<�����!Xg":��Cu�p�,�@)�r����2$���)��:� .��11L�v��.�M�Q��d!>�!Iq�zkf���M���gF�M2�t7.'QtR��$R}L��x��q�(@���!
@*@�Hx����+P8.�嬄�0�9��yޗZ�I�6H�*BM�����hGԻ��_KQX�P�!�$2aX)
`̚�����,�����HX��d�(B����\�!&��.X��n��R�C\��q��a*b1�"PzLfg'��2@��F
��RWK��A��~����4}ܔ����saYpgS!H,H��'~V�~�i���_pr+��S�k���3��!������d���j��a)w��
���`�F2ńd)�#�q���Mƫ~����w��Ao�4�B�
8B|����9���d�0�3#d1�8�>b�Q��%	��3���#���u0O�/���ZJ�ɦ�˧$�H�II1�Lc��	ԅrB�(Hg�(te`R%��R,HX\\��'��[�0�c.c��m����"T�R V+����X��\��s������Yߦ�R��*�Z�I�����c�kyO��M�0����Y>a�1��<���q
�(|٘Ёc]������7�C;�٬19�!0t�H�d1݆7�e�3�js5��I��X�"D(Ƅ)�b8�edC+R�1�����j��P� �8�5\�9[ԡ�h��Ma�.�i�"@��g����>P�̸����!�Y�w�B|�Yfq��4Hj�i�
jB�@��R�\����$��T��p̌��\$��e�.n����H�N��&��]�2�#�V1��
a��6�$p��)�^͛a�L��2❎2G8� \2�	�ã��i�rN�\�Z��!pM7%ɝٍ�f�		�)(�5�����p'Ί�?�W�L�﫯��ڮ;�{�wǌ�����U;^�D�T���,��}���=?��}>��              �� �               -��                                         ��  �`              �|                  �      	�8            h    k    h$  �n��� hk6`��u���`� ��o3���m�(m��lꫥP��fwe�6n�7c���v�s�N�$�g�y�
�`6U�����s� �E�l�i6 7m�R�TK\n�{MKu�j�"�ץ1�"M��klwN�aU�Uj���+iyUz�sI��D�م�M�`
��[T�Q����jBj��Mtf`x��K.�� �u���n�lIA�g�e0�s��%K0a7c��	�ƹѸ��Z@ܰ-e�-+r�T�+q�eU�'��?/�UT���Z����Y��熯 �����ĂI [a�[Amm��r�@[Dk����V�[���KW�6٭f�� �` ��[ ��]�ݗ;�RY]�bRU����gj�8 p�f�[2��$�J�UU[G/��m����Uڀ�����v�@�v��I:HK/ �i l pR���m;t��"A�X�݀[Cl�LH�Lo[R��C�fR��n��v��E�Ud�[@6��%[+*���V�eZ=��]�6pe�0�sWF��0�P�`Y�
��^y55@WUU ��[�	KY�v 2I��	�ɵą�fݰ��D�j۲$�b��tkd��$�̍��ij�I��T��j�ٹ�'̍�$m� H�km��G/IZCZzI,� u�����V��j�1�)ɍUԫW��LP��
�����ڦ�'�^��;l`�2���:�Y<^N����W�Sy�M#[Sx��Ճ�C�9�bM�#Z��d�&�4sZH JZ�]]]Ep��j�$DM�/[!��gF��I��[�S��V1YKT���3��[V���%�Ւb
�m��l��[���iX	�ldY6煷jٶ�x� h6[��EH�� 2������)6�5\����]�"�M�-Qz�c��y8q�*pm]���Qh÷QZB� ���2��{j [SFڎ��i�@ kM���m}'K��-� 9m��\.*U���V�<�6�ڶ������k�ܘp�k�$Y6 �ְ��� n˳n���m��si9�m��zCE^�� $�v�$�mR����hkZ��!4�4��:ɳ%��W�@�$���ll��Y��,�m�`X�#
��Ҕ �VV"e�}W�7nJU�m�;eU�0CD��F&��[U&Ic(e@j����A�[�n�*�t8��UK�����a��ʹ�$�M*�Wn6v�4��j�i��¬#<��i��O:2�+U%lQ@
���Hm�Z1�Acm�n2r��b�m�r;U۴�@m�TK��ʫU�s T��K5����kz��j��2Td�m�U�M�ݒ����m �k��n���p	��-���O������	����d�V�	]䭲Cm��v�v�ܶ��t�-��6ؔ�z�`=�I��sUuT�MʽuUK媥Z��VT�X�\]6�� qb��  �m[ӭl�p�L� pғ��B��6�e��.���� [@�-�� �[UV��`BeZ�vh}>��h�X�i0�	��� e�W�����`� vкY�d����v�t��FD��+���nԌ��RS���c���Qä[PY�v�=	���1^�N^
���a.6��}bf+cj�� 㪃���$X�nvn��t�<�P $�Im����m!�\X��c�kf�	8R��Nq�6�4�Y%[@��k����7	  �E�K] 崖��8kn��M�mUU.��j��;t�V���hr�(i��䀐��K(�t�m��$�gYL�2�6�  �^��X���6*��F����cdYd�n`���`���������URt�N�����7ql�J�)-*�g�r��9j���m�X4`k@�9�m{��9�k�bt�,NXRu�
�T�#mZΠ�5j��8�8u���V=�`��SWU۔gm�myg� m�Mۧ��[��quUL��G]R�ŷp�u�]��)��9�(���m�[\�����m:C�1Эu@���x�(�;t�8�-�ڪ���'Hq!�khm��դ�$4�^qm"[ۭ`��Z��N�@�/L�WD�ۛ&��oh�A�A&�J Eh�ɛl pd�R`�f�(��-�����) �e� [G�m�8�Ѯ�P[@h��d�����#m]68 ��$�m@WYEJЪ�մ�RU*�UWM����O@��K-����l�Xd���# �\��֗ﾑm} ���m��f��v�	��ְ$��   6� -�l��d� 8'Mz�vؐ���x �Ͷ n�u��n�8$�-�mm��[���� rK��Wm���Z�6����ש����mΐ	�U�Sk-��vy�VV�[\�6�� u���l� -��.�ջ$o  ����8�����` ��^����ZZ� ��lN&� ���N6��Ѭ�Klt��(�V��������ۉ�v}R�um{h����:u���ce�l�,2���.)���+)
��k�(b9�6��2,Ԥ�JN0Ia*�v�;N��f�UR�n��E�V�U��0p+2�1�j������c���[T����l䲶� %�Ël�f\�Hq@Z�b6Z�\UR��ey\�5l�=z�MK�{[�h����O*��Q�m�F^�����7Hl�����6�Pye�p�WK�k�t��W@Q���++uJ��H,0��	8H��Iݰ	h$[@IK����f�' ��H *U�]�Z���(J��sO�}gN��h  -�m ��n��8  HNI� ��[�lh7U�h $ 9��M�`-��lv����j�ت(R|���}�m�t
]m�rR�I!z�-���3��	�l�i*��6imؒW���۪y��t!a�e���^{b֩IN�K�"�fT�	"n^{U�4�M�]�X�:��m+�E� #��R��Y$&��P���K)�A�uP�(�UO+O-�%��[�k�V�3���i�J\��4!6�]W;J�U&[��~P>�u�8�ek�*��V��V�w-]+*QJw��a~�j5�H�Z����9�
��h�/�ؽ/X|߀� �    ��@�VͶ ��,�n-����f mZ��ܛQ6��$� �6�i:�l���ط^�[��8�u)̲�uf��  ��;l�E�է
��l�DK����k3p퓯_�Y3�@�pH�n6� 	8� l�@��iͤ�d ��$ ����� �!K�l����wP"탁�y��.^�*�	(�8  ����m�7e�[@   h� ۑu���a�l:YN�m�� m�Eʓ�'��h�`�t�$�M�������H[tP�k� M��H�W�m� ��R���A2�Vie�M:m���nqW�� ��Y����ԛul!$�t�I!��Ӡ�nհ(��J�� jj�X��3�9K���M�Q5]R
(�\���<l����+�UU]*nr��r�T�.��J�U�U/.�k:H�m�Ŵ2BI��dr�@M�-ի8<fj��2�u�u�^���H i�]��0z�]�3����j�ܻl4]T+��h8.�.��h 8����4��zق�[����` []�-�q<p��+Q�m��U��cn�a�mm�8�n�R ,�2[D9k�R��  ְ�f�֬^�՚�7_T��:$
��T�n<P�am 4Iյl�8  m��ԉ$[zt kn�i $<�]6��*.���L��d[@��_L	�m�ڷjR��m�(t��z�� ��oY-�+`�n�C��n����}���'+U@غ�q�:����L�@	g/7:K��wU0r��>]�*N�ڷ�g� ^@�Z���(�@����v�i5�f��lp��m��.�     �cn�d�m��� -��ж����UUW[JK[YD�U
� �T�@]klWZ���I�z�ě M�lx\�� m�@�m3R�mn��l �@4Sd0IJ�l����<U��  HP]�ygb�R��91�eh�L�kh�u�m�8�r,�$�6�{e�ڶ'%���!"%v�7$�۶k͇
���iЭ�0U*�[��n�$��h��#t��@�K���\��2l�ӭ�ʻ��X�^R������J/AT.5$���m9v�i����**��
A�D y���\�v /��!�|�P �`0I���0+�"*��S]b�RV���@�?"ȭ>�hQ��Q�ڇ�lSb? C"�U"�Cj�E�T�DH hD���M.�_� �E�� �$:|�|*�:��ņD��3�P6�? <
��ʯ��G_(;�~P"���B&�B�`�	�S�k�'�S�x���T��*!A�ʈmP>�" �"A@b�!6���*t�`��B�At&Q `	u]
�@ �' �/G*�Q0�A�*mU�@8! T>U6�� ��qP4*PQ;t"�;  X��(iM+�Cy����:Dl��*�6��P��S��(!���=@p��#�P�v ��`�� �a$A����[*��"� 8!�(�qT�P80J(� `^	0 ������>D�C���	 A �D �H:�*]�L���� � !��=C@�>� 	q����T�H!f+���D���
%�A�8�a
�^
��tT�6�EH��耊�D�O�O�(�j�@��1AR, )C D�D��T�~h(UNo�s�m[[R�  6�`     � �  6�   [@�Ѷ�m�� �l�k)�L.�liK���A㉪ŷ�6�N�V����ݣ'-Q�/5`��@�;vR���r�sl�UY�� ��MJ����l��ۢ�J�����u)��j8&�죖5��x�gl�d��>)E���H��Q�T�;5����nJl��,݈�'l����T(\��K0��B:+Q�(�Á�6�6c��r��$�G��Ke�R״�+;0/]I��py��鬹�7ˍ��vXV&Ch�ÝO����)q+�.��#��t����O+�+�{p�`��4g]�H�6�  ���v�b�����K+hz��\Rf�@9t��� �*s�u�lx�D|!�.�
@`�e��Y�^�F��Hlh�1�6��`uڸx�T��q� Yku���clq�k`!9���Eā7�t��pW��mYdK1b�4ĥ�O4�����r�9*�d�֞��fFC�ҰiU]�<��T�fڕfR�r���v
@GrWl�m1�S�X�Idӗ�$���JV+%-��(�b��#��n�N^��ќܜ���t�u��������] �AC�=�\���;X�H��]�Ȓ��Rx���29���4
Ev(��Q��M.c����������#�ˮ�-��YR���n	̏����W*�HMIu��O3�����n&��Ut��[Ke������������q�R�GB�[A�v�Љm�����˅�	;{psl,��`M(Yc��[3`� ��^�rrrbz7\>zB�Lz��.��}d��6��;����.y�nl��=c����6��apm�@%�3�1�X��Z<��1� ��v{쮃�v*OX�OiJ��4��Y�P��(Eu'1�l �79�Us�ݗ��J$&�2e@?Q!�v��@ 	b�,B(�S�A6��S
��@�<v�|�2�9��?Nrr�NI7~��[UUV,�2�ʄ]�g�)�Y|�;���4�[��ۊѹ7@��3�����0r��M='cщ�=�B����v�q��U��^]�qWf7�ݲ�+�X�e���:�=v�&tz��rP�8.8�d�c���x7]R��A���"�ڕ�6
xj͠�o�I`��n�ӧ[#X0�/�Gf�X��/''s��ȳ�K�rY�.��M�Ļ�[��BXM���(M!���Z[�Mv�7ryx�t�:����X�KbH�o��j	 �o�g!����LD�,N{�ޓq,K�糉�c8�3�8�ŷ9�L��X�%��}��I�xA�"b%�g;��5ı,N{�ޓq,K���є�Kı;�{m)Lw4GA.Wu���/!y�_�z��^B�,O���I��%�`����j%�bX��{ۤ�Kı8p�K.pZf��8��s��5ı,N��ޓq,K���є�Kı;���I��%�bY�;���X�%����JI1����an3��Kİ~�te5ı,N�=��n%�bX�}��)��%��)$�8�8���&qI�r���W/����E�=i�e6%|O,�*4t&�����Rg7�8+P�]��uy�^B��s��&�X�%�g��r��bX�'{��I��%�`����j%�bX�o|����(��ݔ듻�^B���s��j�d�h��R�(��,#�:p�>~���&�߶i7ı,p�X�%��羝rwy�^B�y��C{ hSA�s��Kı;��f�q,K���te5��C1�Ͻt��bX�)�=wŇ8���/�G�B�E�*�7�n2i7ı,�wFSQ,K��s��&�X�%�g��r��bX�*I>Y����&q1s��WV�Һ]�&2e5ı,N�=��n%�bX�}��)��%�bw���&�X�%����j%�bX�W���%�3�9w<=�KǞt�W\ۭ9�ק�S-�$�н<�^4+n�8B-A e;��y
�%�g;��5ı,Ns�٤�Kİ~��MD�,K}�{t��g!y���ր�"cE��^N�!ı9�wf�q,K���te5ı,M�=��n%�bX�}��)��E�LD�>9�II&6ۜ���1��Mı,K�=�)��%�bo��n�q,b8�a���� ��X�VH��E�X����ɘ��fy��5ı,Ns�٤�Kı99I٪یً.1s3�2��bX�&����7ı,K>�s��Kı9�wf�q,K���te5ı,Nc��8�1sl�f&f1��&�X�%�g��r��bX�';���n%�bX?p�X�%��r<���g8���-y_��]�������ZƜK���bM��- Jm�F�@U��<ԋaB�fK!���M*�wy�^B'}�l�n%�bX?p�X�%��罺Mı,KϹ��5ı-��zy���^m�P�듻�^B�~��MD�,K��{t��bX�%�s��j%�bX��{�I��%�d��]}��(,�y:���/!��{t��bX�%�s��j%��������I��%�`�e5ķ���x�!=mG8@�u���/!ĳ�w9MD�,K��vi7ı,�wFSQ,KI�9�B�RAB	E	�}8�{�M�B������δ����	�^MD�,K��vi7ı,�wFSQ,K��s��&�X�%�g��r��bX�'��{ř�[mɛ-��p�mp�gqۮ��=��=;�;wiӇ 4n[8ٻs-���7
k�;��y�^B�s��e5ı,Nw=��n%�bX�}��)��%�bs���&�X�%��𞓣��b�Vf<�^B���9���I��%�bY�;���X�%����4��bX����j%�bX���'��a
<��e:�������g9��5ı,Nw�٤�Kİ~�ufSQ,K��s��&�X�%����y.;D��+�|�<��S��%S��Vq|q3��L\�{ �R< ����{T)ut*�M7Cuk �� �R< ����b�:�	+��BV�Ph��Z�H!��ߩ��w�~����m��/*���X�q�����h#�n�ݑ�v�����q���\�4�;/1�,V�M�A��Cx\�óf�.�3�9�5�۔��u+4!]���@ڱ��b�;kzQ8j4l����}�Ӎ����n���΢0Ѳ��WFR Ě�L�1iD�D�\!�]����]T�&|K�#T��D�d���D��eVs!u��?�8ru0�Ja[��M��(���K�9�]���U���3��ӣk�ִl����v�t��@��G�v^�LX��l�����ݗ���d��� ���ʑ�ժ�RuJ��&�����LX��f��x7e�.�;�S���쪵��ğ��_,z��v^�\0�j5��ղ�UE��Z�6T� &�d�`�``\��<�z�]N�v�+�T;���ɞ�E3|1SP"�e�$fh�̕�k-�s��][���o��^�\0	�0=Ē_0��y�b�bN�2��@�� �.��ğ9�5���T�VP� �[Y���ߵ>5$���n����x�=���U&���[�'d��6T� &�eH�	�tJ��j�E�mӻ.qs�z���׀l�;&�D���;.�����ݗ�yO_����``*G��/S�@�k4q���]k��Pe��唵���]�X@m��!a�r��/�5��*G�NɁ�l� M�x˲F��:��.���`g�l��y����*G�vkB�q��)Ӫ,�vʑ�ݗ�.P�&��8�Ԕ�\]쪼xͷ׺�wWT�]� I%�*G�NɁ�l���$茱��;���6T� �� �R< �����`�e�G.�r.�Ghz�0ny���p�O~���o��v׍ĹZ�Q��*m�\�6Ё������{ �R< ����#�'e�*����]ln��0rJ��q����z��NɁ�k�6��b��v�Wo &�eH�	�00�#�7�S�{��V�r��/~~������RNw�ԝ�ej$��Go}��?�����
�5eʢ��w�f�O_�� ���eH��K ir(4,��C2�%���T�z�|�Ӡ۰(uۗd��ݮC�V�6Y+leH�n��6T� �ٌ�:�Wmsuu���6[���^�w{x��f��x�[���,m����*G�N��`*G�v^�j�.��UI��wV�	ݘ�eH�n��6T� ��DuumUr�]��]�0�#�	�/ �R<wf3 ��{��ߛ/�]�� �v�5yN�� ���uX���C�&a���m�uj��r]������͢�F�A쬙���ke�1�P��
��4ک���`W4�1����ŜM!.��]���n-�1"�ᒴ��kX�F�l���p��l�Y�ö��㵎��b���m�{Am@mi����x���ǩ�K�̺c1��M���q�d�q�`��$��I9Χ99����IF�(;D�6T�	�21e�B<6����/8�G��k�5��,4eYt����]� �g� �R<wf3 ��������^�v�n��*�eH�	ݘ�eH�n��>]؆��)�uWv][�'vc0�#���l���z��٭
�N��N�Qe][0���ݗ�l�� �ٌ�>{�7uuN�n����`ݗ�l�� �ٌ�6VǀlQ�����V�����sy��i��2\u�=s̞XNv�cGZ�qR�L��5��݁��{�����LX�����s�0='� ��B�۶��i�ݼwU�:��8s�..]�*c�	ݗ�l�� ��Dt��U�UWM��V`+c�	ݗ�l�;��k�FGI�eҺ��� N�eH�	ݲ<eH�ժ�Ruv��;uww�l�;�G�l� N�x�O<��w��
��J�l�Fmpp�{p���kbV뷭�7W��Q�����˧��v�u�v�UݗV��,��6T� 'v<�������=�冻mS(���y�.s����^=^��'v��������\�[m|�M���{��=�;۩��Se�`�l�� ���B�0�
�ϐ(������%�,�Ç%x�WK��g����ߜ|�օ<d4	ID�A�j�:� $0�`�3�p#�c���֒�R�#*S�C	a��˥]���Ґ%W���Wc 7�&l`F!69a�t�Δ�eXT���	�v>�B�8��2�h�.@"N/����*�$�2ac	���~�Y�1��� �2��64Hi4���"��{BM����=����p���ۏ��b(o��2!!7��@at��²�� b���'��GsƲ�` qQ�hD�m8*�*&O
� ���0rH@t�.DG}80�D؆:*.�t���9����A�8�5=t �666<�}�pA�I��I��I�5��^�hZ�z�pA�A�A�A��];������O];����}�z�A�ll?+�q����;�������k�W$Ƅ��u9';��p��ll}��z�A�lll{���B��`�`�`�}��:w�>�Ѓ���?���?��f�,��X�-�z�ڒ��kY+��(\�l�G�q��a���;N���.��@��_�� 'v^����>�������]+�4n�e� �헞\\l��y��g���y�.$�;���_�2��jܫ�;����;�ԏ �R< ��x˻у��;M�ݕV�	�WeH�we�b��� �!�HA�bԊ#A9�G �Z"4G��?{�s�ROs��%�:�uJ�8�����O<�*���	����Ui`o˭���\�ͳjV�s�ת�Ix���[�u���`�;�33Q�:�tR�͒l�v����xʑ���ʑ�b��2]6X۪���6T� ��p�6T� ;�޼��_v7k[e�f���#�6T� 'v^��x�P��ت��U�n��xʑ����6T� ��#�5�F�t��ҥn�
�x;���#�'v��rJ�:���,�$�I�^sz���UUbͶ���bP�.a����#���{j��zX�v�'7J��z��@#���;u�l\M�����Hn��<׌%m�7���u��ז�*,�ȅI�m`�#.�����v��(��sD /��m��g��teh^����T�4�<�y�m��H]��k�:�kd���xݰ��4� �mŃ�nYe�F��Xku�q�����rͼ��~��G�3��v�K6��V6U�p���;��μӃgo;sX�S"�UsI�x���ݪ��N�]����x����x;���d��)�n�쪷�N��*G��/ �R<�ZĝՕN�E�췀k�V N�eH�z������]\4��f˗pwe�*G�N��䕀u�c8�t�c)�www�l�;�G�k���{׀��N͢�anb�f�R�ݸ��a1�YS��\���:��m	p���]�(��C.�7���>����pwe�.$���	�������N�)Z*�۫����x��%mq&$���X{g� ��y�v�y���_�Ī�?�o�ҹ���������w���K����=g�{�~��ժ�RuJ��*v����'=~��=��<eH�>�߽�� �=���]欷*l�;��l� N�eH��Oe�,0�o�q�kh�����OhJڃ	������Ma3%rmqp��p�#�	ݗ�l�;�G�}��]��Wa6[���� ����wl� �R<�[ʩUUb��7wyΤ��;۩'~�gn���XB*�b�U�$ $V &�8�$��s�I}�+�< ����j����UuN���dxʑ�����w��w�\v�Xh�\��eH���==^��'v�����݋��9w<=�ү�`p��66��octume�)�V�"ʥ�CACR����n�ex;���#�'vc0�#�7�c�{��V�r� �������O���f=^��	�/<���έ���u�v�WJ����f%H���l�������G�W:�	\Ӂ�{���RI���ԓ}�{5".�x#Q#�('���s�jI�c�=sst��UE�Wo &��.��f�[��K��������"���iF[��l�x-%JB���kcasb�Vԋ-%	�yZ��U_�������yLv�< ����j�����UwWV`�1��lx7e�Ip�;��;uY�4a�nQ���� ���.�����p���;��	�/ �K�;�Ł��//w{���vV����[��ʼ��p�<��>_�� ���Y�M1��� �-#1D��BD���B%F)i!$���$?{������ �W+��um��g�3�C�A��M�g�'!�qcK����v.�Sy^����w`đt#�M$=F&n���s:��l8b��ܛOB���n����.��+�����e6�4\<���q��7ml�Iqm�+vB��*�hjD�Ό#(a�0\y#=3�W;pvu���F��;O�2k\$�����SK�[1��#�'�M�z�� ��0Uֽq��]4������ݧ�6�yjϖ�v��r����vh�b�5���	�/ �K�٭
�N��b�E����kݕ��8��l='� �~0	݆,������J�a��w ;�x���N�1`���4-���TS���������xŀn�ǀk�V�F�;�m;���� ٰŀn�ǀk�V%lxɨ�1�->�gg�y%8A�����8�8{sʼ�\WX��m2�q�F��qeц��Fp��<\��	+c�6l1`�67
N���Pv�rJϹϗ�s�.�. �b�z��b���ҙA\[�m}��;$�X���.�[nRuJ��*v�]�%lx�%b�ˋ���<���V���4cn�ݱ�ҷv��JŀG6V�IX���lhS:����N��`Vǀ{�JW���=�� �d�X ���aWL�݊�Q5ҠlOl&3�l�k*jXB� �!�J�2��k��a�.]�=��v��<풱`���>�M8�8��@�;��ely�$���V,?On��{�����pıҫ�[�>�+�l�+�����/���1�%`����{޸��qeц�r�pse`䕀l�� �d�X����I�]*Vꀫ��k�V��<풱`+c��YC�j�5J�Z�jB��(�v9S��b��Ac� э��Ȅ����m�j˗p{����{���6Vǀk�V���4cn�ݱ�Օv��Jŀl�� �$�elx�Î��b�EӪ�X���rJ�6Vǀ}�V,����wN�]*���k�V��<풱`]�AW8�%�ŒֲB�*H� HE�H�R� c� �5s�|O�� ���q�q�U���wwX���.qv{���	�x�%`Y��HTe��Tn�Z�7$--.����`���y��r`n	^F����*�.���WUWo�;=�ŀl�� �$��q|�{w��;��>���0�.\��w�y��d~�� ���}�V,���d{��~4�tѻ��߾�p{����9��qUo�~�X��~��ժ��eR��J��Wu���y���b�5͕��$��}����|�����L��}�V,�.%+����ެelxٝiz�pε��]�@��-�AM�D��`A�b@�0�Ήq�$I��$��~]���X�P������h �bd1�4���dX�b1�4�?JІQ�w[�3�ˆ	F�����ʇuV�c(�	�̦�&t�X�" @���{vo�f���>s��6�#M3_}��XD� �1Ɲ������9@��h� m�q�F`�1�a���˜���� �Q���b?LN��Xm3CB��b�K�c��I4�X Dv�8Q"�L'��B7�%0�B�U�A�2J���� ���]>%6A�`]�ĺ0`��O� Ń�$ �6&C�>��a��$`B,�jg��|k#O��db�3�r!1!�#G�@6�Y���@��B2E�	ix�0��]���� 	��h  I�     m        �����m��@�㭫z�i�N3��=�NrEܬ�(F2�ي8����<��o�>~���۪�7]Y��9�J,b�n%\�cԩ�MueA{C����V��=���"�(Ī��&���Ww׭�hGb5s!R* Zs��Q��<�����#[\c�y+���8���rmp;+����'unM�+dC6�J�by/9����Z�.��is��u�r:U�0����zܜ��RS�V�$�;��jc�hS���+qe�`�^@��R�.k��[���6�*�U Ŵ�����b�R�pJ�6*��p6�E�8�I�6!��6�Xca ה��6�Ѵ�`Ajj
�Tn�չ��!�e%6[e\Ѷh[��W-���i	���L��˪\��mU�e8@ՍMV�0y���a&���oS���HF9*ə�
�6#���[r�\n�ڌ9�d
�:t��d�%�N7U�T-ӱL(h�g��{c	�Z�b�^r��h��1������khGjV�Ȅ�6^��`*�7`��4��Y�������4�7=���.�c6l�cc<�vۡ\*=��j���;#SW/2f�d����'6�V�5�Umt�m�[���G�\ݖ!x�jxU^�E3���L9�Z��'٦��`���+2%.�Fu��5�mc2/B�'�KR-�K�ۚ�8�T�W]P
�D�ӮV��.�����ؑ�tSE�<�DF����8|���C�����Q�T��.gC���,f�Th(Ì� ��!tM�ư�ݳm���Ov�֎�9�b�v6(/�붶[Z4�c\���u�RQ�pm���^1����gYS��m�x$,v96Z1��ޛT�[�&N3k2�;^��7ej  �s�۳�pGnĹZ�[��ק^n�А ��s�'d�H�n:�Ns� EK�Ä#5�EZ=�pR�I������&Ƞ<@�E
��Q>E"� L�P7wgn1�� րnջ]6��K�H�u��˹;B�B�'F�\�"�[s�L�y�c6��V�A�JɃ��fjJ�v�5��˳<;gs�ù�G8��e�3��?�վ��3 ����LK����	�Z�Z,����Aɞ�N+�<����r!����{B�YW;���f��*�IdQ��)���]����b��7��:!q���XD�w��NH�K^�V�is�J2��5��c��*'6M�˹�����l9�v�4��ﷆ�nGH�߽�ޟ� �$�v�?/�v{Ջ ݩK�v�+��ir���{��'�y��������=����l���l���8���@�;��m{� �&��q~��T��n���������tՉc�s�W��ē���_�� �$�.qq�~����7ƫ�.@�7e�����R��W�M�y�$������3(Sm�4�-l*�֘��ͣv(�yLiF l͸�#�Ӝ���P���P����G�z��H��`~�?s����o���=��$���h��V\��~�;۬!�"$X� 1T"M2h'� 8�?};�{A�n׼�rJ����US���1�bn���ʻx�~���nԏq���V��y�lhWuwC�VS�9=�0��V vIx�ĿW�~���$�R�GjһPΆ��=��w �I}����0ڑ�nac�)]�T�ދ�C�N��xY��2%��sG�S��rִ�V��$����yy[�0]*����|��``�#��q/˝�����`�W���f&��Zj� ����y疝��� ���`d���I&��Z��tRt���U�`z�`䕆�Iji%��qs�\�/���'��_`�p�]X�n1%��ԟ���~��I'~��I6I�������`uj�&�5T��U��� ;�V�Kd��o�~0o{��=��; �Ip�.�ĺ�R>��{�W��9������W�
�Df�n�ѝi�%�n��j�����O{��`���߾�����~��6��\� ݗ��d~�� 7���$��;��R�e��S
�EU��%`d������0	=~0��N3�;umP:N���I/�US��׀{����`s���*�����3�߾Ƥ�~�g�d3�l�Ux��x��{�x���V vIx�����ʻ�4��K�<u��:�����=�9.=�#�c}�m���%��ә��3[����}��\���K�_0���0��M��;,j�P7V`䕟˜���.*���~�߿~��7e�<�\l��,c�J�]�Iբ�� 7���$���I7'��v��ۀ~�{٥�(�Q�nj�s�s����I��k�V���{׀~���J�m)�F�8����?��/ˋ���������$��/�B�.1B�� "��3��.:g9�rm���k��C��GS����<�=�Ẳ�)KK�����f��Ӫ���A,�;:��yv��om��ح�u�ku���vk	���127b��)2�)J�36�OW<9�l��6t孊s'���M���J<�j���f�.�Z6ف�Ƣ%�����(�Y��B��[��m�F�(�ڲm\�_=���[�E�ܙ��쓓�r3�NN����6�ۦT�1K�d�ۗ��Jr�[�r-ú������͘��Ӊ�&uun����>�����/ �&���$���;)4��?;tY@�;�� ��͓��;���=��w ���wm�Cf���l� ݗ?&���X��� ��sY�4f�5���~�� ���V vIxI$�� �|4ߊC��-�uf�IX���~�����������.We��U	�(�#�f�<�ٮn�|����	�uآ�.:��I望�k�Q�Ն]� ��x�00�p����#��X��׸r$��f��=�{����BxH0�A�S靈���I��}�I'��s��(�bsߩ�q��I�+-Ն�W�� �$�=�$�پ�� ��}���OSN���8�l.o��\r��V o���6I���~�{߾�`�M?�����e����K�6I��nԏ �$�{Ȯ'l
�hm��.�mK����=���h�cb�Ǟ�����$�tB��'�[�8mc�!�MU������`����}�^=�T��q�њ��(p}�ӟ�y��y<�����`����$��qq.6G�o�"�,vꁺ� ���`d��qq�C�<*��}�jMI>�;�&�8�;�ш�j�.�}��O<�߾�����R<��9�*�����	��5��&s]��x��x��y;���G�z��K�?-�oޢ��+W/�Ҏ�f7G�)6s���14"�3C˄���ZM3�*�i�nC�{���rJ��/�\\��'��uK)y�V�e[[�5�+<��M��޼{���7jG���_�*��&��q�v貁�wwX?~�x�00��rW��߾�p}�zmc3�l�Uxy�s����I^��5�+�\]�..|������}��>��i�k�.�5��C�{�H�rJ��/ �&�s��7T:��2�mf����n&����4CQ,<��V�Hk4Q�9)H�?��������`uV���߫ ;$�d��>a%{׀~�u(}�ш�j�.����>���%{� ײVy$ٱy5��j�sU����﻽�?��O��Uy����~����QLZvR�mՆ���%�� �{Հ�^�'�~�=M;`�:��4����{��8��޿��{��H��8���$���'�{�;��PUUX�m�j�B �#E�Vx.�j���Y����'���i�,�.sm�7���mp,'I�u�m<l����T
���<b|/��!Pj0e�!u�6�d{bS��ɚyx�3�
;T��@���j����hy��������ri�˹�0.^�kYe΃v�h�4��Y�i.�ȭ������ׇtS��ve��l
��be��Ϻ�:��Dů.`F,��Q!�F�tv��,�=��M�Ǝ�����XB,��!�kX�յ@�:�������dx�I~��v��ۀw�W�k�Cf���;6��͒W���ެ ���kN����vL���������=�����7}o� ��@p�j����;��5�J��/ �e��?�I9_w��=�u(}�ш�j�]�{�\���=�>?OVײVتD�
 ,	s���V:�a�[)A<r��Cn��	�yS��Ym�^z=��6\}$���f�l��d�.|�����/+��ӱS�[*�����%Ĺ|:hXL(��U3�#P�@F�T��"� $�i<'{9y��Ԑ��� ���g��q6n�e/0��T튪۫��5�z�f�������%U=������V�i����յ@�:�� ٲ���f�l�qs��ڞ�`�����Cf���?{�yN��Nq)^����=���/ �5�����g�ȼ�� ����s��Eg���� ����fI5Ԏv��'��mɧ0�Xh��*���=X^�X�e�\��8�h'���y�~��tS������u앀�/ ���`ڑ��.q/ˋ���/����F#�fUw ;����?{�yMJ���q��0�`2FCА�����1C�A�D��.0��&�Z���"&��O��W�d�7��lp��Ę��*+����
���Wɑ6���9�����C$SEb�&�_�>��!ˤ�r������B3�@~Cf�ch\�� �\�ʟ(�I	P˰��� c q���H�^!���1�Id& �� 4u��4~CNA
@F�Cb��t~ț�T�\��`��+��4&���@�W �|��:&SJ'Ca�;�8���������;MN˷we��U�������~m�����m���_|�gvb�m��E�L��X��-�VϾm��LOm��J���;���}ݟ3�>��$�{~�[�R��e(�MBjD8��N����Ko&��Hϙ�����`�2i�k��^l�� ￿�}������o���{�����3m���b���UX�'Wu�Ͷ��,��}ݟ3�o�s���[%}�m͏0�j�ƭ���S��m�v|Ͼm���f7���\����W݀{�M� ��M=�ͥѷgAP������cm���_|�o�2�m�����i!�����<�_m=�:�`n�ٍ��[%}�m���1��wg�������cm�q%ʑy��*�L�0�}��K��fU@�a��#��;���ݳ^5nD��]��&Z���+�~ <�����=��|�}ۘ�m���+�n(��m,��-� ���^� ���E� ��J���}ٖcm��(�&*�E��"�Ul������cm���_|�o�2�m���=����7OKE�+͘/@|��U[sޯ�m���f6�����|�}۝��g�K�_vٳZhe�� ~�ܳm�����=����۞���m���+��m�dA!!,�jRД�Z�KB���iB%��@2$1X0� �����on�~~�� [@v�iyU�A�1��4Hn,��76�Rݥ����i.�g�ڷw(<�yVm]��-����zb;E�^��m�rgP]L�ià]ϵ]��c��� �����vP�l�4'AI�^:4�t��<�u�`m�3����[��۶d����H1U�N��a,'�;n���]\d���4gۙ�m)��m\.��1t+#���5�H��T�H�����s.L��-�(�*/)))��(����'^�gS[X&�C\��Pg��Y:��ZJ�.��
y���/}���LOm��J���;��m�Ɋ��f��3gAR���7�C���`�{���l��W����>g�yr��~���놩�%�y����`������_ș�}�~ݛݶ������n�pճ�gU���.���z�@�y�e�v�'��q%ʪ�{��ͷ���0*ڻ�]�f= y罗��>��瞿w�m�����;��m�P�@����"���gXo1�b�3G�XK61�4-ڒ�M��5Y�&afͩ1�m�/}�~�{�1���������~�����$�����枷O�E�W�03������⣵"�b0"DQB� W)���@=�Y��ѝ[m�������������Mo��UUb����������x�nI>g�?$��r��W�>����|�z�-t	E�/}�K��߽����^������l�NNM��{�ހ|���������n��ͷݩ��m�&���������r{�e�
{<=n���͌�©Tj��f#qi�f�+�&i�J�-�:�Z7B9�}�I�u� utu�W%�v }��}�~�޺�6ےO��s�w���^���b�0��WZ�r���=�z =��{/}�}ژ�6�rl���K�T�����[Ws+�L����u�w��7�C�y�u�R�U��V0)��p\��Ow��{|����uս {��n�l�ٍh�P�������ۓe��m�f`co˜U^���� �O[�Ħj�Là(��|�~\����6����o�o�s����{�h�t���.�i�L�eҥ��sG�S����9n*ۤ<0�e@�����6�v^#m�27�ͷݹ��I9��s�������?��:��L��%j�� ��^�}��'6Ǟ��� ���������cm�ي��v��\�Uu!�`�_C� ��={���rM����/@�}���`oR�ۣ�j�:��o~�IUW�=|�{=x�m�$���m�F�1"��U��^�Z�@�'�R�pL�u��r���=z�V�|*���߾��w9����{�w;ݡ�7�m��PHe���#؝�8�`9�v0ux-��4��D5~����B3�^��g;4Y{ =��� ��� f�������cm��E_6���ʪp;����u�99���N*��=�=���od���~����ݸ�z���ue6_�wc��o߽������01��ɞ�}�~�>Ӡ�g���5�������q*��m�=��|�}ڸ<�rI����=���Wbe��(�v�o�27�ͷ��K�/<�Ͷ�g�{ݶ�Ή�m��*E���"g$9$��/���oUUU]6ʪ�Gm9X��Ud֜���6Q�B�V;=mn�m@�F��ɝ���n�����C�/ �.�c���ܥrnݸf�em�Ր�!�n,��[�]�s�q�4S��gcK�3�|}��/9�s����6�5q�0]q\Y�d6C�Ur�ks�������ʮ�!�� ��S)�Y�FNt��$��K���&h��M�b1[�bM[4sW�s����k���Y��Ik��c5������s��̥bf<�b\2�߹�������)�$�@멧Yn�F܍r� ��'@6��/�ov^#m�fF����Kc!���nu�*t ��}���8����#�������6�ݸ^yqUP����&Z����{��~z���}��w����� ;��^� �y�/V̋3��,���o~����`��'@߾�;ݷ��=���M[m��n��ͳmk�.;� ���t ��}�~�����L������e�ӻ)n�\�C#A�Ɠ����۳V!��f"� �ny������N�Zf��S� ���=�6����od�O���s�v�n{�Y��g���m[�j*���=z���&��m\ov�_k��ݶ߻�fj�m�}�￹'6���u�ؙk�J,�Yz��������ve���q%ʪ}��|�{>z����'������d��;��[=���m�����m�e�1��*��}�}m��4�ƕ�9���3���� ���wfx�	�_��wf,E���ݛ���ȕ&獲E���`)�7�1�CXU<�7%��CVG�p��l�,�%2��?l��r��vb����j��@��3����=�^�ϥ��{�' ?{޼���<�6yyV6���U��RO��hԒo��u6$��4����R�7�g�ԓ�c��5$�]�Q�.�U2��.�`yq~⪓���6W�� �[R�?%Ğ��� �-���UQe�����R<���^��ݞŀ엀k��Z��S��xU�%��u(����73e����u�C�,5��Ӝ��8mfQ��\�ٿ���}�� ����`{%�v�x��R[�E&�Z*ꮮ���f,�����U��^��~x}����N�V�gl� ~�%�v�xys���T�V�=� �R��̢��L��'�y/�_������ԓ����2te�b"� ���M���]��&�����f̙�ȭ��{�����"���%�=���~�xݩة좍��k]����n�๳'d{tG���ɳ����I�GggIu�����{K?��ŀ엀}ڑ�q%�ϘzT��ֶR��]�T�㰺��vK�s�qq&��{� ����ً?q$�:Ű�_�v��.*� �����;������8�{�ذ��^���U5V��SC������q?K���7g�`ݒ�?��y����^�t�9�hMgg-��ˆ }�/ �jG�M��X�q�T��J�F���P��b�
B٠2+���x��E_�5�M������M�R?&�Sh�]���tiG��q���X�R���R&�0�2`�D���\ (UPδ��Uq��'1��p�:M���V&B�b�2XĨ}��  �m�l  ��     � v�l      hm��� ��kX�%hëT��"q����� ��[eI��#kv��g�^2_"�{"���˺c�
�@��m���|tl�`ȓ�BJ�*�˦�j��p`��ڱX���T�s���F�Kqa�k�S`^�^�Э�-�9*9.�@�z�F�8 ��z��6$�<:���ԅ=GSg�P3�\�l�.;^�� �h oZr�l�9��ΒD� �jKmv��X������;s�HV
�#��1t���& �]E!u��ޘ�)V2bs�6�5;*�p�v1����w[��>��p�˭uj�V��G	B�`�X���.q�.@u!���ZU��;5c`���)�5l.��B<R�E4w�m��P�J������
��
��f����g %�3TF��>2G  ���qŖ�9�m��KVŭE�cs���㫋y�W�F��uu�ukn¡5\�����	J�Y��r�v�3<Fd�&�����&tB�R�%6�N^U�m�]eY�%�8��5=�x��E$p	**�=�vS��7�)��vȚr\�qK�@����Z�s��V�dm��a'R�+�b6
�����C�؏+��h���'DO@�*�!�+*��hKգ#�PI��Z.���՗j�1�!S�Ű�Y:�:�oH�C�=�8ST��cg�:���R)e�8rśI�t��V������aI):ѱ[��J�:�` �il�R���]Lv��kr�3.�c!����+�wn��Y̠ZA҅����"�d.Vj�,yN*��P�6���沕+a�,��B��m���2�� Ɖ�8l�c)�d�ʨc#�.�e��yl��ͤwmK�a�ɞv��Bk�J�IR�af�`:of�;�,<����m��66n��&�[�e����k��KY��$��#��*��@�	@�0qj��=X����Av�6�TD;�gRrry�NOy'9��u��{UV,��U˱(g1��݋A��BdmW@y�n
*�7-n'��囬!#���p�K�q��F�#AαU�q�+���i�wdx,�u6�69u��%�ð�&,��vw��GV�B�wkiV��LN���X��ٻ���ɜ����ha1��țs�h d��;�q�M���Oh��v)Ǘ�L󎬼[�nD!�l\V5gs�nM:�A��n�b�H�l����Zys�oX���1&��R2�R�����^nKo+s3����~������keג\_0����;��z�Uv]�U����;ڑ�ke��ˆ �w�?��O<�c���|?�6d�vF���^�u�w��vK�;ڑ�����͐l����O<�_}�� ��׀w�#���~�=u�u����vU;bv���%��H�	��� �e� ���U��+�Vƭ;EQ,����h�³�7�Ɍ����ˢf��X�$��Ô𪪶��黻���׼�	��� �v��%���^6�QE]�I�<��1��'y�w8�vE�gS���Ow�����v�y����m&��wAH��S��wu��׀vK���I;�� ���;�{�FS���9���]�~�o��^�^��&�ˬ�\I7�|��O���ح\)���n������므7}���%��l� upd�p����nY8%F�K	�5�#h[U�z�
��qtn��sfe� ��`{������q.%�����}�?��d5��rn ~��^%�û�^ݯy�}����ě:�����Tڲ�����~���n����w�i�B"� z)�s�Y�Ơ�^�t�8S�i���n������I��<9��X{&, ��^����1��k
�ټ��ޛ�}�{�����x{R<&��ݖ��4��]����&,��	�Ą�Y��J�8�4`ĵ3n��5kT����� >���>�H�ľaݯxx��L�`�fq������y��Z~��� ���<��ŀwT����ݻ�E+����>��0�������{�, ����=��C��g;%S��{�Ϧ��s�ѩ$���u'�J�F!U��Ы�O�D��=��P$��xڪ�X����� ��b�����n��p�?s��T<�YfԚ�جeS�ˏ2u�.�bMJ�� ;>"\�kGJ�䅜�����iP�? l���;ݸ`wU� ��b�:��s�r@v�r�[{����������&��+�`=� }ݗ�ots
(���6�v����#ŀ}ݘ��9�&��y�����=�w��4�Tg ��1`�%�wn��8��x�`{��|iXE�\ms8���x��.wfx��� �ً ėW"9���$ 8��h׶�f�]��gM�	�4�U�S�j�7a��j�t�]��3�8}y
K&�Oj�^���U	���[<��7M�f�Zl�V�����θkX��p��^SZr�5�Y�@�V��Hf�fYG���Ë5�/9,�Y<^�.6v�l����'s�I6�{Y���roI�8���N'�6��ͻg�VS���Ml�EY��I��9�N��v~n��B�`��s�p􈜽(��ۢ�����{f��f�lu;��ZZ{=%]�l�vC;��%�.$��@{����;;����2g;%S�~��ş��ě&�b�	���M�g��������Uh��AV�N�6{ od�"I��B����`kv�T�2��+%����K�;�~0��ً ��t�9E[M�UM�]��ۆ�ų�/���ذ{%�(�ϱ�.;Aqn6�쏎�N����۩�gw�u#�9a��mcuS�]5�\*����ŀ}�1`�K��8���9�	=��B���v���)�����>옳�/�9ľG9�b\\Y��%��p�;�<�NrNNsk��������]K�:�=?~�{.vG� �ً �m�:j�ˡ��W���K�~�� �ﾼ��f, �d�)��(������՘d��s�}=���޼{.���:Z\:>s)*`��1�o7D�=[N����V��z�9�6�玁n�]Sui�-`�1`�%��p�9Ϙ{߾98����d�Q
��p��^~���l��� ���	�1g��/&Ǵ�|y��3e��[Ux��?� ���ѩ	 �EO�A8 |�&�C��o���I&���RM��z�ŗe�mS*�����{�� ��ذ��?'�3���ti�Iҷv쵀Nɋ ���z��_��t������b��-���g���#�C��y^.\�۶��vN�v�g>�;sؠ�cY�]ݗt*uk 7�^ٷ�C�$�P�߾����P�Ύ˦��W�wv៸��&���b�;=�X����/�<�c���|?�	�9�5N���� �dŀ�/ ��� ��X۫N�mաӵ��$�}��� $��w�ѩ0/���z!QB��>��v�|����M��`���<��%�{���y��7�b�;�7�	P4��J�����j��-�0=Runyh��sۣ����t��n�ܓ��.P��n�X�#ŀNɋ�s�|��=x}���v6��2�����`�b��e�v៸�����J��B����YSK�Qk8���8��޼?�8��{�{�;-6�J�X�쫡S�X�\M�O^��� �d1`~��{��� ��R�ƨ�M-u�xf�0%����~�utO߱`۲�'T�F� � @圼�%�n��UU@UV���8���-�jƢ#p7��[��,��r./��7,�Lj.�ŭ͹�=A�c�1J�b�K�잘�vޞ��:+�\�<�o<�M΅�J=k��	n�Ag��Н���ӡ��a��4]
W[v��ت7]��
�h��6�]y]	�2򱌥�f�c��il](M�ɢ��LV!l�1nD-�X�34̱��䜓�s��䓟rN�����m��j+[��NF9�;N�v�n8Vx-���յ�:�k��L���T�~�NN���' >ݗ�q/�zOb�&�y5���:�N�Xf�Y�s�6�׀M��`l�,��ٯe/> �ջ���������7�b�>�Xf�X�M5�8��ۥUuT�� �ɋ ���͘�=���׀{��1�.�ch�C*�`vCٳ w�/ �dŀu�����)�Ũ��������>��m��� P�6��_���֬��+��@���X����v�	�i�
WE�we]�����ϗRX)"����W��	)ė�!��ŀl�1`ݘ��q&��X��UV]�7t:��;=�X��b���=� 7g� �j/�
.�����n�`wa� ��ŀ|���?s��[�ߺ�	?/ɬn�ۺn���:-`ݘ�˜I.��W�v{ذ�� �Ⓣ���i�.Hˠ���_붅����j0�l�@�V ���֝���Mݮ����>�1`v+��Ϙl�ŀl��?'m6�U]:uu�odŞ��Q���?{�,�vV�T1e�vSERWk �b�`�1a�9�uE�e*�Bi(�,1���(0��%�����;n�� ���C�W{�p5�ӈ�!���� N�O���� ���ؙ��S:CⲒC�b|�1!"E$��!����|*
T�XV���fp!{r?;p$W$	A�5AI��5Dv0F�%��g8�Ld�$�&#4���1$dB�&2���'ū���'A.i�MT�D��C9s�VfL�/��qN/� &�C�O�P�x���? ���B
!��A< w��q���
i5�\�ԓ��tpl:{��,ɥѫfN���}���`��`l���.�ۅ+�ڻ���UZ�:�e`\�9���ߺ���_� ��ŀlQ�����MVDiw>; tD���cI�x��Gh�Gs����kd�jX7m����;���y8���wf,�vV�lD
.�����n�`lW��͓ذrz��LX�(����:�M]�wf,��+ �dŀ}خ_e(�!ݪj�i���u�e`l����:�z�H�V�	Eb�L�L "R �CB;�Du;/V�����L��J��ӫ�����wvb�:���%�z��y;�e!L�S3\V.ZML�Rǔ����g��vȝm~k�4Ը�@f%2����x���ً ����>�1`h�ʺ��T[�ʳ ��şɳ^�V��b�>�\3�q���M��N˻*�eU�^�V�ɋ�&��_�d�,�lh��[��nʪ����q>�{�w�/�6LX����`O"�x(���۪V���� ��./O{�'/{�jI�w�5$�8b�P� � ��8�V+�)��X���� m�k�]:��.��l�y��:��u#ۆ͙�����B�N����n��V��<a�f�/n��$���6��ԭ�9Zǝq=/8�{���\a��3�N܊�;0#8h���qAn�݆Q^Ga��9�-�t�n}i}<mj�be��m��m=(�����E\���ԭ��մ��jB�����\b�4̹����z���(�E��쭖�6����1��&!�.�)����Lite��;8�aM�:�����&��cU����g�X^�l���+���J>wj��mݕV���X�1`lWl������TE�o§�;i�J���U��߿b�>خ~I.7��b�5���7M���;)��	����ĸ�<����b�:�e`dŀ{a���AfM6�sx}�y8�%{ޯ����`H����1�EƓ93����$�aۓ%��`�ɘ5���V�X�4(��FQ5詜�po{+ �&,b��q|���ŀI-�x�j�@n��[}��z�~�ܓ���F��B1H�"��?�K��߮��s�ѩ'/{�jB)�@Uuc��T�լb��&,<��&���X��,{x2���7LeYEݼ�\��{�,?{Հnɋ���_��{�^|��4���Z�5�+ ��qrO{���^��;$��	�ӽ�d��X��Eΰ��؍��M1�y�G5pv풢���l����!ng��U]:���7dŀHT� ��IX�ye�N�h�Buv���xd��rJ�7dş�#G�껶Z,��[�:��o��X�%a�\�\\�qqUIs:�G�N�M�S-]+�*�mլ9^�� ��ŀlU#���$��}�s�o����W4���1`H��1`ݗ�{�$��{���\��d!����0�2���	�!#h[U��,����C�	��[T�ծ��*���ݘ�n��>�1`uG�.�ʦ�L�����ݘ��M������,uT�?.$ٯ}Kπ;�m;c��`����1a��q�j�y�=�X�M�T��6�U]Sww�wdŀ}
��ݘ�;�~�9�ƒp�ڢ �T@U��F�e~EL|���W���u$�r�V���T���`B�x��͓�/�='� �dŀ~�9��J?xC�·��8Qcx9�n8�n^ݷ7A��;Fׇ�!k��c���D�Qغ����ܜ �e�l��ĹĿs����~� �?���Euq����޼��{��'j9Xwf,�s˜�Q%͍US���UX��,{F���q`�e�v����ӻ�T�լv���wvb�	6^��O���`�y�˫�TӠ��e�`ݘ�n��>�1`��w �O$����or�UUX�m�����*�r�n5łtT��K��[lj�ku��(z�og��m�A!�nj�Tu�ţ�-Wi�X�����۞���#t��(��cN틗�y78e�˸�K��J+**��������Knrl���"[G�ూ�Yt���cqN�V�*nɖv���k�y,k81I�yxۮr����օ�v@|�y<�y9�F��!�v��uCǏcnndlEW[ٹ)�������h�@~�y
�#��[L��C�] ����;D��wvb�5Jn
��mҪ���� �dŀN�%`ݘ�n��.Z}�����6��g ��}���� M�xݓ:l��E��T2��?%���O|��z��LXc�����^�F:+��l� M�x�&,�l� ��ŀ�9c����Bt78�	\�ū�D۞�]FwvG#�x�woN�⇙���\�_l}�b�;6����X�����@Uwi�۪V��ٶG���ÝK�V��$��9l�3 n�x�&,n��7wj�:AV��o �ɋ 7�^I���,},��:�)�uj�2�-V�=�q$��z���,�l� �ɋ ��oE.���t������;�b�;6���1`�K�7�\��ع����\�M�,��i��hp���.��]Q �Ĭ�����m�Yݷ�K<��1`�K�7dŀF��*��i�n�uV跀vI� 'd�vw��w�S��w�ZKۨ�G8q��Ԓw��:�s��Me�H(A�U��B��V*�"����S�U\E�(:�w�������?~����\۝�]��\�I9=��,��;$ŀ�^�ރ�ЙYU�F�p��v������|��� ݓ%�v�Zz�ح�'<j�ö�t��7WA��Mն1�\�� J��cj���@�*7�~�{� ��vL^��_0��y��ԏ
�v�-;WUk ����l��ŀzK<��1g���5z���[M�UWAwf'�� ��G��$޿{Հ{}~0	��Ȯ�4U �]�n��$�v\0���s�p�p��W.���>�׻8l:w���GE�8���p�`�b�>�w�\����܅jαsr���DVVj �<��� �i)l��P	s
&�+�\�~�vLXݎ��Ϙk��X�X��'umӺl�� ݓ�c�`rJ�7��\l����x]�wvꕺ��w|���$�{.옰	�;g
����2���������� �ɋ�}�<�k�R< *���Z���{.�LXݎ�u͕�%xDS�0h�	��cD�f�bψ4HR4�f�3������M�R��(m���) p�B(a�|�̌X0b�s�� ��#0����|�m��% ��=GCv�wو�`J�a!b��[譡�	��*�9�R��w1�!(�1�D≷���4���o�Ү�'��slI�C�7QmY6��������I����A0B�A���%I$@��eH٣C��iB;��۵r)߄�f�w<�;���l��/bl��4a�ZP6� > h�$չ�� �hm�`  ]6      -���     mi���`m�gl��m�WѬcc^kK��Q�+	+u@c�L�y@׭�3-Ɩ�CE������Ʈ�s<���l<���s��w<�q���Z�Z�M$�Ɩ�wQ�86k��aldrˎ+ۆcjV@�n8�d�h�%Pù��j��L�#����%e��;` �+�rev��Ħ�mH 챮�ûA������ۣ��1���W<����[��uҮ���`��7I1�s7�ՇY�&,8z�/]��� ��gS�x�q����dFGi�	7T��h�Z�ݧ6^�]��S(b`̱���cG:����0�jM��ܶ�W�x�;Ju�ec�-m1�U5ʲ�C��s*���I�T���q�B�ty�7cm[�EC�-���F��*݌�P����y�	�ER���o8�.qۀR���=�����3c2�YEDbکZM��ɺ-���x�nx	�D6^�[��w6���(��K'�֢���',.�T9��a.͢ ^t, �Г+�̋Ҷ�5mg@���U�q��|�0 <Ԛ���2;���=��t�+�p<n�ހk��EY��vWY�,�9��%V�֎^7i�M��i�	`5��!%�SW.�146��"E�a��p�J��O���\�^X��p�S�c��CCZ�ԂZx���=���$���s��3���\���TNcvӭ�n]s@*�)*��S��N!֛�㒖uj63Gg��j�4�<Ӧ�	��魢ʭ ��:gj��fٌ���q�Q�Y�Ʈ ���Ѻ{�as��N��dɩ@��Hkp�.bv��m';mD�bUryAcB��J�m����6�r;���ۑ�}���e]�VJ2v)��xjݽ��ý�Ih���<n��u��1�Ve-dz�P���Q�8V֒� 5m	h.�p	-R2�L���
�r����r~�q
9���T� P�5 ����DW69h���!P��5��?@� :���6�؄՘8�t&6��$�N�t�5��u-#�!YK[lx� �����]J�ucl����nZ^m��Znk�60�/Qk�ċƹ@���0v��<����G����P=�ǩ�k�Ã�WU-!�Q�2�Y�"�[e�{l��w3yA��b6�v���Fdܠsq�`�����;��m*��Hs����8�S����q4��9�s�Iɧ9:�?k��� ��@��v�د5p4S�geu�!9���'p�/D��8�v� �1`v;��6W�%��v����0��@����4U �]���p�:���7��odŞl��l���jӢꋥv��_�� �ˆ����ק ���V���r���y�s}�0	��,��p�:���;�XԤ�t]�]ـodŀ}��\�X�\0��"ݱ:����N�x�J���vs�Ih�c�
����s�'�5OM��	��crU������=�����p�>�1`u.햅U@�1s��'/��5�U.4�D��n�LXݎ�kݤC�����h�WwX�\0͘��� ��+ ��oDKi�TU��� �ً ���0}���`MH�[T�T��Xݎ�{��ޯ����w����}$�Ϸ~>��� �1Q�:��M�� 9�RY��w���B���tyai�B��*ݣq]]��׿�ۀ{��Nٳ�����;����Iڶ�쫡�U����f,��p�5�J�;5XԤ�t]�]ـvlŀ}��٩�w`�N*�����q%���J�6m� �@����N�[����Is���0�ެ{.�茶X�G��wl�*�aN��5�J�$ۆٳ��I�}�0B������h;e�� ���v�c{��m�9ݵ��s��`������\�����f,�%���#�z�Jn6��-��*��n��;6b�qq.q��޿{�V�����D���EP��`^���5�J��\�M�/���ŀk�c��XZt;�u˺� ��+ �ۆٳW).uq|�'�NY���p�����V��Wgp��0͘��̳ ��+ ص�HU�blkm�yA
�W_1$$K�ת�wd��;����m\�8��l:v+5��f,�,�5�J��O_���|Yb�����������<������==~0͘���?U���wv����Wf�?~�l�a���7����?}߸���<&Wh������� �Ob�>�2�./�럿V�����aM6�WV;� �ً ��s�w��Y���`e� �\�y��v 7m�m[��bE.�ajӰ󃨖xl�N�/3/�T��讃�݀-�mPv�{�E*u�`�â�uc��A���N�`B�YJ܃R�h6��c�2�m>�mY%/_�ݳ���5̘[��6Q^!�����9k(��i�t��ж�M/98�mӲ�G�0\V(6��<��B@��#�QBQ�k�U��$e��I��	(�8n�f�u�^]�s�<�dŘ�JK�MD��y�͹[w/��@��C�\������Y�k���&ˇ��;��X�=�ul��wN�]�ـk���$�鳓����8��YKۨ�EL��$�`n�Xy$�}�V,�����cR���캢��ݘ۳���`mlx����0�ȿ5wv��[�n�����`���	%� �l��?����ǿQ)B�	sT�;+Dٸ��1˨cR�F�1�&Ǝ4Z�r6�LL�l��)
���Uk�#���$���$�a�{Ջ �JG�
���j�Ƥ��s٬�D��"��os��b�>�V,{[��zږ�n�Uumݘ�f,�%b��\Mͩ�{޿����(*�uuk �IX��lx��}6b�5�i��[-5NۺWwV��lx���/{���;��X�Jŀjk�`����)��ϩ<��p<�;[�y�hʉ�Z�3�(��t�򕦌��v���^���{��>�V,��+ �m��I��wn�wt���ً?~��UF����`��� �_N���zYb���r���{�9$���n�3�V -DZ$BB�@H,(^��et���ܒ�0�&,T�	�[�AUL�UU�.qq$�l�`����ً �IX�{��pUwuH��;��Ip�>�1`I+��+ zln�˔�6�4�Ů���� +�k���8w6�۲V��N�.�n�_��s�Ht��@l�.π隣`I+��+ �\0	�R��AT��X�Jő{�%�Ty�;����7�j�6oi4�n�MS���լ=�� �\0��X�Jŀ}��H�+UeP�uwX\�����߷�jI����RM��ƍI���I��'8��GV���6�+6�� �lŀ}$�X��<Ip�?%��w�x���P����Bl-3 ^�@��:�[y�3J��c]��$���z��T�]�t������� ��ǀnˇ�>a�Ob�<�^Y\n�tU;
�� ��ǀnˆ�ً ��e����l�JG�
���j��z�`M���&Y�okc�>f�j�i�|���0?q>�{�w}� ��ǁ���I���{H�5�"��WV��&Y�okc�7e� �lŀ���˜ q�����kf��v��p��^-���=-��<Z�B��;+��7Sٰ`%wmc���
ʺ\��V��y�es�,ܜiɌ��On�(��;�؜{�$����	 F�2��g�������{=����(=���k��>����c�U���) 3Aֶ2�s�)�4]\[A�k|��PԱ�Jf\ �¢K�T�n��6rs���gg]�F��4��p�,�pZM�hA�u[I��k_+)(�#���dt�p�Aq�ڧ}�����7e� �m���_������e���?�Ҿ]���*���.�nݓ,�7���专g|��������P�v`��ݓ,���_���w}�x�?� ���3�m������ɖ`����p�>�p�"�S
�wuM2���Uـokc�=�q%'���w��`wfY�ut�`ݖʅ��,l�s�k����h�C���L�ѻ`��V:Pm�+�V.o ���0��0��,�7���3u�e4۾U]"����|�B�8��N+E(� E�� ��h��xT9�����5e{� ݗ���&�i���PU �����e���<<���ܞ���p��/��Fdn��U8�y�q9�<�	=~0��0�&Y�}�|c�Ҿ]���*���.�nݒ�`�p�	�9enݍ�US�!����qTZx8y�[Z�ט.��yj�X�f�>��N%9�VU�����|�p���`�p�;��E�E�Ъ�Z�V�۪� ��+���.ӯN}���%�ӽ�^[e�6΅ٜI~0�aK�|ԗE�IW�P��HV�A�A���cR�3��� B��?:>ND Sc��Dç��*��$�PJ�a�Bd��m��A �# �"%���l�JH��S�(�����ʁ�.��� �A
��Ȕz(�D�(t6���y�g�RNw�5!�v���wv��h���}ݸ`Ip�>]ً˜�8��y�x��Lw�wAwf���ݘ����/�7��[��z}���Vh���h����Df���Ν����br g@��L��k���U�V@:���E�~ŀn�� �jG�s���s�v�~���Roߛ�v��tʻN������͕�<����:�LXݗ�8�W�eP������ �K��Iq����`K�H��JUwi�t�wf��>��� ��{s��f����b����榤�=�3�	��X�[�p����p���?�=�}��z��\0		dݲd�͂nh.1K�l�B�VZ��s�V�n�F&�tljPV���6g �v�w�p�>�#�>]��v��	��+N���NI�y�M��_�<T��X��3���g��g�N��|�tv`�{� �wf,=ė�_��/�:D����PU ���������`K�w�p�>�#�;/��{kd�Z�2�ﾽ8���w^��}�{�RM�s�5$���XAj�*-"�J�F����s��rm'4%��z�ڪ��f�5U��9]���f���Z]��E�q���0rWv2�]�z:�J��&��8����V��"�Q��q��kXwZ�a�V�s�AB�Վո�5�ùs�3�<����ȪqOg���5&�-�Pθ��f��0�4s��6��.Gs��mia�v�$޶�61ۜ��dn;m�1�%��;���Y��]@�N�X�ϟ\�^q�O��D麖�^.�VֲW+��g�^#[s-����[CB�T�
.e(����k������p�w{x˻1s�/�I/��/X�R��N��v˻0�H��vb�7v�}ݸ`n��Ъ�Z�Vʱռ��1`�p��.&�e��;����ceݲ��U�V�?�8��<��Ҥx˻1`�i
UwuH-;E]���� �����ճذ������{��-t��c�ٷ&�8+�\��/F'��Ӥ���3h�8�2�R�gtv`J��.�ŀn������0���yy �VS�Uv��vh�rè�	�Tj�~�(~EķL�g^���}*G�D�7����YuM��*�`���wn~�M���<�g�`vZbq����T�wo��I/ˋ�U��~0�_�<�ݘ��lx�X�J��:.��.��>ڑ�.�ŀwkc�>��0�ˀ;�p��i���nzD��>y�$�[n!u�ŅQ4JF��������޺�&�1b\۫>�g�`mlx�ۇ�|�J�x���cc�*����v��H�ˋ�&���<��vb�.~�9�T~s�B�]�2���{��po�����HB�9�Y�\�,v��Fw[P�SLw�wAwf��=��:�{�.�ۆ����tT7wX˻1`�9�o��>�/��d������oF��̣ŚWQ,��4��2(ńBw��x���3�N

�6���*�t	���0��^�X�ً ��LN2���J�*uv`wn��/��<���`=��.���^���Wv�@�v`�z�������ק �{�=,�\1c6.��y%������ߺ�	���0����0��E��A8C�'{��[�os�'��+�k��eui�.�q.���� �vb�>���u��F$2Fb.u�Q�#t�K���\Ų4t�
�L-r��w���BK:�4����π�� ײV��ŀvK���-7MP����^�X۳�.۷Y	j��
n��f,�\0��Ĺ�.*��{��_��� 쿋}�Y�m\�����}����#�>ݘ�ݴ��)_��Ҫ�� �kc�?.%�s�����I�{��I>�s٩&�7�
(�
��Q�0�0 B	Vӽ�I����ߞ������K��!�3�ۢ�{W����Z�ҳΛrT$�p�U��d�q�v�jݡqZ�n����Lɛ���CTK�4X�����6��R�yڞ�9N*FEH،�b�=��jg�qj��Г�x��ma1�Ѻۍ�7kh��'vt��G�^��@��.�'f�:ֺ�lk�b�u���@sKheH�faW,�糚~���wݔcʓk4ڐ�&�Mh��,�mZK��QٶK�޳w5�V-���`�Uwl�t�Wo�>����>ݘ��~��9��ʞx���5N�Wj�Pꮰ�f,�9�/�$������7��� ��+ �uF����0�uv��Xv\0��<�d��ً �!�j���e��n��>�������f,.'��� �5y��i��N�*��{%`ݘ��`J����v�5��5J���:cP�74�Jk[,�T�{~3�|{g^�]�y퇶B���=� �ˆ�����5�z�K�o~��2m���8����鼜�qg9�vWc�>rJ�7�1g�8��;#)/����Mt�)�?}����}����I��ذ	���(�]�)��U���ē���`g�`�p����y���ך:-]�UCwu�ovb�7��}+c�:���<�8��U�#X��qb�Xw�]%.wv�#��ɵ��v�T�^pj6�98L�����pw�k&�4�tO���>���seu|�vZ�$ֈ`�we�e��n��>�����v��LX�\3˜I�3W��l��|��e]�_�� ��Ň���8����R�:>T�k��ԓ�㽺�ݢq+t������X�\0�lx�\K�\�������~n�̛j�j���8����=�����z���XMu�1�E�;n��)v�w;=�\��sn���ry�3A/�+2�]�D�T`'l�|�T�Ҫ�� �Vǀu͕�ovb�7��n�c%*��S�l���u͕��I�l�,o�����?/%�����XMpŌصw ����oe� >�/ �+ �H�X:�
ES��;���.$��g� 璘 �+R~D� )6)�C�U��@���%�GJ.���������X�f,{. �67UcT��Bʴ�`�k	e Щ@`6K�c�-�����V��mF��W�]�W�~����ovb�7����q.��߯ ���~��t�H)��`ݘ��`�e��}����}�+d�W#Vp{� �l�=Ēn?OV6{��'J�t�'I��0��se`ݘ��p�7T���]�)��7wx�����X͸`�e��O�!]�>U>H�$FF�d� L% ��$��R� ����>bC�u�!��a> ��ٚ�p�
��2.�209P�5��:x����mѨ@��A��3.�	��a~P�8�8�����\����VC��y�B"HH�FbH�6����8�U0C�\W(CFY� 0H��FW�qn���2J|.�@:ȐH��XX�Ss=��� ���հ  -      h�i0      $�5�m�h< k��d!ݶ5ή��� ��5�����}�4"\(��url�=1d^t�S��j��ív����`���dX��(b��
����*:LfM���ب�B�d����e�,�l*�glċ�u2��8��TL+�D�b��cQq��&��e�v ����u0r��+�x���q���U���cet�U�4i�R��ʠGir9r0���@���|�+�k\t+���5� 1C;�i�yݒ�'�|�R����y�8�Y4֡�r��J(���-fը�.���ÔK��u/�ɽ��v�rgգ��9F�gL�A9��:�,e�
��r�!�+-�@�ʀ-�@.؎�+���P�s��v	x����|p��9* ^{�CGnٕ��m<�焠z&֩2p�7.Tp�t�n�sá9Ͳ[ͥ���S,is:�;���P�b4��2�	�]U����SxY2����ɑ�j�e����^3<��XQe��%��T����jJ�; S�+)��j�s֭���U�$�	��m����Ɏj�G>��ůl�^tnln�
�=���U�m�����練d-��@��/]�e�i��q�;�i 6Ѷ�
�l�v�n�uJ��:'BEr�T�[eB�n�ΰA6��Nn�V�޽��b���fwdzp�g��=�^-b��@��	�B<�l�i����ٶ 
<�-�ȼ�S`�%-�Թ���{!/n���J�6��=Õgd8��w�4�W�3�
�J���Bgg���s/�m�F�N��A�A�pr�&�I��v����Yw�r�l�`K��	q Y`�SR��m�Ϭ9�2e�ڲ)�M���lZ"����g�Iہ��q�^{c�{e�Uhu�(�z@t�����e$���7nݏ���Ξ�[�M"�eaTՔ`h�.ʮ��w6d�{���׹S���|�|*�
 8#��{��d����y?I�9$y�y���1L�UU��US�'���.5a[�<�����&ĉaٗK�{X���y�2�.��#��R�����`�Pt�����V��:ց�/Uk*݂	c��6P\XԆ^u�Y�"�he������n�:W6�e'����B�ڔMLP<��Fy�cՌ�K5ֱ��k�ـvv�u��=1�V{����<�F	G	��^���Y��*�w/U�q�Wd��Z�ͪ�H̄,&XZi�.�{�1s�
��@�����x��cB�E�jӠwo@���,f�0�����Ikt6N����6m� >�/ �[�ً?���ɱ������YTt��UN {����6VǇ�s����X��:�p�SLw�j꛻�elx۳�n�M�O^�/x�` ���x۳���zg��;'� �[�}7z�F��4��`����--�m�[x--�9�+p<XQXY�����͕&���lۆ }�/ �[��ŀ}�m��`˜�n3��$�9��*Ȩ P�D�	����s��W�<�߱`6្�8�g����vZ�t7t����<��f,f�0��x�[a:-]�U@���.*�{�V�޿� }�/�Nz���y6�n�e�*��wk ٷ �v^��<�ً ��l�;-���]=�F9���ǃ�ɨ�����p&a�m�v�gg!������$��t��UN ��� ��c�>ݘ��s�����`�7��SM��R���� �[~��l�ŀOK�n��5�N� ��x���ԓ��{5>r����� #O+�Z���8��z�xޯG�D�͍ڻUeU]v����9�*��}����^��<�ً �v��J�t�'I��0��x�s�O\����X͸`uk�P�E�0��j�qt�㔊�ЗM�όM�ʆ��
�J������K����k�4v�O<�ً ٷ�+ �V�N4*t]��U!ݼ�ً ٷ�+ �[�6�w@��*��wk ٷ�+.$��O<�{;��,��t��9N��y<���~ܒs�ﮤ��;�RaO���W��/���wy�^B�}=�\@mq��I��%�bs�ﮓq,K�{��f�q,K���צ�q,K��{�듻�^B��李�u�m�h����b�!u��g��Z�<3l�6t͒�p۫�2�m��r�rwy�^B�~��٤�Kı=�k�I��%�b}����n%�bX��{��Kı<o�o�n�0(,듻�^B���{^�M���LD�9�{�4��bX�'�g߮�q,K�����&�6%�b}��_cs��!�g3I��%�b}����n%�bX��{��K��19�~٤�Kı?w��M&�!y�^O��uK��k�4u��Kı=���I��%�b}��f�q,K��=�M&�X�%��;�cI��^B�����>%�Ջ�
uɸ�%�b}��f�q,K���צ�q,K��ﱤ�Kı;���I��%�bh0�J��{����s�9 ��m%mlһ.��-P�U�2O-\�pnVZ��V��&��r��+k;���3�˓<�%��,Нt�n��a}��mUpq�nmY�1A[����D������v裪yem@�	:��e��H�$8u��ݫ[Z �������ƕ��]��u�%F���Ŵ��b�I���I�4�'"�;�m�}vN� ,�9����I.���'9�N��w[h��%�n�s�9�8���5�VI�=��ƭ�-�lnD�]mB�g@�)j�Qg��T�,K�k�I��%�b}�w��n%�bX��{��Kı;��f�s����/'�zK>��P�p췮N�X�%��=�cI�����b{����Kı=�~٤�Kı>��듻���My�}����G\g8�n%�bX��}��7ı,N�٤�Kı>���Kı>ǻ�i7ı,Nbzy/���%�����n%�bX�w�٤�Kı>���Kı/{�gI��%��f"{=��Mı,K�;g����31�f������n%�bX��u��Kı/{�gI��%�bw����Kı>���I��%�b{;|�ɜf�w�N���nx��E���R�{���ݶ��cGlP.xZ;<Xhiv����/!y��ﳤ�Kı;�{��n%�bX�{�٤�Kı9���I��%�o'�Ϻ��j�Q�%r����/!y��=�i7
"y�bb%����4��bX�'=�zi7ı,K����;���/!y?y>�k�!1�ջ\��7ı,Os�٤�Kı9���I��?�������:Mı,K�����n%�bX�=���8-��rb\��n%�`؜�u��Kı/��gI��%�bw����Kı=�{f�q,K��ݤ=�S�Ͱ�qsq��&�X�%�}��:Mı,K}����'�,K���߶i7ı,N{���n%�bX���}���%.d�͓���F{{;j�5��[���r��;k��8{��������ڹz�����bw����Kı>���I��%�bs�צ���&"X�%���:M������_���J��1Q�듻�D�,O��l�n%�bX��u��Kı/{�gI��%�bw����Ky�^O&�ۦ�f��ι;��%�bs�צ�q,KĽ�}�&�X�2Z���bX�`�
~z E��M����wMı,K�w��&�X�%��{M��˜��1���&�X��{��:Mı,K�罍&�X�%����Mı,K���8�8���&qz/`�Uv�wM�s8�t��bX�'q�{Mı,K�{�4��bX�'=�zi7ı,K$���8���.����*�-�j�ݫ���p]���g�;r�%�ԛ)����iηS�n�)6Qٛ\�듻�^B�>���I��%�bs�ﮓq,KĽ�}�&�X�%��9�cI��%�/'�ﾁ;��T4X]��N�!y
�'9���7ı,K����n%�bX�c��4��bX�%���t��bY�^O�zK>��P�p�'\��B�,K����n%�bX�c��4��`ؖ%���t��bX�'9���7ķ������}SXͣ�r����/!?$D�{��4��bX�%��߳��Kı9���I��%��z$]��V&���:Mı,K�C��|f�ɋ�3q��I��%�b_��gI��%�bs�ﮓq,KĽ�}�&�X�%��9�cI��%�b~�ߧ�rH0�qu[����� !�/E���(��[v�~_}���-&KKc�ۦfn�0"e����bX�'���ˤ�Kı/;�gI��%�b}�{��n%�bX�����n0���/'�2��Y�4�ru���,K��t��bX�'9�z�7ı,K�}��7ı,Ns>��n'���&�������R�i���+��N�X�%������Kı/�����K�,Ns>��n%�bX��ﳤ�������z��i3�9�EN�n%�bX�����n%�bX��}��Kı/;�gI��%��&"w����7ı,N��~-7npb�ۃ9,��t��bX�'9�z�7ı,K����n%�bX��}��Kı��~�듻�^B�����~�ʭ��[@v�O�o�O�i/L�+f�m��J ��C�Ϊ�59����ug��5=��u�cR M�kBf.ݮ`�bhLE�ck�l�p�M(%3d &��Lֶ�JT�nWRh��W	,VRn�X�U�X�}�7��\�ց�����J+���� 1M��ck�p��܁G�/���o��aFe�Է����rrgѴm�f0��M2?�s��ܑ���;��hV$5S'j.s��u�ֹxS�7T�<�b{s�%�w�s-ĭl&Z���*u���/!y����{:Mı,K�{��n%�bX�����n%�bX��{��Kı=�_g�mW`��&r����/!y��=��7�q,K�~��&�X�%���߮�q,Kļ�}�&�6%�bw��_�2b�˛��7ı,K�}��7ı,Ns=��n%�bX��ﳤ�Kı>罽&�X�%��x_n.�f�&^�;���/��䡈�����Mı,K����&�X�%��{��n%�bX�����n%�c��́~�ۋ4Ɣ�޹;���/%�y�{:Mı,K�����Kı/;�gI��%�bs�צ�q,K�C�?v}y�
���bi�e6�x�K�\���8��lvm��T�<�^%䗦�7a֋�ݲ�����8�}���q�;�^��	�ܦ�z%�b^w�Γq-�/!y=����]fɳ�'w��bX������:����B"����@�*i�Mı;�k�I��%�b_w�Γq,K��3�]3��^B�����N����n%�bX����Kı/;�gI��%�bs����q,Kļ���rwy�^B�~��_�v-B�Å�Mı,K���t��bX�'9�z�7ı,K����7ı,Ns��듻�^B�����}���lM�g9�n%�bX��}��Kı>���I��%�bs�צ�q,KĽ�|����/!y��O~"�hfUq*���;����=�n��^NN���Un��g}���;���&nd�\��O�X�%�����I��%�bs�צ�q,KĽ�}�&�X�%��g޺Mı,K�9gpR�nڈ���'w����/'�}�פ�Kı/y�gI��%�bs�ﮓq,K�����&�X�%��d-��k�1q�q.s4��bX�%�;��7ı,Ns=��n%���t^�}�&� �l<B�>$��a(�?&����)�B"k�2#��&�@����Z�D�� �҅w�h���=��p9�B N0�$��j\9	�21G�M�!�e$Y\�;��$A��
�.!	������HiR@֤��E��P��?K�k�u5
��d�*�2�t�`�b%(P���� d�R�M�KR�vg&Љ+��G �@�ZX�J2�#�Va�p��Ʀ�R���.�ϒ,�eK�ܐO��Ô�X�|�??�JE�� gr1Wy���	���w����@��B2�Je�f.p�W[�hM� 0���D�F|�<D��6(db��J��@�U (*jN'UL�hDr�u��-!��;���4��bX�'$�����&q3�ڽ�=T]�v]6���9�n%�g� b'{�~�Mı,K���f�q,K���צ�q,K�31���t��bX�'�~Է��4V%�ru���/!y���~�u���bX�'���4��bX�%�;��7ı,Ns=��n%�bX��x�2Р��H��"peELB�P��=�Ry���t���:l��kc�����-�{�[�bX�'���4��bX�%�;��7ı,Ns=��~T},K�����'w����/'�|K�{��j.g3I��%�b^�Γq,K��3�]&�X�%����Mı,K�{��\��O��1ɯ!y<���E6؛��s��Kı;����n%�bX�{�٤�Kı>���Kı/y�gI��%�bw��_%̖�˜g7I��%�b}��f�q,K���צ�q,KĽ�}�&�X���j��0��W��� �0 ���%�@�0&)! ZU��#�?�M�&�w\�Mı,K�9|����UC*�U����g8����x�n%�bX��ﳤ�Kı9���I��%�b}��f�q,K��'Fv��R����M�ԣ�CB�䍋^4�;s�î�6K{EWTݤ�Nz�pf�O[)�\�m>�bX�%�}�:Mı,K��}t��bX�'��h?(�蘉bX���~�Mı,K�Oƥ��3�ٛ�[sfq��7ı,Nc��4���Qc���bs��l�n%�bX���~�Mı,K���t��� LT�Kǟ�ԛEa�\�w\��B����{��&�X�%��=�M&�X�%�{��:Mı,K��}�&�X�%�ý���cl�pc8s�d�n%�bX�s���n%�bX��ﳤ�Kı9�w��n%�bX�{�٤�Kı9ޒ�{��j.-듻�^B�����t��bX�'1��Mı,K��i7ı,O��zi7ı,L��(�(� ������s��9�j�UR��孡��Zv��{q¼�m ��:nŮs����N._`����=�V]�a�K&�m���f��pâ��y�8%�4hs�w51�0�u�2����l�U��Xݵmi�H��c���Vᎄ⺤�;Ef3�qŝ%��v�79̻Lk)
W +���r��Ɗ��x�CWW��ke��@gR���Rcs�NrM�]��"�YC�i9tB���ÔW5$5��,!�� 4ĳ%q5�	\5�bl�9}�����b{��i7ı,N{�٤�Kı>���Kı/y�gI��%�bw��_f[s%����8�n%�bX��}�I��%�b}�k�I��%�b^��Γq,K��9�cI���^My��ޟm,7����ٝrwy
�%������Kı/y�gI��?�a����w߱��Kı;�߶i;���/!y=��/�'���'\�ı,K���t��bX�'q��Mı,K��i7ı,O����7y�^B�}��uO���U^�;�bX�'q��Mı,K��i7ı,O����7ı,K�{��n�����>�}�n���4v3P����%Ŭ
@۶�2�\v�N�N,z�	��l�e��'w����/'�{�s��Kı>�{��Kı/y�gI��%�b^�Γq,K���B[{l�S;��듻�^B���Ͽ&�� �#1���U6�q,K����7ı,K�;��7ı,N{�٤�Kı9��z�a6eB.��'w����/!�|�7ı,K�w��n%�bX��}�I��%�b}���I��%�b}�N�a��͢e^�;���/!y|��I��%�bs���&�X�%����]&�X�%�{�{:Mı,K���Y�hb�W�N�!y�^O>���q,K���ﮓq,KĽ罝&�X�%�{��:Mı,K�);�~�!Q�6i�����l+��@2�B�Ɩ���a��cObl�u
�Ḳ����2m>�bX�'?g߮�q,KĽ罝&�X�%�{��:Mı,K��i7ı,N��Y�f����8��n%�bX������Kı/y�gI��%�bs���&�X�%����]&�X�%��5/��6f���g9Γq,KĽ�}�&�X�%��w�4��c>
E�*�("���M{?z�7ı,K�{��n%���/'�ߺ����l�ʯ\��Kı9��f�q,K���ﮓq,KĽ罝&�X�%�{��:Mı,K����cl���p�ɤ�Kı>�{��Kİ��G����}ı,K���t��bX�'=�l�'w����/'���W�h�\	).m�f�Jr�֩ l:k.a�m�^�v�vI���:���mԫ��u���/!y�{�Γq,KĽ�}�&�X�%����Mı,K�g��Mı,K�z{>Ç4f�3��N�!y�^C�;��7ı,O��l�n%�bX�{=��n%�bX��ﳤ�Kı9�>��4�Ţ�\��B�������4��bX�'��}t��bX�%�{��7ı,K�w��n%�bX�1����}�B��rwy�^B�~�ﮓq,KĽ�}�&�X�%�{��:Mı,�,Q,�Q���M(�����{\4��!y�^O}��b��::��v��ı,K���t��bX���=�~Γ�%�bs���4��bX�'��}t��bX�'��|z��Ĥ����/B��-�����/<3f�ax�f�W��5���H�ь�n��A���'��^B�/����n%�bX�{�٤�Kı>���Ϣb%�b_{߳��K����}����a�c*�rwy�ı>���I��%�b}�k�I��%�b^��Γq,Kļ�}�&�~E����'O~�JI7�JS8�sq�I��%�bs���i7ı,K����n%�bX��ﳤ�Kı9�{g\��B����{�/׳��җ��Mı,�(��L{߿gI��%�b^�߳��Kı9�{f�q,K���צ�q,K��=:{8�9�ܸ����9�n%�bX��ﳤ�Kı9�{f�q,K���צ�q,KĽ�}�&�X�%���������\Yw� q��26����{7*����y�v���z.��e[G`���M����U[�G'��D�㱭dՋ�2�-c&#���i�K�`��ڞw�8�6���0��,m�͌%94�' ;��xg����s�40P68�3ZZ�Rf��{Xx&΢�am��2bs���й�����V�2�����d����u�b�2�8�s����D<�xC�9'';�s�߫Fۦ�֎*^0e�&�t,dM�-ٸ���5��`��DEeZ�	�IS6\�n,�9�z��bX�'~��I��%�b}�k�I��%�b^��Γq,Kļ�}�&�X�%��^�.<g.1�q�I��%�b}�k�I��%�b^��Γq,Kļ�}�&�X�%��{�4��bX�'y���̎��pf�޹;���/!y}��N�X�%�y��:Mı�D�N���f�q,K��k��n%�bX��g��]*8���rwy�^B�y�Γq,K���Mı,K�w^�Mı,K���t��bX�'��|@���ʯ\��B����}�ݚMı,K�w^�Mı,K���t��bX�%�;��7ı,O�������U��T|!��m5�q�����ř���8�[bW��6�iP���%�l���ɴ�%�bX���~�Mı,K���t��bX�%�;��?
Ϣb%�bw���4��bX�'}�O�u��m�,��f3���Kı/{�gI�x4*C�ρ����D�/��gI��%�bw���&�X�%����M&�X������}��b&U듻�^%�{��:Mı,K���i7ı,O��zi7ı,K����n%�/!y=�}�d>�F�Ţ�\��B�,N{�٤�Kı>���Kı/{�gI��%�b_��gI��0����7��K�t�B��rwy�ı>�u��Kı/{�gI��%�b_��gI��%�bs���&�X��������\�2�,GBm.zõ%�.k�f��r�(2�ha�8%�KKnfp-���8�9�34��bX�%�{��7ı,K�;��7ı,O��l�n%�bX�s���n%�bX��}e��T�⺹z�������?y��\��B%�b}�{f�q,K���צ�q,KĽ�}�&�X�%�ӹ�e�L����3��I��%�b}�{f�q,K���צ�q,p�BU�
_D�%Ϲ�t��bX�%�}��7ı,N��I&�e���3q�I��%�b}���I��%�b^��Γq,KĿs�Γq,K�����&�X�%��v��t��2[1s�\�i7ı,K�{��7ı,K�;��7ı,O��l�n%�bX�s���n%�bX��y����f�IJ��6KsuCe��gmF�X�eu�Z�:��`�X�N\�Z�&[8������[�d�,K���t��bX�'��i7ı,O��zi7ı,K�{��7�B���gޖC�hSA�����*X�'��i7�G1��}��I��%�b^{߳��Kı9�w��n������ov�}�5�`�3:��%�bX�s���n%�bX��w��n%�bX��ﳤ�Kı>�}�I��^B���>�_��GS8f�ɸ�%����w߳��Kı/{���n%�bX�{�٤�K��p Ґ� ��H)��'�SX��g煉q,K��s�,��-b:�^�;���/!y|��N�X�%��w��n%�bX�{���n%�bX������Kı:w�ܒ\��9��ݛ��ڶ�;M�0��WK�l\-\Rg:�����U��Kı9��zMı,K�{^�Mı,K���t�I�LD�,K���t��bX�'{���ce�3�a�c:Mı,K�{^�M��q,K����&�X�%�{�~Γq,K����7򘩈�'}�C��s���9��f�q,Kľ����n%�bX��ﳤ�Kı9��zMı,K��i7ı,O���ع��3,�qL�gΓq,KĿ{�Γq,K�������bX�'y�l�n%�bX��ﳤ�Kı9�w�ǋne��9�t��bX�'�﷤�Kİ�~J���|hI�=�~�j	 ���В	"_�"*��*��DUj "��_���� "�� C�袊DA" �E�*�"� *�"Ȃ�� �� �H��A�*�"ŀ* �H����Q_�"*��U� "�Q]�����DU� "���_����@EW��_�_�1AY&SY������ـpP��3'� ax? 
  (      (�   P ـ ��
�x   ��UT�"�*� ��@�R Q@R��UR��
U ����
�RR�EB�      *�  �6 �|.N��,�-9e���,�� t��'B�U� ՝����P{�=�J!�  
� : 
      �    
 �     M�s:�q5JU��:� ^�Jҷ����� bu@�,��  x8      �� ΩT���AB�.�A���)ӝ�*�p �����Ƕ.���sh��� 4��n��R������Ǻ�{����|S��/T���o�/=΅˹f�� <��\c�d�ֱ��^�ϷUW� �|    P  ��U��ښ��cӽ��}3�*������N��w��6\۷�v����6鯾|P>��R�o������ y׏�n�ϯg�>�=��\v��.����wy�t�� c�ۓ���^�ŕ�w<��� ��@ P   V;� �ۛ�Ʈm���׼��&�{� ��������{�zWq��[�P;��\w|�t�k�/v��.�[y�����Uq����ĸ����������P4w���¦\��<��[�v�o |   �   �� ��|������>Zyyy5��Ƕ�� {ޓs�cN]�嗓O[�}��zW\w}�����  /O-�=�������Oyzn.�=O&�=�z^^��� }���-*�c�[�o;�z�x ��̔��F�S�H��R�� �<z�TOT@  Ob�R<�R4  ?BSd�� RԔ� ��t�����O�O�������	Oe�{=���{��PU�f���@AAW`�
*� ���`AAW�YAENw��?ю���/����0��тh7)�:L�&B��D��M&�7������4����y��ly��TGk��A�xgņ�0�a$h��P�R�a�a�4Z��Q4DP�&�82�F0Ł8N:e$�#I;P�a�f{o8i�U�Zx�{�o6�S]���?$}��
-&��7�<�y���@c�1##D�a��5�s���3��\���h�,���WG���8A�0K�j�Ra�qu����pvn0�����p7��4N�+4��F�b;�ہ�
|��Id� pB>���L�ZI!�I.�6a���1u�����g C�F����'L��[H�B�0��@�JC$��R�F$HPI$cf��߿}�8�&a����u��4}�|l4]��VkC�J�g[Af������2�0��o^l�Ca�����1PDs[ٛ�e�ă	q�2��t�(�ێ�u�Zc�κ��Li�(*J���h~q+�>u��˶��x�j����XLρ�UĐ�J���l�<��Y�U���1��������k�h���7���8��r4��4F�E��(��N�f�&k~��kE�j0,�0Y��:J��_p�_<��ic�k�^����=|���f�֩ޝa�z�� ���p!�'\��3��k�Yd��hޏ<q�,���ya��8Fp7����<�\H��SǄZwPi�4C�h�X�F�<	�����j��i>��M�p� +,��@f���Tç��z`h	�4�a�ֽ�g�٣�ְ��q5��ލ��>)8��.�&�'!0ߧ�e�<F(6m�)�m����$�jX�n5����Z��y���R��"I�;6�8Q�����M��[�3z:��fq�&$�$����v{�y�{��sO��8:xx٣o)��y��ow��<>X�X�14���M+8F1��X!'���'t\�6�!$"8�<<�CN��2�[c�9�k��3�p�z����NL٤�wRճ�F3Z���4j��sz��ȹ:7h9Î���#V{����
����9����&��$M$�V�Q{�㎻�>��DM���!Y��������A;sV�6q�@r�E����2����1��v�w��8q�9���ױ�6F���l����-uG�=
$����.I|���40�@a�{g���d�u���Ը��ي�N�QX�+�`��e����~<��?n0l���La$��$��& ��&=�v�1�֮�k_ZY
8�N͘�ŗJ��1�A�M{�쵳A�����X�fi�M,C��<9͇I���G[�QrCD7\|>��HR���Y�����v����;�1(YJEQ0����8�e�e�x����8��:�����R<�@���L�I��z��}��ϓ�Ϸ�$�|�C�l��_0Ѱ�����^1i�&C�pbh���g���v��|0L7��4����s�I���MM�G��Ʌ�6k���A��}�#��s|z���g4�;�2����6FLB�l�Z�5��x�x3�L�`���	h' �a��9�s�{3c���"3&L��ַ�_�1�[�m�f�9�͜��=��Ed�%Td�Y��tPI��y�9�puȕa2�@��v2��r�y�/�^��sv:�5��ѾT�a�a���Pa���	�
"31�����w����q�w:ݯ���G*��5� ��"�̠�m�^��|��3�v��F�N��	pI��H\Hj��#A��6�`�a��]uÜ�,*$�`�67��1��{Dg�؈�F����5��8x������l�vfyK���r'
`d'�1���ƒrH0�H52D�\�h<|:���$�1�2&	f��upČ(�ߏņtݚ�N:�Z���IC
��� &X_��"�`�s ͓�l5����=u�����D�3���텭�X�l��z���e;ʽ���]�������9G�}$�~z�	���y���ӿM��m���aefe��0��K�l�Q���������m\Ձ�q�#H��2p�1��X%��+Q�j�?<Pؑ��F]���9�g6�������;ߙŜц��1�ny������r�f��Ϛ�sRl���Fq�'lp�3[�ǊA	��d����l�[#a�Ʒ���[��ɭ�8I�8f�٭��85�R8'22�#�I���I(�(hvp�3|�:#�ڰa�r0������כ���X�\�ϋ����{�ך,���[1�����v�,ٲRL'9�Ȱ��VS�9��M�f_f�oY�VI�Fk4oϼ��p�~70�he�r(Ƶ%�cl���}阮�l5a�0
��p��5���H�ή�y�^��e3\$���F$F�$s^����Fь0�0�f��if�ⶣ�|P-NH+]P�O�q���b{漰��m���{������ ��t#����fg�3[�4K���ݰ$�����Gʿ2�0>�e JI��PzZ��D��X�	����G�`>�/g��M/�1oa��9���8{�'��g6F)k�0���!ߜÛ�aş\��m�y���>`�2�����'5m)��z8�����7p;V+�4!#mp��L&(Dk�-9�x�`ǁ��%�D8�8E����Nh"6D2�F&����Ѿ34
L�����f�6a�o��,a$�eP��;��|#�c�1�9-�lf��ۜN�&Tf�a�4Fh#`҄�8.�q#� xzo��S��A���` �Y�hL<58� 
c<ms���`q�Ű#3�hC��s��M���Ѡ'��(����b��.xn1�)���������r�.�YJ̜��>��IW��*�NQ�U5�CNa��+#�6�E!5|��?��+�>�J$��R�g�Fy��%��y.���<�$½���+��+5���z!0�%���L��!A����S��>fc���412a�3
`�2Is̸fe֝Z9_9�6�����蹾h��$a�8CY������a�%��c��q�LA���3�� x��q����H`����'���Vy��9�90l�JRA��a&�Se�l���淛��䬂��'g�\���0ס9���S��"4?F�7�i�F��̆ц��I�bFi�����V�x��W�B�.��t�R&�|I�I�3���<+�5^�l_���9�����>��@F$@�i�i36sK���4Î�fr��b�j��H�<���V����3��9T��\�ݧ#�y��g�6h��N#�٣
H2�����$�%�|�)ȟ��vou��3��,Ѽ����TJ������)X�/�)���4Y�0�bc�Ѡ�ż�6x�y��z�}�����#���V�U�n��1}:���r3���$�p#���F�y��l���}�®��v��c�`:��А��	�0���+�i`����q�5�l�Ѹ�6p�Ff�'[,\0��mzl���#��d&����J��8p�K6�vm,�`�f��2ͧ\0Գ�
Z�c�c�oz׾}�Z��Z3~ٳ�9��F\}$�Uɚ]��k^m���v�Fm���(\m���
W�!�??ڸ�q/���*��W�ve�-��'>���н<eVٯz^�~w��${#sG����e/�i�f�Fh#	=�5��N!!��p�#Q�gǬa�LR��G�N��BSV�dԪmmތ�[���ӄ`�kϪ�F�"/#S�A� ������C=]�$7Τ�$�`�!9jG.#�Y1Q4&'7pN>�p���-3p3|<��5���9 �5ߗms�� ��9@��'?@                          m�       �      �              ���            h�  %�                             ��h k�� ���    @H-�                        	   H  lA� ��� -�j��`��6�m��3�ҮC< [m*�V�U���%�BےG�E�����\CV8�`���h�⶞��AJ��ҭU׃�.�:UH����+�U�K���� ��[���m�}U��1[F�A{V�H���Bj� ����n�]
�toQ���V��8�B՗-�m*f��m��q:M�h�l��8ඳn��8�-�t�S�˷0m�`�$��Q/t�[�yU	�UWŭ5gf���}��R�ׯX�v�C���H�UwI�-�]jn1�cX�����q���u��l� ���d�Amd���!�Kع`ݱ"ڃm��� dlq�$S�ۗ���(���i�h:Uj��U���%���7f�YZ�V`���IUfդٶ� ��6�A���H��nם��F�ls�z�~�m���V���J�?Ϥ�ۭ����3����&�kn�Wfٶ� [v�I��j�` m�ז��lm[ �  �ۑ��4��-�@��[A"Z�ꪞYAܛPkcf�ɺٝ�N�ۡ���� ��Uժ��|���kd� �����l.If��\�ն��[�iUV������IKۥK��ltѳi�v�˅�2HE]�mg\��t��q�5oɝ���X��X��d�P�Rmy�c^��#$	�	&�wX�ذ�u��[\:�-��Ev��mV^ۀ�H���A��iU�n�i-6 YE�V�r�&�WUO)v-���w�i�P�/5�>y����{j�h*S$8��Q�3M��Ӝ��zM��TD�ʶN�3&��J&��kI6�h�F9�z�k�n�x�LZmQ@$ 5� m.Y�Ҁeۮ�l��V֍[,�S����5RH4�έ��j�v0���̉���lݶ �@��<�5WOh���j�h�X�Gҭ ��Ug`Ej�`�%��*�ԫZ�I�U�*�v�\$Yi���� q��^�UV�O�/0��vmÖS;�-U�u�m�-�T̎46�GY��k8G6��*��M=g�:z�-�x˝s+�)�+S��6�gI�
���6�	�ۅ.�.�n��J��SiVB s0�DW�UP�Vq��nŘkj�]�8ے.��@6���tݚ�Cd�\-Y��n��̴�"��ڭ�����W��(!���Vl�KװJ�l�i�m؁J+F�nݥ�
�깩N�m� $E����[@JP�.ٶpl�B��n;\�m�,b�2,���va8�jVV���UJ��P-�3m��8 �m���l��X�Kz�d�"�i�۶��d���j�`��m~����h�յ����$[s� �c����aη^��mJw�U���G/X���-)�\. �Mm����-�/M�%�*U6����|��K.�6iKF��� s����n��^�ɦ5J�(� Q��mc�k
��[�I��y�8a��n�oP۶R��t��и�ʪ�檩X9���V��\��M���`����`ۮ9YN�i�\��0]:ۈ^A�l7��T�X%Z�UZ���%��mS�-m6d�2v�4L�㦪���uca	T��UVV�j�P����̴��-� [���7E�kn-��O��k�\I�:GH� ��]�ַ�Ĥ����F�ܐ-�� 8ݶ�G�!��[v� 8i����lm�mo]mZ�� F�{ =!n�s��e�8�ƵAݕj�nY��hH�mN�r��Q-f`�j�_-Yvظ&��; �][g�j�%�bċn�@E.]C�]�˱UU�B��mjկ'�%�c$��Yj^���� m�qml �n�6�6�r��AQ��=U��U#���Q�m�mt�i�[dm�m�86�� ��m�@춁���kl��$ٴH�� �$k�B@q-6�7G��  $$�ku�u��5�Ѷ�n�	$[N�h�  	m�[� $m��UQ��%U%����,����Uڪ�AU��z�5�� ��m��m�ۗ����ml�*�V��pJ�P!+UMf�v[D���m�2�&�L  �  d��]�V�j�&�PƲ\ �m�S�Vݶ ������^�� pt��a���)��I�}��$q,� �Rɛl6�h�ª�jWU�Ca@j���ll	� �ȓ�d eU��*���r�k�e��[a��	6ۀ۰-��$	 ,\�U*���ك���[j�[h�ód�r�-�(��	�jv����\IJ� ��y7n�d(
�j��1T�[T��@��Ѷ��Uyz�^`��+��Ą�m]�9�3N�[I�t�'n�hU�m��gNj����|����7�wj�j�R%�{'-��
T�=ja���\�`�he6T�G�L�*��qW$M]T� �V�@]��Ɉ�mm�	l!���I����m5���D��1�Öݶ 
ڄ�����/Hz�vM�[�� 
���l; � u��F�V�$��l�5�INe�Iyʷ[�)ً���z��D�8	z�tLgo0p$rޤ۩�hm�6� HᲀJ�*g�y��y`B��m� ��h��Q�Ѭ�p�� ݶ m���-I2e�v��3��+`'B	,�m�W�]��u��,rBD��\F��	��6�m� 8HHH    q�m�@�:]���6��[KN6��'�^��yc[AÂ�5�M�l]2�H�I�i�Ӏ m#�j���jU�Yej�X 0���`I����m�۶m6���*��J�����U�u�R��I�Ͷ[mɰm[q�м��F1hb]�9��n��4ݯ�m6�� 5����!�	�m��5YZ���/::�8�6��-���7iٕj���L�f�U���*��j�Y���+
v�w7$�����N)1��iEW@UU�]�I��i��5HMh������R8�D�uIn��u��4���5�� ��Z��f��;_Z��ˬ�Bt8����˕]�nx `*�@j�Nb�	�j�Ur�6�ګq�U�ҙ�A�����P8���Y �c�8��AZ�`�'9q;�z��c,�쭬�Y$��8m�i��gT�zYCn͚M�e8m���������;m�[m��5��r�[����U��GYm��[�<�,�UUl�����eU��Kl� �s�`H 6Y�Z���_��Hh���4P��9�M�K�m+6�md
Z[V�P�uR�S`*y[`�`�ls����ZmKm�-�~�}����[�������2��ST���    �i  �cl����[  :���G��햀X+iPU�d�(���&�8,�X닖�U���UU��(   �Ʀ�5\V�>۰6�0��X`$�],�!�m�Ö�^Z�U�8�ny��c�m�� -��#lIз��:$k�ԛ�#  �[%�I��[  -�m�N��m�N;Z�>����f۳m�B� ���/Y,� k��PH-��P�j����U/ 0m3d�d�[�9�m���ޞYeeV�j�����ﾓ�[M�f��8� �� m�-�;e��N����@�Z�-���[rͶ�	�I'4P  �E����� ���'�`�� -� �'@ ^�f�[Km6�B@qn�m�� �[%� ��:@s��%�l�I�z� ٫` ��v,��M��Ç[R�r�WC/gث`$q�-6���L��6���;J�R\t���v4�`S���'n^���q���Y�̈́�	���ۈسi��nԑ��s�F^�Jp/-�\b�Q�P<d�`� $	:�b@�G �!���UW[i	�-�a�
� �����   ������J5��[Nkղm� 6��Ko�md��UUU+Fv�g���v�m��5� ��¦�]�^Ɖ�t��t���H^3ݴ�<:�|}\}e�㊠��ZS�l[v�.�$�T�6[@U�Ų�xa��;����@̆�m� [@ m��p-�mt-��H  "M���'!�l��@�-)�m����5J���`�nom��!�m�nĀ ��JCe��kYb�γ�ֳ��� �0�m���$��ǻ��w{��{���P,�'��> *�&�O��0�?�C�T�"�*����z�1!��<}@�D<(&�x@����:h� {�TODM �5�� O�@�<W�P<|@��pzB����^��BH2�>�S�z��(����0o�|U:+�6�22��!�<6z��LW}�� mDN��,*> ��]����1��@�}T��~T��/UҀ���+�;=T`OR�"iN�����Y,$��tF�1I>O��P�N� � ��|�!k`b���H�� �N��O|A���@
z��;�LUsϔD��:�(b��'P< ����<z"`"t`�A�U=P:���0�\Y�� p<D����T=OP8 � T��.Հ>bt�i�b2�C'2���1^�A ���!��x��+�	�WM�"(i6�m>E�F%�^��]���]��}<�E��!0�+!,�J'��,
$,�#�C@�
�� >�D~�v `!�A b��_�_6(�+��}Q�p�J � H���\AWL�0�$���
�d �S ���t�w^�������o��    6�n��  �  [@     �]� $ݖ�   �k�ķE���MXէ�����Ŝ]R�X����i�)X�O�9嗎��v�:["6�<���K�)���6;sCn�^�f��d�*�cGu����鋠�&ډ)�d`T�"^:�,���+��pܓa'�	J�i�{�:kM*pgaF�k�ݛB���Qk�w�f�Zb�TNt���l�ź3�2�]L�=�X�o6�:R�1[�\dװ�Nr�{N'P;O#@����nnv��.x������pr�n;C�6��3���U�*�$��=�	�'��$N��l8h�p:v;V�ݭ�v�:,��yn��a�v�K{Y�z"c�2�9�%n��e�ɹ�n:�d^r�M��s��N�JŽ��	4U�cGUX�m��^��"�n�e�i;!7,�r�8���6�oi���R��
��Q�،�ʁ���1��#��+I��p����dW`������rh�H���r*�mU{�1OZTz9 �'GMNHAœq�Pn%A�1�&�nD㎺�sǖ�pڱ�j�I�v�����b�oSY�2J�a�s�u��^�z�|qN���zz8��]���m>�c�Z]�8�VYZ��4eeL�m̓�ƶ�RS1��$�C�i,�]�r�WX�U�v܎�w��a�rr�W�b�qrgOn{���ˣ�v��l�m�(���V��ŭ��δ���ն�:삗m��Z��A��n	�{vv7MaRΰ�$��U��Az�mV��^�)[�̩/M�RI�g�ϫd6⨠��I��{f��%��]Ek������� gj��Cn�d�H�.wh�K��� ��v��шخ݊�<�]�r�et)$l��S̵�U��L�MX�9��]�	=F��	M��F4Z�:����0�f4���3�c�I=X
a{kZ�_ퟀ����bP�	Y���(����h@v �x�&������| �/�����_��5������@a�L�ێ�'�h΍ѮN`�k��ɒ�]md��s��@]M�G�M�R����O`���KS�0��՞����i�������S���5ǵ��vy��ك�{m�Q>Xq�"��l���0��5��9dS
�ñ֝Î{%��^�I��u��Y7Tl:�{Xk]e�od�b0�{�ǽ��{������m��(����1����g܋���dy�\�wg�l/+�����P�ݺ�;ܕ �ɇ�s�_ ��v��~��*e�'@��j��ffڿB�M�����|y���V�ѭ��GV$��� ���K`wtt�����
+�%/
V,���Ж��������d�IP2��J��-���������0=�V�ܮR���H�EL (���l���$���^��nԒ�͊.�Ӭɺ�V�@8�P�Jd�NHQ$����]Xn�,���`ff�X�mk5&�)Jq���`}�X^�jh��P64%�k8ͩ��l{v���ݺ�
�w]k"R&�9p�;�V�36��W������Ł�LZS5H�	8�#�33n��2Ձ�eaa��9�́���Y�j�^e,
̻̯$���d�$�fmՁ�����:�Y�4��Ӧ$�`��i��'j9'+�[�0�{;:.h
@�ў�L��2"��nW�wޞ,������遽��������(Ax�x0=��wGL� �����3v��DA$I�(C����]X����H�E%d��@,J��LuH�	� �RE4���T�(l5}$�����v����%2T'$(�U�����d]R[����cMrTmFSnU������en�36���n�X��^��L�ԕ)0R���E�N��حq���G�f�� Q�m+���ɺ��H��*r6�����`ff�X�:`zL�J�B�����3�u�����遽#���07�GL���Xz�&���nJ���Ձ����(M��36Հp�d̬�D���%w������t�������:�ZF��ԡ���J�o}�X�:�.���*GL�0=&A����_�o�[�r��:�aX�ш�6wn�888��0�6.���OY�y������[�^ex	'Θ�0=&A��05wkc�u	P���IVs6���vi`}��u`ff�X�mc56�)�FS��`zL��R:g�U��RO�0:O�Xv����G"J�#p��9�]���U�����R������)>���<��;�Wt�����-��f��g�)=����R������)>�;�JR�}w�8�)K�@~�lt��`���=�w��{76́a��2lu�NN�����e��m�:�4��y����7h��.M����X���4��#i�4��*\��X����ժ����}}�]o:�7B�!�e���ݞ��ې����ꍌucm���N�	����e���n��$d��19�]Q��z'��r�l3.��V'C�!:��q>��8.q���s�%$!6O�WL�e�*S��IV�o���;.n'q��Z7]X��V���h�
�'�NEAv�e�' ��j�8D �[�z��*R��s���)��{ÊR�����y)J^�.�Z;��[�ՙ���)JR}�w�<��	�����8�)I�����R��߻ÊR��w3��˺���ox�kzJR��}�R���ﻵ�)�w��)<���y)Jw�˼+f�oVn�og���'{��^JR����8�)I���C�JS�o�ÊR�����ӽ�n۽Ž�y)Jy����)JO.��JR��}�R���ﻵ�)��������Y�k -%�����j�Żu@m�2�����&��=��n�t���u�-kg�R��߿~��R�����┥'�}ݏ�To%)O~��R�s+<�zD� !�7r�r����������C�K?'�m��I »�4l�G��ͦ����)��C��)9����)�~�ÊR��]�t<��3)�
�I!(���I*��r����a�)�w��)=���y)Js�r�� �A�碢��RU' ���p�)_��	�xqJR�����%)O}��)JR}�u�y)J^،��������Ҹ�!scQr����w��)>���<��<��q"B�,o&�Ni6�Ĳ����m���x1����m����bg���5�G�5���b��qeox٭��R�����┥'�w]�������R�������R����xV�ެ�Z��)JR}�u�y�C%=���qJR�����%)O}��)JRv�:wN�ճv�m����JS�~�)JR{��py!�"f:��xnS5w�8�)I���a�)yv��gr�l̵�-kg�)=�w�<��=���8�)I���a�)�w��A��JyT�u@ɩ�4�Y�!s����)JO��%)O=��8�(��1��!B��S�T�T�S�@R��q���t@�V�'��˱<�kY�t�^wA��c!�R�)6�%_9A�Pr�5�<��<���┥'�������;��!B]�5��ʒ�9U55����w��$�'߳��JR�}w�)JR}�u�y)J{�.���F�n�ֵ��R�������R�����┥'�w]�������R�����f�.�[�U��f���J��}���R���k�<��<����&H���R{��py)Jw1#n��TM(�����(9Y��JP�'߻�ÊR��~�߰y*���W�!.��njDʙnJ���n�}�tZ�{�Sf�v.�g�������Pڐ|���BS�i¹g9A�W�ͺ�%)I۽����w��);���R���Gڌ�f�ڵ��R�����C���!��}w�)JR~��_��)�w��)|>�������Z�Z��<��=���8�)I��]�������R���{ݏ.r����)�zG!�JM�IW�Ps�I��]�������R�����C�JS�o�ÊR�������h͛ٚ�{���|��=���qJR��{�%)O}��)JRw��a�)��O�1P���9��f���Z����# �n��?��y�i��g���a��ױ�ͻ9l����%�֭�gGV��9�:�7
m���t�(�i�R[��ʙL^W�������)��5c(�����Yˡ֌�u��QTsmԓ�ece#n]�[n��nL�\k%��] ��IC�cŝV��-h2�z}�5'��G8N.F����z;a�I�3�;��];�����6�s6p�o�z��p�v�V��4�b݉�ܸ�k�]�g�V�z'/8ζ5���"�������Ȅ!x���������┥'{�vJR�{�x�!B\���s�JIe
���BR���w��);���R���ÊR�����y)Jw�.��o7���og�);���R���ÊS�@d��߿hy)J}�s�)JR}{�;�yZ�n٭��nJR�}�xqJR��{�%)O}�;ÊR���u�y)J^G^���jنkv�kg�);w���R��3����R������C�JSϾ�)JRw���lE�:�q=�.*����z�f�Ξ��c)������sv<\�L0f��ַ��)�gxqJR���%)O>��8�\���~��C�J�Y�YS:L��I��:�q"B˽�zk���Х7��ÊR���;�JR���w��)>���V��UI�*���G�B���iq�����R��gxqJR��ﻡ�)�t����T�۫-k{��)I�s���)�~��┥'��wC�JS�~�n)JR{�ϳEfk]ޣ2�kz��y)Jw߳�8�)I�����R��߷ۊR��w;�JR���������6x����]L\EN��&ǫ���Ysҙ��-����&�6Ʈ�.���Y��)JRv�hy)J{����)JO;��%)N��w��)=��;�yZ�n٭��oC�JS�~�n�@'%)=���`�R���s�)JB�s�J,��
�G��l���Ӛ�Y��R������y)Jw߳�8�'3��e�	��c�y�<C@Ĕ�h�C�9��jb	`�??��?:x�F>���kI`��ޏ<S�����]��b�N{�H��u��onq��kIR��kH:њ�wl�b����n�jM�~A|�y�Mԇ�a
F*~��fl8����"�_���>xQ0��pq'!� �j4ʸ~����u+��t<v(@!�+����'�/��q<R&R0X�� X�L�_�A�L+Y�a8�srV<>��6������xy�e�hM_Ys���1JO-�;�D��"&[ 0�`�H�����s`wB~qP8�!�	����1P���] z*D �|(	�D�
�H_(!�T4 b��h`�����R���n)JR�w��o5�3[,�oy�nJR����8�)I��wc�JS�u���?"!d����E�"u*v�f��H�R�UJ�
R�Ͼ�ǒ�����)JRy���<��<���8��J��(L���(J!(J��30J��(O�������z��l��`�]v�t�̶nϮ�[�c�]�Y�a䃋��e�d�8ꓛ�w�N�I�BP��	BP�%	�%	BP��%	BP�$BP�%	B}��g�	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP������(J��(J��"��(J3�(J��J��(O~�����(J?���H��(J��`�%	BP�	BP�%	��P�%	B}���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	D P�B��=31�HTH�ji��	(J��J��(L���(J!(J��30J��(O{���	BP�%	�`��"ː�%	�%	BP����(J!(J��>������(J��J��(L���(J!(J��30J��(O�~���(J��<���(J!(J��30J��(H��(J������x%	BP�$BP�%	A���X%	BP�$BP�%	B6� P�B-�z�s>�#e���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'����x%	BP�$BP�%	Bf`�%	BP�	BP�%	��P�%	B{����(J��<���(J!(J��30J��(H��(J�����<�J��(H��(J���(J��"��(J3�(J�����8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	BP��v��ްѭ���7Z����(J��"��(J3�(J��J��(L���(J���	BP�%	�`�%	BP�	BP�%	��P�%	BD%	BP�'�����P�%	BD%	BP�&f	BP�%	�%	BP��%	BP�'��a�(J��<���(J!(J��30J��%P�_>�$��� d�`0�$�0BXY?�����(J����吏	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	�~�k����f�٬��P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP���g�	BP�%	BP�%	Bf`�%	BP�%	BP�&f	HJ�*���؃�4>���À�@�B�}݈<����;�r���'��F��,�c�x���h�]���қ7;gV������]�͝1���(J��(J��30J��(J��(J3�(J�������%	BP�f	BP�%	BP�%	Bf`�%	BP�%	BP�'�w?xy��%	BP�%	BP�&f	BP�%	BP�%	Bf`�%	BP�����(J��<���(J��(J���(J��(J��(O{�߳��(J��(J��30J��(J��(J3�(J!qnJ{T�&�\�74�B*��0J��(J��(J3�(J��(J��=������(J��(J��30J��(J��(J3�(J�����	BP�%	�`�%	BP�%	BP�&f	BP�%	BP�%	B{����x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'��g�(J��0J��(J��(J3�(J��(J��;�v�j����l��Y�����(J��(J��(L���(J��(J���(J��=�s�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP���g�	BP�%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	�u���(J��<���(J��(J���(J��(J��(O~�~���(J��(J��(L���(J��(J���(J��>�����Yl���ַ��J��(O3�(J��(J��30J��(J��(J������(J��(J��(L���(J��(J���(J��=��8%	BP�'��P�%	BP�%	BP��%	BP�%	BP�%	����x%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�'���pJ��(O3�(J��(J��30J��(J�@��
N�ff6@R9��|���(J��(J���(J��(J��(L���(J�뿳�P�%	By�%	BP�%	BP�%	��P�%	BP�%	BP������P�%	BP�%	BP��%	BP�%	BP�%	��P�%	B{����(J��0J��(J��(J3�(J��(J��=��~�<��(J��(J���(J��(J��(L���(HP�b����@�RNmU*�������v��s�����u��6��n�g86�0��������jѮ��&�+m���qp<��":Ж��9��ӳ6�a�^vM=O6�/��� Z���Q�c`��8[��!nZ�݇�� =�qi�y�+ٸ�'���q8�X{�ݐ�ۣ$�W@;��\��	�����7b6��F��x��+��U�� ��Lk��S����w���duP�t`��tz��[�x�c�3��0\mr�wc�]Z2���ЪY��nj�kZ���%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B{��xy��%	BP�	BP�%	��P�%	BD%	BP�&f	BP�%	�{���(J��0J��(H��(J���(J��"��(J������(J��"��(J3�(J��J��(L���(J�뿰��%	BP�f	BP�%	�%	BP��%	BP�$BP�%	B~�����z�F��7��k7���(J��J��(L���(J!(J��30J��(O{��8%	BP�'��P�%	BD%	BP�&f	BP�%	�%	HR���g�	BP�%	�%	BP��%	BP�$BP�%	Bf`�%	BP��]���(J��0J��(H��(J���(J��"��(J߻��<�J��(H��(J���(J��"��(J3�(J��?t���7���5�Y���(J��<���(J!(J��30J��(H��(J�����<�J��(H��(J���(J��"��(J3�(J�����8%	BP�'��P�%	BD%	I�I��&��(J��J��(O��?�<�J��]��(�!B8-��=RR*�*k8�)I���py)Jy���R���ﻱ�)���s�R���Fw[�o2��Y��3[��)�gxqJR���{�c�)�u��qJR�ϳ���^������W�h�N:��v��+r)��̮f�;�.�r8$&��s���v���原��j�l���f�{<R�������)���s�R��}�w�U�s�JS���W�!,����n����Qr���k���AM+�
�Qx�R����py)J}�s�)JRy����O��D0u)���/�kO��5[uk7���)>����y)Jy���R���R}���ǒ������\R�Pr��ƓM���SnE\����W8B{�s���)=�ly)Jy�w��'�O{����JS��s�[֍��޳u���)JRy����R��>뿿k�R���;���������)h+��ޒ)E `�P)GNJ��$��i���{u���F�uؒ4�܎Ǐ�|'����f�k3{%)Os��k�R��}�w��������)JO>��JR�����JCD�4��D ��_q���Hd��w?p┥'���%)On��(9�s��t���C�4�I�\�)�����)JO>��HhP�iXH>!$�%�eRXbQ��4�~�Jo>��qJR��g`�R��߰޻�ַ�y���Y�[��)*A�{����R�����8�)I���py)A�De�ߕ� �A�
v�)UC�U3UJ9)Jy�}�┥��"c������)������)<���y)J}����r/=�Y�Y@�#�W[vW����Y�&��a�s@R��=����;�{y�����)JO�g��JR�}}�R���ﻴ��)��w�qJR����̶K�ڂJ��5D �_t�Z�����JO�~���R��?�k�R��u��!l$(dB��{h��R�i:�F���)JR{����R��;�u�)��{���JR����R���t�D�JTR&�n�E�4P�;�7�JO{����JSϯ�ÊP��P����| �Q?}�7��y)L#����)��i�M� �A��JR�}}�R���ﻱ�)����B���If�=TU�����g�n���e�ӭ�������3:n�ڌ#i\����x�`���=����o{�����8�)I��wc�JSϵ���#�񙮹g9A�WsG��!(�����R��}�v<��<�]�qJR�ϳ���R�����┥'��ֻ�ݬ���ַ��%)O>�{�R������<��>ϳ��R��}�v<��=kXwD��սo8�)I���py)J}�g���)<���y)Ij���V븄!f7�2�.gj	�ַ�JR�g��w�)J?"���폒�������)JN��w���Q$_-
�(N(+%*��������m�m D�l6���ά��q{lv���փqli�ҾM�f9u&ծ.h�H�'!x��'mb�m)�/-7g�ԃ�]3�3Q��G�mԷ�����.�m&JeMγ">�a��G<0m���82V����x����-צ�[Ûb�LLs�W�srd��;d�LY�=5��u�m�o�����=[��ˋmr��W;.��]�������W��܎��v ����LGl�n�M�ײc�VB9:RR�$n�N�ICQӤ�(�NL�(9�W����JR�}��8�)I߳������^<ڸ�oql�$�E"iT�ҎJR�}��8���:�������y)J~����|R����ǒ~!�K��l���D�h���q"B�y�E�R�g��w�)�@d����c�JS���|�9A�mn:Z�q!�r$⧒�����	������)I����%)O>�{�R��Y'��`�R�Vn�Oԩ��DNK�(9�V����R����w��qJR���hy0�!u��*�D ��ɓ&F�&L�E/n�ƹ�F��N���mv����rxԪȒ����*&j�|D �\��|R�������R��>ϻ��rP!gwiE�"vZ6\�e!Q$�5�R�������<qC�;3GK�8�." uU�@߈rSy����JR���ݏ%)O>�{�T!s��̶Ks�(M�T��!'��}��JR��{ݏ%)O>�{�R�������R��߳�-f�h�[7�ݚ�o|R�����c�JSϵ���)=��t<��>ϳ��R�?{���-[7l��zֶ<��<�]�qJR��g��h|��;�����)>�vW,�(9���TIJBn	�Sub6�B�5ۛԆ�vlH�&�=���n��>y���u����6[-nַ���)=��t<��>ϳ��R��{��y)Jy�����Ps�[����H�q�\����+��>���'%);���JR��_�g�)=��t<��=����L5���l���[�o|R���wc�JSϵ���ŀy�D8'o;�C�JS��}�|R������7k7�5F���c�JSϵ���)>���JR�g��w�)JO;�v<��=��wD��սo8�)I�����R��>����)<����R���w��{���ow��߁��p����A$l�:ˍŵig.��ւ�����YS"d�J��f��2�fk{��R��>����)<����R���w��)JO�~��aܴ7R�5TS�����!y߻��)���s�R��^��%"!u��*�D Qެ�TK(�E"i7���R���w��)JO�~�������)<����R���_�]5��l��Z���R�������R��=��┥'���JPm�>�hH`��,��a�Hb㎖ۡdTz ��f����#��)�Ӛi���UT��!B�{�u�)J? ������)J{���qJR��{ݏ%)O~���{�[�Y���ݨ��\�8�<�r̨E˳�I��h��ƺV�<n�H��)X.ղi������{߻��)�w��R�?{��?'�B����q"B�E���D���mS��QdB�����K�2!���'���s����)=����O�9*ǐl��*�I�U7�!���(�)�{�u�)�V$��ly)L.=͛�A�z�\��o*���9���R�`�����qJR��߿�<��w&�(^��3���ȄV���f�h�f�kvk{��)=����R����w���)I��ߴ<��>�]�qJR�C���e�:�HdCJ�,Ͷ�����Xc�`y�o��{�}-�I'R$�-fb �0|�oxX�B����;����t���3|�l�p[s�;2�Iy�{���xx0`iIng�0��sɌGM�}(�����6������1<6����	`��@<�HO�Ǐ��f���Zh&��h�	�7�����<��&	)�Gc�l��-�2���O�T�۳c��N
$!I�P>@��]{�L�$b�c8�����}��<]m�qLT�F�4뇫A$�|��|�4��Bb���5IL�9^b�FB���     m�ݰ�     �     %�j�� u�h    H�H
*�%�W��s�b�.%�Ms����1��{Na�ѭ`ZMY�2Lslܒ�=�rh@xk��D�ci*ֲkfɳ�Ϸa3ujU}�Ny�G�f�ko �ti0,��A]W�] �'��$l+h�Y��8��;d��w'���_4�͉yc;DF^��"h�:4� `,���h�5@�h�wGOU�u�vnT:uh;YG;�l�i6�+�� dܾ�7e�q��G����%����h�c����T�$�蛫I.��iB5���QM�ct
 ����YR4̥��B�iA��a��ɻ&�g��eb��E�Å��v1w��ݓ��N��N��)92�B��3/j��݋����/1!2.�b��.���&ĥ�k�v�P�LJ;pśZ:P	����Z
G6�a͕��T���E��]�q�6���h�N39z���^��
Mb��̇euN��h"����$t��{snr$�X���B�1m���+;q�;�zx��S*AY��o�b���O���:�vk�[���UP=�'Qru�8T�-�n��=q�6����L����|�n*�iMOI�T�Tz�����T�4а@�Qru��s�[6�J�{n"[;�I��R]1��ېS�m�ic���f��ؗ�ځ86Ypg�۫=8Œ�v�)�H���es��uU��x/I�F�u�;<�7N��=v
ق���ec.����$gX�Yg�-b�u�c�j�%Ms۶�5�J9j�Eir�c;�$C׹�ҝKLR]Ӊڶ���d�c�B�u�a��0�ԝtڎٺ;�@g�L��t��vgg���s��m
�)[r�q�����(!UkM������]up7�ļޣ
��{V%ն�5F��D��]�����ulD8��� ��:�O� z� @��(lM�| 
0 x�D �US@���T���w�{��������9�l�t�<tcIxΒN�7M���7D�9*+�+�W|N�vM�{V�-�b��N��}[kW`�i(�v���'nxWW=����w�n�1�r�,h�L��nܾ0�9�����!�7u�q��RȾ�3���U(c-Ŋ�V��@ԇ3��]��_���+%�m��a�"���c��l�Z��q��GvM繹��n�w{���>��i�X�DDk��'d9[��g�ۛ�J��x��0=p�v��3�Mk�vnއ��������)>��t<��>�]�p?�\������JR�����J
N������!t�d��~Q�!�O����┥'���%)�����B�M� ��ܔ�jf��Rs4��zJR��]��R�����py!����jS������)?]����R��g���3JYJ��T�!F�������<��>�߿k�R��^��L KT(DFen��A�:-��͒��5f�f���)~���┥ȡ=���C�)����8�)I�s����Ps��Xm[Db�8�H��1�q9:����!)ٝ�ļ�<ը����s��_������k9�6e�v����)I��ߴ<��;���┥'�ϻ������R��ޫ�A��z�Krߪ�����Jy)Jw�w��! �ʄsk&!�A�Y@� �z m؆�P���JRw���JR����|R�������O�Jt�~��37�F7�[���8�)I����JR�w�W�5BLQ�ݥD �[��w	JP����v�������kx<����g�����)C߿~��R���s�P����jN�g��JR�c��W����fkv���|R�������R�Ԓ#{[��D ��y�E�"��U��+��n
(9*T�ʑ���Xds�.���]Y��M�SZ��[��*��������ҷp��6�$����Ps��{�|����>�%)K����?��DBZg�*,�A���S���S�R�,�淜R�����py���K{�W�!,;�*,�A���w���DB��������%�'#j�����JR�?�┥'׽Tـ/����%7���8�)I����JR�|뱚��F��j3Z���S�UI���������u��8�)I�s���R�C�������-li4ߧB�n:�s>̕U��9Ý���?�)O���qJR����C�Jy[��+c�A���Jm��R��&� S�y��uy�"B^;a��js�}�:��v	玍���k{��)>�����JS�}�qJR��{ݏἔ�?}�߳�R�Fun�D�@J&�s4�Y�!g;�h?,�'~��k�JS����┥B�>�Qd-�(dB:v3i�e�RsCz���)I߿k�<��;��qJ�}�;�������R�����O&��J��355SB�"y$��Bj�����)JN�g��JR����P���/��N*� >d���_��R��?Ο�QID�(�W�Ps����C�J�N~����)JN��_��)�u�s�R��G~�˦aoV��l�Vd�f�����2ЖהlT O]��ְ�$[�S��(�����sI�ڧ.����K�����)JO��%)N���ʡ.JR}�;�����:����6e�v���JR��{����O�ԧ�~����);����y)J�ʸ��
�A1��%�s;PIBs��<��?g�ߵ�)JO{�w�����~��|R���ߵ�JR��-ԩN������A�����py)J_�����)I���ג��"6svn!Bջ4K����M&�[��)���8�)G��������R������qJR������)��&C��<�iT�!w����m��k�f�n@bzW���n���uuiP�v��kç��f���e����lR����'�g2AS���-F�\����\��+�]����]�[l��"��[c�lV����n@ٸsz7�˗-nk��v�;��z�v���\c%�
�o\5U�I��V˺�g=�|ˍ�4g�u��}!�n�'<�3�<s��h]=�g��a���wy����w�>?��j��ڒw�C�<xW�9��-�ͷ�ɦM�����F?�������
u��n�=�)>��)�����)=�}��BO�B����\B�^�M���$�¹g9AUZ�u��4�77n���/�\H^�)"h� 69��36��3�����wkK^ń�g몲�)T9�>B����VwkKs&�RJfޖ2'D��J����`s2��?DB��	z{���=���`nn�X��ѦI#c&{]��m<��[u�K�p4iu�qx�y]��^�
��UW*��Q�bi��
M8|�����r��3���"%��֖-7ln�JtB�������B\� KqR��	B����������ɿDD%�$�Cq{�D���)J�j���Z�9�XY�BI�y�6f֖�v;��2�*Nhs3J�a%�����7f��r��Ԣ���Xչ)�{4ԗ������K`wL�t��6i`b�J����T%R8�)$��ۑ˗�R��h;��;rs�j�Ϋ�P�����e��hr&��!H�w�Ł��u`wvi�/�k���购�sV�iR��C���73m_�ID~��&{�����zl�+�
9�:)���I�!�+�߷��]�~�h�����C��r�ߧ������Z�M���pd)˚,5D$�=�ݛ3kK;�����D'����Ŧ펦T�T��47U6{����B��ͽ>�������`~^�7�Q�H���I6��"��>��/O\h��F�D��)������ݙ5�I5*��>skK��������
_0���`V׏(�� '܅��٥�Jlכ�`fmi`gr�����_�J�
���Βk��Lr�q��`/�����٥��R^�O��Ł��f�9E1���M��	�m�`nmi`gr���Q6�D*��j���7f���ź�nT�%PM��=��,͚X�u��4�?���X���b�6�p�6PT˺��m��u7�n�h��=����@���{��ؤ��T�"sTpo�Ł�3&��٧����|�Ƽ�4��AL�����dޥ��ZX����V��6j�m��)�UB�MM�������q���
g��Z�:��M�g�D$P�Fܫs��-پV��:`yI-�:GL���J���+�7TX��V��99�?��j���4�.�+�G(�s�G73�HHҒIl �ͅ�e�&��9�5�FK����	7����+SR�ˀ�͉%�u�e8�%��3����?���&�?I=Y�N���w[:�����9V�7���Gj����{t��3��-�pC��q��Xw]g#�x��6����IH��kkl$)j2�H;/7/v���<�<à.֍f�⫷$�q�zmF��ݮz(�S�Tg9�\��� �P��ơvD�c�wb��#Џ\�k`gN��]k�hr��g��8�&��Lr�r&��_��7;�����aB���m�{#�eMS�SPK&jl��؄�g3+Kw5�˺[{�F���N�J�W�^�����ܵg�$�f́��j���8)'$�&H9�,5%	����<͛3�j��B��)���,�~�2L�>�"������rlP�w7��͞,�۫�{���Iʊ�E������<�	�v5�nY�tq�ړl=�Ӄ���ҩR࣏�=��Ձ�d����Z�D/�q�l��4S(��4��kg*��۞��5�U3 �f	���0��'�� $	<+H`�r����@L^��r��V����Z�I6,Zz4�d��)���]X,�v~�W�DL���Vwkŀ,Y�C%��RM$�RJ�>Y���۫�ɥ��ʮR���U��f�r(�IH�`n�ڰ6!(�f^���j����6�ʜ� �[�u�4:A�`�7��o���2�Xu���6v�G�Ğ������?��������R���Ł�ܵ`|�ܟ�~�����Ձ܉�"�H	�L���,�������k�v��(�K�Dɻ/ΛC|���2IV-��`grieօ��G6g��'�x��
h ��a�Y������6%R�(H�>=%}�4����sBR��>7���#�̼�?��_*�4�����8�~	��$�`pw���+
��>�� ���Ñ�O=0��(zB������>v�Z��vδG�����.#�cZICh#F��`oB:	�A����@Uߕ�|���~V>TP�P�1�Mb��2�u����_M @��U莀�D�
*!F�&�wvՁ���ۗR�5*B�q�ynm��;�<XnmՁ��k���ph��J�����ri`o77��}͛��a`y(]ݷ�S�/e�����Bq��{��ͥ�"v��MZ{-�m�<��?��[��Mo�m�o�X>w&��;Xy%�̭,q{]�:���'�U����`gri`}�4�>�۫z�zȢ"��3S`w��,���͈J|��Vf�������e�R��D��wvx�����ʼϾ�@�
���>���`j��*˖*��Я0`ztt���rl󵅁�{XXP��Z��M��l�Z(��3�Íӳ:��K�\����X�nT���9D������gU�ͷ�~~~�;�K1��w��՞��t�VVaW���`v�A��}ӣ���/��C���J�����=�`}��Vkf��Xܭ,��T�r�iRr�TӰ�J!z{���{��XܚX�uX}[����F2P�R�XfeX���^��;���;��/B����`�KH��=�K׽����~~?@��6���8�Փ;UWI%K��f����=�v���;R�ϴx���;<p�����!����;j������k3x�`Xn���f���k�!�ع���S�b�Z�eB��!�{���ۂ�1��]۩& 9�F�;j%����u���c��I�ڠ���t�O<�[a���Ӆ��΀%�!uq�ধ��Kv{��1���ww����{�{ky�٬ތ�ʷ��"ʵU����	Z!3٫kQn��G�r��4D)�RO��~�,ۑ0=::`I����V�yYV6��M�;���9���wv���&μ�%��0�r��S�9���32���&w6�X�����e�
eP�����k3)�I&0;{ ���L5BI�s~V��͹u*S��ӧUVy���Ԣ!n���nm� �̫�����0�8ӰV�zsh���Ż=�;qr�H�^=�@�Ѧ�y��m��mvnx0$�ӣ�$����UU^A:O�է��:nT�H�7��Wf�^K(�����*(i����C2�~��|��o�ʷ^�
���׭����(rK �ݫ9���I(���gu��6lqOgZM(ۈR���^�9\�S�߈����t�B��feX�M����nT�%Q8�������s]�n��7&�ݬ6�їirJ�i��&�WΕ[i�JO�mî��rޅ�Ⱦ�����{�o��WtR	�7$]���; �ݖnM6����vd�ҝ:ln�Ҧ9�`I��0$���o�߫�G՞��l	
qE$�7��u�X#l�q���&:Ĳ��+�i�(��9�پ~�*��߷ʯ{�k�%H��IIV��V-�v��V�O77�`j�h��LҠr�TӰ:�6������f�ڰ3'uX�kv(�C��%F��l�d�h�:v-�5�֬e5��r�m	N.ǋ�W�˫�̢�
���c�GL	.E�W�^Q������v}#&��LuA*]UX���
f���̀ffU��j���i�nT�%Q9%|���`b����I$ٻ�Vnm�;9)�P5T�?(�BP�}��{ޫ�ܵ`�$��1
��v{/�S�M��&����`��`lDBY��/�ݝ�`f��Xwu�ƜRG#�d�z=P�f�� f��H��p�����j{����v�8�B�QI>}���7^�:tt�$�΢^ef�^RJ�X����$��)�}��`��Vs�j�	zB��z�NT�*)�M&��:`I��0$� �T�I=L���8���=�U%�{���o��׺�=���o��2��15C�	R���w-X�
�n���͵u]�{�U��d �
�������������m[� �n�Z����\�N�c��v��c�$��ggn�v"�S�ъ�]v�����]�e��vL�moCA�]QƎzM���x^ˢ�ݴ[`F|0�Y�а�(i�[�e��u�:7����۫�qm��T��Z��=��Gj�'n�ژ�WX�U�Dv�.�:�ȥq��V۵:���	Ƹ�A�c]�1uٴl=v��"�yi^��{���6����39��[ճE9�[5��ٹ��=̴�]�5hSW�̻���2�6����喥��%!(��������۫ �ݖnmՁ�����H�7$Vs�j�/��{��X���2sꄑ����(���eD��`��,܎�\��ӣ���ڼ�t^aSN�UXjI<�ߕ��;���w-Xz!(�B�������Jh*��U!��`Ir&�0	$��06IwOQr8
K��"j8�Z�|��ٴub���
j��գj�<~���wړN狊���j�33*���Z���$=����.��MϦUL�R&���`��s��q.�P�E�9v�d���ܺ�s�����d��� :jI`{��2s�IBI���V��V�ƫ�ue�2����_��������j�33*�a������4RMH�:�����m�����o�(��zWͶ���/�m��4V�K��qI#����%���:��g��V�V1gr4�΋գ��9>/��)�9rWz�G�<KI%�����$�\�ZI-�߫�Kk6ݧ�Re(��*�m�w>_}�f^�֎�m�������٤�r�i,��u)�$P����&��ҭ��w���狊"��%!BI8!bȄ�����d�YV�os����?��Ԙgs������w����=�����=��V�o���}�m���[m�_V뤞�Dt��B9+�HݚKI'�,��8�f�ګm���|�����.e.'onJN��&Vy+H��Fފ��sgMb�1�6�Jp�~������JR1[<��<$���{�$�G�I%����I%2i-$�٪�W��e��HJ'$��$�͵W�#�(��o}��}�m���U���w>��I-{ɥ1�Shs�"�������������U��	%3;��/�m�smU��[�m5#@�✉9+�^�s��߷�[m��ߗ�6ٝ�Um�p�B"�a�<:��8�������33>;��q�u*Te(�rKI%�����$�UB�BJ�}�\m���|������U��y�k�tݎ1΍r+f�F��G]n�<;GG:�k�]�T��������7;s�#��uK�l�媶�y����m��UlDD.Wͤ������$/y�$t9Lt�$�ʫm���|��aB�Jf[{�Um����/�i#sn���Wi.�kB�%&���}�m���V�o9������̛�j�$��}�}�I*�y��4�����~Jg{���Ͷnm���y����~���߷�ZI.�_����ȉHJ9$��$��α������$�S�cI%6OW��3Յ�6� �		f@������^�F�Z�m�d]��@�1m����ևcy�:�i�'����LlG��Y��7�dz9��tzi0=\{�d��p����}����b��$o|N'L;�|a��6�����5�j|D`|2��nѮ����     m��L      �      mӀ:魸    �@@Pu��+�n�˄��d�U�\��X�u/.��z+��`ll�q��Y�ૃ���VgN����N�]�[�����N�3�5�#U>�#\j"�Y���X3���[DU�6�	vm�!݈l�v}�s֭�*�{J�s�qv/n�n7���3�T����Zθ݋�t���v�Mog{)� C�ŘG0���9wHt΍�ظ'�� ul�J�cc�.8����q��ڶHo3*�A�;J8zmun�)V6�7i۶��Ļs+s��jqO4n��4s �$�	P뇩@�Mف��3�Ӓ��p��"�cltu��ݷ":w/++ѫ���ny�W��yd����];���<q�4�:��̎m�� �N������]GTY�>��6��MMr�c��ʾ҆�*�L�Z�b�0�	2Z��ۃj������m�T� `�Ij6.j�@ܫ�/�[;�k�T�Ke˳-:$:U�N����Xu�\"�ȏG]f-�OR�&�{B�y�ѻ:�ѷ;Ћ��6`3�e�]\Y����'�NM�|N�;9ݫsl�S]]�Nׅm�����87j�g�̫en%�җe��b��(iG���ԩS���Vu����O
�k��2;6�y�_`�|��&I���'C�v�Aݶ�z�fS35�9K�q�L���ek��V�㜅&�jRYk�e���j�M���tXՇ;��Y�qح3��N�EP�Wn5��6W���T&
�k�����+/<�v@+( �VڻN뢰�t�sS�����^F��q�kN8�^�WY8Cc.��HWlu�U����p7E�T�`�ssr⸦;g��f6wP��e�tV�@J-;�v�:@B
�{�F�
�5���� �9E�Al�f�(�zm�������X����*GH�cλ�ٙ��$��о"�8�|?($�!�t�G���Q_TM#��E�N��(��������m� d��۴.���v��)6.B�Թ����n��V�p��{u�燳m�u.�s�=�j�b�a��B���s�Û��0�y�n��O9R"�m�&[�t�ӫ'��3�S�vgi�]֞v�n���a!��l����t/���Du&-è�v��6�g�ݞ���ȝ�ݜ����[Q���UGN� q��Ԋ6��ʪ*�U|]��ĩ-v�g���T˺�N�vݔ�n5e�f�����roo�������w)��Q]_6����������U���f|�"9�m�����I{���jP4��"NJ��Krf4�Sd�{�$N���������UU������;�]5*���:����m�����y$���4�S�z��Jt�i$��2U*�UH�@��6�(�/s~Um����/�m��Um�Q	)���/�m����#��c�9$�T��[�߫�I-͕m��ϗ�6ٝ�Um��	-��ꢉ�	X# W�B�����GL\g�Ps�M���49���?�ww�ɇ���	v��.�������m�{�/�m�;���>�m�=��IV��Tn8҈R�r�K;�������j�����sY~��Um���ߗ�6��5~��3-���o�7n�I���U.q��o�U���f|���ID)���[m��ߗ�6�N%XD�1M������Jl��y$�:^4�S�y}�oaBJw7��m��5K�H�u檗�6��5m��D([��\�m�m�ZI-�����$u�z�$�
 DPJ4F�n7<N������;dm�9���.�t�H���FR����]�߫�Ksn��m���-���r[c�٫m��t�T��JjpRW�$��݅�6������I1�lն�9�j��P��ݝ��R�HӨ��4X���ɱ�BR����G4�8��{Õ}���ʯ�X�*QJS�H��R��K��׷�`f{֬󵅇�!>�w�`���jcJ!HG��wn���76�|f����nk�7��&H�t�TD�2E�/Mt�����^� �$-�ycs��;]��#�{6�'�N�\�����J��OŁ���X<�O�0�wmXR�"gY.j�4X�r��Q2u�}6g�j��;X_���H|S�9%X^�;�ݺ�b��D��׋3޵`c1��˦��#)D���9ř�}V��{�ua����D���Bh?%�K��0�=Pz��%�~��6��ʥJ�P���X��`n���:[vGL��U]ߟ��nH�
��g���4�����됎ٴ��Oiq�n��nKl��1�wy����s�.�W��'����l�0;{ �>�քǪSaNR�rU�������z"&L�zՁ�����3-X���USN4���q���Ձ�ɥ��9If{�VW����Jط�;�r"RII$��ܭ,s2Ձ����z!$�{��1^ҙ�qD����wn����ݺ�3�4�'9�q�,�$��6�m D�l6����4Ǻ�WowR$=��R�	���L���\7��u�X��倮黝��m��gۯ6��[$�:0���K��ͅ�\7oֺ\�3U�ga�2�ۓ��E��QƸ@�b����͌b�j�ú����zC�3�7E��·gX�Bv�7E����<�3&k��4�cl<-x@�|�fd+�#"�6!BJ�\o�M����`[4���u�������������f�.�`�*JNAP�✉�+@Ş�;��Vy���Q脡.Hf{֬3��隖�B�����wn��W9T���Ł��j���2oСCa��ʪ
U@R�P,�`wL�`n����Z�,vGL��B`R���A�C�3>Vsf�ղ[w����V�,�B3���`yl��ղ[w��07���p�'���ڄ.-��ɷK�ka�W1��T:�/��h���e�����1���쎿����]����+�~N�I)$�I$�͞,�VW)50���J%E{�Z�8��6�fU��I����C�5 ɚ,�vՁ�[ ݓ��`
�J�E��9�U���מ��zX�M,�v���j׭ƙ HR���w�����쎘[%�>����x�\kk]$Ji��͛��ݟN�噹}��0�b�t�M(G�R)�M9'�fl�����d���0&�me�YR5IS�4X�V��Bl����w},�&��$^֒�rD&�5��{�~��U}�{�_ Df d_ć������?y�nQ�d�`�l�Ԍ	I�qH�32�s�������S��vl�m?y�k3��YY���;�|06L��dv��,�a����+)�鑵#u��*��n�R{h�T�e|��[йvs��)��y��'8n���`|���3vX�M,�Vm'**m>9ȣp�>]ݛ�IBl37j��r��9�X^�Cf�W���2@��R; ���������2-���%���*�U��s���������2l.""1B$!C��	K̼��w$�u)�R5Ib�x06L��d��&07{ ���b�4:��BTn�鲔%9{G:p�W%v7V��Z����ҕb�x�\�i0�e����-�wI���06L��W��'R0%'����`w��,fVϙ�{
M���{�nԑ�JT�O����X�۫?s�K�=�`���1[��Np�,�0<�K`�c�W�˺?��=JB*m>HTQ�V˻��37e��~�nU�{����I%+
�{���ɶl�t�x�å���鑗����:��Q�^N��r<1s�7Z�=�ȥ�S��i�s����Ym���r��jJܼ��Tv����D�Џc�Z���N5(rm'b�����Z��t�k��s[K+$�, \͗�Wm����[�[vvx�E�;n�r��Ng�����j��O5;s>y�NBP��34��4��$���P�����L��i\�]5b�vz�m&�:��bGW8���#V[Zv�iXdsv��%?m���cw��:`yl��=!.���NK�ɥ���H�zx�:�|�3vX�����)T��'d�0<�K`�c{��д���J��U����`����d�����X}��"u#Rpr6�&07� ��#��Il)?��u�m�����u�u�l�F�&�4T���ø�"�o,m9����m���φ�0<�K`�cȣ��v��kme�n�^����~@���$ z���('Duɯd�7�07� �6�/*�W�0�,�`yt��;���d$u`j7[��Lr�
Q7#���`ovA��GL.���%�RX`R�R9��9���B��ߗ�q���f�=�Y�߉����q�HC�P/Pp�I<l��m�V�ڮ�g��جl��qu��9�)(�U*����3��Ձ���`��ܯ�f��`�ѡ����P�x0<�K`I���0$�^�ű'"h%)�#���`w2ig��&��)��z��&�~�u��T��Mh�G�D%��F���ZL�I���� g�p"BH%�<h��:�w�j!�!���`gݲ�%�&0$N��|>��3��n�����ă,@�� ��1aB��kC��>D8FV!�N��t o�hl`)�)iCGˮ��&�C�9�Ł�� $��~��o#�ݡ��Q�8H�7�'�����^>b����W����p��:x���΀�eW�^�|����m:�.�
�f_+����d�釭�wnj�I��:���ОnߋwkK�ޖ�$������y�w�fV��'3g��ڰ>�k�׿?21T��7lܼzDւ��� ��]�\��;:.������unQ�n�,�f� �ݖٓO�{ޞ,k^�J&���m�`���W)#��Ł�zx�>Y����[����<��1���I�`ywK`I�	,邺J�YU��^	&A���5ʮ���+����#I1$�a!�0HP=U̛�X�thhz�i(B
IV�2[ �L`{� ��GL	���e�����VȌ��q����,�M�6gnKtreS���٤z���l�?m�����vA�$��]���?ƫ�ڼ�e$�R���&|0$��˺[ �̫���%�)5"�� ���}��t�$���vA�HWL�B�O���`|�5���>̚XlC���X��s��r�"t�f��33*�؈K����n�ڰ>}̛�� �A�С� ؗӽ��I�w���{�ޞ� 86�k �j�v���[$L�mOF�΅vxwmL<E��u\��c�j����>Sv8�k���y1�im�v �Wi�9 0��L�ƌ�[��'�]ؐ:�϶���gm�p7+�mձ��-���6�֖��0M�潎��7e��Zt�J]�pl��:�,/l˱�hL+�g�\�+�Ձ#�{UtvNx�Z����9���@�(iD|��Z���e�Y�և�zik���p���4v���J����gC�t�\T&F���	D�'&��l���GL.��t����0WI]��*��+���GL.��t��������hh~q�(�$��}�`�eY�$�s+K��j��Gr�G)�������������Ł�ݺ�>Y���O�U�v����R��|s+K����|ǹw��`s2���+:�.��X�*ļQv��^f3�
h�	�vH��3�{�nuݡ��E���GL.��t��~�^A�g� ��*�ɘ�A.iX>�M�������Ќ��"�i%p}J������2�:`N�q%�ԢB�M��3vX̚Y��,��u`uo������0%1�,?qBP�s/K��j���2l<�y��`nɻC��Ț��:sE��̵`yBK�{�?�7}�`w2i`w2-�A�&���+�M�6v6e,t#�uϞX������Z�Y]�0`�RcCC�6�����n��&07�!�U���� ��O�,YV�)f��[ �ݐ`l�����~��������ӑ�JT�O����`s;��q	D|�B�o��`�e0<���U,W��J���0<�K`�c{�aK��0���b?�V�7]��Uʥ��O��������}�������_��n��8���I�p:��i�%���WZ���n�=�	a���B�M�� �����ɥ��ͺ�>Y���[��)D`J$crX�۫gGL.��l����r��Wb��X�)�����Il�L`oM���4hhz�i*�A9*����u_{��{�{Õ����B��@a(F�bB4*:q��8!��$�p�6�]V �Q��ӥ,2�`^^e��1��#�Ύ��u���f��Bd�GI�Td��2_�������[�jۍ=���=�+u].�lo�;�R��*����߭X������%	|���Ձ�F��:sPKr�X�05t��;d�􎟿~H6�����������׀{{�0=��V��I�J6��rG`�����gGLRK`*KYI`e��^Yw����gGLRK`���}$�������O�>CZ�ER�BH�ڵ�8�,�]̅c�d�<�lN��]�K�Z��k����3Ş��R�A���hƻT��{:�n��t��v�7V�*�z�d� G�d7g`t�r%��u��7N�p�mn	i���>��pv�.�� \t/61�Q���J �q�x��-c$,�&`�u��Gk+�%�A��`:�©w���{���}�7&�q�T,u�F�ڬjԻyͥ�"z8�ݗ�ܖ���nw�~��]�g�1ZY��o��L)%��1���� �t-v�̴�f*�0<���;d�wGL�?�
�D�bŕh%)�#��zX�5����o��^�;;���;-ȇI%*I'������ߦ��o�Xyܛ �3*����"eR�yE�Uy���09N��;d� �͖mj�J�)FATd�Nd��	ผ�7=��,�V�3c.��`9��kw͌��o�#r�W���3����f�;��VkX�֔mJ$)D��;�ʿ�b�脞»%��6n��3]�wktr�R�P����f�`l���T�.�[ �������,JdaQE4�l6"!yD��V=�M�gwe����`sH�ڊF�p�M+��ɰ=�����u�6w�j���������e#��� x/#V�[�\�/�;��� h��VG��f!�6������������-�;����lʼ�"$)R9>�=�ܪ�������[ �&0<���*�+�KM�U6w�j���rlR�CW�Xd �'��6��\��(8*of�z��*�OL��<�|��V=!��"9�V�(J}�͛ ��Ձ�Nc�9�۫u�I�J7)ԅ(���wvX��$�wo�|=��`q��6{���'��Ia�����S�s9���ӗ���v�ɰ�i���3�����mvg-Xy�63�j�����Q
>`gwj���?TbM���nH��m���W5{�v��K��RA����"���hC�V=ݛ �3*�$�$�=�����]XfQ��q�iJ�#$��;zc����0�~���C*9R��RI��TD(��؄���͛^d��ם��C��$�|�{���sn�Y��;�,U�+}pVP������:諬�y��@��PUVr�Jw-�M���o>RU9CT���]X�u�w6z|��̀sE���IL�T�4�]%��1��Il�?�RG�j	�%�$)D܎�3��`un�>�۫n� �ktr�R�P����IlI09t����I>��??T�$�Jp�I���v��ś�ʾ���{��uʸw����C@�I�4��Q�WM�ˮ���pA���S����|�}���.B��4?��^A�]�i���ͩ꤁���8��� fp�H	��"B�	�q��% b�S�N��f�C�Cf��zS25C}��8����خoN���!@�4서��0��+6�J��e���Ѥ�5����gx�
��1hWHz���Q��y�GH�!�=T����i:N	@>1�KF���P��$���{���w�������     m��L6�     �H     mw]5�    �p��.���lΓj�Z���u����"�6h��N��[nT"a��R�hZ���'4H�Ўl�9RTU�-���n:���vva�AMT��uN�ʅ��d�{b��M�e���UT�����'1�u��v�����n4��J���;AWpP$ʷ�vX�ȸ��tmۭ��yر2�m��Z�2�6f�T��u��q���53��m[<�+D�q�0cn�k��X���$D[�;��d9f��:����LJ�#��Q�[�H�=�wN6�8}^�ܮ34ր�Sm��A�3vˁ3����ݭ�J�,�vz�G/B�x%�V�˴qV�f`p�I7�mV�&��ge㴠i�l`4��&�'H�4ۋ���r�a�Y�;l��ByPx�[m�&M�L�J��ΎrtѦ$�M�ɖ�$�^\ae��VY��3��ZE�U�U���(�2��1.ʣu=T��X�İtۘ�^R����vn�c.����Fݭ�s��f[�91:���$�op�$ ��1�b	���b��e����'G����[,��Kg;Hn�'9ѹrku���(ʵS���RN!�ҫ�.�GU+ slCB����uF��_S�S���9���ڎ���T���1�y����-ۇ/H�v��4�A�!m�l�w �դq�f�s�{PA� @��ta���<�]Rd��p�6��G1�i;��򬵼R���cs3���m/n��nԹ+��[%�y�b�Z�;N۳�՗gi(S�&����x5)�c�v��K���L���#�*B�Wb�:7d N.��˱s�#�y[�Ӎ5�
Gm�L;s��Nd\-�t'3�T�b��۫�(OL�sEq�v)8�G�QBw�iw=��'zY-'E�{U�Zv�R-��z�),��_��v���!�^��q] ��8+���聡�"mW���C�Pv"|���'���G>uUUU��W+�s�v��IPm��$���F��<uMU]$�)&�1�+]i���.:���O<d��f�ށ˞��B���6��\�z�B���O���t��g�gm�T,,�g̏	6�"��4�ջ���b�ۄ��c�;%B'n:�4�1��;fwF�-�L3�s��ۡ-f�G�rx�蓗.Л�Q.���p[OU���շ�NvV
�������{��������۵�/�u۬����&��U5��;7J.����Z29Q�t�s]�ff��w'�G��}�Z����t�ԍҪ
��-�wt��%�=$t���[�"<�S��M�5I�ꪪ���>�˦.��wL`y�KR�2�)Z��MM��Q	�w~V<ݛ �{�a�g}�`���U%L��"r�Y����05I-��#���(Z�Y��;��-�Lv���^�U<�$s�y�k��-�s�Z����q��(������fM��fZ�/�c�ٰj׮��J�V�[խ�|���{�x �x�
*0��,�� �͗��=���ě)N	9�w���1f���`un��4����iG"RKfM�w�ʰ8�2l5&���`03d��Mʐ#��37e�����{v��̛a(Q��oAKT�9�*�1���#��X8��9�M[t���:�54�t��8��*�ݧ%)B�I�~_����>�ʰ:�2%�36�25d�H*f��K���&09I-�wt�)%�����*��DP5�-�v��w|�vC��S�CBa���\�S�v�n�z�$����4�f��aDBM���`q����̫f� ͭZ�50%1�,��lvL`r��7d���fe_I��<3ƣ)h�/I.v��t"���˛kl�,2V��u�˺�������*���rl�̭I$�aǻ�`��)8�b�Dܖ,�w��*���f{��������,�6�C�5+02˼��&0<���6I�]���]?ʼ�Ӓ��
H���{��9��`u��6qBk�B��}����;Z=�DnSj�G�wwe��3]�ff�廮���f�8����j����$N�P-a�ٍn3rt��4�5�΋�F(1�g��$8�
���ř��37e����`��`oZĞ��q�!NG$v��U�5���wv���v�v��MT��5��ջ��;��ͅ����v��Vs)�ɑTM1���o��V�� �s*�T/�����6��j"���&�I�`n��`z""f�|�ݛ �fU���$�������V����t���e�zm���[<�0��6� �a�r�����V:���q�)4����v�\�V�]�Kӹ�;&^�=�:� #>���.Pܜ�Aprf.�-k�
�v�۷jCq���F�\ԁ�	Rl.4�N$�B���l��Ŗ�
tT��ۂ�y[��hw];f��ۤ:,ܙ����a�j�l�ҷ�����?|\�-�A�=�'ar�w/n����g�/\�ۜ�m�pZ�U�T���l�@ȗV�}�w��c)%��cK�09t���yݧ"%$)#��<��; ���5� �ݗ�#�紧�F�6��q�wv���;?Cff�X�vl:�:2B���PE�k�V��,[��=�q,��,cZ��j7♘�t���$��L`r�[����~��/��l���Sp+�+;�2��A�����]��=���!��\�����.�[��r|�{��;���Ż��r��wޖ�����8�I9�wwe���� �ܷ���W�w���u��k4j"�����#��ř�`�eY�	G�I)�~���3��XfQ�J!ƚ� FI�fn��ld���$�.�W�*��W����USU��vl$�}�����v��,݌��JA�RR(�ʌM�eu�۰v#���\���=��� ���&����ƍ�mQ���3^���`b��`�ǣ$8�
����{��y(S!���_��`s2�쾹���q�!N)$V����.�W0@����$� �	�=�1]�� g�|��^�w\���3��U(�	DQ�,=�r���o��{7��Ź��7����k4�Hl��Jy�oL`j�-�M��L`{�δ���u҅vB�h�L�`�pa�ϮX���dls�hw<������{�����'$�j���1{|�{�,]�v�� ����QDܩ2H�{�/+RI%2ݚ_sf���]y�2T��;��D��$�|��ߝ��������`��`|�n��&�F����~����P�՛�5�}6��U�D.�F��*�U(�݀ok�(��2"�G2��K`zc��l���?�W��������X:��I�F��gq�t�	���8��ء�6�ղ�۵ɇ���{�>�&�B�NH����X�5����q/�c�ٰ;���hT��*
n����[�������L߿~��#�?"q!��)$�5f��[���͖.� ��5��D�!qIV�I�w6l��V_3&��	�w},�(�Ti5r��#��6X�K`�1��t����̬�˻�;m�%�ݭm�;��]�g|���NmnnR�pV�N��0�qy,A�6;0ۭ��e3�L��<�� K�glD:��nrl�t��8^m�*��Q�ԲU���M��K9ٝ�	���aW���e�6��qл��9VK��71�H�:8��XobFm٧�8�<q��pnh�<g���جs��� ��Bry�V�cm�M��(w�{߽�����?Ć�Kٍۡ�s��鯮���8I�ьV���֎,� ���C�K�5��n�9)!G$��o���}�ʰ8�?�P���K�f���<��$�]�e�0��`�1��t������;K5H��TȊ��������̫=�
&u�6������7�GD�8���ٻ,]�v�͖V�;��wEJ$p�)%���ɰ=��w}\��`feX����>���ufj�;]l��Wbf��t@�'�v�켉r[g�;�c^��:�/-�wt��������[ �+u�e5�S�1�,��w9�r��H�p�FQ����A�Nz	�D���W}���WVff��T�Ve�1�r���; ��Ձ��ɳb!Bl�ͫ���`|������ԑ����W*�c������`rޖ�=$����j~7)EJG`�����k��vX�ݖ�Z��ҡJJP�t)�I��S{BC�+T�E�[S�M�D��ZG���{��r�R
*J�@�r|,���}���;��`�����Z��ģ�B�M�[ ����;�cV�oꪯԑ��^j�T�@'��Xg�,>���îM��@���e��Lϧ�l"Lq���5�^;�C�&�
"&�m>6�Rm��y��Ӟ��N!�����c3V���ka��SV����ON"�� �}|)���\@��M �T~O��;��_}��u�N46T�%	9,36X|̛ �3*�R�I��v��-�U"�X��yj˼�������7d���,����n*r��8���Ϫ��=��GP7O3��SID�nu3.�gt�T��v��� �we���O�$����!�=�:�Ҥ��7n�I�Ȝ� f{���#wg�{��>��`|�mk[��r�T�9%���K���g�J6s7j�;�ڰ�y��:�5%1 �Qa�g��`�ڰs2��P�D	8;�&��;�O\�9�Ԣ�SNf�l��U���P�3ޝ}���:����u]8�(�Ƥ�Ym������<d��z9�nGǵ���e���3�T��@'��X{�,̚X�K`�cK�ş�eg�2�����{X_����)�{�`��V����ă�y�cAr�j�p�1f��ٙVj�	��ݫ3+K \�;�eG(r��#��\����zXg����05l����ud��O-I��W���X��3/O�������wʽE��~օo�`b���T��6�HSr������{��h�sa��.�15�������1���;]��x�e��Ŷ�!euԸ�=�rÈ�Ӝt�&P�γӤ��H�D�$v���X���&��KwVz��uF�rK��,Q\E�울�=�n��.�tX�iM�I�1ֹ�ua�g�m��j�6���	\��{$6}�:9�m�e���Ҙm�ղ���Gg��=���o-��k-��@�D���s������ҏf�-U��x�C��1P1R�|��C��6�RGR��JqQQ�4��3&�>����%��ݫ �Ou�VZ��(�������7d�fM,������B�M���L`�c>���w\�09}>�ޥ�].J�	�����Uķ=�`f=�5N��=�ct�����C�W���,���s�������K ������~/ءLZ�Ԏ�eNbv�C��NͶ8m������6n{Y.�s���ɡ��ZJ�T�l�&0�3����_��1Ve�2����2H���w�l�"T�0ɒK�x�������{�`unk�>Y������%$)��5g����?�ʪK���;���>GĶ��T�r;r��B���;��`s2��fM�IJEy��*�@��LS��l���[v�&�"B���-P�vD{c�Ѳ������O/S.6���p�v;k����0sܮWe��a!J'$ w=���:[v�&)��z���eH����-�w��U\��ǾV�f̀}�ʽQТ"d��ĹA*S.���2w�����ؒ\K�@&�O�FEٗ�V��̀p�̚%˦�R�i&��,~�; �{��Ź���^j�
�ћR��� FI�}�ʰ<�B��͟��g5�yܛz�m��'TݖƇ��kzٕ�ٔ�Yڭ�V��K��t�������7�.�13��.��`n�D��:[ ��x�� η�ڥ4�D�M��Oq��P�~�J"d������j���dߒ��ul�R7@���+���3��X�������58&(萧�;(����lՁ���`s��vK�(oҎX�c+ߐz��=�=Ձ�m-j�J�	CJ8偋����ʪ�ɾ_���`��,;��"�z�G�v��<֗gbBI�w�0�yV�0-N���w��7�=���sv�;�|��K`�/�K`uH��%&FH�M�`unk��k�.��y��+��6����2J� �;�V^w&�D(��	D�d��ߝ�������妡)!Gs�5f��9ܫ�;�a�y�٫��Lz�SR�4Q5S`�r�������x����:��6�����
O2�$�V�Lg��k�ȃ����nl.�˞�c��m�.�d��;v��5UDB�҆���n۵���7"�݆�atػv��Q��f����#2{Wk��W���,�vJ�7��M/5v�([j�,8�v��;;�;��Q�ܳ1¾V6W$Xs[���1��]���-tFxz!M�j]ˉ��g`�F:L[�H�W>g�8{':4h�dZ6f�ky��+����̼�T\���W;�5a0�lk�ɘÓ���Ί�H�ymR��:7m#_�|����M����䒈��y�6{�<�tH8�����wW�UG�2k��l۾��;�`w:�K�Ȩ�	C"�U��s]�nf��Ζ�:KJ�RW@�Ve	^[ ���K`l�n�}_�����`J��R�RI�չ���滫w]�nf�s"�lJATI�)NDZP{>���B��Y����F�
�pQ��
��c� �RRr@��;���]�v��V�B��^�́�;�����r��ܹ�_���}_D%q��33�`|�ܛ�ܛW��l� ��*jUKN���^f́ǝɳ�$�}�ٵ`c����kң)
�@�q�~�qc����ٵ`u�rl6!��ڰ3t�\��Q� �$vw5�X�5��5��5��Ur�}��*H6ت*��@�H�te9��9љM��Y�i药Y:�R�>�w���m] � �E����ߝ�nd�)��^A�,�t��Ҥ������[ ���5v��=�[�)��߹��A�׼��%*q����������^*{�����bLL!b��ʧ����]���Fv���'�NAH��k��1nl�w�V�P��DN׷�`{��:����7"i�_�=�`r�K۾����`ws]Ձ���ةH2J#�ƌ��M�ey:�l�.՝�7h��GV]�I�D�����G`������`ws]Ձ����ū^�$T���H�<�M��P��s5ڰ1�l�w�W��\H�x���b��9#�=��t��:[ ���K`t�RӤb��
D�t�Xz$�N�́�3f�����y$�|���D(�+�:���^�(�������[��&)��:'V-�vw"ڄ�%$�7%�Yy3r�לp�g�6����Ϟ�Wr��nv��d	)S���$��Ź����WV-�z��DrC�w�`q���U��f[gKt��:[ ���K`M�ە�X�ӎ	D�MJ�^�; �̫=�=͛s5ڰ>�i��NVay����[��l	��-���kң���@�G�չ��������`c�rl�ITD*��i�(l�\=�Q�(���C�L���%M��ҼM������ �9�6�m��\rfxp��@�.�� ��.�CD:=O$���H[� S��Z��@�ϯ�������$��r@0CF�-
�:6L�G�]d>��� 1��}�$S<̾���8kBw�?@    [@@�      :�     ��� $ݖ�   ��/o� uj��I<�[�D�l箨)IklX�v�C�\�G��@�Ű�e�{vp�aă�zX9��:.9�j�ت�m�ّҮ�R��<l��[���j�|ղ��kQ�sg+�K�{M�n�z�wdC���nr��m�qI���#�c.�����a�����H�6"�ݬu��ثm6�]����E���Ea�Lp�Js���e�kW7E��R���rzRg��n0�x�۵��n^&�1��;�w]"`�5m��e��5��s,@���n��f�,�pQ_?}�7�S� ���a��m��v���ðL]p�7G10v( �˛'��� +*뮫<S�Jy���ڌ�S����g�Mӄ�(BS�,�H�>ϟ�9α8�Ȳe̪��ݠɅ)��P)��%M��AsLc+lK����؝S�Q�y@�X.DG\f�/.;+mUyԼ�Z��9��#�<X�vB�j9We^p�T��4k42D�'2I9%rb��wQæ�r5a�+k�Cu���M�p�c�M]���۝�]��\��ƀC�C:bƍ���낪�),�\��`2��!�c�����RA�0�D,Y�V�7C��=�{wq��;.�u�\�&��TĮ^ή�sm�8��܍�Σ����6�&�r!�+�k�Xr��]��X�yen6)�	~~~����uH��:�ܹ�cv����b�v�����*���
��zy�T���ez�0�.t��\I�&6��<�\f�9�:c�[k`j[YSh�P���n�t #���-��I��]�$2`���� <N'�2����,�.\�'�-\���CF�Y��wS�^�"�U\h��xT�L�״4���'S˵�vw:fw$8Iæ5�F��[#gFM\U�j���7oz3F�k6P�>P�!�l8 Uʤ	� {�v'>U:�:��4������}��~��m�ְ�����9��8���r���Ɠ��z�<We�u��v�`��(���OP�λ\�Dv�O&gh�
v"��	��ƌ�
�s��#J�i@s�ΣœBb�n�F�m�\�+l�C�LF�66��[nv��݂�:��qc���ӎ�7X�9�,�ǖ.�<m��pե��]��-�q����YOY9\��ֻ����wt�߷���c�O]'��XM1la����-uu��Fh�v�a�=�խ���V#�e��������l���5N���Ե��*@%%�w]�nf��;�`g{�����2{|���S.R�� ��������Q�f�V�o��t���I�8��rI,[�6w��Xyܛ$���l�ΆmD
D�NB8���u`~Y����o�������r=j'T�J
*8s����ݯ�˹kYo,��鴊�SmiQ3�d��Y$��Y.ӎ	D�M�����`|�5��K`I��0=-U�~
�u����y����W��⟈4��	��ƖT?"�}��~���W=�V��U�"I���M9%HW�e�"ﾶ�-� ݓS��;�CS��R
.7#��9\�\����V��U�����y$�=ݛ���WH*T�JQ�,�ݖ�s]����`��Xfj�q9LJ	S��)��/�������m)ٸ]�����$f�g�w;��'H��)$�>[���� ��Ml(�Ir@����1��s>@S�C�;����W9ă��9`���>[���u�*$�H�#��7�w[�W�������!�X�S�3��1�@�+�g���*�=��Vm<|��jAĔM9#��s������09}�l[%�	:^0=-U.��WXQYy���-��d�Ӣ��͖�Z��ҡJQ�J	ȐG�a{�Iw�b35�e�6�kQ=��1���>~�H����2)�j�y�nj��͖��U���50I'EHC����E�gL`z_D��[v��AR�P�n)`��`}�5Yꤱ�vl75Ձ���!�eªM��Xz(|��v>�̀w;��%(�HD�����y�{��^�rֻ���F�Q8�]�v�U/{�s��zX׺���v�qGHQN%Q�s�֥�.�h7������c��J8�nt37��&jTI$�)�G�f�`��>׺���6�֫����NH���ڿЛ9���}ݛ ��M_��l����S�BMUX��v_3&�B��fnk� ��Հf,�(��.�3�`fb`r�-�t豀nɌ����j`�N��(qI�f檰<�{�_͜�`q�2l	��	���;�{�w�??�`-�ET��A�7^7G-����iɌ���%rq�M�z�[VM�=��m7Y��E�;�wOr���[u�W�u�և<8�s�&j�O+�5�3��ҚExe��R�˹�5�$�'F�>'+[�b�k@s@rԷj����o��]����z6�{tnzx����)ٮ<�zp�7j��]�P�'#Mp�$���ǐ:��U?}��߽��{����?�Cd�p�%\ݺ�1��N��l���X��ܼ���z2�W�۱��u`�-e�,�N���05l���,�`n��:@�2�RRI�`f���_��1�6�����̫�BI��ըo̢��4�R+{���^�v�͖q� �:��G$r9	56ٔ��3�V;=�a�D%��~�7�u�~���M�nh�> ���z�&mȘ��09WrU>�c�0�����|G=J��kv*��N��_%9����U)���n��u
*9'�f��`v܉��� ��J��,RSPUS�:��6�$�%��z��z/���w���d���k��EE8����v-V˻���������{�`w�n��
� �Q�+��-���v�&�dI�$R��$�ʐ��vٓK��9Y�|�����w]���[�HƩġ#M��w6�z�����:wf�q��qfiM���qu۞'\��"��u4G!`uw5�f�J���2uG�!���`g�4蚩��S�e�=�"L-����05oK`f�1����ԃ�TJI�������o�/G��񃴋B�a�m6��>Q��!�ٝ��\��dԬ��������B�I��dс�z[��`yl��:R�a���ׁA�y�V����v���-��d���j7F�R ӕS�s�g5��5ؐ^j61��&^{k��`��������(�����w��X.��ɧ��,�;=���tJ�*RtG�<�K`{� �ս-��2Z`I�t$�"�R����2i`uw5��.���XY�; 鵨m�'"u4G!a��{�67ke�>fM�D,Q�HR���k����0�
��Y�(9�)�G����-0<�K`{� �ս-�������?vN��Qr��<%�s��\���gs��d
�n8���u��7�����������5�j���>̚X]�v۳Z�>ָ��D�2H��&�Ws]������w]�s�����J	q����,Y�v��[����]Y�;��Ł��&	ku(j(qI��$V���-������u��������*T�R���N��wu�fM,���k�>����BIrH��5M���{[�H��uʲ9�d��mтբx���9�O[a	��w]sp��e;t�;t�,�k�c6��k��8^չ�ض�X�7��v/`�d�p�W!���68��mě�?߻��&N����Y6fҽ���臛vҦ��-��`z�u�y�GY��at]vGd䳗��u�AŬ	a�1���4�hg1aP��]�Y@9��	%Ԕ$�$��rg�S�N&):xǋڍk��I�c�b���]<Qv�'L�*:S5):N�9R��@�l�X��L)	l-���Qr�-eeը�!`w�5_�:������y�̚_�q ��<�҃��������;�d��d��0:U�����Y��Q���\���~vn�z�]��N�`se�-��
��%UM��ɥ���7��;���`|�����q��$����e��z�N�j����عv�,�s��]�4&;�<1�yѻ'f��w\0�˭�{��n�F�Cy2���5N��'M�$�	!� !z�� x����}�uʼ����L�ID:�����бe�<�K`ovA��}����K�I�/�!I8��M,���x�l=	'����Zɝ�Kt���e���R�[%�7� �����ʲ:�<����y��D�N����sk�2vI�8(�WJ�*�e��K[s���0<�%�<�K`ovA��}6���ǜ���TD8G�Y�;����L)	lK�T")�+�FI��ɥ�޼�f_9XrsUs{B�n.��ξc��z��h6���<$�e�'8僪`�2b�����	��7��D�	�`��Jb��I����z>�_64F'�S����C$-4�������vȗ��#>�yB�y�^�X�ꇬ#%��JI!�i�%��|�&������!'����vIE����T� � ���xn<|6I,��T�o`�ppmGH`o��4�F�`0a�o6�AT�4�B��5!�y�$���,	(B�h�4��=O�m/�bC�x|��+b�ǧ):JA7*���sv��oǣ��=�1D�n�t�T| ��;E����D6 �Tv���
ȁ��&�̀H,N�:��
'E@�����g���U��k��Y��J�@��X��V�0ɰ>|̛$�$�s/K6^LВ�BQC�Ȭ����wu�̚X��V�cz�S��TQJmΠ��e9����cd����2�]s�5�OI	�<(�@@�%'IB;���`w2i`s��z�$����`k�����)U�I^[{���R�[#��U�oxڔ�8!�X��V�B[�z[{���K���k0*�1^&��-��-�����/�/CJ��Щ���8&US7Ｌv�P���-88�5����������-�������~�8���1�v��%�Ny^M�@���S�un\ѻE��uӓٞ;����t����<Xw&���k�W9_ ����-�*�dQR��!`}ܚ_���I��:�l>�́����I$�f=��%� Hg��;���`|�����0=��`l�J!�YYJ�X��[��ݐ`{{ �����"�`���2��-������q��r{���r�S
%	�g�m[��u�`x�M4�-W���U��<��R
%��{ū��vg[3u� v�շ=���6�ڑ����r���狎�;
��;Q�q�O:����[s�m���	��g�Ӥ�/9p�q/i9�k��4-�*%����r.MP�n���zv᭶��q��W�ȹ��r�]����/�8�S����p1ݭ��5�c�藒yݝ��w��}K�"b�t疕�
�h�]u.�ݼ:6:ٴ��΁��ԛ�vtS ���jR��C��>��Ł�!-�����^�%��f^b�
�ŗ��B[�}{���&�f֎��nZpp��G�׾v{���D(P�3+K�V��d���[AQ6rA���۫�ɥ���u�c�V�k�!S�����`{� ���K`ywK`wtt��G�೹c��g��q���$�\C��F��JuC�K�	�cgxk0=,��]���0=$t��Ԟ2�
�*T���S`u��7�;	(Ũ`	p��'Q�@��<�遲GLK$�]�t��*�
K2��0=::`zY%�9nk���C�SjR��Cr��6����K`rޖ����W��p�X�#�)��`}��v.�36���sn�r�����Q8H���P$L�#�/�_m����#;.Їi�����J�O;��r�:�-88R��G�~^����mՁ���Xk3]���UѵQA�H7����ӣ���-��z[ �W-*B�ƓnU����Xk3]�ʣh���C�^gy�U����}��V	)xP����S�T���-����GL�ID�efayIT��|�M���37����V�dٷ������s��jf�V��E��������؉���te��s�+hy�{kΕ%�l�0<�Il[����!�j�)A�!�Vۛu`|���-�l{h�Tfff`U�^fS�T���-��}ӣ�3k]+����p���G��|쯾���U�~�W˵�ҐK a(c�&(��2�����������1֣��|�n;1��\�ߗ�q�ݛ��ɰ5(K3�{~��N��c�]��$��N������#�Z��%�9�ƃ=�u�F�9fb�����T���/��	.|�^���(@�ʰ>[[����������w-^�	&��&��aR�	(C���{�`f<�`}��V���`j�z�.$�'
E`f_D�����d����x�ȹ�]�����������*K`v�E`f<�`uP��]Y�IRH�rI%!5T؏����^@�u�����0/6xx�:�fã��ع����J�v@U���;F��'h�k[�imi��t�7.	�aH}"c
�mI�ccb1�-����f��)�;���C����y�˷Gn�vW[ŢSj4"��Ku����GNܸc���5e�`��d�g�� �'�.$s����{Wk����H&m��9�'�-o7�f���U�>s�ּ��v��7��e��[��6�+��R�L�Of:���T�����E�):��$�H�rJ�:�^�;o�`w_D����һ.ϊ��0�)Z.�/�E��`w_D����嵺��J�A��Q�aR�`f=�`}��Vy$��ջ6>�̀p�d�%���EX��������-��s]���U��E���P����*K`rޖ���}I,O�l���
W]75�c�*vo3�|���ŉ�s�^;b�=p�!���.6�j��������u�LN�0<�Il�\O���'%#�3j��yڨ�딎U~0S2[R[����W"��Ve+/,Ff&�dR��m�Lǚ����YD�G(�#��T�����r&�d*��+�v�	
M������y���rA��*K`j��}�<��*��&z�k�<K$�t�5��Y�-9�a�۔�r�IN2JL*F�_�����ri`yJ����0%Ւ��1iR�������*K`v�D���
+)xP����)��*K`v�u� ��OAֵ����^w���^�RZ��T�A�J�vw6���y������-�K��/����x�,̦��lN�0<���oGL�{��������'�u �㇬h��O[f[�`;7n3ڳř�6nv�Eŵ��uɘ'�)yee�_�ߦ|0<���oGL]5�v�����5"9p�:��]ꈆ��m��7f��'���/%����0�)Z.�/�N�:`j�-��r+�+u��iH�N4���nJ��(�}�͛�;����fM���8I4��:�8��1"Je%~ L�w|9U���'V��̶��0<���wGL]ߏ�o���7��F*.q7F"9���W�x�!j�-�`��rev�	uiG�y�C�	�"��ǋvl��j���ruD$�A�zx�3v�%x HP����Z���gs6Ձ�������&�"5g��Jd�NHQ$�w޺�>ݚX���0*U�V�ee��RW������-�������]��eE$n!S���k�'�G{�ޞ���ٺ�����_������

�����������"

��(*�� ���� ���H�	��
�@��$�����PU��PU��AAW� ������� ��� ����

��(*�� ���@����

��

������)��ؑ���,�8( ���0���    P          
    
  ���� �zT��h
���ӻ�(� � iM
�wnu�� "P
UPY�AE����h4�PU��^     {��z�`jMd�A݄���q��	9��/y{{����6+o�����=��==�s�k������7��� {�S���}Ϫ)�p� ��
 
�� P﻾	<���>�n��� }�q�{���;�P�  �T�ET�l� jU(s�uT��������u����w�o�|�=w|�Ҕw��R�g��@��:R�wX)F��)��R�;w4��� J-e({b����N�ܥ�� �� QL�� 6e��n�R�]`R��ܥ
R�(F�tPP =�z(��UD%T@�[�ܯn������r� ��R���R���R�3���zS����>�z���`f�|��v|os��8 }]���w}-iw۾vy�oOl���o6���[�s|=��h����G��X  �{f"$�b��T�(+÷-n��
[��e}������qһ�:=�ѫm�������}`��}�J��>���}ϐ>��v�����T�Z�'�w����}7��y���}5� ـ��!�}���� ��ᢩ�
�E-�h�'.��������ϰ��y���/>�|���@��}�t��}��#��{���   �|����S�z�������{�z������ik��|���;�����;��'�m�IR&  4"{J��mRh 4 i�T�����hL�"~MU)'�P  ��5J��A�F�))M" <S����������g������O_{X��{^�B���7�Et("����
���PE�@U��(*������1�	"ۙ���4Bsr4e�y��\�	t���'!.i�1�kyh�,��M���r��]-a4Ac�2���.voWv��f�cF�)�nGf���� ��!0ޮki���ą\�c\CN��X���n�&m�_�F�} dKO7t�ĉBt�����WFI��I���@�2Rɒa�4F:F���CD@�@�a���w�O��%�{����l�Ą�jq���+!3����'��}�4�H�eL��N�Ԑ��d#H!BG�cB�.�7,���%��I(BJ�$#elP�V�Bw]ۆ��H�#
�茉$a���r��d�,Μia�Ia�J�\�V)��C4�XD��#e�)��h�6��gġkD�B.||�a�)��F�799�a���5cV0!qd������t @�e�D�2�l�	BT8�if��n�f�ʑ�)4St� U��paVH�"P���\��:��H3MW�s5��P1��NB�aBiH� T�	H\�	7���0�S	+%��
V5�p�0C	ffe�\%�1-H�
rF&�]R�xlbR%0�>�̏f��h�῵�}��$�|d�w�wG>Ԇo6K��&���5�
ڔ�;�&�dY�ܹMD�	��ePrI��4��3(¤+
���< f�}�٩�w��J`��1l�0�`��i�YR�H���J�JJ�j���;/�&�~����J�������ܤːx[�2Ie,�$m��
m�t�����-��s����}��ɭ3��s]!��w�6���Z��P�R50�.�_�2�&ᬡ$4R��.}~o�K4�^�:=�ץ0��7 Is	��[~5�U�1ԫ.�f����oC��u!Ä<�KjMo�c����g2a�ĉ� ��W7p��^��	ha��Ѹ\=�z#�&I$��B6ȱӉ(ŀai`A�oZ��@�Sۺ6K�Hg��z�{��2���vp��Nk{ٰ�8Js7��ˈ}��bH�]!*F��L��K��, p`P�]!F�.J8H�k��5��V10�k�
H��Xl�,��׻�7���h�F���LHS�FPaaM�ko �P.� ��>:�a.K�0���|l8)���0 Ip$�6r�Y��C$!H��"Q��|��X0�:6���u�M�JD�NͲ�5�S��,�\$���%YK���T�91��1��e�nZs$�$��$���X�Jc.��c!°a�##�!��>5M���c7�n�����Г��!26[����Nq���t���$&a��&)J�be0%�$�0��_q�	��	S�D)���jI
�!�\#PaX#@�|G��%	a��SI��jH߶N���d������'İ�6�5sR0�3�eC�'�0��%�k��$��L
V4�.���8G9XY��7��JI
ߡ$d�B:�}r���.����}��$�C���eLLޠN�H5��X�(��qH�#�������C���y�Mg�ww���N�V&�BP�H$>ַ��)�IaR��.e�%�N�t)H+�hB���J��˘�$'��I���$jd�pn���\w
�����&r��(`ofްJ��q"@���s��~����B0���X�2O}�¦�:(0$r�0t�C�������aP�,@���X�QK$��jN���Ӻ��`oЗ\N7����`�!rb@Ħh�.��a*²�,�hb���;�����0�l�	�re,���.��oI4c)�a��B� ���+>ݛ>�)�c
9&1Hp����d�²[�\��@��R+3
D�q�D�!L# ��4�h��N
�+�o&�BR&:w�U���I�:���0�,����J�,-�S$$!p�!�dѕ&�d
8a�n�@��B�hH�%��!`�7	�!XRfS�	LcLYRP�%ĂSRM܎jHyY��s�y�RR�_ A�?}&��:j$�h�w��J|�+
0�F�5!X�!X�L����� ���¸�#�$����V1I\�q�1cH�1�XT�f��K�J�I�����䅔�����xBq��8a~~ܞ�d>�A<q!�!����#f��;ss;��2��B�藖o6�&kA��H�I�"����A��{�!Ldq���4l�ӎ7L��!tM�dk&�jX��7
a
c
&:.ko|7�B����;>)Lvs�5�ςBR�Y����f����Xgӷ����e���2c��X]����3Z�&C�	T�1�u���(B;nC��~!\d5$'���$�3#';�����p&N$���!d�!R$4�0��0���c|?^�$��d)�@��¡�4�ă "S�)LߒXU�p�F4Di�e��̲�)���Nk}�})D��BZJCni�!u��bR�nM�ؓqa
���4B����YnɟrPɽt��k|�D �"�����\�2Lif���	0B����S	@�`�P0�ŮeR"Q1�seM��ȳHB0 ��,�#%��L~6������+�
8��8$�[ �V!���&%�4�$!,t˖��&!̦8�Ir�,1ŕ��$���L��\�d;�Q����r66CN�����t�n�!RL5���PWۂ��z�:��H���
��.e����8u�Za�d$�E�(A����jV���F3)�;��ԓE$�4���e�&�T�#H0cL]�ϡ�Idٶv�4m"I�
���l�E�b��L����>)p�%@����.M�c)����ם6P�d��6|Ô��!�|'��\��.�IS_l�Ӊ�
�������]o���L��CL��o hH�w���s���&k��O��k�d,4hs�kn��OB��	��I!�$@�
�1��Ͼ|;��5qd`Mp�"C��"�,��:�HD�R,H ���a$#0tsf�Xf��u�m$"]>~b:F��b�JF��[�)����cLgx���l�GXi�#B$IRT�Ys�)�y��au��>����4��yNgr��>^S��Y������m$�BB��2�.�p�4!ԑ�G	CC1�F��.�[���=��˹�fͰ�3s���	�L-�A����.���p�d���S�&�d2����S.�:֌"� m"ĈK"��]L��hA��j��������74c'���.h�1��B�V5���5�'XAiXF#i!#0�"Mʴ�6��	���C��$a*�$*B R����c�0�"�dj��Ht}��z�%�]��7�;��O���d���O�:ѢF�53�����9�	�4@��捒���z�le��(���)��5f���ށP  ��4H�m��X��rf�H�'��я�f�a���S �4Cp�t�$�4��B�&�VYH�::���C�\�)��$H� B�),�K4af�Yp��d	�n_����0(ʤIH� D�%�ޘFjC�sL��І�l��ޙ���dL~ P"R�BL��$��u���z7H]���L��X���	I.1{q������!F6\�K��\�4kA.��{��_u߹�u�R�%��ã�m�7�80'M�4� �%޷{�ua�,XQ���$�'o@���B��D�6;�Xh6�H�P����Qt��R����T]�I�����O��L��B3fDi�>F��F����j�@ C�~��sZ������F��I�#��\��9i��nHBI����K�0�Ѹj%H�#`FFjݛ��,Ӱ��d\ܛ�	`kD��I�0w�M�!�M��2HP� � E�!!H� �$[q�A��f$���.<�|�HG��Wϝp���&��0Ѥ7o�SZ�Ɖ1e�q�F�����+�*��	&�`Ŏ�Ѯ�Ml�\���S}�C���o�&�VVL�3D��k���F�!8B�B�@&��K��]c��Y�ˆ3�P��6���,��	X�u�M�f�]F�Y4h������3�A�JR�	#9���є�[��W��3�=w��'yx]Ó� 9<`�L	chIul�[�Y��v=	�Sa%�ʚ9�tiH�,��H$R�8�0��Ɂ�<f���]��B᠋L�B�G#dX�M#���*d��ģ$'^Q���G��0M)��� �ŮkB���35N=$��\T��BbA�ԉ��%IV�p��ٽkUR�UUUUUUWU\J������UUX��j���ݕj�����h	W�RZ�]=�[\�;g���t�*�@����^V��Uumm��gl֯FU���Tb�AV����>�FX骇��D�rqAs1v[�u�J�^��-f�UZ�tP���+�w��@섓�.x�H-]Tp�����,��UUZ�j�r&�$�J���׵v��`�`���tt�t]Wg�0f��j��ʤ�]V5�����"d�y�y��U�b	���UH�V;e��b�`�vwI��M��U^�v��eAj�m����k�Od�ƪ�V	�7SD�$�&A��G$vyvn�vx�t�9f����9������^�B�z�:�
���j�i�e��`*�e�9I�k(5.���j�+ez^j��`���EQV��Tp�/m�Uȵ-AKPUV�vj�@�j�j�L��er�VV
���7��+E(\����]�k�MJn^gEv�UVʵU �6ڪ�݃z.V�YT
ycT�����UH*��V�W�f�U,�^z�Y@j��ej�v�0��T�8�Z�$��L�ll�j�P*�#/�j�`� U� +*�d��P���J�L�]W[~���U�U�t��UЈ��m��T�Ξ�Q�y`[���\��U�J�ʼ���`CU�=�T��cs2���lU�J�pU��UN��6��W(�&:m�1r�U*�UUUTP
�U�u@����������� jV�����r����Թv&݃mB��WP0T�tº`1�U��WUU�H*0���t��^�H�5��V�S��Mul�(�y�Vz�������Q�ݫ�WhؔmmUUUUGU[U�R���j ���:v�5AJ����j���T깝��[7J���+q�+vwS�8�s������P��)we�U�vk�@Ke�Z�UC�V�@j�ԅ-Utz[UU@R�UUU@��=�8���q,q��HҭJ��Uc�-UUP Y!V��v��<���!KͰnUPUUg	KWU�T��UR�UTݪu�Q��T�:�iZ���*�����j����깪�7%mU*ʺ�UUUT,m�VP�3����/ ����3�����+ȝG	.#�+;gDb�TA��q��<!&�m�W+�c�W�]�4�1�����!�͵.�*�UmT�����/+]7j�-�ݕb�[�{my�A��d&۪ԛ���l�UAī�e(*�-��X)�j��9��UU7L�UUAUh��AV�5�MR,������	l=��!ZUla��j궩Vڪ�������Ug�j��j�����T�H'kF�Zǯ)���J���Z��U]UM��k�mThV��f�.���v���UUJ�U��k&A�{G��V��yTH�^�a����	kjy@��p����MT�W^��:�ue;f
`S��C��h�m2
j؄˩6��I�2]v��x3�PS��������ԗ��� ��T��PhJ�3��T�0�gۥJ� �=E��3@&��G%n�j���v�a]9�v��ի�9iv]��q�:8���T���)�Y'�+db���V�ۤ�5]Q�OW<��99v��j�j����+]J��U_G��m�յt�5AƩU�
yU%�;�5T*�UJKUUUUUWUm���PK�{R���h܏7[TW�_U*���U[�j�
����*��U�
��r�@u,UU]m]uJH3�ڪJ�W]ݢ���WTP]Q��j���+����X%Kq(媺��f�P"U-n)`�
U��U�ZT� n�����
Z�b�V���]����(��yU�������\ ](UR�U�UJ�*���Qj��F,UV;(r�@j�mV��We`ON`�j�������U �%-UUP\�UhaV+UP���oUWUUmR�Ke���۶٪�����t�	��&�6i�^`���:��6�1��W�������6�UV��U�T�̫�[UU�D�UT�]UUU*����&z^�%j���讎��U����X�NZ�˰��sm�p�\�]�i­����H�U�U΋.�\P!5X�T
�T�\q�
�"�5v�zy�m���#b��
�wc�\�]�h՚B������)"�u�2�b�,r��Ep�s�����Z��䖺�Ʀ� ��Lb��ꪪ����AV���t��)�4�^�Z�j���ĵ�wgA�дJ�UUV�Pr2֮���aY��%]�\&8����芋�m]Tڨ@����*B���@b��i�9�q�T��U1\�1V��^�[��AWh�scVH�U�i�F�tJzd�� s@[�#�sV�R�%j����
Y	���f�Fݮ��u���U��g�mj����?iN���yVyy���j��ݠ�s���	A5I]Euu�0�U�s�Q�S�@�E�R�[sI닩׉.X���˜*��OpK�*Ӣ���( 5U���Uʵj�:�ʁq!u�h�iΨ�Q5[mI*��n��t
�:��V(^��-0UUUv�|�������
 ��[; #������l͵UP�����se�t|L�UU�(�U�����ŌU B8�f�"�|���V�ں�r֊+��y]�Y`��U%�nK�+Y����ړ-��4Җ�UTpU[NMU���6�ɸ��XX�!-b��P�5=mUV�hx�F�g������r>�iIj��^j�ZW������Z������ *
������]WT�e����tTP�B�J�� @�*�UV�UڪlZ�@,�/��8��
j���+ny�U��W�۵J��b�ZÆ ��:�J�*�(�Wc�jk���*���\���������eU�������U�8������) Kl���Mvƶ����
�'mAU@���R��KV�٨	v%����U�*����
�j�j��h6:���Y�;5!;��,�UR9��]Z�!�6�p4�M*ꫨ8���
�V���`E��j���ʃT�HQT��y�����c����еU�F�d3U�e	���UU[J�ҭ*�R�2m�C�i`��UWR�+UPUT��֪���������P��
�UU�mUUUU�UU/�j��UPl@@U[�]Z��6�V����(*�5UUr��  �@UV
i�UUeX	V��vuU,UU*ԫ+�j�����U���;c���{gf�j�Z��ObUڪ��j
]�6�p5 �j��Rn�F!i�[�m0Ŵ*��UX�Tev�V�v[��������[PT�UJ�u+UUZvC��Ͷ����ꥹ�J��UW]AAtqu�4��j���������t@��F���\�x%�9�ͩV+��5MP
�U�F�@�\R�Ō�UV�O~����>���tAʩ-N9&wGKҽWOb�����ź��@W*�Y�Dl0umn�[E���	�=�+�&���Uj�v�N�v�*�!���ꂂ�8i��i@[�U�ј��U&�<K�R�P���pG[�Ƞ5@U\��*�@m�aeD�B*��f�5��һ�%&#��*����R��+eZ��V�����2}�v�T������ +;,/�ru.�UԪ�S��5UWTUUS��UU���U� �IiUUUV.��Yt8Ң�	e�UV7-.����
�NM���*��1�-/;��R�UJԭ/5�]t�<�T���u@V�U*�U�UuUm<�UUt�R��(���UU!J �Uz8*ڥV쬒���f` j���t�޵V1W]*յUJ���"�*�UUv�*��Z*�Pb��<f~��!���MUT���^X*���GR�U*�UWAKuUR�����h������j�����V�wR��F���;\ʶ�U��ˁ��TUA*ͺT�kq�b�!���O+�KJWU�UT�mUm$3�5m�j��e{�����UU N�	�]-UJ��JHci�U����m���[�mU)�]mYF�����H�۪�ET�J�Ԩ=��Z 	vW������Z��4��Q`�J˝�qĜշ��������km��DЪ�P
� �
�
���5Z@UQ���ڠ��⺪�t:{3UmB�5UUU*�� �������%W���-suR�/V�6Q��UUUUKЃ*��sFꪪ�(�\���W9p5[V�Ul��8�mU[N�ڪy�ay�'�j���UJ�Uv�'�Y�vy�ԭ� H���'� }WP��UUUUUu�Ee��2��-p��TK���}J�uTUPUej����j�({���2�m���
y��UJ�p��z��9� �V
����n��V��Q���vg���j��hڗ�vœ( +�=�mk4��b6t���/JT�%���{�\�D&[]�P^Ӟ��;T�mU]U����O2����W��UU[UUU@V�V ��,�R�cê��cst�-�-UUl]Z�����a܀�@T�6j��
�j�e����f���6;!��UUJ��+���Um{$�y��uB��UUUX����*��������RT���V��;@�UUUUUUUUUUUU�JY\�n�=G	�<k5��O��GU��Z���=r���� ����Uc���UR�ln�h�j�V�O��qbP&
U���5[UU@U�������@	�&�ҭ+l�r�6�G)�l����t��O� `EN���t��Ƃ(_��@��.0X*���`� �O�H�1�G P�)��(��t;� � lBH$bt8l6���~P~Dv������ �P�����1گ�(T � ث�SN�a B H+�t��N�� qQ~�"T���!�j <��G�*i>��R�Wg����N�)��	(?
 :U��8��
!�]��@#��t���1�UW��
�D>PR�ΑP���T��
�F# " D"�H�HH H$`�M)��q+�E]"=H�G@��`�AW�|�	�:c��b��Aҭ��`����#����@*��h����m
�=US_P������P�  ,�#|��L����!@'M���<'���*i ��Ⱦ�(�(�!
� 0BQ��YD�P6)�U��Z��� ��u*[���~"pH��V�"(`Zl�X?/���� �3j'O(�ρ�%R� �Ҩ�����!������Ł�>����O��Ӣ��MQxi�H�@�@H1B"��*��G�
��uD:���8 (qU�z��C��@:�j$���Q^��? ��bDʐ�&�3DdMEa�aPB����޵3.�L�`i�dim4�.S.��:+4�/�����ECt�iÓn�t���J��C����ڊ���粆�a���U��,���Jw:B�˒wA���H�]#���9����l�g1�zҏ'�;Lt�%a�A$�r���9�8$�/n�m��!��Nk�\�7uZ�ݴnj4y�J� <sЃ&ؘ-�Q�хbʂB�P����W�㶌��Y㗓jU�]nz�&Q�yoC���j��S)��81[���\:vns���O.�ك&�̰@�ڒ��%�.,�*�j�Z�Ra�;v:);��|s�0���{I[G�vm���ނ2^�:n	������(Φ��\���/Ò �q*E�sn�'
�ܚv\eӇ=�r�IQͻ�t=-�o���HU�6t#��	G[���tR`h��&�:bs5�%D��)ŷ3��;7A
��ׂ8�6�����-�kk��	��Q�!�5�.�Z��dm���%a�^���[^��p6��LÒ\Ae�ݧ���D�/<H�mɆ$��"J�lΥ�y[�Z	�b�m�ŷaەM�&�U��e-`��=̭��m`���9z&�-ێJݬH=�2�,�ł5���l������mr�&)�a�x�U���C�']�l�<Yicld�Pi0�Y��8О�#vm\G���E+3��w`�����R�R8pf�9Y�L⸲ˣg����Նa�¢=N-E��'2��^��It�W>V��BR�y��ډ��1::js��I�E�l��:^�8��U�Y۶eyS=uҮ͒8XQT�X��݋ �D��E���SųB�lgF��z�[/.J�&�%�u�	]��g��&�K�.�"b�>Ў�r���uŜ�^ɡ89VM�v1M���\:��z����u̖u:$o!s��:�n��]�Q�:-�6m��d׆����������ԩ�%���5N����e��3lOE�dI���՘oI;�����@��FH��H
�U�'��)�����QQ�� �x"��Yx>D��Ν'�t��ۤ�l�?�P���MZNunSF;$Eh��Ғ�5e�R:�`B�b7c�iH�ĭ�Z'�B!�|�	�'R�<�� �%{�;����Ħ�j�����/�����l�t�9��/]�x9"�*���)cz���ye}T'd��^�"R^&�1��n��윖;7C�� 7i�sOkk��`�^!�Ʋj�I�0��hGzܶ[M逥�-�!�-���i�q��3�7��q�ñ�3�+�Uf�\0�����z�*���X����ݴ�V�ƕـ}Ş�*�I}~0	�y`�p�;݉��j˻E�CI��7��o^ŀvm� �=� ޲�'wm5Cj�6�ـo^ŀvm� �=� �ˆ���.�Ю�mYi���vm� �=� �ˆ�{�V���i�M�$��$�gm�n}�D� a:ܜ�ŕ��]ϓ��P�с�i���cV+h���;�<��`ױ`�`�Q��M��t�wwrO���7�CDL��H�`���b�%�Y�]�>���ܓ��ŀv5ĥTC�M��n�z�,��<�|����wv�ak��w@�n��ˆ�{�ˆ�۞X����ݴ�V��+� �=� �e� ޽� �^ŀ{���s�Ԡ�����Ҳ�{�� �4ö%5��R!{1�+B�J`R]]HuƉ�(�!�����ߌz�,�{�{�Y[�����n�n��7�b�;ױ`G�`>���g���}�qk
�m*7e�	��]�9���6 iC��b���ā@X1�F��Ř(���0H$�(�}�ח ;�-4�WB��][Wwk �=� ���|�c�;ױ`���۠Wv��.�v<�{��� �+�c���	���z�		�\�{'.�q�]cFG�ۺN8� g�$��7cE�>�O<�{��� ���wv�Z�V;շo �^Ş�r�;��;���v<�*��Zi�We�Wk �^ŀ}�p��\K�O<u�,��1�Yv];��v��.�v<�{_9Ty$#�D��2#�t�����t�NQo-�},������%v`-���2���Xd�`����;�Ӿ��ŉtK+_���q��"ru�����qc%g����%n3$�Z�.�n��ӻ}���+ �^ŀvK��ݏ ;���wB��][���{�.�v<vL� ޕJ4�X5wt
���.�v<?%'���v9�wZ�[U�Sv4[��T����$�����Xd�`݅*�E��N�um��7d��>ױ`��'/{�ܓX`�Ø�@��&�H"�"0� �H�Pq"H�#!�``8��	E�B,��}���Ұ�2P�2����&A워�O�6��N���=����n��6��M��/N�zg����n�a���C�7Qf���Sr-%N�1ѳ���y�u
X�n���Q�Y��^c�*�8�(;'9���+0(R�STn;��j����U�>s6���d�U�Ɇ��O.��
\��N��s����4t�$�e�(�[����s<�];g��̩zE��5�P����S���i
�;)�ے8#&t��r�U�m7�y`��|�c�7d��;�`՗eӾ'k ��ʪH�� ����>ױ`�ʄ`;t�J�$����&V��� �wTu��Ю�LV[N��yI�}Xc�Xd�`-����[i7t*�*�ؕ�`kذ�p�>[���e`��}［Oq4@��4�e�&Ik\\�hicfLd5�;���k1v�GK�LH�l�wHWv�O_���&W���9��<�	渔��
nƋv`-ٛ�4AJD"����3��2�1٣ �1F;�渡��Ug+�\�}���z�`��}$)V:,�v�n��&V�n�`�"�;"�dv�E���v��=Uʪ���� ��� ��&V��1�4��];�]�0�p�=U�l�y|����&ˆ޳SQ�en�zK�8��l�l����n 5�[@^�
�5����G�5ֺ[T�����>�2�	��nˆ���Ь�1Ytӵ�vI���)#��� ��� ��X�ȭ���]ڢ��`eɹ'{�zni�	� �^�?+���:��XݙX�R�J&���v�J��7e� ��Xd�X�p�65Ķ�!�c�"ݘ�"�;$��&ˆ�.�(!t��a�n����m�����^g���s�Z^��pGb��%��D� 8V���y8u��7e� ��XdUl�դ���˷wu�M��+���=~0G�,�L��"c�b�l�w��v`��Mr,�L�l�`�ʑ�+N�Ҷ��0=�/K������	%�j����6(�  o;��nI���z5��]i�e�N��&V�{���$���$r,�V�-1���	[O�'Ae�瞭�I��;;\�p�Q�;����-6õ§e��+��$�v\0	� �+ ;
Q	D�X4���0�p�r����?y`�{+ �\0�q-��|�H�f#�`�e`K��.��R�v.X�h-�v��2�	%� ݗG"�;"�q��CmZ�.���$�`��H�[�}�{f��?D�I�vf��[�N�p6y�7i�tk4����Nδ�C�.j�\��U��QeJ��+3lL.܊�j��hk�x����� !"���nQ���*l@vEǢ7W/V��;tV:�B�o��.((``*��pg\�q�!M�(4ZEr��=p�n���N*�v:���X��1=Ps�ϊ�=��;�v���u�Y}�]5:�Nw2�ph�)�q��S'2�L��9nI��]2tv�7m3���p��1�ws�;A�i�Z�m�4MQY���'�;��Ӏw��Xd�X��wFT�
؝	�m%v`9�&V$�`��w���ۺ�J˦���L�Ip��9II��{��X�ȭ�7t&Z���ݘ��}��H�Xwn�R�J&���wHـ}��{��z���%��$�jZ ���u�*%�^C�y|��!��]�̻��]rZ�q����F��-�����wn����*�A���wg�U���\նk&���'��7��h�bE]!H����G"�;"�n[��M��˻n�Ip�>�p�"��ۆ�ؘ𦬻�]�շf�ˆ����0	��ob��GIZ��ݘ�E�wv�I.�ק ��<�b^�@�)e�6U�̤�kq�� 8/C&��A���o1%����Sm�5l�J˦����/�$�`l�`9 w�+lM�	��-�wf$�g��r�;=~0y�� ���=U�H7�/!/&���wHـvz�`9Otl6W�;� ��ۡN�Q0|�O��dB3(�X\��/�?vQ�B?3��S�d��F���F�S�ޓ�B�
�]1���4�Q��T�!�_�j��$��uLrl�t辏���W��(�\b�c�	(ŊC"R����t���6m��\���%Js]{�D4p��-�R�&$��`�}�>6��HX͇Ú�Y��@���pz��+�c�a��A�"<�� @�D���[v|'># ��0��c
��!��g �M�"~϶"����E�H��U"��y�+�`#UR��Ϙ���iE8��� @��(�� .Հ�4���V䗆�ۆ�k�mTC��bE�0	� ��� �\0=\�Wg��ݜ�V*�WhCeݬ��Ip�>�p�$r,�U�W;.'M4������u�a�Yj�
"c��Ol	z{b��{7T�6\��Q]����Ӏ}��lr/W>A�_����2����m�0�\3�\H�~��6K��?w�N{$���jK=ŭ6�0	��,��Ip�>�p�;�Q�m�%v�b��k ��� �\0w��ܛ&���
(� �؁H�a*��à�C�)���o���V�~���Йj�LWv`K��z�=�>�~��;�u`�G��:�l�����8���'ptk�ϧ�3q�L��s�9�lmXw�:^R�]�h�e
��=ﯧ �Ȱ��=_ ��~0��(�y���!�0	�<��_�����>�p�߹�l��~T`Y˻�Cc�0	�_� ��,=UIvz�`�_��
<����j�ݘ�9K�����Nˆ�ɞ0�ǚyE�ݗe4���}��Nˆ�ۆ5�X��Kd�u�/Hi�߹��bQe
�Ps�e��������)�/��[���M�V��]��b���f�$�k���­Ϊnx�W�&�g���N���&|O.�F�3��H�;Ra��s��{m���=k��;2v;tʡ��Ő�N.�]Q�7sD�<g�]g���\S&ur;����	��� l��r�0�fW^�v�Ď��;GU�	��i�ش�,��M�'�I�;�e��4��Hآqf���g����D�z��M�"]@A��)βs�I�����z9�wv�M{�ˆ��<-����LV]4�`ݸ`^ŀ}��N�~�Hվ�n�j�n�Yi�����,�v\?�666=���lA�lllo����\�&�]f��Z�؃� � � � ����6 �666?����A������M�<�����k߮�A����ڭ�G��L���ff��A����o�؃� � � ء� �_~���� � � � �~����A�A�A�A�߷�lA�lllgo�.e�����fm�nȻOc�i��4{s��w$�s�s](<�[[ʶ�[��;�'kll{�o�؃� � � � �����A�lll~���� ?�T�A �`�`�����M�<�����R_�5Y�و��'I�,�;Y�v����׿]�<������z<V�x(r:���}��b �`�`�`�����b �`�`�`��{��@S�P�������\�	�ֳSZ�[sWb �`�`�`������y����b �b�!r9~����A�A�A�A�����b �`�`�`��~�cL�̗2Y�MkSb �`�``�����lA�lll{�o�؃� � � � �����A�llA����Aä�gI�Γ�����:�L\� ݈<����}���y_�׿]�<��������b �`�`�`�����lA�lll���O��{Y���\����9t�n�p�&�a9����'��#R��-�~\y�c2�R8�Z�؃�lll�k��؃� � � � ����6 �666?��߮�^A������M�<������ߵߌ�r7\��t��Γ��'X � ����6 �
�66?��߮�A������M�<�����k߮�AV����ڭ�G��&\�\�3Sb �`�`�`�����lA�lll{�o�؃� ؃�uC�P�O#r(1��>��*{�;����k�]�<�������M�<����}��'%���Z�˗Z�y����yߵ��b �`�`�`��}��b �`�`#`�����lA�lllw�iw�V`vZU��;�'k8ߵ��b �`�`�b�������� � � � �{��b �`�`�`��}��b �`�`�`����$$�ro��Rb{�ӧW:x�.	a�V��b�"�>$�-��4����YEV-��w���666=���M�<�
9�%����6K�ꯐz9�u{���Ҷ�b-Qwf;.��%��=��>�p�ԑ$^u�ձ[�m+.�v`%��&��R]����� �쉺i����v&;�0	�b�>�p�O}�znO�_��DBZ���!">��҇˵8���nnI=�}e�&�V�؅wk �e� ����kذ�\�Uy��]$�$�V츘�Y)9���&�q�]i	�zN<]��gY<6r����47g�{��`ݸ`=� �e� ���*ąeYwaV�v`ݸ`^ŀ}��Nˆ݊���wc��vݘױ`l�a佾���z�p����)U�.�ڭ�l�`��wv��r������#��I؋\.��'e� �+�͞���'�g�]�9�k�rN ��(J�P!V%J�T!(�%P�@�U��IA1RЩD+7t��M�Ov���&*;-�
�ȷ[-�nT9aTG++L�s�ۉ�u!�PMX�Ӕ\�9^�u��~��w��ɂ��y�7�����E��<`��Gc]r�Z��Ц=�� ���u�@����b��U�v��h�ᷫ"]��n&4	��0h��`��3u�%�Q�U��LD�Bb��kXH����%ص�y�ZI�Xe�XnM�����$�����w�L����Kh�@h����ͯE�[r�h�o]���$;Yܐƨ��ODN*�k]6�����`ve`l�`��uvD�4���]�ݘݙY��W9ʤ��_����wv�� ���/�V�V�Bn� ����$ۆ�Kd�V�Oe`F����`�v���9��O��}��'��+ �fV��T�=�0�U�X���.�*�Wf�ٕ�z���������p�>�
	t�Fmً^'#u)+c��,<�`�q'u�M�v�u���8��*rπ{�}��>�p�$ۆ�ٕ�}4��WwtkXk35��s�צ�Ҋ��Q(�b5b0Z1��"CHm�+��̪�2�_Ll�X�2����Dĕ�"��0	6�wvea���I{��`�����b��4Yt�� ����$ۆ�ˆ&�0�ț���;�bc�u�I����x�z_���+ ��j&�!U�l�$�`ؖ��l�jB�m��@��9S�x�]�|Y��M���ٜ��8{���+ �fV����9ht�v�� �n��*���{+ �����\0����VU�vi�� ����'��l�?=~�
��7�S�� ���wb�c�v�;��n�����=�`���`yl����ǅ�$����Վ�� �e� �����6Oe`ve`��҃b���Z�k�1s�^�h�v�x/qӹ�n����uݢ�[I+lE�v`��wve`ve{������+V�wbh��f�ٕ���I���� �n�?{�GMuafZ�����y8͗?s�_����_�{߲�	)đJ2�������R��x�=�u� ��ٹ4�'Bz���4��(��`��a���9	Zf�WJ�|������}�ڭ���4ݦ���'e�0��+������?{߲��\0Ԡ��aq[����<�px�o
�\�s�7���s�-(_3Dq=�l�BV�wv�����XݙX�/����y'��޳��������Q]�����&̬�+�I���.�`��'=�KO����Kk���������0	6�z�Il���=���")hJ�k�ݘ�\��\�{��`����I�+�9U���}����~��V����h��7V`ݙX�Ur�U~��ݮ�����7$����rMH1rb���C�*��Gf*o>���`"D�2R�!����� �h���.i�7���\�V��$ ��2�-��]8�A�h8t0H$�����Hr2"ed�ɲ�H,`@#9#!	$CIͺ\�K��\Ѣ\Mh"U��j��X4H�e�*�+@�u�)���"ϱB0a��1���	�;�'��@��@�H�����d��$F	#�	g\aq'
*l MJ��n�{T7�oُXh���K�R�L[�h��a*J�P �"1�D"D��o� F,C�la����H\dILXP\d���c���6hw� h��;&����XvU�`�K^�t� f��7	ILB:�vU��,�u�8�d֍X� �X�!L����II� JT��P�>��XK�˚t����~z|P(��}�@9�%!�.l:!$9��n0&�9�,gܕ�tVYчYzI~Z���R43l��q�� �Z�s!���2[e�\�@��P�bU��ݬ������Ѐ'�[F����>6�K�<�Mz�	���t��Э�6�4#�v�^����<*�l�s�$�!d%�
6�3�bv�嶏\[vx1xBs,�U��\0�ZBV��ͩu�d`k���:�>��RI�[/��]��x��w�h�G�w.��cdɊ�܂�V�D��MSR�֜n
�\8�rnK�<�`�ې�]UW;�y%\]��ӂ-Š��T�<a"���은keMvΙ�#s���PGl�O�%�j��yGq9��r�d��:]�57[�f8��r
eaԬ�A/V�R
3uNA�M6�՘��:�3�(����P�.i(�)�+�U��U��m̯ 2l�ql�Zv��%�Q�&��ӻ9sx��1�����u)��M�ZvZ��	u���P#��O� �N8^�g.��7��I��'[�u��Cc{c/�^,;7&v�9�L m�n-SX�mv��64\
�MyѮQ��O\�3� «�-МlCPl�@�d֝%=�8V�	x�q����km�z ��A���:x]9d��y��	�m�bm�ؠW� ���nέͳ��8z^U*+m�g�r�n��y^C��6��i:�6rܽBUr����qGJv��R�c��f�AWR�d�e��=�ѷg��4q;�qb�7\Y朻 �	�6�1�q���y�r��aM�j��B�gu����ۃm��ø�,�U<�VvBⴷ��uV�8	Fۡ����]X1��"���+Sh��y���nx	���ul�˞c]���-�ȕ�2m{T�v9����Nt�ɕG=u��z�D3	������y^=:�v%�C̴#����u��(���YuE(s�8��5υx5��MQ�Yss2�͓ġ��1�\��YW�e}$d����c���`l����Ԅ�SZ�mŶfv���zr~V�EE�|D�<
0�����#��� TS� ��1D *�Ԝ�ٛ���7V��F�3��^#i@��9��3���c��`���j�RbÅ;5p�L���K�'N��y�59F�!.Ktd�mۜ�\IG;���#[���#�q#���Ã���=�{s>�4\�Ǜ�/l�x�۶[��s��i����8��5�/VCp�F�Å�D"�w�x<���F�N��Cp��ZN{U�5�h�"�o�K95�̦�[ |��
�,hQ��q��x�u�\6�R+Z��r��O&�x:k�2Ը�g�w��ܜ�ˆ&�C�Uϐl���=�~I�+5f�sW%�ѹ';�zo�E�2~��`����I�+=U\�����꫱��,�7f�K�wfV�U�����߲����`wUEX������WV`{�ʥ�{��=���s�\^���~�=�j���떬����pg+����x�z]x�;�2���Q6�������r�M%��rQ��nC;[!�ͤiu�~��e��7l��V|�����$ۨ`ݙ_���UW:���~��?_���f�����;����2L�D��J}�H, z��vi�7��w���;�~ٹ';.��RF�y�vƝ[E�MS��l���;6eaꪤ�=~0	����kvab�.3���y{�~N�����ԋ�9��\s���O��$�_�J�v��&��\0s�n���%��;6e`P(�%Q�m�4];�@�C�����qV���*-&��R�J͛=�H�	/�C��j�ݟ5׼���0͛?�_�G쓿���7$����7r�]B�k\h��Xwn��*������;=~0��{���wt���������(�T��֦�����rNw������C�\���{�l�� ��AeZT���ɚ֍����� ������~���rN��0%z�ʧ'���ǼS�"�E�v`*�V���>}=��}��}�� J^�eVْ:F����@i��6�hf�Y�*�b�a�O�A��v��=�
r=&��t�|�~0͙X�.�ԋ ;6馮�WvX����;6eg�;=~0	���wv��$o��G�n���;LM�`���ԋr���~0��V����9ht6�Z��+�~����'�~��ܓ�w�7'��?�v^�Ⱥ��ٹ'��?����5���%uv���0ߪ�US��v����0���N�n%i�I��ں�p�����;�2o.�^&�
�aR���/��Ӽ/����-�:�����N��^���R/s��s�%��;��
ۦ�LwwX�.�����W8�����Oz�f̬�9��GW����t�m���0	���wvᇹ��%����;=~0�����V�v�T�`z�T�L�o����\0=UT��{� 7�ź.�WvX����;6e`��W�UW�g�/������ܓ��7$�+���1����弛w\�VĤX���C�j����2@z�fɊhB[X���ժ��h[��9.���OX�Y殳��6|��!�q��Pf꜍�����i�г�,�bC@�V[LVw:�l�BB�^-�ڲ�����g�P��ۦƔ�����;��,˫ja���.5����F\��/���͉Z�۫lcA����Z���dԲJ[���
iU���ȅ3�ek����f9=f�3��L�
ۧk�;&�����?�U�38[�������n�����'�~��=?Z���]&�իCv`��ԋ9_,K�ｽH��bX�'��m9ı,�^�M���2%��x�Nla�Z�w�>^��צ�=�����Kı>�}�iȖ?� ���M&�X�%������9ı,N��}�V;e�����5��d/���ND�,Kߵ�i7ı,N��޻ND�,³"{���q,Kzk����۷�됀ֆVy���MR�����n%�bX �5����iؖ%�b~���X��bX�'��m9ı,O����H]h�,ճZu�n�C�I�����@�N~��Ĕ 9��mt�ko߽�������d5wUk��zk�^����?��ӑ,K��u�X��bX�'��l?*��İ{�_��q,Kޟ}��;�X�D�u�y���MzX�pÄbF,��"��B&lO��yQ,N����"X�%����4��bX�'~��]�"�����^����$�Yr�p�]q,K�����ND�,K�k�I��?�"{�?~�ND�,K�:���צ�5���>ݶ�4G..fh�r%�g� d����Kı=��]�"X�%���ڱ7İ?��������iȖ%�bzMB���C9����צ�5����}�t�Kı;�{V&�X�%����ND�,K�k�I��%�b{>�ɗ}�GU���j�YGt�n9h����.��Ҙ��J����NY˶H�TMt[�>�bX�'��ڱ7ı,O��p�r%�bX?{^�ȓ�2%�b{���y���Mzk���M�x�7;5�X��bX�'��m9�C��������4��bX�'�h���ND�,K�׵bn'�@ʙ������7l��42�Ο/Mzk�Y�?���X�%�ߴ{�iȖ8`����S��"�5"{���q,K���~��Kı,�wՅ�٬�5Y�ji7ĳ� 2'�����Kı=�~Չ��%�b}���ӑ,K�*̃���4��bX�'}���c�U��O���5�O�_j��Kİ� 1��~��}ı,����Kı;��z�9ı��_ŧoL�1.3,.���Ơ:��|fۅNe�z�m6;x:lX��l��f��Z�7ı,O���m9ı,��M&�X�%�ߴ{�a�'�2%�b{���q,K���_���fu�o�>^��צ��޾ק�~A#�2%������9ı,O{_�bn%�bX�{���r'�!���MN����V��^f �A�O/Mzkŉ��?��ӑ,K��u�X��c�B"w߿p�r%�bX=���I���צ�>��t��lcU�)y���bY�H���X��bX�'}���"X�%�����K�]��*?'5^���iȖ%�b~�����@ss�5]zyzk�^������"X�%�����Kı>�z�9ı,N�^Չ��%�by����C�R;,�%�)nZƷP��7n��nc	D�FR�%j�BI�%���5������v%�bX>����n%�bX�wG�v��bX�'{�j��9"X�'}���"X�%�d�Vf�,�f����Kı>���9��"dK���X��bX�'����ӑ,K�����n'�?���K�����c�3��.���^���?~���Mı,K���m9��D���j���4��bX�'�h��v��5�Mz}���&
�(4j.�<�bY�P��>���ND�,K���i7ı,O����ND�,K�׮�<�5�Mz|�>���:�P�3Fӑ,K�����n%�bX~Tc�l���%�bX���j��Kı9�{�ӑ,KĊ��b@$����6�j1r�nu��4�.�<R^��BѺ�y9�	�1ˎn�6s��щ;��6ƛh#���|MN�g��:���4�Ν���y����8X�q����Ƹ�s�JL�x��Ju M�Nnb,�×�K!��d1s�v�x��a���+�s�Y�3�W�ҡ�������l��eh鐍��9�ln{�yq�wd=:��!6�΄'�I�{��}��}�܈����aa�����4nח�jSy���9�.��pGC�_�ӟ���0v
z�Mı>�����r%�bX�q,K��}���İ{�_����Mzk�����O��b�% �8�Kı;�{V&���L�b}�߸m9ı,����Kı>�}�t�zk�^���}�o|R�����bn%�bX�w���Kİ~��4��c�!�2'���ٴ�Kı=�~Չ��%�b}���y�-՘f�S33Z6��bY� d����Kı=��~ͧ"X�%���{*n%�`��]D����M�"X�%�d�����%�̳U�֦�q,K����iȖ%�a����?eND�,K��~��Kİ{�zi7ı,O�{�v��[%�0e�76��H�v�#,���9�6�����t�<�4��y�NNY�ӱ,K������7ı,O��p�r%�bX=��4��2%�b{~<���צ�5��=?0V�A�nf���X�%����NC�D�)�	tS��;Z`��6;v�h��j�Eҿ�� 4�&�X;��f�q,K��þ�ͧ"X�%���{*n'�Tʙ�����A�r��g�>^��צ���t��bX�'p｛ND�� ?�A��j'�~�쩸�%�b_ki��zk�^�o��z^f� ��^�%�bw�ٴ�Kı=��eMı,K��{[ND�,�(L��^���^��צ�=����ͅ�[��6��bX�'��쩸�%�a��~����,K����t��bX�'p｛ND�,K�d$��)��%�ݷ/R;�62燖 7ckI��\w2���I:Wͯ���kG`UM���bX�%��ߵ��Kİ}���n%�bX�þ�l?�?�[ؚ�bX�����<�5�Mz}����|�e3i�kiȖ%�`�;��Kı;�}��r%�bX��粦�X�%�~����"?��5Ĳ~��X\-�̳Uֵ���Kı?a���6��bX�'��쩸�0�vEM���@�+$`D �h� ��;�[�L��I�@��$�i�5�빴�T�B�-~]���@	���w� q6}ń������0� @ �b1#�G u�:���@�o�:��n��@���Z�I6&����4�	>R�o�a�Ϗ�>�18D�	6������gzm�0ޙ�"��!6���1��$dc�ۥ4kH[�V�!!!'��z����u@(򢩂G�t��(�)�;�4Q�"t��0Q�C�*UQ�T�vq�@��(/�]AQ�/?�Q5��;��"X�%��?~�O/Mzk�^�?�o��j��]����'"X�~P��?k��*n%�bX���~�ӑ,K��w�I��%�bw'�}<���צ�5��==1pV�A�.f���X�%����ND�,K����~�ND�,K�{߳iȖ%�b{;�ʛ�bX�'���~������X�
BE{l�S\�7ln7=��ې��${	n�З?�>E�y�u�������bX?����7ı,N���6��bX�'�������&�X�'���<���צ�5��n����0l8 \�%�bw�ٴ�Kı=��eMı,K���m9ı,g}t�/O���^���~���[�&ӑ,K�����Sq,K�����"X����Q5�?]&�X�%�����ٴ�Kı=;l��k֮�j��kZ�T�K��2'�����Kİg�]&�X�%��;�fӑ,K�P  i*:���=�7�צ�=���鏒쵀L��:|�5�bX>���7ı,? ���{�m>�bX�'��~ʛ�bX�'=�p�r%�bX�ȧ������IrSR�4h���;��x�̡��h�X�\
���l3W��O5u���.�٪Y�jb}ı,O�~���ND�,K���T�Kı9�{����ı;?k���Kı?�}����i�]����t�zk�^��s�쩸�%�bs���"X�%����17ı,N���6���C*��=/��n�n�^��bX�~���ӑ,K��{^���c�a�2'���fӑ,K��{?eMΚ�צ�>}��opb�T-y��K���P���������bX�'�?~�ͧ"X�%���{*n%�bX����iȖ%�`�/��ڍ�33SY�kZ���bX�'p�}�ND�,K��Z����ʟD�,K����6��bX�'�����Kı?���B�ղ��JA�mJ��耉Q�5t���� �T�=	���s�϶��%����*�SJ��y+P�Ek����v�2���E�� ���5G
��^�p�.V�)hd�*��Gx6͋��30&%y�܄�
�#Q���a�;RT���<B��!�q�t��یqBv�ۂ��r��Rt��6_U���_v�h����z���΋���N86�g��8���!�%`�+%��)�k4%5]��È���K�p"��҈��%�3$�H�c��h��qu�]��y�\t]��Ai{[`��RŎ�wwd��y�y�V�@O�?צ�5�O���%Mı,K���m9ı,O��鉸�%�bw�ٴ�Kı;;���X.h�
��yzk�^�����]�!�X�L�bv~�鉸�%�b{{�m9ı,N�s�Sq? eB�ק�l����.�Xɇy���K�����q,K���iȖ?��)MD�O��?���X�%���]�"X�%�d�}X\��[�Y�ji7ı,N���6��bX�'s�쩸�%�bs���ӑ,K�)2o�zyzk�^������-0We)�kY��Kı;��eMı,Kʌ~��߮��%�`���M&�X�%��;�fӑ,K���̅�ƲTZ�wm�g��G#C;���竓8��v g�׶��if�b����������5�bs���ӑ,K�����n%�bX�ý�l?�>��,K����7�Mzk���}��LƸV�w�>T�,K�k�I�P0P��8��&��T ��Q>�b{��6��bX�'��~ʛ�bX�'=�z�9ı,e�2�&���L�kY�&�X�%��;�fӑ,K��w=�7��,2&D���~�ND�,K��oI��%�bs�����֝�֦�fk6��bY � �C"{��MA$����ؒ	 ���@���Oh��fӑ,K���/�޵���UM���^��ק�_}�t�Rı,O�}���bX�'p�}�ND�,K�׵bn%�bX��M�r{B�ڦfYc�*֊�㗇�c��C!qk��9U����w@���y5�tl�W��Kı?~��Sq,K���iȖ%�b{�����9"X�'ߵ���r%�bX�N��X\��[�I�����%�bw�ٴ�Kı=�{V&�X�%��k޻ND�,K޾�M��
eL�b{�?S�f��fj٭d�f��ND�,K��~Չ��%�bs���ӑ,uMZ)� ) T(�P�C �����E�x�/�
X�����֦�X�%��O��<���צ�5����� �˩�fkV&�X�%��k޻ND�,K��z��Kı;�{��r%�`~T����Չ��%�b}�^��r�a��
ڮ���^��ק���t���,Kʑ��{�m>�bX�'���dMı,K�׽v��bX�'Ǥ%��=;7nn��W���&ζ�� rO$i!�v���yc�>F�Zv�X�%�N���ӑ,K��{�ț�bX�'=�z�?��R�&�X�3��m���^��ק�������h�K��m9ı,N罬��~�L�b}�_�]�"X�%������bX�%;��[ND�,K��]ffx�ar�Zњ�����%�bs���ӑ,K��^�17���ș���kiȖ%�bw?~�D�Kı=�w���m֦��-��]�"X�!� D����17ı,J~���[ND�,K����q,KI���G�^D׾�.ӑ,K�������ZL����Kı)����r%�bX~@u���r%�bX�~���iȖ%�bw/}���bX�':tܑ��X���m�����f�Z����\h�6����l�,k����wM��i壒��R�
���%�`�?~�Mı,K�׽v��bX�'r�ف�NDȖ%�O{ߟ:|�5�Mz}/��B�h
�]�]&�X�%��k޻NC��(�MD�?e�����bX�%?~����"X�%��{�I���� ��5���_��	��
ڮ���^��ק�~��Mı,K��}��"X�%��{�I��%�bs���ӑ,Kĳ���=�cl9C����5�;�IdȘ{����"X�%����4��bX�'=�z�9İ?"�Ȟ�����Mzk�^���~���i	�|����,K��]&�X�%��G�����>�bX�'�����bX�%;��[ND�,K� 9�[J����H�C10z��0��Z�55����D���I��@�a�Kpuť���I�;Ne"٬v(�;���Z�9�f�Ŗ�c`͡\*rb;`�+��Ѷ�M�s��.�#D![m,�D��v�pj��)�丱�v�&@h�K��u�ɩ0���r]6،d��:ŇbPnض�^^kk�8����W�f.7qn^"y��h���J�ƪ3���)���n�.e�r�0��.��z�L�Fh^#)��-�\t�sة: �Ԯ"����˦CGt�^��צ�=�׿�ӑ,K��^�17ı,Jw�����bX�'�����Kı=�i}�$�0�an�j�9ı,N��p����j%�O߿kiȖ%�bzk�bn%�bX�����OӤ7B�ק�����Y�TҘC��,Kħ����r%�bX�Ok�q,K���]�"X�%�ܽ�bn�צ�5����{��Gf�s,|�,K?+"vk�뉸�%�b}�_�]�"X�%�ܽ�bn%�` !�]D�����m9ı,O���3%����ӧ���5�O������bX���f&�X�%�N���ӑ,K��g�q7ı,K���x��%%�e���6�ط���g����N������`��R���]�mW|��Kı=�߳q,Kħ{�kiȖ%�b}3޸����~���%���]�"X�%�g���\�rۚ��k5���bX�%;��[NC��y�� |!^DȖ'fo�q,K��u�]�"X�%�ܽ�bn'�L�^������ ^#H(L�O���,K�?~���bX�'=�z�9��P!�2'���bn%�bX����[g��^��ק���&b�q��%���hj'���v��bX�'쿿�q,Kħ{�kiȖ%�b}3޸��bX�'��/��MKtS5������Kı;���Mı,K�R8{�����,K���߮&�X�%��k޻ND�,K��>$�d�I�Ф�]թp�u��n��9��]\p9�{f�x�������Y�\�)�:|�5�X����[ND�,K��l���%�bs���ӑ,K��/}���b[�^��g��v`;W2�WΟ/Mx�,O�}�����DȖ'ߵ���r%�bX���ى��%�bS�ﵴ�g��t/Mz{����TAf�q,K���~�v��bX�'�{���K���eJуE�J�"6a"�M��"r%?k���Kı>���Sq,K��M{��.�2�����צ����45ۿ��q,Kħ�����r%�bX�v�Ҧ�X��"~��~�ND���5鯻�~惶\�P���X�%=��[ND�,K����ND�,K�u���r%�bX�e���Mzk�����1�5�
���Lɺ�q��c�T���3g�J�i@����N�|�i��$&���zk�^������Sq,K�����ӑ,K��/}��NDȖ%�O���m9ı-���L���`[�yzk�^�'=�z�9���uQ,Oe�����bX�%?~����"X�%��o�T�O쩑,O��/�^j�kusWiȖ%�bw/�f&�X�%�N���ӑ,�HdL��_�*n%�bX�~���iȖ%�`�wՖd.��R�.����bY�P dL=�~�ӑ,K���7ı,N{^��r%�`i�!+�P�$B06��&<:��
~���o3����5�O}���e]X
fX��"X�%��o�T�Kİ�C�k��]�bX�%�쿿�q,Kħ{�kiȖ%�bR{�Қ�O'f��ܭ�d⧒ |�I{����Ħ�G��&���ױB�����k�w��d�,N{^��r%�bX�e�q,Kħ{�ka�I�L�bX�����yzk�^���{ߌ1v�uv��bX�'�{���?������%?~����"X�%����eMı,K�׽v��� �L�bY�C7����s�C����5�M=��ϝ9ı,O�}���X��"dO�k���Kı;�߳q,K���=Ne�i���\�fk[ND�,K��l���%�bs���ӑ,K��/}���bX��{ߵ��Kĳ���2l��AfA�����5�s���ӑ,K��/}���bX�%;��[ND�,K��l���%�bUoTXBe�9�}T �}��H&���t���wZ�e�9�h��Gg�89�m��+�e�|7DHA����� `Fh4�Ԧ#�X/F,��{k����B�I��1r���Dd*�!!(��@RP�=X��*|>(B'���H�	��7H� ������ӄ����HB�_��@O�Ǐ�'L��~دM i�0H�@0B(4�!�"ss�!�$�b}���Er�u���;R��i-V�4J��-��HNw>�S���;�����" ݌�ɮ5®�6e8Y���=�����4.���T��]��l�gh+n��Y��X(��[l�|2uE"��-���7EY`�1�x��2f��#���\U�o��3n�J��]+ݢ���^T׋r��)�Þ�)����]��2��J"��f4�`Ω\`����`�W2m�$�z3T�q�����ؚ M���U��:'���F�=M�Κ͇�b9�Md��R�}#�f+�ܖ�*Q�v��/6��`�IS;�]����ð����g���p���m݊��j�L7���k�Mν#��4�d�A�Ԧ��:����4.�y%]+�v��7`ˍ� �������b����#�Zí8܏�W���Fp��e�努���7���:H�0�����qg�a�J��aD�i��֖��z�r�:덮�����	,=�v��l�vtK�����,"Ũp!)E�8q�+y��$-ћ$��ڹ\'Vz�L�M��a�Oh�$\:,(p%�7��in�^�U���!������^�k#n1�6�m٢{Z��AR��q9�Lз;�<m\9Y枒��s�G
Risn�6��G���yD6�ge��l8���t�.t��H�TY�5��E��b�(.��Q�e#䶱՘n��U�S��C�����E�+�Z-u�/W,��۔���Z���iIʓ��Ta���jY�G�B���̳m���:W�T9�6KnWm�6�D�:�z�A�t�C�ɕκ��6��v�j[��<��i�GnYkAh�Nz#��Eh7[;nx�b�uX�.�`�e�H��۳�Ie&�F�p��%���ݤ8{l��t9$�V�|C84b*�x�J��*��Ɔk�h	�6�4��UEӰ5Uz�sY�w-��X*ۮ��b�&R8����;��t��B��p�T���X=U>�@�A^��F+�M
i_U_����(��vJ�43�kU�r[��b���h3=3 =�M{e�v���D-�٧�kJ!�{�:_9��/,v;t[�Fó9wH����=�L�Y<٬p�JҤ&�vH76��B�F�B�ur)юڙ6�݆�6h׌��.�iNm+�
����{]x��Ѷ!�g�Y.��T4 �H���\�s��vM73�r]��[��%�i��t���e�ݧ���rG�w5����c�r���SK+`�.ŀ�)E�{�q�4n�2�I��|���5�K�}�17ı,Jw�����bX�'ݾ�C���MD�,N�k���9ı,����̅�����u���Kı)����r%�bX�v�Ҧ�X�%��k޻ND�,K��bn'�ӿ���ޚ��������
���]�"X�%���_Ҧ�X�%��k޻ND�,K��bn%�bX��{�Ο/Mzk�^�a�� 5C jT�K��2'߷���r%�bX���ى��%�bS�ﵴ�K���2'}w�T�Kı>�߲�e�1�����:|�5�Mz������X�%;��[ND�,K��zT�Kı9�{�iȖ%�bw-��̚�Ns��y��m/�P��v���=.�m���a�ω|x`^g��7�Ѧ�v\eP���ץ�bS���m9ı,O�u�Sq,K���]��O�dK��_~�M�k�^���}�~���k���Ο/%�b}ۯJ������V�: �N?D�Kߵ�ݧ"X�%�����7ı,Jw�������2�׻�%���2-�<�5�'ߵ���r%�bX?g}t��c��ș���kiȖ%�bw�_�Mı,K�v���MItS5������K������Kı)�{����bX�'ݺ����%��ȟ~���iȖ%�`���X\�������]&�X�%�N���ӑ,K����J��bX�'߿o��r%�bX?g}t��bX�'�O�r��MK�E����δ[��:�"y��F�8A5�;t���.�++�\�_:|�5�Mz��۸�Kı9�o�iȖ%�`����"?�_�j%�bS�����r%�b[��?���`j
��7t��צ�,N{���r��"dK����n%�bX����[ND�,K���ߥNr��s�.�^�H��0.�7a��92�Ḍ�~�t��L��S"a���fӑ3+DM@5��!��sj�D,L�N��ҧ9S"fTȟ{��ND̩�3*d��9}�ے�j�f����*dL�������~��m92�D̩������Tș�2'��9&ӑ3*dLʟM{����3*dN�OY~a9��n%<���нt��oҧ9S"fT�~c�~��6�D̩�3*vk���Tș�2&k��m92�/@�=�z�]�5��r�f6z1Nr��\,��i��fx��z1�.��Gv�@X�����нt/O��y��t�x̩�3*}5�\Nr�D̩�0��f���&�S"fT���J��L��S"~���y~�3A&�����н���������Wq7�������r&eL��S���S���3*dO���ݧ��7B�8����cM�.n�.z|�L��S"a�w�ͧ"fTș�;ۿJ��L���S{��������r&eL��G����Nr�D̩�;��sD�\�����>^���u�wO}�?\��L��S"w���ݧ"fTș�>���'9S"fP��>�#(j"p���i�iy�v�< �(�S�'��Șs��ͧ"fTș�?��ِAP��>n���z���m�r&eL��G�{�I�Tș�2&�}��r&eL��S�����Tș����;�I����7�gM�HH�c᭸��O�@�+�v�uhY#�<)n��Dn�z���QU�aU������z������>Tș�2&�}��r&eL��S���S���3*dO���ݧ"fTș�}w���^ٻ.\���t/@����m9�?��u72�����Nr�D̩�=���[��Lʙ2�������нt/O��{��'2`�	A�m92�D̩��p��Tș�2'���nӑ3+�j&�G����9ʙ7B�'���Ο/@��7w����+��3Z5��*s�2&eL����[��Lʙ2��������3*dL;��Y��Lʙ�5�����S���3*��i��|l��	6p��O��n�L�?k޺Nr�D̩������Y��&eL��S޿�T�*dLʙ�o~�iș�2&eJ���Cȑ �)��exuf���Rsa�Ҽ]@  �7k�6��R���J�㵄dsc�͋<�9�pCs���@�<D���ܼPaP�s��ph�l\8�N�;t4sBU�����S�D���5�q�-]v؟Kҁ��ۛ*��{`p�m��xH�wFMٻt$Xq(�x/;��]�=gut�]�������ʹ�.�d�$�$�����D��4�,vwn��u�pel�v8x�̡��`�Z��͗\�[�9�|jd�jdLʙ=�~�m92�D̩��p��Tș�2'���n���obou2&eOM\Nr�D̩�?~��\ÉrkH�*y����z������>r�ȨGQ5�������92�D̩ٯ߮'9S"fTș�w�ͧ"~�t�ǧ��n�����C@T6�9ʙ2�D����nӑ3*dLʟM{�����a�2's��Mı,JUn����r�T���BIRt���r�^{��/�I%��I%�����$��bI.��bp8��]��ݯ�@��X{�+ �\� ��E�}P)�ƈ�;@S2��Kv�K�ؤ����0�ix����R��mcc��#��7�}������"�>�~�s�ϐls� �[��LɭY�7$�s޻�>qj��L̟c�`W^ŀw�2���9Ib�V/YB�T��V��u�� �kذ�fV��պB�MRVP�\���WԹ�n��X��Xz�X��\r�+t�ժj�`�X��Xz�Xk^ŀuT�I�t� E�w˾Xz��Fc:�C���L�A��Mr�5�&�UHj&�m۶�n��Ȱ�Ȱֽ��}���p�w�v����vT��r,�+��s�Q�,w���>�"�s�i����i�iWm����ﷀ}���s���B1@�	"1جC�*������5�,�j�-�����n��ɕ�}�E�}�"��Rڗ<�	��4ݪlNˢۺ�>�"�>�`�{����>�J�Ө��[WJ��xr]�Ls �1�ڵ������c���ভs�g�b�(WJ��Jӳ ��E�v��X{�+ �e� ��!E"�e
��+��w^Ş�s�T��=��vz�`uȳ��&����[�T��Wk ݞ��>�p�>�`ױ`�"����m۶�n��Ȱ��Xu�X9Ϲ\+��W+��̬�Schm�WV[wvv���Xu�X{�+ �\�~�m�}�zKy��&��t�Cj��DK:��<��攌v�z肴;��	c��rՓ���w^ŀw�2��Ȱ��X�j(վ[9we����;ݙX��X�r,��,�Ur�&���v�;.�n� �~��>�a�Kc�X��V�v�ZD��t�ۤ��X�r,��,�ٕ���+�]���R(vP�LB�Xu�X{�+ �eɹ'>�z�I��bd��B��C�M@�;�r�*��FYDL��vŶ��J��\و�R�鸙�Ƒ�]9bZ���gN�.%��:wZ�c��sM�O;J�8b \�VG;�ǆ�9y�x��h�3��ڸTƐ�[ظ�U�C�<�E�=M�l�eZ2.A֍ۋ�^��(2���y���94{q4�'�@������P���q��1�R6�@�7��Š�JZ:�'N�}�N�'�:?&���um%W�k�5��8X�-��>�A��m����R��\�m�n�ֺ�e`l�`uȰ�ذԑ`��V6��m7wX�.�$w_���y`�̬�]���n��-��v`uȰ�ذ�fV�ˆ���*�t�ݴ��`��0�nݗ��ڊ5o��]��lN��ۆ�\� ��E�w�p�'���C�R�]�g�1��a��ct���9�;q�R��^I��$l����l��ـv=� ��E�oe� �ve`nҫH��uv�;X�r,��NW+�`�E�� �4�lr�UU̮s�2�\0�fV��,�t���+�����ٕ�uM� ��E�N���wJحҧV�ݘ{�+ ��\��W�g�j{�5cmݴ�wu�uM� �\�s�����M���;ݙX���ݴ��y+y��p��:(\������]tPpGGN��y?�IH��j
��i�����`�̯�U_ �����13�B�.�N�����I��X�O<��5o��]��m'srO��7$�����/�K��X!����H�6E�٭�L�|�A΅��S �l��G�$4$ ,#�bċ�x���٭2ŋ/6Tn��ϕظT�r �ak	B!�[��||��!��$!
x�6m�!r|ЯD�D��j�$��a[]z�o���S�S_r�HkM��H BX�@ٲ��(��<����L��1�:�f2.؟!bR� �!4Sn����m�VT�v��6ki<&�)c�a1�BM�����byO"��>D��� O�𦟕���(���.�k7� �.�P[��I��v`~�r���y���,{.{�{���R�.�nw ��w��{'�O;������`Sc�7eԠ�Z���gEO\mnq,b��s��@���]ֱ�� ��ml��YE"�e
��+��}��ۆ�6<��m9@�
�aj���n���#W���~��7�e`���`�Um��7wXT����X�L��ٕ�F��T�����ݼ����+ �ve`*�"��P$ p܂�`�`���'n��ܒ{��r\��WE�i���7�e`�̬�lx˲<�"i:fSB����V�mV��Y�,���Мk�zg��Cq��ͽc�uv�J��fV�6<����+ ��-�K.�ݧE�u�uM� �vG�od��;ݙY��RD�EZG��]+-�i]��}�od��;ݙXT����R(vP��Wo �ɕ�w�2����{��}�uQ�J~�4�n� �ve`��s_��ğ^����w�{f��Fs� )��0Ģ�2�lM1@��^�������cV1�)�Axes`!�&ѻv��Og��i乸'�Z�k��Y�θOd�A=���9�������j�'{;Lu�`lK�*�q�Vv68z�]A����8�)4ң+���{mF�N�%1���Y�Ug%՛qv�	�J<]�"9����L⋡�i������{<=��\
�=n�qj�����5��	��L��R߅^�҈�>T�ٰ&�4-a6�lw�<�+ ��uנӭ�����iZ޺պ�D�A����/H��dx�2���~0��m5WJ�n����>]��l��;ݸ`M�=\��|��ת�t]�����Oe`��0�r�����:��xѕ�Ek��]��m]��r���Հyzy�.��	6e`ݤ[hr��ݺv����s��^���=���ٕ�mm SPJ�N�,UWv�t��%v��Q�5rg�"R�,X�8�r0�И��un��i]���&̬�ٕ��\�����C���B�Li]��=��f�+�|��� ��AH�K  px'���}�r���>]��*:VӜ��I�M�`�̬)��.��	6e`�B�SI�m'lm��?Us���� �y`l����g�� �'�M6��ݶ��]�xT���^����{�XSc�;R	���Ch����n�����;m(��4�8�F�n�:�72�P��2�ݷo �+ ݓ+ ղ?���{� ��'l���H�n�g ���������#�$ٕ��==H���wE&���wX����$x\*�s�«�0�$@B!=��f��{�rO����
�Fh�w�<��������y8�`M� �����:i�[��I�+ �ʒ���^�xT���<�����n��_Y[�,����j�v�W ���i�ӷH����x��w�����s��d�$�ց����XSc�:�� �fV�6�j�I�bv��Ǟ�*������=��uȰ�dm�۫�jۻ��v��#�$ٕ��\��~��<�<��GLN�Ql.�vݼM�X�`M��s�*��9UU���5����@Y�lZ Eb�ҧȠhx�������|�'l���x�n�g ��w��I�~�����$ٕ�~�s����Z�y�=8�N�9�\����g�7m�up!�\Pl���}�G6SmL�%��ew�=����>�#�$ٕ�W*�����<����$�EX��]
�����v�l��I�+ �dxScϹ�r�����8�ĊT�v�=��j�V�^ ow׀N��PЭ�Ln� �dxSc�	�^����� �zx����Ю�hN���l��I�+ ��X���	b$A��K�Y�W
�n3�f������0e�	�j\.��Y7l;]06G�'�\�GHe]�N�N8�n/`9���y��MA�*�8ඪ,]�r��vƯ�gq��G�
qvedݵ�CrbѨ�nb5m�d���q�NB1zi-88�*MHYZ�;%!�8�Y����tM0JV��\�m�� �٭`����2<�p</me8���s�ﻗ���M�^۪���kG.�n�s�e�ku�3;@�[e������+灃b�n��ۀ'� �fV5Ȱ�ǀ�A���n���[��$ٕ�Mr,)���/=I�**^��VUݖ6�� �~��${�U�RG���}＜���7[���gy�o�UT��X���&̬k�`�R�t+�wC�J�`l� �fV5Ȱ�ǀj��i���ҾH8�6���p�ՙC�.��ט��5G]�/���b�j����z{+ �dxSc�"�:�U@�hn�`�f��={�f��
���c�.O���f�uOy�l��%M�4�������)��l�ԗ�=��yOy�4�����-��t�'�N?�߿<��~��&����(1K���.�.ݼM�X�r�s��������~x[#�?Uv���JH�[t]��i^�݋���6<���>n:ғ(\q������c��T��ڬ����xo��p���ve`��[r�Rn����"�?r�����y���X�E�vij�t+�wC�-��"�<ṋ�
�J)`��G�@b���D�1,z�R�b$�?��>E�5���]�"����� @;,WMS�Wk�*��W��ՀyI�E�:�X먪�+Cv���`nǀ{���~��r����Ϡ~���Mٕ�E�&�ڎ��r<�lE�1��%m(ɓ�ƮL����8�D����ڛ;4�[��;~���N�7fW��s���z9�uBy4��(�.cs�������%��＜G<��#�W*�7�T�~8p�E�jӷ�zOe`ױa��ʮ%���:����**R�]YV�m]��{/��nI��{7$1dG(�2$`|D�,� �[iP �s��Ov��H-�ߝ*M�㻻X]��-��ve`ױ`鴭��Y㔳$^��f�Σ�q�s�լ��xg�g5�b� g�K��p�Z� �-��ve`ױ{������ ճ�e��cc�xݙXu�X]��-�窸��u�^t+M;iІ��y`vG��%�=�zOe`�S���lN�����/=���=�Mٕ�������"��m�wWiݻ�N���7fV�{I=~��rJ|+��H�� Y��X����hmc��l<#��B M�x�IB�0	ZY���3:���!FeK�&K$�B����d���4^:$��@�D���>t�"`@1H9�MF� D�R��6�XMړE�D�"J�E�UO��z6��dCo�8x^���) ���� dXY���D̓�c	�(:���.���JE������Mq�u֐uj4�S S�������!�aaX�`YrVH����_�:ma�<)���"U�̞
�w�g4S����<� D� ������#	!��������a��|"��4�Ԅ$Bc�� �	���"u�`�@�2) B9�Xߩv'����P,2�Q�C�!	 P�+E3���jf\�eؗ���K����v�XQuU�$q�,FДt��H6��+pK���z�6$ �H(�# �J�eUSf �L���s&��U��m�v�ե#L��kD;*ewE4�[9�����v�7Az�C]�{�����jLN
��[6���EeB�;b�����8rV][�ٻY.��0����ur7 kt�*P��=�<������9tzP��pV��o`�ް:���B�GG7o&�:ԩr��@Ru�pv��*۵ְ�)���d��H�x�ۋ�pҤ���D]͌i[%49�n���Wof	̦ȾwH�p����x�c����m:2h\�����]l�ʽN�[���C`s`�Pn��]�����NCv\�)U�5e�(jz^����)�Zz���;1H�v8�h���d-��������ɸ�^850�
4%S���X����]��K]�sҷ�hh��Mn��u�0�d�;�A&�Eu����֝�\�8���k���f �*��-`ú��j#��A.�ʱ��Jf{7�4NTEVfV;x+���ܑ��Umr�;N�A���IZ��T�1Ø��Y�-N���1���#��؀GT�oTݎ�\J��Hl��P�Σ{kX2v�N�@��]+�sn:&:�+��6�؃h����#O��6L�f̓e���0��2�G5a��"܄����x���R�����b�r��mk����7\��)�	Y�Kl:�m�biF�@�JP�O	��ya@���H\������!ْۈ����:蓵�K�ޖL!��2�WNºN�WI���Yay�mI�:˷�j�H֨ۅ������{Iy7�A]%]X��vm]%�k���ӊyB��v�3��GN�)ѩc�s5�����v�.��r�ӭ��gS�Ơ����MUV�5UPngn�9v�v8̈́)���z�d�V���[���ꃁ�&���|��|�bQM��L_"��Ġ���4( �pG��!L�A����ׅ����R��ep��Msڋ7*1�V�tPV�4��A�̴E)���KFc�p)���£�::+p��!�F�k+���mJ�2�yŌr���dF{\fp�l�+�(N����t\��B�5��7Dj6�W�㎱�9v�A������=j����&xж*kXʉf�u����n<l�,����l��Z��������f�L̳t��.d*ۍ��9�Ф�&��9��6�׫�a�f�e.Hx:uvw ���y8�ذ�#�\�~�+�5~������J��9vU��Wu�n�� ��<�$xݙY�$wg[I�:T���wv�-���<n�0ױ`�Z��*�#����y<�w�������7^Ł�����y��x �鶩��xݸ`�K�_���>RG�{����!����mk�OK��G۷g����Ekv(<�����w�}�lJ2:�΁�?~X]��)#�U�I~0	�^Yi�7m��6��`vG�
�(�hPO���ܓ��7$�w��I������n���s��>�{� ��u�X]���U��(�n��շo ��V�x]��{<��~�}�p��l,���G)6�8����#�>RG�Mۆ��\�{���~��m�f4�e�D��#�����Q�
:0�B[��Zn^�����!>��-�7wo�~S��|�� ��ܪ�|�^���?~�6S�0�1�#��>^�� ��+ ջdy���U$j��JdFm��]�=�}���oݼ�"X�(�;AB�Ef0q�*�%��=��v����=���h�؝��CwX�\��� ��y�-��?s��qzO}X�y��m��cv���]��-��	�2��n��Oн�f,�8�`ԅnͬ�^� w2��>Mt,�X���D@ۭ���Q� cQV�;�'�7fV����s���<��x�x��窋t]���xݸg�\��H�� ��y�-���W*�#��e���)����{�Ӏv��w �nǀMۆ�w����T�7o��� ��<�7fVҕr�q�UW=����p߽����*�e��p��xݸ`n�0�#�;*Q��
t�[�=E�n�+C��G}]�8�8���k�����m�S�DX�s�?`='���.Ǳ~�U|�u�,k���wJ���wf�e�?��<����n��I��e�ln�.�i�f<��ݏ��9�RS��`{�Ӏ|����Kt���9�o׳� ��� ��b��r��+�߳ߖ���V�|�T+�էo ٷ�UW+�s��'���>[�����s�\�FED�=�?Z~�ۗZչ��Z��td����W�I��.tj��cT��Md���m$Zzg��6�G��.���=9ن+��!����\B]�K͝�^�v� ��m�Q��BS,�hp�v���;ql�(ܦ�N��"�NG�����d�6:�m2�a��=Y�@<���Q�qn^��y��>7��}��!vY�u�\��=r\	Þ'v
�@�t���N<`b����iZS\B����tv��z��.�pY��V$��4z��vSi��>��� ��,��*����XvqR���T��|�XǱ`-���2���X{*�""�We�Ң���>[��6ea�r�.�~0	�<���Ie�-��j���n۷cذ=\�.�<�	���&�:���ۆ��X�v<f�0�UW)W}��"ӴՇn$8�m�^�U�3;����ti$��z�8%���c�V�;
˵�'�;�ﷀ|[��6��~�s���_� 4���r�Z�h������}���Cɼ��W�qr�F�}0�\0�b�$����*�t]��;x͸`wn~�\�8߿?~X��� �v�%JY˲�ݔ�v`wnǱ`.�x͸`�qRƕ��wW�]ـl{�W9U]{<�z_���� �� ��$�
LT,w5-[(fabX6��ɞ:N.n]����cMe⹬e�V������n�ۆ��X]�$�2Ֆ�n�wo ٷ�r��RGv_�y�,��u��&�:����znI�g}w)�M���kXB�Q�D�1T�'T�	@0���s��'{�znI߽��U5*�0�-��;�M�����oT�xf�0�n�ݍ N��˴�۷�|�c�;6�}�b�5vC�o��]��49��c������u�g�6��i�l��E����N��m扱g�
��5m������,Wdx�v<��bU�]�n�ӳ �^ŝ�UUr��"�VT�x����\H���K�R��_wf�g�n��;6e`n�0�U�D�j�wWN�ݼ��*��"fw���nI����7$�{�Mȝ�X�2�?�����'/����0�e���]���2��n������x��O���/�m4J���=��<mX����A��2�����;�����w{���26�:�ց??�� �� }�/��\��{+ ��<uv�ݶ]�&�n���< �v^ٳ+ �^ş���h}?w�h]��)�w >���ٳ+ �^ŀj� �*��*U
��;m��~[�0�<�]��~�O$��{��?tž���V&�' �v�j� >ݗ�vm� ��jSNk��5qB�U�SL��n��]��N�8WknKs��tkv�5�K��6a��]�6�\p=���u�!9G������8ֈ���Ʉ}JkQYݭ �u��UFk(�&α�m�,������l`��&�٤����&Y�)��=m��Y�آV�ѻI���J�r�]�
u�,g�����k����x��kyp���	�H��e�[�L�e-j���l�����vbo\8k�ynJ�<	�&�WR��>mQЯ�T�w��\�a��UO�v�����v^ٷ��Ur��=�O�j��U�M��;��we��p�>��0]���-�Bj�M5Bww�o���>��0��s�IE�������\�v��B��>��0]��.�xf̬���.��˻��iـj� �s��u������ۆ���C{��qP�U���,m� L�m$!��]x��m�`VmRX*z����|����p�>��0]��EV�eJ�X]��;xf�1�*��8D��0j.�%L@���m4eF��1��1��8�7��yOy�.�y��6K���vU�Ս�fݞ��5vG����).��x�_�waIbiڥM]_n������S�g�� �=��ݸ`wfV�ʵHQ���J�`.�xwn�ٕ�o\� ��M����VV2����h�e��`E�P�K�gˮF�=ѵ�}�y�^Ҙj7]e�w�?{�� ��p�7�E�|����\��`Ӵ�wf�v�o\� �wc�;6��s�T���其���7cm�fI=����I��}��5�=gp��@uEp�)������0�L!a�GN1��t	�
m~3���R)��{xbp�������!
%����f�`��M��O�6�����G�M!�D:t�Q�:C��ʅt|V
&¬P� xP�qy��d�`��m$�.��.��X˻ٷ����\�qM�y`��[I�
�mZv�͸`wn�Ȱ�v<�9�Ԡ��:U���'\�2�u���[o,����ZYz� n�,���x���
G"mr|���ذ�v?Ur��+�\�	����?O~)cI�t�������7�E����:�y��~0����j��Bun��]��ݏ �ۆ����Gvz�	��X]�$�2Ֆ�j�wo��L���[�w��������T�)��{�nI����nۤ�i:�� ��/ �*�s��W�~����� �ۆ��&�����7Pޏdz�{.N�x3w(�R�5*]��a�@A+ll+`�ջ`�q�lm��~����>]��͸`u�X�I'Vi�v�ݬ�ݏ?W+�+��6O޿�����7�E�����yU��^���t�;x�_�W9UIM~��:�y�щA���-�ciف��������&�y`�ذ͸`�8�!ݺ)������7�E�~��W7ny|�_�$���]�'�a�����jC�]zuӻ��X{��LU�]���	&p�4#��M���w}���AȳJ��u&i5 �F7�>�al��Tpu�um��JM�@�ۉvq�y��X:8�ɰ�'�q���"PB�Yf2�`�
Yt+�m筁�sl&�:�dcv�{r�Q���E��ݧv4�E�e��*Z��9ږ���eXb��c8�'��veӳ��^An�E8^1Z�@u�`L�)����N�N��w����k�ۇ����jLB�M*:����t�k����V �g��ӠF��@�?y`�p�>�s��|�k����HMU�-4�6��ٷ��r,�{޺9��av�Bـ}�"�7�E���T��X�_���]4���7V�m����9Jm�� �s� �ۆ�\� >7ci$��պWv�n�޽� �\�V�g���y`�"�;Z5���j��v� �b�c��ۄj�����8���z2���x)�ҧhம�)[��vm� ��E�o\��9ʪ��X��x~|.ʶ�njnIϳ޻��4D�]%D���U]s�*��?j�7\��;6�od�X�v�RWW����o\� ��b��+�K}/��s� ����%�cNӫ�5v�=\�����+�f{��'�_� ��b�7�E�E݂HMU�-���Xf�0��,z�X�{�i�QV�H馮jأ"(k�r�k4�Y�k�(0c ���*�Y�i/�ӻ�e�x�ŪR]Fπ��o\� ��b�;6�w�G�M��cum�ݬz�Y����;�y`�~0��,�W*��s�UM������ut5I݉[v��ߖٷ3�\��\����`�y`EVҨZ�WWi�-���Uqo�x�;�y`�"�>�ذ�Ġ��)$��>�ذ�\�rm���;�y`�p�?W*��_��'�Q �,jݸfxz�FP�����p<7�m&��m�%v�F����k_5�� ��b�;6�}ױ`vRM}��Fje�[~���?wN����������6?~X�ȳ�+�[<$��Z�h����7��`u�X�Ȱ��,�tr)m�av�Bف����.��,k���^Ł\ʕ�+�#�hM&	�h:��6����}0�Q��n����[i�k ޹���v��o���>�ذ�KS��͹���e����s<�X���>MzK��v�r]�oW���w&~�P�kѥ����vm� ��b�7�e`EVҨZ�WWm��k �ٕ�unǀod��>�"�;�D�P���X�wXV�x�L�?Ur���S{����'�~��'d�X��)RWW�����2��Ȱ͙X�K\�xw�n��]���WHwwX��X�U_��~���@����$�����?����{aA �CJU� ����G ���0��9�����\�@��C�6�i�R�8����3ڂ�g\�����6�� Z�� �&-�h@�X֝AJ����DjE���r��ͅ�[��>-�wWX�댬@�q��V��ˠ��,� ��Jʻ6�Ƭ��n��`���
��6	����ԝ�Fӳ܌:.����l&����D'�����rk'|�;�Ye��[��F�j�ۅ4$]I����6^�c��"-�{m���' ۱$&���B|�_�߯��:�c�7�eUs���;���G<����펄;� �ݏ=U\���O߲����`�p�;أ˦�7v�ui���{&V��ٷ�v< ��En�utWuh�wX��Xf�0���=�R��}X����V�][lE�Xf�0����X��X��)�>.0-���hzq(]ZW����1>�t'u�!�<���̈B���-Э �����X��^����_���q,Vݔ�[/����7�ef�|�*��r,�nV�y���q#��H=Wi7c��;����� �ۆ��%�O<o���uw`�U�����X�K}3��O<{&V�e�� �ts���l.��C�0����X��X��zpd�y�����m����|#4:sn]Y�T�6�"z�tc6$�z� E+[�~����m�i�ݶӫM���O߲��Ȱ͸m|�V�`��mН]J�]���V��� ���+=Uʤ���6��[�؋v���V�ٹ�:&�#)V UX,F	+A"��M=A]��ٹ'��XtbH�
�[�Wfջ��+ �l��UW9���q����~��q#-ۦ:v˦���ݙX��s�{��;�~0���� �t:%>+n,O��xK�֞Vg;��S�L�����nB �:m(�m�:3,�/��p��� �ݏ �����
6;Uj�!�����ٕ����F�<�	��X�dy��;��y?7M��n� �'��ٕ�|�G�}6e`I�ӡ�cmզ�v�?W*��� ���>�2�O�PȂ�����\��ܒ{��n�ut+��;wX�dx�fVջ�ٕ�n�M�5O�Cm�O���,0�7NW���(]��blv�g�qI�<vȬ�\��i��>�2�����̯U~�r��W�~x�bH�_��[�N� �ݏ ����>[#�>�2�	�8��n�;e�wv��̬�<=U\K����5I�}�J�Te�V��]1���>[#�>�p�:�c�7�2�킍��Z�6P���>�p�:����;�}�rN^�ٹ'N �H �@w�����@��P�A�a������!D�$0�:]�K����:|�6z������P�=vcT ��]��|��b|eI�ӷ������
�  X��KBĤq_��(/Mc�;�^1J$� R��+f��2*T~��@�BbHō�î!��]�QЬ�8lN��D4#���:6�1Hu�8�v@�(&�~da��!BH�PY��mX�L�]2ƙn[j�UA\U�h��j��Q(m�CEdk��*�탋���n\��\�b��v��tͅ��i�s�HM�-!�<�����FH��&T�V亞�e-���"��̹��;&5�]�`��u���"h�"��l�9v���Ip�e��Ds�;�O�ɘ��:�p���b�=�q.n���G0�H�5�؞Y�/V�&�[���{)tn��n����)ã[]�q�r�������5�VxK������8Q����6(ɖ��-ۙ��#��g�Lr�X�ݑ����(�,�m��W��r����a�=�G\F�vaC�����q�jp96Jԍ����WfL�$�1�@�)m�(3�Sv�s�9Z���:��Г�0\u�XW�i�E��t�=��ݝɧa��R��=Z��I<2L�u�+�kx�a�Or����{�X��r�Rm/"nWէ1��:Gp�'吞�v8���#��R��p�9R�ɘ�+��GgA�Q�MEd�p6LM�Ek�\��ڄ,Ys��`	̕=��V���,]VWP%Z.GsR��\tC;*D\�Q�P���Z�6imӳΝ��^t�'F�:�Z�i��X؋$Z��RH��p5�7cc�`��h��v,�(
.2� rjE��h�e�m�v]�&�zl��]O����݋�ԋD��=x�:\�c�]��G,���v����[Ep�(:���k�ݜ�vWK"�by�}�����h�b�ʕ,v���TV�����l!eT��f�[q�Þ��� �����gGI��)���,e0�NӋqw;�i�U`�Ö��k�
�֣Kʶ*�,>NMV�� ���U�DK\ù�tr~Zx�ݰOVl����ŵ�q�����Xcg���u�u�G6�A�7�)��qf�0X���ITU1%i���h����q��E^5J+E�R�U\E�cF�*�� ��5�ޭ�4MC2au&�EO���S���B���3��H"� ����jQ ���=W>D�� p��ۢ}>ə�k5�2랻&�%n���I�u!���K$GO��#�l:�[�U�4�]ftʶX��\R�)68�&X��q+*����\���fz����Z�XQYĳsn��F�˂�Y`�Ps��o2$js���%2��\���Ӭ,��u�ɞ��9��La�v콬�U���ڋ����yyUwe��t���Q��.Snm�h:3��m��;��$�ylCy��j�s35g˼�p_"�T_j�9.z�q�a��s����w{?v�?/6lt!ݚ��ߞ�ٕ�|�G�}6�}$yui�wV�ui���{�+ �l� �m� �ݏ?��U����߿$ĝ]I�hv�^���M�X~�s�Ij�� �=���#IB�pv�m��>�2�����̬�]s�x`ė��t�ē��:�c�?s�g������>�2�	R��UҩK�^K2\�`�K�-��Pwq\9��Nqt�;��R��"�h
�[~���������̬�v<��UiK�cXk35�rN^�ٽ�'� `� !R]2*$�І���['�e`_���ٕ���\�$��,��ة�����Oe`[��ݙX�dx�tr'��펄7u�����~x��e`-��~�+���� ���-�n鶝Zm'o ����>[#�>�2�����Km�Zn��܏��c���I�:��8�zU�U@ݵ��5l�6��0X������w �6e`[���r��==�+ '<�SU�k�J�b���M�Y���Uq#T��6{+ ��y#�e%��Bt�ē��N�~���w��f��8��4�P��P�"�ɉ���H@a�U_\��ܓ���f�>�w������v��~��� �=�}6e`[#�>�b#�bN������dx�fVղ<{�+ մh�"�"G7M����#n�n<lp�'�c��r��f�mzkHl�V��˼
آP4ڊ|��Oe`]���p�>]���G"��*uv�B��:�����|�#�;$��>�'��I2�U�i�x�`.���*��{�X��x_o{kK��F�����O%��{�����f䓝ﵹ>ބ0I"i��W>[�����ST�9t�+N��&V���'��$���>[��]
r�i�7����RP�<[ɋ7!���c7��6.,���c�p�!]w���v\0��xd�X��)c�%ٖ�^��^���I->����?{����e�ꤎ�U��jĝ[��+v`Ry��ea��U\KV�<O_� ��Q�ʻv�ڤ�v��2���x�`.��룑Kn�:�c��`]��ܓ���:��xd�nI��O��?z~�K���̚��ԦL]�y�t
y�p�ۥl�ns�،P�:�w���z�\j��Sl�NAg���� .��gm���v����q4��������ݲ�ήxf��c=\r��֢{wW7e{#�Z^�p�i�]�o@ù��Sd��t�&�G3���%B9�������&ׁ���Kf|�C�]&��X�r��h�jr!mҥ����w�I��D`R����#e_%2D�W%�r��.GW&t���[�M�N���m��:Kb�V�v��e�0�dxd�XWv< �dJН]�|�N���~�USd���V��nˆ~��A9<Ʃy�v��o �z�`]���p�>]����Q�
�Wj�Wf�ݏ ݗ�����s�*����� ������UXK�.�w ���N�vG�vI��uwc���M�R�HKI׭�y��LiNݓ������`�)attr���9.â��N���w ���0��X�`݄m�S�lm�ٚ�nI���M�B! *yUO�&a-��I��|�#�;��*6�t�ݷI��;ױ`����][�<}��}$n���N�تնݬ��'��վ��;%� �^ŀ|��t��
t��uv��˲<�W+��g��ճ� ݗ�8m��uWm��+iX�{)�1�����/�	��}v ��ō��=�Ҡ���m�Zv��2���x�{�:�T��������HWj���`]���p�>]����N�)7�wn�M�&���7d��>]��U<^�E��\@�oi�!4�I���H�4��/�~��~�����ꗻ9+�Ee��/׾��==~0��X�2���6�)۶6�$;��M��{6L����O��ⅪT�Un�nꚻ�*�E���r'c��قШ�Q�0���k6�ЩݷJ��>u�,l�X˲?������{��[����U�m�X�2��dx�p�;ױ`-�lI��:��]]���>]��e��n��z{�X����UӶح;x�%��߸nI��~��=�{f���,-��%ms��w���x����D:��Wu�|���d��>]��	�e`��O��v�ƳL��2�`%M(��4"�XY�2hM.y�tk8�`t���+x#T��`wo�6{�X˻ݓ+ ��b�>�V4�ն�]�m]���ǀwd��>�ذ�Yꪤ����:���`�B��l�����,�&V��ǀltiݎ�;��Rn� ��b�;�e`.�x�W)l���}�'�����[m��;�e`����=�7$�����8l?:$J�J���xe�aی4T�7P4�[X�]�3���G��S�ԖجJ�\ܦ���UK�3`ؑ:���ң��\ֈ�^�z� ^��q�m��md�x�-��%q���ekA����7k2s 8d`	L��K�]W��#�5Ǆ��K����A�l1�Xzy��t\��A`�܎%��<C>8�ۣ��.�P���������\�(��[aGkZ�p�<(>��������3&�s��Ί�k���Jrk���Z��ݴ�GF�Ѱ���um��e��@��XvL��ݏ �ɕ��Q�%�N�b.�`�2��)#�g�����>]����Ky�+��&�� �wc�;�e`.�xvL�l�Kwn�M�Cn��z��������xd�X�9�]{<�Ȭi��i[-]�M]���ǀvI��|����e`
�����"H,�-c�-�*��cK�9�6�:bV0Dp4���%mm��[�g86!M�������V��Ձ����7]�v:T�Y���7$���]��@�  B4�hP8&��lܓ׽� �+ �e�L��J�[m��7d��>�ذ�2��v< �d-�:�Vګ㻺�>�ذ�2��v<�O{��	ȼĒ�r��lEݬ�L���u���	=� �H]�6M6��y尉r)�$qx��_+��)
m>;���\��.�.����w�>�v<vL� �+ �'2��Іˢۻx�X�{�&V��ǀ}�V$�ն�]�M]��_}w$�����Z�#a
aT�y�P!JԂ���v��`��#�$tW1�iN:���	�:Cq@�d$��.��!�K~ ���7ݢj�>S�VX��"�VT�$�ȒI�'v�O��@o�s�z$XF���Ӵ�	GSoF�5�FaPx��X�S�@�� ��IB�!D�HmYC�D�$��ZCH�m<R����]����!�Ƿ�u	��%�K;$����<�> ���q;�f�1/�,�to@��`A�0�M�AI���1�r�, !!��VE���|b��nHM���m��	$H@!�V��aX}������ϒ����'�����l���BQ�CsH']�@�P�V/U���E����"p��D>�Uy � �Vt �6&Ê�TM�E~:��z����=���rI�Ș��n��vP���z�������x�X�r��׳� ��<��bC�n�M�`.�x�X˲<�w��|����x��� 5�3j������n�>���D��zpC	[�̌5lP�V������|�#�;$��*����5l���x�$��v&���ـ|�#�;$��:����G�Z(���˧m�Vݼ�L����dx˲<WZ���I���5wXWwٹ'=�znI������5B��C�!�� 4*�������}��ȻB�fWe��z��dx��0��x�U^��{�2ғ�r�oH1��]��<#���t�\�sn���+bysXy[��ή2+Sd����w �ۆ�ݏ�U���� ;��c�Wv���;��n��=��URF��x}��|�#�UUr��7Y^+�ۦ���T���5l��>��|�#�7v�|���ʹ�[��vw �޽8������ }$Vĝ]ĝJӳ ��E�n�� ��ǀ}%ɹ'��hD$J�"D �{}�r�TB1@�Y�U�)wg��P�\�f.����NM��`n�rX�
���7AF<dq�W-�^�\v!u{ɂ͚���%:
ո^�b�i��1�-��Q�ұ�#A�q�ݎK�k,nA�3(��8����Z*K�==,���^�]yâ��p�sI�Wn6v��9B���r��V,\��eLuɘu��I�ZF�k�PAĖ	 CUB���t�9�y��e.)Hp��:��0��M�۞:�y������o]�[]�v��7�{�_�}�G�}%���;��X��K�~M_.��N����������${}�*YV��C�t����w޿�r,=�W*��_�V�< �uSq�v�c��b�0��X��0��x�\0�c�Wv������7v�uwc�>��w�E�|�+SJP�X}��݂_�:N��NI������n�y�m��FT�U4�1��eO�~���p��`�`�p�>݉�wI]��]Me��nI�{^������"iLP������ܓ��7$���f�;�n��t۱�ӳ �\� �ۆ���� �)D!(av�1[��n�� �� �K�޹��%8�j�[��ӳ �� �K�޹���s��PC:�=؅�2,�pbѓ��;��7"���M�:��DvM�啍t��2�.��}}8z�X��0�����M��ZM�˱���;�"�7v�uvG�}%� �l+�v��e���n��	>�{ٸ"�>@�Z
l�\��Uq�k����=�"�;�Uj�65C��ݘ��x�\0�ذݸ`n��wB�M1YbWw�}%� �+��Is��$�� >�^�ډ\9M��	 �E#��K[�I��ny�J�Z ]�h�	���n���hm��b�7v�I/ �K� HRԕ(���ݬwn�����`�b�;�R�!�m	�f }$��.�ذݸ`�8�e��$:wI&����`�b�7v�ܟ�I�jB��k�b8FUD�	�n���$�z*mK�m6;.�+� �{�I3����x�\0Ur���xM0�`�Ctܐqq�Sn��p�zf1����#�Q� c����c5�dV��ڭ�{�ӀuvG�}%����7_���UO;M�Pƨ�wf�����r,~zs���y%���ێ-aV늎�; �~0�Ȱ�9�q)%��5o�����4�Ю��M����U-���$�Wdx�\0kR������i[��n�� ��ǀ}%� ��޻�w���E`tݾ35�5�.��wb��O{F�/fa�!6i�e�ˊ��S@�����]E	kJsq6����!� �e�c�sk�	Vz'�$�юi툜Ju�[ur5g��m�)8�w��ݷH3v�vu����ez ���f�g+A	.K�n�U-(�d-R�4r&="`��������i�uƯ�4ph�ѶJ�<�;}�hͱ�,�nwkyP��_	�lCg$s)�H��m���y�J��y��XC)�*t���.��۪�[\I�Zvؚv|�w� �K��\� �ۆ;',���I:�wo �K��\� �ۆ�ݏ >�Tڗj�lv]�Wf�\� �ۆ��u�,����>���X5eݫV�M]�wn�{�� �YZF]�*�Ҧ�� �K��^ŀn�� �i�Q"S�H\��zzܷC�qF�An��s1dJ=u�=�8�=���m���Zmj7l��zp�w����r�� ��u{�i�M]
�/2j�SrN}���p�4�1!
@kP��U�\�9`�n��X�\0V�D�����4���7v�}ױ`Ip�>�ذƸ���|�ӳ ��b�>��}ױ`�p�'v�e�e$�����X�\0��,wn�{7EV�|�H����\r�v��#�{Ʋl|i1X4H����+�vTڻ�m'N˱���>�ذݸ`u�X�\0��1�YwjժWk �ۆ�^ŀ}%� ��ǀw��#.ؕv�Swf�\� �K��F+	�@~S�o�^�nI�s޻���eں�M�e�ݬ�����ˆ�\� ;�-��wB�j�l�v`]���\0��X{._-��t�}����H��*d��ƴN@Fu�g���GVnxZX"Pt��f��C���2����_���ˆ�ݏ �k�J����n��{�H����5l��;�p�7�
T��e4�����X{.Wv<������{f�˝n�T�S����$��y����r,��+�k��I�%����bDȠo��� �"c����vP�v��\0�`�`�b�=U]ھJ(+�6��VC-Ʋ���1��q����xx��v�1�P/$��X8D��2@�-��?y`�`�b�+����$�x]��]���Vݬ���+���s� ����7�E��W�z�M�t+�[V��|��ˆ�r,�� �"�6��&����ˆ�r,�ncذ�q)U�Rv�-ـo\� �UUo��:��`w��
�����TW��@U��@U����
��� *��� *��Ң��"��H� �b(* ���T��X� �* ���"�0� �(�"("(
)@A_�
��E�@U� *��TW���+����
��� *��Ȁ�+�B���E~E�1AY&SYC�R c0_�PY��?�������`O>�(|]�_ o�  �l�DB!��@&����h}ۼ�
��������>���0������:w��v�����s�z�/�����������dϺ�������w���w�.������ݟ=l=� w糬@P��7����%�@,�y�u�H��B
i�Bh�Q���&�@�CF�"l�R�� `�0 ��UUQ�  L   d`Jz"P4��&� 2h  @��&��=H�4��b56��
�)����Dz!��4z�=C&�N	�z+�'V��
Y�{�T�(��QAN*{�ȤA.!����'����c"���P�t�i()�+��
�)"�7�7�����M~���~��{������������������������������������������������������������������������������N���������������������������������������������������������":@ t���$�yBT�"M�����������������������������ffff�������������������wwwwy��������������������UUU�������;��p�&�(w�=2�+��qG�#���j+!�&SP�f14�`�M���Ւ�8�(����N@˜e�[9q�$��LE��� ��
P�U0�]�&]�:�*2U藹M���v.M6m��!��]	 ���"kKa����U��K�0Ӣ�ع�z6���$ѱ6Ì�BS�`�$hcE��Je�<�Q�����i)�Cw��|9w`|ς�H[��}��zIL{�9��/`z!A
.V%���C�֓7v��Z�u��L�q+���bڧJ��=x^K�*s�D�ǡ��Q'rM���=Jx�YA�0����0��7��XU��)��'�Gǌ����������|�>N����e�k۹F�\1��x��4���K*9����^��� �9�0z)9���oG�]��rC���|��r���Z��"	)4�!�/��͹y��� S��K@E��$X�*1c��Qblf�ӆVª���٪���6;;-�s3-r<�f�5m�v�ީ�N[2��vs���"˶��'�0��=��n�j��Ʋ�Y��ZΐٓN�;J79�J�Ia�lve.��t`�se뛭Ilh�I��t�t�i��Y�Vm��k�J�)l��Zj��Iw3�@�O���/}��'�`0Q��9mr�$c�rz.r9b���k��                                 �                                                                            ��                             	q�7r��d��]��f6vlv�uƃK;t�:I�h�Ŋ��$[GFc"a���l���P�.��7jl[�s5�TV;lR��
�!�T�m!�p�o
yGa���f��T�)W8���U���s:�Z�R]�����t�a|�N;-�/6��fa�Gi1��fN݊�h�c�+���v٦I$מ�yw��|�vK
i��#��:��"�U���5۵٥�;�V�kQλOh���N؄�5܄��	v�Ԓd�iG�*�K�U˶�0J��ԫRdj��Nݎ��nN9���U��V����ڝ�M[m�L2I ��$Iv���.��B ����E�� �&�]TYZ�Jא�p�V��)P%jN�������I^̠4�j�[��Wj�-�՝n-�j��U�7kR�RŶ�&l� 2H ����L `�� ��f�UU��fX-���Um��UҮ���P��&�y�ivX-��iZ�i�T�4�l�]R��Z�U{Ե_�6�ڏ�C�ő	|:� >�<(ƷW���וQ^E;���EPxA�QO��tN�Ax^U�E�Ex�x^U���JJ)(��)!JR����UUU{�U^�UW�UU�U{�UQUUUUUUUUUUUQUUUUUUUUUUUUUUUUUQUQUUUUUUUUUUUUUUUUUUEEUETUQUEUTUQUEPUU^Q�UUUUU^�UmG�6�HF�� {��=�G�h�N!&�9Da�PS��0�,V� �͕(D�K�����M@�!�)d�nC1%tt��F���$�u:�ZQ�t!�dM��f�;��Ndm���J��G2��N��n�GrwϿ~�V�q[a�m�S��Qʪ�������������������������     vE�[m�[a�m�p~q�p� `�'���
/����m���Uf6ݶ��mn�8���'wwpY
�=�#�v�:��u�%��(�c�7�����      [h              ��    �e�w�,���u�N�m͑��r��ݤ.���\IJ:�m����O�.:KPcr�b�q��YZh��Z������f�u�l�]���C\S�ܯm�ۈ���<ũ�B���J7 n����M�#��̓}[�@[h  [j�g6�u/�r�[�wlɣ�ҝ�����T�ZZ_?l?=���=U�r���>�|�=�US��wzx���HK�-9�(�Ini0��.�j��r�+.�ˢ\���DVw[l8m\��J�f���)QZ9�V\�*#9�T��:y�U�|m�%�)9s1&U��|�.�f<�b�sG0eY�(00D\��.T��_;��ne��M6��/������0�]Z�X�us{|\[��DA��[m��m��`  j�̮6TdMcf�%�R�dkS�3��]	�L��iL����,Pt���SKF�[�E	��R��y���m�@	I��o:"�C�zT t 2r��Z��a- T�}�т�`MD��m�B�m���
j��ywIM�M9�@@T4CT����Z�b�s<�m�L�A�ZS/w�Y�x�I�����ZB�kf`�������3��>�5I�n�%���˫y��ʦXsz��榸8d0��h���ǯ`    G�F�S4ɪwWg�dצgp��ͻqr۞�O^��Til�n�c��k�nf�:j��m�fQ-M�-5[�kFUP��Zf�uJ����gj�mL�+�� ���m�-��r�*%"o7.��xĵyT�t���=�٦�����ϐ����ɞ�379�>�Z�"yt�$�x�+c�{=��ۗ�&�a�$���㡙���s��0�c*c>����ڱ�b #�#y"G�V�l2L�$�(^r0�.��{Y9��,��5�"^>�ځ�<�2��X�8h�!�����Z��$V!���ܐ,���ےSM)2��r��uML�oɌ0͘�=�w��W'L��p{����Iw1ט]�u��ݴKp���a"�D�"f�7s��7ϛ�    ���,��JC[@��ض�u�����>=��罶2ȪNJi!z� YH���Ӆ8x@�6@�^NV��G���_�H�`�|<��N�cg��Ͷ��)�ԫ�ށ޿UMpP�ȓ��ؚ�K��w�Ei�i��H����C�����6@������E-�-)���7�!��&8x@��ӆ�m&5`h��*����O���<0�l�)/�� ]HF E�D@��[nK��)������	�t�&�TI/��сD7�mT�(s�
GUT�wRH��F�$z��:H۬�]%�w���D���n���X~�":*�Ͷ���JX��m�b\+{|y�jhR��m�VgD��ౘ����3;��9���3��/�   �����4qv�����gt� ^��j�s�͐�/��I��o�U���<ߠDq�ު�p '|��ڵh���iH(&�Je�������GEō]�U�w�]V��� :�j�ko^��2�)�)-M�]O�^c��X�`8��S��O;т�N<��[m��M2 �Uo,W{]���ٚ��*�8��`L!�>}R��@n{��$%!��RZS/&��Rg4�o�1Q���uj�{�\���~�[m��m�磌1��m����m���A �0,��b�KaeEK���IV؞a�VF${!�QK�D���Aq%.X-�V�UKUC�}���EQ�yx�r��&z2�                            K��r\Y�)�R�v��Kt�Fms��9�d^��a��il����l�s�7n�URiq�&�j=LX�4�=��a&6�Ŷ��xxp2���c��\k�'\�X��C�KԪ�}�	1b���b�&�s��@⼁���b"�0�؈q��m��`  �Y����^��GGY0�d���n�@S_<Ͱ�D�l�����o���"-H�Z�R�'n� �oX0� W�|���3���-"Mp��,7���O�N:������G��[��V �ݶ�be�Дٖ�{��^?x���sX��b񿀒���#9������B�{�M�H,L�e�2�3s�@z �6&��������k�U| j ��1�"��&�k�w����kk��`�i�KA�&�(�؛��� �F
�>�Me���_d�7~m����  ��2I)�hڮW�x��q�n1Ŭ���3��e�9���"ś[�y,\=z�����W9"�~9��w::�M�*C!���J��g���yNM���jU�Z�UU�x��g�=�W�GU��.,\���M�ʔ�)�)�ҹ��SB� ���+� �3Dw^f�| ������^c]S]m�岥9M9i[2y��/�]| �k�o^��<����> �� KC-���[m�)ɓ-��X�Ļ��
����'��)�
�KT�{z�E��D�卶�m�   ,�ni�ܭN��]�e ��]k%�s)�ܹ%��K��9SO��w��������pv!Ƕ>;�؁����rKl�l��Ā�ԫ�(��� Dd���]E��v��oDW}�}�!`��m��3%�R-)�+Cr��ڑy�����~|z�� >{���ϐ����m��/���xB#ʪ!�=�Q�� �i�nDq/$��p� x`aiC�xߟ|c9�mU\�m�^W7��`�JT�)q;�=]F��9G�c�rĹ] H  ��v�� ��6�E!(J-�w����os*[��M��@����Iҟ�$�`G���    B�g�ӎ��T�N"=;j�u�L�n>��8�_<�b0k�{�|}���=3bkCM�p^\i���3� e'w� ��>m6ܔٖ�m�[WU�y��ּ���u���bD�My�A�_Yrj" �s�9�"Z�q F�i+ C�/�m�&R-&�"m�̸��#�����t��9�@�=Q F�y��n��y)��r�Gj��a')��2��U�֜�����RY/��
� 8'<� ~�ճ���m�\���.s-�gf�S�ќ�x&�_T���r�^x@���>t    �E@W\��H;[�itNs�3`��Ź<_���x�r�w��\;w^l�H���ۉIKF[)�|�.�{�U��. M���xe�X%���m�Wy.{N�lK	)L&e�T��y�Y���n��+�׳�W�(*s�R�fC��o�*��e4�8�:̰�����������ts��ne�f���)�NSs6�Ū���.).�����f�4*ep{qz�l�߽�|� |�{ހ�3�o376"Bq8eXE�`�YV�j��'r�d���`Y�xU�NxVnr�2�n�nf�O��@                          U�È{ez�7@�c���s�Q�%Hn��^��mOP��vJh��a�.-n��gY�N�v�Bi]aV���vdۗd�hC�v�.\,[��w&��ƺ�맵v����t-�,�h�\����}�>����sq��4�T0)0hQM��̌���)��}s�/@3�''� �*p�7�~s�����     p@Le��VT;S�n��6M�m,l�\�Yuj�?�ۗ��7�S�pe��v�������BЊ}<�-���[l̴&Rbzt�+�3x ��aq��8@A������මK>��9x�",1d�#C>��]��d�
R�++88�dH��n�seOg>��/���r{-Wݗ=Ϡx8���M����ۙb��� �{C�9X񎎌
�Ǽ��91�� 9��Tʛ������R��J�`��`k�WT�ޭ�k�mP��v�L�Z3*ǡ�,D	 F�"oɶ�m�   9[�ڗvl����R��@�z喛m��12��6�Y���W��Ѽ[��q��ʓN��Q8�����Aq޳Uuw"�	 �%�TN=|�ǧ��/�"p�}z�[m/K�[&/��/�8S�$8j-����E�5�"�[]��j��o��OiiΙ���9���Q��U�V1Ij7��H��+����z�#����bZ%A��Y/ڨI�I1*	 ��A$LD�$�cfս]Ilsc
�Q�0�Qls�#5�S�8S��>m���]��Y8�8ިMU	 �&bTLD�$�H$����H�{�9�-E�͌W�IF*-E��:���Q�a��ߛ�:��Z�Qlf�,j�(���e��q�Z�c���ּ��h��*%A$�BH$�������[���b7Qj8�j*��b��Z�Qlj�*-q�>7�m��+s��S��
p�{��p�Qj-E���*-F�X$���,��H$b�A$MD�+Q�0�dZ������4�-E���*-G8�-E�͌TZ���Ɲ���5Qlb��-E�ŌTZ����������Q�wߘֶ�Qlu�#6E��a�Z�x��N*p��8S��z���kf��qf��q�p��)��"�Q�0�QlgX��Z����H��1Qj5�j-�,b��!�P�M��\�m��LCn5�M��S���j��ogh�>��     [���cqYS�uͷ+���RD�!3�̹��@���,ML2���.��ӤE�y1͟ �H�Eޤ�Dtً�ݺ��da�h�6+�!�!n=m�m�&[	!Lٲ7Suט�f�va��������4���0�#��,�1f��bȄG�#g���s!$�F[.B2���"��]���E��1ש.�0��� ��u�?~������z��<ffsVP�C`�����s=��N�#(j�`�IJ}s�������Uu�m��L	�Mӻ d��̠B@��U�$/���y%�ǨS�.�/��x���vH6sa��k����e�حٛ�Y��t��y�9�t�`���������YI�I�^H��a�?��d��`�B1���m��-&2�0���(�Z4!�a� <1�:`U�B��R�$�:���ũB���m�Т#24����2�- �_�f0� s��aF�(�$�u�F$���c��,��G{�����fs7~_�   UUU�gu�e�mXY�F���n8��U�5U���ۛb�'|�2��Mrhf$��F(�\\	� 2 ȃ�q��ek��k�0��T+�>|&���h}ra��"�Q3�Y�@��C,����PG���\�%)aZ�"0�1��"L2#���(�~Q LF��,�%Lr�H`(�G�@9\�m�
h�l4�L38l��Jb�M�q�� I��ѩ�(��ˋ���SD�<�u��2L��r]���8D��
��N���]y�\T��+=��ݛ�k>{�;����g���~s���     �v�K���t��u����2LM�-K!�6�A��f1f���
��{_��<z=�O�t0�Dg�\�f(�"6YR2 ���m�%	��(dY*Fn���Dwh![1d �ԇ�4G�"�?�H�}0�KW[l�JH��Je��bȅ��������jǶ����!�f!Q�	���+���8q�`��0Gyۦ�����*Mɋ wR�C"=>� �cV�3f� H1c"B*E�H�b1 �@��:x�OT	��~��e���j�h�ӄQ�=������ds�B,�<�̷Mы�Y��xuS[���R��7����� ��{�>@�����
�b�-G�0Sr7��5E��l�F)"���	
�#UD��z���H�Ӟ�p����w��x;�                           ,��w^�<c�y�/`0�k�5.�S=�ˮ��vN,�F��K��XI�=�4�a-MY5���X똺q�Ŷ��=�.l&14˗u��l���:���F�:�ݲg[S[��X��8�M!2�!�:�<�fs���<�s|���  UUUm%���.��s1Ƙ�M���шj�,��-�.' bLqj&��.DO�fdF���b�LV����0��gi��m�l�J��='Ǹ_Z��㏀8�䈲(梢�� 1uj+���I�0�����B�G�a�w^m�Crٖ�	XY0�@�M� F/_6E`����j���|nXsA֦�1
9��n���m�4��6M�m�H|'�fC�����ݦ�(�8Dm��a��@��(���ܩd&%Ke̩�Is��u���N�KX�@F�P�FF��|�
�`v��
�O�@    4u��b��UɲH��;XĒ���s3)@ݪ%\D���0��^}���L" z��� '1�h�و����"�Q����s2Bl-�2�hY�@s�ܘ��� �:�{���EF7yLA1DI����h�E��ۆe�2�X1�D��:{A�؈ Y,�ِȊ �=��Bޡ��Y r +����Lb������-�� )QV �p��!�'bh�Ōa�C{bl��� ��7���1$x�O+[m�2��Z�Lc�{�Q�1O5�1f!�ax�dE�F�r��B	�Q��p���`   Wi�dųrk��ь��\9ZKck.�j��g[&���C�C��g�����#�w&���"�Yq�b�tc@����q(�2���i�`t�0�x���jr^4"A�04�X�grb�x%��d �O9ζ�E$����b�bH�L��A1D#���c��j���m��|�z����m��U��Z�sĥ��I�b�J�ݳ��e��#�Y���;��,η�5�=����}N7Χ��̓.�.��T�v`p�k�p��x�i;�0��wȣ��u,�����8D]�|�cm��[�������'���~������aӞ��#Z���"9��gw������c��g��:     ��m�ԙ$��97YpX��*I.�d��X̗�6ۇ2�M(�Dx�w}a����SF�1ˑZ���0:h�sR�<84c��q��L̖X�l��FԌ> Ac��%�D#���=#*@�P0�LN_F-H͗M�"fS'ԛ$���#�]bψd ��(f�� 0�?V�4t�T�Et!�#}��$H��b��x�<���&���`�2`����l����4Fvt���p� �D���(��4���l$'%I���M4��o�>7wm=���Q]}7��j�z������Ͷ�l   w&�Ul�:y!�0���J��mX��&�m�.eJ�˓(w�����0g�O}Wv��z���:�ͮ��m��,�*S- �X�aw�n�x�w�D+T�A勹瞚�|\���(�A̦�R�W$�N�+]�DEW�k<Dr��^���_�T�8ۻ'׾m��I�˕&Xɵ�m���٭<�̩�{� @�%� �b#���v���ߛn\�R%0��9\H��JdU;��vȈ|�*ř5�P���W�� }���=z {�{ޅ�9�6[*���T���tXX�a,`��Q� 4�'�fEId	gG�D^@�"/(��",�ΐ�T��>m��m�                        ���7rE�2\7.��%U��m�qm�`�p;]�/a��cdpC�n���3�{}#��X0aɰ�D��R�ӷ1�����7.�⍤�r��5�TX��n^�2���&2M������s��s3�g�s���s1����    �r-��uےo{v^�.���-i���i�~�i]vQ��W�b�0�z�.��mp����n��)%�ZR�ɼ:U�?LQ?��x��������c���U����l��%0�2�n����CǑ 
ӵ'� Ȁbqs�9�/�/�i5�s��eJ)	�Hd�ϫ��r����V#�'���W;�n�.��~m�B	��mKK�k�����͊�]���|������|�������ߠ    	���ȍܗc57IWQ*�Sr[m[��WCsY�T�Sd�\��7m?+���|2�i��M�m���撶����J�m�dɔ̴A川�
��Z��7s�UT�qmg�o�{u��fZM e������h��,�_X��' @��~Uuڿ�r�n8�[m��̂ӓ2���7n�q�Z�w�2����w�
��
�s_[l��f[)�������N�e=���oGvy��>����1��   UT�D^KW=�ny�w^Acr�h	�dj�p�"e��L�é�W�ɛs���l��d�P����z�rK$ӗ2��q5�}>q�g/� �}�s���&�Zy�r�%��ٜI[W)��/�����Gg��m���ߝ�^� }g=󛹜͋!�H���Ӎ������� �*F�8�] G6"4�t���=>]�|ϠZ��K�\���m�SfRm�y�"Z��ۤ��Ug@1�-X�o� 3�^���;\m����r�X��8��b���=�}cq1���]�;���϶:`b _x�m��   v^$�� �:�e�d����B6���z�b[+#/�ry���|e������Vi���KV��ܹ�ʙE����_5��g>A�q��>�n���W9�W-V�y޶ؙ	0Ҕ���;"hUS�cu�^�������]�;�+��mA�Rl���/w+�w�y��޽SvQ�z�_�yP�K��{�m�e(4C2�7�`~���s��̷=��7�d����9���D �����    ��uTY�v���/{�c��.\�bV�l˒�����m��JSD�E�����ߎ�r�Û��!����f��%�v��N�6�l�EJl�6���uM���Ϸ>��W�" �}Z�w��"����e�k�}m����m̴�.d���2�s)W7}{���yU�}�M�o/[lL�NL�XKy��nU*\�9S\�զ�Ϩ<>��ʛ�km��f�����τW�ᙗ*{�J�g(W��˵o���>�W����d#'L�FHB
�)T�b��~�~��'���U@�0�|���J��P`ز�U�Z(b킅
$B �UZ���H���'UT������dT���R�#[�M��%�C�F�tI�����V-I2aHD�dDV��e4�h�Q$Q�+q�yal[���xr"���PI���n?���vD}^��Jubؒ5�� ��	a~�D������q	�?X��?	������ i?�����}&�i�ߕ��L>n���x� AOh�t�8|�O�5T?���
�)䔌�Ϗ�C֝'����v%'�\X��˰�>�8����I# �P�⇟U�K	!�+*Rh�>�m��I#����T}Y>��ƍ7� E�9z L��I"�l��I�%�*��	AH�"�PO "�*A*XHCUt$�-ZUZ�YVU��KdK,B�E,��"X�s�$�	�x��t�����i��k�W�~���$�C��9��I�ſy�����>��D����rvrz2}>�O�P🯠<�*�)�����������~��>���B�+��}}����w�ì�a�q��Y�ߴUN� ��:���N����<��w7���#��`�;N�T>���4a׃�ĕK�X��7M� �2?D{1 ��>�-�tʫ�?��V		J��|0�Z1��%�Cz*�������;���%�CFEP�i�e^p�@S����W8s���O�}��v>'���GAEC����za�1̤���~�
�)�� �=��*��Ap^�����vsp_���O��c��J̊}�n*����ʵ޷�}���;�ܞ��m�0k�B�
_�qK��574
�]�;��5�t�������)�������=B*�)�`y��-��H-��o�T:�Aq��qC��!��ơp�!�_=��! �$����H�
�\K 