BZh91AY&SY����_�pp��b� ����a` �P        @  �      �}��  �  D�IR�P PH(( *��DB�)"�)B�(

%T   	E   "��  @��B@(�
(d i��qhVl�f����ZS���zZQ�}��y4����O�y}�ťv�7� N}�_An��@���^��8C�q �`(u�=�
����q �H  <@(P(AT�i�P��9��}��rӖR�eO}� �|�W����ݵ����seK�(�R���w> m^l�bҜ�� w���髛/�>�u+R� ������MNM/�v��som�� �� ���*���`�z��}m�7N�ɮڽ��Mo<����J�n6��T˗V��ﾔ��y���������y��+�x �����d���ε����]�Nz���J�v��^�iWq�J� �x)TJ��P
ŀ�O�9o��}�^��R��R����U���������OW��]�� :��'�3�3���m;mw�ޚ�=�$��Ҭ��}��]n,��x��i�� <��nm\���ֽ�����t�x �}E

$ 
(�� �զ�n�nm>޻�˴��]��P�;�*ru���{�ye;{��=S�x i���q���ם��  �^M*��{�j���^���Z�&���[����u��甠7�m���)�{�����wr�Ɣ    J=H�m�R�?T� �C�i�FFO�l�T� @�� Ǫ�PȦ�     تR��j�  F@ S�
)�*��4�   ������hCF�)�� i�6����O��������y�?���|:���� ��������UW`**�dQUW�PEU\H� ����|�DUU��I�"����t*����������I�YG�5���9�[��|�	NLY	F�)�l�7����.byN~!(<r�r��s_�=
/�4o/���%&%�7k� �����ǱN	Ic�,p�<�h0��j͘�t���7��g#��i�Qfb~4ţs�0O����G\Y�I^������#��Q�?����|r<�7xp��x?�Uyf�_z36>߲��L�|�it�i���MI�d���N��,wύV��iލV�F����ȃ4���o^����[���y��py�ằ���NӖ���>S�����l�����X4�����:9����f�g<7���3�W�;{�"J��^LED\Q�ܵ>�ۓ�j�>�^p���$$���8}��6T�	By`&�pٮf�#z����,��;�h�R!(�l�%���X��/5̝f0�K4n���S��p܆R��X:��c��� ����FXbE�����7��>k=C1������7hoMh?Vp̃[�5�k3E��k4c�̸K\�Q�NG���O��t~�m7�h����k3�Y�a�+���u���f����NRjl�G'5��q�'��q}����5�&�p�J0��K�k5����|���y�Y�y����k�`?/��	@~2B2�͜��尝f�8c�F���p�F��~۷���'���h��(�#�q���(J����.BP��c�?n���<ggN�ѷ����Cp��泈V�Թ	���%8�����Q��%����Fd�Ѽ�x�	F�q&��9��9K��#�Ƶ&o���E�Ra>kD�Q�<��̖Ȩ��ћ8�X�D��fÛ���tn�5	O�BP�&�|*C�b�7�f���o\#t%/!���zƍV��퇅^��<�e��I�`���P�d'��eS���,�m���	_��5x�F��	�bi7q��%���}�s������6Ѱ�<�1ѩĊ���D8TJ	�	�t�dG�`�d%	By	��%	BR��2!2�&Bd&�)y���|ϯ��O�����������X�`�Z�?X^�{����ub�a͉BP�	T	�)��nBP���%	��$�(MBP�����/�i�o4�RPy.QTN�� �a�𩭚)9&&�/$0�
��6H����pʚ5��ߢϵ�������Fy�NK#�	�x�P�`�~3�����ЙhjR�qͿ.I�oX�}~wY�<��� ��`�J����F��޲)��]BP�bE��Dd�&���<y����ddm#Y~#�j\����yA�㪃$�dՖ&�_sF�L�Σ2�#��gTS�����r��f�$� ¦8y��a�C��?�dC�ꊲ�l�>iʎ���r��0�p�}�`�\q��4d��kn��F�֟jq�<�Q~=��,�h�����-��4`9^��rU��Px��2O��6aE���l��l�I��&;5	A�~�8	��K�MM	Pp,��AY8�&De�S�:7�y壛ɏ��oD!� �$�>ާӨN@h�x&�<��F2�>�C�dZ�K�`G�`�%	K�'��� ƌ��?��*����5�^��$}^�98q<�\�f���e���y�mߙa��9g�w`[5���&Z��8ލ.�I��D��z_5o4��}uI���y	BPe��#/�~�
��I�d%���}��2N'��(tm8��ZM�m�m�璮U��L"T$�>��Y��w*~�q������p�א�O0O$�d��A�_�a��<�y�q�9��q9�4٭\��9��O��B�X�:�C-7��&g�dE�<H
��7s�����3ۚ�"4~m[v��f���o<���۹��.;u�~�m���8�F�P�l�翼�g���K��~5��#!+`Y8Ay�	Bn|$�L�%	@a�!����6�RI�4Bn��9j]:�\�� 7	�L��(J���e�9T�21��M�P�&�(J��(NBR��d�faj��\���Q��;5�ky$�L�4��M>p´�r㖒4}���A��<Ǒ�Ց�ӫZF�Q%�%5���"�,�Z��6n��<���kXBP����d%	BV����Ǒ���a!yi��z[��π5P�	�A&��'!�Zw�a��F���^؄�&X��4��\ѥ7fs,�������&�:�̍1�����zI�G�x%��kr1���h��(�1呭�� 绀�!5:\�q?&���5�I�a�V��OJl5�\0�F����W^��{�Cu����;�]����s|9�9h�s��Q���!��>�,�$��y�3[��M�33Z Յ�5ZY1�Z
%�����J��(J��J�7syfk�k�����o�̼&�+�d%	q|r\k��NF�!����#_�y��ח<Ks/8�$�sa����	F�����2���r<�d�c%�J��<��/�C��R�����J=�ѨJ���2C��f�2�bi�*�J4�WƵ[�	������dК��Hdm<ub!(k�(J��s��^f�ώ�+�f�׻|5�/��u}��r���CBd��%b	@G�4Q�g�}h�\/+���G���4d�'�f��3 �C2L�<�i�r�e�Y'�ͳ����&�*���4Χ20c'��Q���լʈb��%	C9BP9�&���jj?9f�����ә[�p�.T���m�3����*4kg�sF�0�jCyp��� ��24ѻ�xm�j��9���� �s�(1,��;�,	7c�Q��%	I��	��(J��(J��.	��(J������R�ַ���A��uB}�	��BRbd���&`a�(0ry�P�%	G �J����Mf	BS(lJ�J�id&f8ε0m�(89b	HfI����O3 �kIP�2�N_��������_S���4���1����)C�A���8��F�P�`q��J���l �8�N��hDF��J�!,�zh7	�0J��BP�%	@l�&�7�m7�!)t��i���%��|�0e��Z$��hա�� �2�̀ٚK��V��O�~�#NZ�'#�kA�.�@a�Y�2s�f����7�f��F����sbS�Hg��(JOp�f�W�NG�����*٘q)�Py���Pl~�+q�8��ݝ۟:��X�q�{���zw��ߎ���w�j�C��\2����#F�;�٬�߮O�oaQ<>5���L��-�f�+ԙj2̊0�s�Ն����zV�C��;l��BS��㐔}d%	Bs0;}}�?�ѭa��׃��A�Vf�5	x���o4��VI9~pס�2##5�v�>��I��[��y�5��sBVhl��u���a��g袱�Nh���˻�^�����}g��E��F��r���3������g����|�<���ww�0�o�<��������z���2��jC2����٠ٸ<�z�{���.X���� 3Fkf����<MF�F��\�O���Ų2\�(J_�BV&��	JP�%	ZC$=�J� ��?'`�~
%�����?{�q�]A��ȥ�����FT��A<"y��%�Ͻw9�J*y�W�R�TA�r�SW?w��B�Y��}�4�F;����r_ӎ�P�f0��=߷߿ڱ�V}�Ca�Z3W,��Z'5f�u�F�)���1toY��y���6��ͻ�ߛ��H���7�	�<vn���oq������?�в�Nj3�9�M�m�34ᠵ�9M5��{��l�&�f��&0�j���J��)J��(J��(J��(J��(J��)J��(J��(J��%	BP�%	��%	JP�%	BP�%!�BP����C!(J��(J��!�ްJ��(�ޟ�x%BV��\�J�DC����ӬѲ(�`Z�Q�6a����`�i����Č�6N�����[9��7���`��A��qr�ٙj+�p��8Pn�$�9	BP�g��J����?>���[�������/��Ͼ�������p�   ��           �      ��|   �
Pa��޼�`           [i@A���` ;���  �   	�      �            A�        >�             
�            d        	(   5�9���o�v�)Rm��d.Sm7   �)� ���C�U
%꫶��`l 6���m��wM�˻\Hm��       �|��T ����ox �[j���Pe2U6��  oi��` � [@ sm��� 8���-�n  �!m �i�h  	 ������e�B4� o͟   � w  �� 8��tٺ
ͯ6�݉���]/-`$I�p擄��JKn�J�U]@B�8H	nLm��ۭ{-��Q�i0-�#mͰm���e�u-�   V�/����O+&��� �x%��*��F�1�gk�Y�m��� ?@� �&� �Tv;J��Ð���Pm��v1����6��
����UW��b]��
�j�l$y��� :[4�� �)�J��Nļ�J�UPm� ��Z�8lҀ�m��9%�5�J�̵���Ő�$:8��[�f��
� ��I��� 6�Zд�m&�I���u�  [RI/n�]s�m&��   �  -�m��}N$���u��uV� �v�jݛkjH�   p�i:m���p [@� ����$m�p6��H�d�ݰ�]6�$ l��-��  �m�d��ސ��  m�ݰl��@[U-�*�;8n�'RH     �i���`  �%%�8Y-[e�Ƶ�Hְ#�����\ 6�6Im��ض�m&ć�j�D�b��K���ت��g��N;���Ⱥ�=��8��6����m$�Z �kl��e�^������� �`6�փ� �ݻ$-�,0-� *��B@�`*]�������I���!�m[m��` $$  � 8 �ٶ� �kn����M�`��86�[@  mUu-mP����:  6�[x[v�۶�6� l �l [@hi� m���ZM��}�kzɾK�� -� �Pn�L 	j���c���[B@���۶�$�m�H 5�L��ŵ     ��  �nP�A��d�;�  ,55�p
4�-���M����   -� p�`        � ���f^��l��Tb�L�+�UT���f���� �l�!��-����R���5p
� m�  lpWR��S<U/(Q*�P��I���@	'����t�� -�?@� 6�� [Ԑ[f�  ��     ���Y.�v�mmL��` ְv��m� �@m����U�P
�+[R�j`k� -��}�o�          �Hq���     p�m�m�� �	 ���v [#Ywitr�m�m ��m�'�I��0 H�]	��C� g$       �    ��-��%�	:I"���9���KR�Q�� 4-�� � �m�� v�-�Xa�8 kn qUR�f��L� 4�M`U�d)��Ur�PR�V�JK+q���h���2[��m���[��N��� ܝ�M����6��)�az���2�!���O�Z��Y]m�),���(,�lѬ�UR�-W@����ďAq� U-��
��B�r2@J�U�U� �ܪ�Hm0WV+bvU`Mҭͭ�n�l�ڤ�2�Ԍr�UUVҎ�`ڂ����-��T�l-�ٶ  �̀��/T���M(��R��[J�
�R�V�V�T��� B���G�}� [�+m�d�kh���p  n�ۀݴ�m����m���*
@�)2B�A&GZ�l���� �` ��vm]B���eU�%��U�l6ۃj�f  ��@  6�@   	      mjm���Zj�Yq���#R��ջI���@		�m�U��L�8�[B��Ij�cIKu��]�&�m��Xh���(�i%��[@Ãl�	 � 6�a���!�kn�[�8��.�Kchm�= Λi�*ඊQǲfJ�H [C�mf�Kd��C��[�M���6�S	e�f� �޴޶t�� $�I  )@ 		6�`  lh��H8� 6�n��5�wK���� �� ��k�k:ʹ���-6m�2�T �khW���>�} ݳ����[t�V���
�bO��}��f���m(�m���5�    �JP IH�e����RK�� �k5��ٛa 
R�5�/;X¬�YZ�]�)Um [@��$a"魸-��0ăF�(
�UU�*�Y��〓�m��ͺM��f�u(	�N��mnl    �            �M��� �ڶ	�$��HI�$9��IW����uT�uʮ�tٶ�	    ��pڥ\Xpf��ammn����Y��l �p�A��m[:mpp�i��/�J�UUuԬ�*�
��U    �-�Em� 6�%�1Ĝ]e�e՛   mY�g+b.�\-��rꀠ�j�P�U�Vm�`6<��Jl
�j�YS�d��#U�E��{e�J�AV�ȴ6��H��# -�5��  UP@�geԄv�MT�m5�mm���   ��{D�m'  m�   ��d(����2�n�Mځ�M�mj��m$z�s�a  6�fa���Y>��O��[�	� R�A2���sO.�j�j�� $ �d���n�*U���h����R��  �@M�q�m�Il�6� m�m�-�k ��ru�f.���( ��  ���6�6��ׯ����}�6��$-���}��MAm5�    � ���5ض���j�4k����\�N$�d8m�m��l�     Am qm$m��m[��nc��v� ImwLmz.l�Ƒ��t�� 6�  ��"���[A���m��f@�H����      ���f�l��`E-�^�n�����e�f�9�h�@@ �����8  ��7ɲ@f� 
V�)] ,I��I�@]3m.� ���������� 6� Ē ��^�	  �[@�I�     �    �cl�$�aM�[UKĻ=�9�aP��ծ�f�n�I��H�   $ sm��hl ��E�n��@  �e�]U���+��@��jU�N )"������u��܊Wh�[�"۶m��)��f�    ��l  @�`8����    Z�n�գv�%�Jʼ�.�*�*p4�m�Sm��M�m�`m��-����� m�8�@  ��   m�   ��        �`m���2�r���B���Ď����m��"��n�� -�   � [D��t-Yq-C�#.s5J��l�_}���睾���^�� �m��� �H�i��j��`6���K(����ݛ6E����   "A8   
������� �l�� 	$ m��v���`   Im��l�[h[BCmm� ݤ��8m�Km�H   ��J �` $l�i8 [Cm�U   �\�`@   h   H 8 m��HH  խ��B@  "iC�k��}�$>�m �  Ӏ������HI-��[@�f����J����:Ŋ��S[�  ����_��^��l  8��ky��� '�uʹ�S��t��n[Lr{v+f�3Ks��UT�m����UIjCR��l�Em$ˣm� ��D��4J2-UAg��2�	�P	$ r�-���Y"���9m�V	 )R ����� ��su�#m�?���r����DU]��������O��������M���
��8��e� ��hiЂ��	����D B?����& �=== ���@�`� �@��>(���TЉ��<@Q��Aq8 /��`���dO�"�T���?&#$�
���6�= ���8	��$��4+ID(� ��A2D-4��(@��-JI�K"��$ �H��C$--"��
z��+� �=�@G��$#C�(�%��]�k�Bك����Q B��'W�C�"f�B!?�����ªz�@l`��+�q�t 	�kH~D���~�0U*�� 8B�(���x�t���~���*
���_���-������G�~�0�(,���B�������ww{����?�}���l   �`J �mq�      m�    8 �mu[iv�e���i*�mSd�� ���ŝÖ
@"]r��NԜU���	V5��л�۩��a�m��83hk69�.��rzYY6���`��l�إ ���@���f�f�t+B��v״V�9��.^���잕3��e�u�Z�R�0���fZ�$f�n� 8�D�ѷT�$���F۲Gk���j	ڣ��uI@J�\�86�0IsK�$�֤��2��ې�,�)�˩�lR�9�M�d�6$�j� ;*�m�YTp�����(gJ*�T�9N[��eI�cvA���[t� �q��a��AU@UYv��{m�#�eՙ�*&�B�@mm�e��u�i�f�����M�s ��[uۢ%�.*�r�Be�ڛ��\G����ks�禬'b�veBn�(:k�3�3����4I�J�v����"ύ��  
�*��q��@\I̻�20Q,��Ynꮛm�u�ܕ��[���i+#e6�f�h4�V�q�m<��.K�����e�q�+(x!����8�l��ʻ]�f\׭�u�`m� �e�eJ5R��P�ۜ&�;j�
��Qp��5��^x�-��P݅te��ZVw�Z����!M0UG���`°qR��۲mp��2R�$�v!���`ƉY�HA6+�s�E��ٷe�4�X5m t#%�[m�1��6�͊���9"a�vV��P��N��LĶ�U���1J�U*�X�Ny�8]��ȵѰU<�@���<���t�KR���T��qaN��1�v�\Imm��cm�B�@(J�p�K<�i`����@@��*�+[J�76�K��=T��R�D��t��m�&��vٶ 	V 
�8�تV{m���K;b��J��u��N�h��F���ꕭJ���x��7e>���wq����h ?�DO����hUO��!�>S�3_y�oVn����t�US���w�6��w�W��%��r��)L:ۮx�V�����Q�h��S�R�n(N�A�̀*e��n��v�d�Bs:937NB�tv��6�m�
e���e�81���v����WN����3���q�r�qv����Mvv��ݮ���b�9y�D'1�C�y�\뭶���雵�÷=��w�������O9˞ݶ�<vW���s�8�]�M˶{>X����X�1 \NO�~��[8�zE���� ��# �@�D���IR$�w���J�(�I!DB����1��p}�8��X�{�f'�ě��+F˖F .J��d`=�.蚰���j��呀��.Y��}�h�B�FE�U]Y3aUq���.Y�0�d`����?�.-c�m=��DG/]l�ǰ���j�v�q�m���<�k(ss٭.�7[M\��˖F �Z0\�0rW�{�1�>�p��6���7�4�;���Dm��DY�# <�^�K# )�Q(�&ੲ�h*��<�d`� �%��.V���*������*������^�K# \��,�}!��A0NN�n�8�}�o���{�d`� �䪰����l*�g��v���!��:2i����Wg>d�n����D��6���n9�'��3�o�i�=ܲ0rW�o%��t��]�M�U?MU���F .J�Id`���>�3s�ɚ���(`�� o��|�Ͼ��-�D�C�P�Da\��p�>��J���# <�
V]QwSW����]����+F��# �x��a��7�cx����� ���0.W�jK# D��TMTK�$��[3eH��OM��k�\�f#l�ۍ�3ƭ���e����vN]�!c�f������^�,�.�`	U\�"����Crg 7}��wwy�w�N�{y����&�jE4`��0Id`	u�����呀	r��ƍ'���ͤ�4���� ����U}��o���>�AT�<�]߳�j����� �"�7�{y� K������F ��#�\���|���� \�g3�����)��Ot3�ݸSt�����Z����}�u�9z�`�e��ӼRY]hqD}�	'����;�X�����8ww��7}�wr���^ܮ&�%_�]E�UEUq�%֌��F %��Id`輱�����cng �>�{���\� ԖF �,� J�.���"䠢��0�d`ͽ���0�߸r�1A������� � ���&���v �[V�ƈ�E��SA�����l�Ij�K��v�RQ��uОf����r쐓�	�ck����.�H-k�y��u�u�i�P�\�y�ke�&n�������7i��n.��52�8��Bj笞0k"nZ��x�Vq�f�nJݹ�F���Y��v����]3[���=z�]#	�����ټ�N�����⁕�q\g��-Ri��mm�w\A��Ӝ5���IW(C]�s<��)��^��vwR�7gf��c��F �,�w,����d`�R5�$��6�x6�p�o3�o�����F ��F ��&�]�7p�\���`�d`	r�����呀tw�E¢�,��f�*�0�d`�d`	r��>]�# <�WsuD\�dU5W�Y\�0ܲ0�d`�?�o�?S��~��Q�]9��m�H�8k&4�Ct�=�����Þ���b�M^���TI5Wi�`�h�呀jK#����L�48,L��=�M8�.�k20$�0�d`	UY6\��EUf �,�RY\�8�� ��4ɭ�D�L0x��5%��%�# ��F �,���B�������L�\`	r���,f��y��0z��Q*����쀰�\C�f�Z�D���vɶ<r<;m���u���Ȝ���#ȱ93�{ޚp�o3�/%��%�#��l�����U]Y3d�J�t�R���G��P�@g��8�}�l�7IɆ(���7��3�}��p�(x���S�D�5��p�o3�{�17�gЏF�$����F ��F �,�RY ��D]MIVLMU��֌.Y���w���{�[�j
6�#PQ��*�\E��kg4�ό6�tv��n��s+ml�E ��1����p��3�n�y��~��;�2kƤP��K�5%��%�# �S�	r�s'*`1���!��$��n�g ���pw�8ww��=��OrF' #ȱ>�P8P�3�����2�TB�#>>�>�6%��p��Q3X�B8%$���^ ��F �,�ur���_�����˧�cw87$��N
J�-�&�֞s'i�鴥�ӅmZLt��������呀.�S�	r��ى�[>�x�&$���7}��\ϱH�'8 �w�/%����
)u5%Y1TU\`���\� ^K# K�����䄂jd`Ɯ\ ���RY\�0��8�E�����&�

��RY\�0��8����U��"������v���k5@ �U��V�s��}���U�=-��+�m�mrEr۷l=�����xY�H0q5�8�d"�P��솈�� �֣;׶&vH��i�,�Gd^��D�h��[�S)��&K-4����B�M�E�3�v��k�i+�N�'�V�X/[.��$�{�$��˞�b��Vi�.Ò�&�L�Zf{g�=5�F�=�]�k�v�c�ة�.�{�m�`zM�ֻ��0�i\XDnےu��\��q:��O@��Vm�n'�	�M������py�.Y�Y.�&�]�5a�M�� ��N �,�y,�.Y��y5��#�P�H�﷙�7�e*6"P�[�J�y�s@g�����詻�j�0�0�d`�����g ��bX�ϙ<��&�p�Y����9�O# ^K# ��6��\�I����vic����Ό�λrǭ���F�Ts�G^���X9rр.�S�%�# ^K# K�F��E ����4����g?|����-���d`����*&��ț**�� ^K# K�F ��N���p�z���$�m���܌ur�.Y�Y�˪��tM�g�zO{Գ�{)8���I?�:Y�ά�e��݂�(��HC�Pn2Y��ݛ���9$Y��۟=m���Dv��GoFzr۪���.�a��!j吗+�]�Y��A
�njn�������Z�d%��{�B\�3߷q'���#yM�f�fo�{y�g��?��$�U~�hO?b8$`A�������)�����B�	&ͣ���b(�(h�%���	.(X�``f`*Tc9ed�.d�fZ�#R����CM�T�@C�㔙�`�&I�����8`f0B�S�J!�j�a���D{h��)b�)Y�	�R/=K;��4c悆���a+9� �4IP��2\�Y�AA����� � mF
LSP$�
)j㉙��J�,���������Ȩ~D�T����DD?9��<�a>@C��=���AZR������җ_s�����l�o0֭kg�T({��w��)���AiJN����� %)���R��h[d$R	1��ffb�s��O��S���8(Ҕ��߻��Q)N���┥~���G�JS��>�?���e� ��wm��Vd�4�M��\�"��[�鹈��;uܵ����]��dꓷf��%)I������JG���8�)C߽��%)N���┥'��Q�ݭ�fm��kZ��JS���8�P����w��8>JR����8�)N_�o3�}��٪�bw$i<�1��8�)C߽��%)N���┥)��ҋ"D&�Ҩ�!b��1��on�[7r�s�%)N���┥'w��|��;߻ÊP�:�� �����" �J2������C���������;���Y�o7�V�k|R��y��QdB�	�>��x�(��gc�����1�H� fFے@x� Ή̽����x�H�I�ۉӵp��8��x9.��ztff��e)N���┥~���|��;߻�)JR{�{�������k.�Y��խl┥����|��{߻�)JR{�{����{�xq��3�hn��jA&4qG9�����{�y�)JO{�{��R��~�)JP��~��JS����tZ����Q�[���)I��s���)Jw�o��(~��w��)���qJR����H��y�o7�3f�{��JS��}��)C����%)N���R����{����`}�nf}��ǭ�$N��	  ��xݬn�[����sLQa9n�X�ۭ��P�{*��ۇ=��ݹ�gX�S��
�Ar�7v��JOO�XC��7T�ʚٸ�p����F8�r��r
t\K�����p��MV�E�'nN�c�����d���n�d`粩��<���8�Zx�Es�3Z#����H�r�dŠ�H�:�%�)��.�b�;R֖z*�r5��Ut�h+��s�2�7:��c�kk�o�|�n8��i�q��}�;��}��n�_�g�JR�����)JOw���)Jw�o��)>=}˽�����l��7�p|��;߻ÊR���w���)Jw�o��(}�����)w�;���Y�o7��o5��R�������JS��}��)C���%)N���┥}���X���#y����O����e��)C���%)N���┥9�����O����/�J���'��cc�┥����|��;߻ÊR��|ۥD �M��B��ޞrN7�ĩH��KW�Wv3������5��@<S�q���v'��^����o��#p97�_|>JR�����)JO߻��|��;�}�┥����|��?z]��E��[�h�޶qJR�����#Ҕ���$2��Cr�����)L Qm�D �M�QR��AkP�{��:��3���D �[�{5�!�{�ҋ!-�u�JJ!/{wiE�"K�\�5��.�g�Q��j �(}�����)����R�������JS����)JR|z{fw��[ۛ���f�����{��qJR�����%)N�_w8�)C���%)�n��ܽ��nX}>���w:9y��x�zy[f�x��n�bxs�v���ڲLMkF�[��)JO߻��|��;�}�┥����|��;߷ۊR��}ޙ���r޴oZ3y���)�����(}�����)����R�������JR��a�]�k4f��kV��┥����|��;߷ۊS�R�	��G�y'=�}��)J~�_w8�)I��uئDۘ�8���}��>�-�ہҔ��w���)Jw��s�R�>��{��R����w�3{���Dh�{ҢD ��ͺQdB��H����BR�?}�����R��{��R����������DS{lGk�Fi�D���tn^�k<U�t�ғ����<��(��&����)���)JP����JS���qJR�����%)O��a��MoV�m޴ao[�)JP����JS���qJR�����%)N�_w8�)I������onn�n��8>JR�����)JO߻��|��;�}�┥����|��.�G{ov�{�[��添�R���w���)Jw����)J}���|���>
��߹ۊR��}ߌ��M�f��h�淾���{���R����~��JS��}��)I����%)K���ֵf�Z����8�]���j{3�su�׶L�V����\��mu��;N�!�9sn�თT}�v��h}�߻��R��~�n)JRy����JS����)JR}}�g{��6o5�l�լ��%)N���┥'����|��;�}�┥���x>JR��.�y�7��n�F�o{��)I����%)N�_w8�)C������{��qJR��O��gw���7��޷����{��8�)C���%)N����)JOw���)J}�}�t����n޴ao[�)JP��~��JS���qJR����x>JR���┥'�_���&���I� �h��{UeM��q�
��r�66�la^W��:�6��R��]���a;br�N��a�v�"DH�q�\��4h��]�N�ے�gTc%SV��*���4z�GY���K���A�Eu����Rʒl��������*��>k��8�\gm���{�y*x�0t��r���sn���fl�x׊x�鱮9�L�d�2��y/��=d5��t�U���Z�8Sm[�t[v;�z�s>'����dk��u���j�G�B���ҢD ��t�Ȅ	�74��A$B���Y�!�����f�����ַ��R����{��l(�BRD-�n�D �@�3^ҋ")��}��)I���Z��kދy���)�����(}��w��)����R����{�������Ž�ַa�[��R�>�߻��R��{��R����{����{���\���4�ծE2&��1��s>���)����R����{����{���R������ ��˒��s;h�oZ��J6��;�"�#1�E�c�'��c,���ocC�Yۥ�n�'T��	���{�!fn�(�!Bo��D �@��mҏ%)N����)JOgj��3{���3F����)���� �J����JS���qJR��{��|��#�a��MoZ�[7kF�z�qJR��{��|��;����D��>�wiE�"�7f�D ���H���z��[7g3[�8>JR����┥'���E�"g1�D P�(I"E��C�):G��Z�����[8�)I��x>JR�����R�����������R����{��a�ú�,�-��l\f͢&�͢���͹�۳��u�˞��M��f�S��}����m���}�┥���x>JR���xqJR����x>JR������bֵf��h���┥���x>G�D	���Ҩ�!}�ݥD �X���B��M�Z�S"i���8��}�����xqJR����x>HuW�¦�ֵ���)=�;�t>JR��_[��޷���F�o[8�)I����%)O���8�)I�߻��R����)JR{��v���7��[s6oz��>JR�w���)JO}��������xqJR����x>JR���Ι�;��7�7���.�l��\IӉn�q�V;=���T�vss��kC��J����xح���{ݤ������)J}����)=�����)�u���)>����u����ٛ7�g7�h|��>�{ÊR����{��R����s�R������%)K��6�!�<R$�6�s�>����o1�R����s�R������%)O���┥'��ܮ��Z�������R����s�R������%)O����&l%� �� �jQ�	=00%A�iXA��X%a��0Yp` %����=~Dy'>�<��)J]os�3]�ZՆ�3z�qJR���߻��R����)JR{�����)�u���):}�gn�7f���F��n� ;Pq6�����7�u��v�4&�D�)�k����.�nÑ�7�{�{ݴB��*�A���ҋ"D,mҤ�\�������C�)����sFoy�ᛣF���R����{���PJH��v�D �A�u�Y�!c}��)JO};��;�7��٣y���)���R����w��|��#D-״�!BX�v�Y�!d���}��Zճvh�f�qJR���߻��R"mҨ�!{<�(�![
���U�!,ń����z�vN���]��|��;����)=�����)���8�)I������)Jl�?z�A!��f0�c1���k�p�x6�n��J�*�$!�6�x�)�I���JR$�1(3�c�h��&!��0P��HAPK# ����D���@�($ڏ3�L�L�)	$��R,Jq���^ГO4i#J��2DZ��[ȴ0��S?���X���M�' �wp����$H�[K!p��iq����0���d�󾫠���2'��đ8�M1K1.f���0)h%�`����R��������A/��qA�	LSB�!��r��G�Z ��LS��!��2A��?��/�MM���    6Ί �m"� ���          dY'E��M�q�Ni����ݥj��m���ؙ�P�ލ�$ii��UTiB��h9en�/!�6% �q"̝�*��3l�ηaьFݬe݃TN�$ �⇳��q^��bڝ
4t��\^�{)Z�1���q��v��;��s������2���2j�A�zU��]mHp��ѰmS&V���qGc'V���$]Gl�N:֐�v���Ԋ���*��%���h��s�(��u���:�ٓ��V@н�xG;��%R�q�x�o.��1e��� �{^f��&Кc��c�%VG��[N���q�lS����G\���)�l"6�6�U��`����0t$���	g-x��`�٬�RN��e��j�=3��x=yLՌ��붝�"*��4�UHKT˜q�u��ݴ�˰�;$NT��%c�sKW;���ZAײ�9�L�؇�&z##M\K�J�s��Vݤض���D�������%��L�
�ܜ^S#n��r�p���-�����	@��ݻu)I�r��	�jeU�UuAؐvu��Γcv�#M����ʘ��ϥ6��` L�h9۷ M�Dj�UV�wB܈H\mF��ʃmUN�됞��������ݧWRe�h�Ur�9�Vj�)�U�����Qb�8�!&�,];5cYXH�ű1N-�`�/:�nf H�ڴ��������V�F� ��
���(-6��T��J�G��7��YH&�1	fڃ���*�UU�Fx����2-t⊪	$�2n�O[�i[�
�}�~�?5I��ݭ��G2�6���$  m����ҀԨ3��0��M��W6@���s�}R���:�����o��I��I+�G�<�F�ۂ���UX݂����#�[y�:�/p�ہ*��N7�wS9��y����n.뮵��'�l�62��O���������w�u�& ���?���*��D�{��w��w�����~߀���k�  4�Nn�:��N�䴮�xK�[���'m��8ۂ�\0l���ޭ�H��\�v���p3^6M��Q�<���!�N����ꭍMӢ�8���ҥ%����_�J��>p9�݂�xD܂�Vk�4��[��x�'f��Nsm�r�utQ[qR{qf�6��7#Sc��:A��AP`�j��7;3O`�rU�T����u���j�ێ�.Ĵ��Eɬ�cwf��I�5� �8K�]��0�km>6�H�\Q�\������y���a�k[?�R��������R��{�R����u�p|��;�{ÊR���N�t��ֵ��F����0�7J�_�(DI���쨲!B���)JR{����JR�}�Y��Z֬5��Y��R����u�p|��;����)JO~����)Jw������<mj�"�N`��'}��>���w��)=�����)�~�)JR~����>JR��.��h���z5�-��qJR�߽�x>JR�����)JO�w_w�JS�}�R����ٶ?v��-�k�U���Dg�y���8�r��`�*H�ԈLr���l���{��JS���8�)I������)	�:U�!/g��(���ӽխo-�h�f�r��k�w^c�  �%!	T�Z����ʾ��{�w��V̙�	��L�]]]��꫖��0\���� �v��PBus5R�,�Hpo��@����ٵt5%:�i@n��F��������`>v�ܭ9�o# �M��p��}�'0n����zٚ�f��-��s������e�!G��`y�N9�s$ݘ�,f��y�otճ �kV�ȚsƘ�8t�y�����ǝe��)��B�3���s�{�p��w��������B�{~�:����e�J�7�&�$��O# �%��O#�|��ͩ��F71dO	���� ��y��m�@��\�=[�JB)"HX�m�,��$j[�����N^��K����"Q�<H�"�8�P&D�'xt��8|��:nprX� jN�������&�0���	�s�{��h+� ��X\�6���I;�/���{��h+f��� p%AT�	�&˒*K��ܖ3@i[0���{��U=��U��\$��	�1�p��� �&�@}I����<�ɋ/�!���m���դ�[mv]�/l���<�́��a�+�"�$.-c�T�7f.��|���'8w,f��[0��T�&ܟ	�r9ށ|���{yN�}���������a#��*���� ���V�|���'<�"ؓ�IL�b�w:��p������;�{���ue]�L�]Tœv`ͽ�Ss�w$�4���ʿ�dO�`��(bD����Ow~/�����YSm�  9L�s���E]ԕ��<�#zU
���R]��y�V��3/�=�����d,��آ:��ޱv�:ٕ W��s�b���9�kP�P�7N��vjG�Xr���C[��� ET���.�D��f��[�^{]
�ksѓ��!�įSE�3�0�vt�H����V{mze��5k�Gk�����1v�wwww{��p�s���=�[���+��#�D�*�V�D����oh�9,)��ã��	�|�G�Ih���\�ݽ΀�:��I+��7v�V��<��r{Ý;"��f����ٓ[�ٻ�`?s�mjגLq���q�g@��N����'8sOc@�Y���wuE�D�Y�w�{�>�� ���4���j�+	��<NG;�/���;����`�ot�VY7K�-��k��t�j��&��@w8�mA��c'����(�|�n8���˭��ڣ��oc@i[0y���np�LĜx���,M��@����f|��l�����74��v�RS#��-�:s��M��L\�ـ{�~���Np�Oc@��N�r��O�����I;�?W�h{��X��(5D�����59|&y��(��x���{�����e���~����z���}��c��@�����sӈKq�{=5dm�l�\�
׎\Jv�i��.�s�$� ���ۜ΁��N�ս�<�9�;�=��D�	���ꋑ]�:P�n�a%�d������k�o�S�w٪���7'�x��w�~t����ƚ�>��V�����Դ�#cd�� �.�z��@�l� ����l�z�h�%���x��]�SW{�l�7ͽ�<�9�;��� �Z7���cq4dX$D�3$Y�չ8���w=m�k��6�[v��<9����Wnf�[�T��ݘ���Γ�����+��w**$�h�$���{W ���4��`����*�f��7D�rED���ܞƀ�<�|���{W �Q��&)��6ns:ء(�x����v��1�_G�;��g@��8�!l��drg ��oz�'8w'��.O# P��dMYu�C�'��z]�1����.���#��۫$��'�Ƙ%!R`�Ƥs��{g ���4��`������]�TUu ]\���4��`����ڸ�x-���"X����<����Γ��<f��"��s&7O"Ng ��oz����m�:�o3�m��*$�#h�$��Γ��<f��<����b>�;�?�ȚU��&  7k����Wn�����@s�R]��:���V�v����>�3ݯ��ܦ��S���/�'[�7m�I1s���*�#�hܶ�h���Ƥ�գ�����5֞�3Z�z�:��c���5PrF��Z�6M�7�v�+��"G.��j�v3�9�nklquX�$�n�5r�p �[�=26%:�!�6�c�s�����s=�{����r�̮�?��q�l�a�Uڞuu�gi 8�k���J��:�:P)�"�g�b�ED�ܠ=���N��<����Γ��F뤘�9�`5���7vS�o6�@�� �V��j%�2]�wQ7 X]]�ͽ�<��;��:��p{5PJ�7ēƤs��v�ܭ9���y������e�E�sQ!ws�w+Ntrw�o6�@�^��?ϳ>�-�7���piLQ .��`�&lF�/m���Z����u�u�*�>և09��	<�b������8}m�@�^��=�W@���r�)��g��~m��L�<=�ݚ����n��6ܫ�|�G�Iށ����w+Ntrw�o6�@9TLӨ&8�ǉHp{f�����;�oz벜�F퐘Lr�����������Γ�ܭ9��C���\��n�Ga陇	��(ET��&����nznoa��:�K�����V)��������<�(���?���G���8�/�K���B7#����pr��@\�F������˲ꊊ����
�0r��@\�F��Gё@u�H��.� %Ѥ�4J�s 4��i]�(@ĲB�5!�K�;���x�?eDB�x��g瘈h ��!(H�	2�,Hʳ�����Dit!"~�[��� ��$�$	2~�1PWH�<^ �@3�(�b
�� �L࿅G��M�zy���z��p�<�br6dCȒ/s'@\�F����[0r��@��1��mH���p��{�?]�`�m΀�<��}�
e��?�gԩ��w5��6��7N5�D�W��v�cl[8s��
cXL�#G�I���w�prx�ry�7� �ʢ���WSuuSus�{��h���=ɽ���p
���0����Js�@\�F�M�歘�<f��D��
G�|d�$���oz�����yN����o��8�*�J�R9�'�Wu{�y�s�{��h���=ɽ�?��ݱ����F����d�:�Z�4�&�wb�3��;q
��<7<N�V�!ZT��5�]������0rot:Npz��Ȝ�ŉ<�Q��@�m�prot:Nprx��pE:�n��j��&�0rot:Nprx�v�g �根&6<�$���{V�o�.O# �M�8r���D͓W$LM���o�.O# �M������ʰ?u���qQԦ)	iY \���7����Uk������Q�%igHů�f(�Ӊ|FN#]q$˦���Zâ�q7z��[k#Y��l\��{.(�C[��F�u��nu>y�ݍ�v��n�ν��!��\D�v�qϣ�B��d(�Nѻ6��܇c;3�gv�����[���v���ї���	��:��sW]X���0)ۚ�x���Mў��W��N��=��{�����~��,J\i-��"���6�ِێ
�8�Q�j�I�mtOg9��#��Wծ�5�˲O�0?��<��7��'8sx���N$H'��g ��������{��}���?~�T�Ԏ$����^�t����4��`ͽ�?VTҲ&�Qc�I ���:�o3�{����ڸ�CQdNF�Ğ$��$�F���Λ���g@�����O��y���ܛ�4k���wH�o]��0�Xƞ=��r ��j�͆��&�,���;�{�y�s�w7�����w7\�G�Iށ��UJ�(J>J�Q�n�,�:T�ۻ �U���8�ddŉ�pz�S�n��pz�ށ��NV�uئ���u�hz%'�`w6�@�W��#�[��ĉ�"|�)&pz�ށ��sx�$�052�j�d�uq�M��vFy�^θ��z3��	5�m��&H92(	LjFLC���@�l���3@I<�����je��T�WdO�7f��3@I<�����e8�CQdNF�Ğ
w�@����^����/t�
�~Q7��wېn����c�	�$pRc���=ͽ�<ݳ �o�	'xj��01��xa$��������@7v��[{�=����J1�F<2,\cnrem:d�aol�󡣗KȊk�mѬB:�#�	�r5#�#�ŉ�pz�S��g �������j7l��c�6]f �w�w6�@�v���f���*�D�q����$�������sx� I;�=�R�e�]�L�W�7u{�>v���f�4��g����dݗ���ʚVD�'!�R��3@N������ ����s]��jVS�Zn����܎��nM/f���)���jz����h�~w�I�����`ͽ�KPe��6�'�)' ����� ���΀[�p�����$���l�;�{ �w�w6�@k�H����MHpz����g ����� �Q�d&�<l
�����0����f����$������_���t���  Mr��.ݎ�,E�[��_��^�F���y����gms�y�̘�sZ��{`iy��:�Nʰ֣=�v�ْv�l3�u�W��j��s�۠�F␊��΅��8�',:x�e�:�rvT��%��۸s���ҍ�[���$���[N�j�"v9���5-��mzۚ��;z'��n�!Iֻ:�'m��SMZ�$�G��8�hv����<��^�]KaaUxu�׊�#D�]IqED��ǀK��۠6��soc@�o3�~���*�q%��s�݌�Ē�37vՁ����6����s�N��RH��JC�{���@�o3�{�oz�)�?]�B��H�<"�i�`ɽ�;f�m�h
^�c�ncny�p{m�@�e8�mڰ�J�؄ޒ��$�9�޲rVջ&�JuH��yF�Kcm��Lb䰦c�FE�L�7�a�r~����� �6�4���;�{�2�����շ3Y�ܫ���|<���Q�	�CǷ�%����0='*w5���QT]^F�4��ɽ�;f��:��Uĉ �c�I8���@|�soc@N�z��E]GP1���@�v��[{���g ����=k|��,�H�1��0Y*쭹�]�ѹs�6��ק��\sq܎�>�rdA�4�2H�2H��m�t���[{�/���?]�Bw$�8��s��'��w6�@}I���������I�<�s8�m�@�{W�%�����/���6�n,�'��%]������3@}I�菣��W=߬Q�-s{����:�����y�3@}I��M������swSE������Wa��%-��t�l�z��U�QG\r�b�y58����� <l'8t�Np�otԜ�汚%#��$���JE�=�m�@��N��yN�|����P��8�K'�Rw�>V���3@s���M��C��w#M'24�E�?z�)�*���=����+E7)������~�3�v�j��LpI��xt
���~��@}I��k��ʨuqSs70���hv��z�g=nN#�4��.������}h�0$G��y"��~�{�/Rs�{��hy:��S����;(Gy�݀��sZ�Of����Ǽ�=��ހ\��Ȥx"d�%\����N��otԜ�zNT�j�w�������ԡN���=۰���?z�)�=���% �h�7�������`�{�N�}���JZ �7s��fJ�PWL��)hu���J�L�)����c��M/8��t��-ZF��� J��a(+�廍!)�yx�pY�h(�h���IH!�e@rJd�B�!$�CT�b9[�D�SG��Q�g�6h��!:yϼ1-p6�EUA�#=_I(}SH���xC�%-42�c~�"Sb�`�&�(H��44�XTC`⤌0dScAcT�fT`8���AUS���S`8��4���/�����M�T% ERKV��+2b+ɚ!�?%�@F	kV���f�kZ��   ��@ i#� kX          �l+^q��[�`*�mxs. �&�J�m�Zض��횕�O]�&��1�iB���m�ݜ�c��B��"['rfN��`�Ԥ�qa%����T�H4����.X{<W/U�����a�WA�q�s�Nd�����t��<OCJ9��ƣ*<;v�6x��$͵�d�l�T���f��3�U�	�g'j=�v�[3��f�W�s]�:��O%��*һ6����.Z�rUմ1�u*%R��/a��H���UUQ$ܲ��n�,�a,�c�J�d�HBب�'�8J$��knW����	:�M{J�4&,��n�6 6�:�@��%�Y�;t�����k*��`Y����6ĵ�U<���RQ�����1��N���+vN�b�&�6��m��x�v�fi�%���-��zY�� ���Jv�ͱ� �n��n�����ҫ�pH{�v���R�y��"�R/��^� �K7�^C�n�W������)�q�3�
[J�muUN3�Z����X-ѧH��(�kBY�`��U"櫶����r�T�]��.WC��^:!�u��0 UU.w��ݝ�Q;nȫJ�A�����nu	���i'n�9�1�ۥ떒f�Vݲ�'l��U��m��qTi���%`�U(,��n۔9�)g�[���g�\��taj�nL�`Ms�!n���)��4�UP�����U�nlޒI";P�]T�չu��*��,�=��7m�6h�x:ٮ��D1�\K�Zp�KJ��U@�iw��EZ�$�PZ�F:�R1n�)Z�����H�P�x��Y�,��n�bE��  nڒ�k���I�B�Im�ݙ0j��� ��$u��Tr���9�OT�<��m�T�u(��T��	��� mmI�Ӓ�n*t�(�U����v�-�m�b�§��g�����k97H�bF��n��^Z��Z2�Y�6� $~D������]�ߛ��e����Z�� FK�/kr��T�ݛPF��s�c���hm���<g7<k'n8�r����X�	����aDֱp��.�����W�YN�u��Ξ�1ٞ��ʣ��+��G�wn�����c�U=\7���AӹR�T��y�Qrd&�\9�n�u;!�����ם �83�qIL���m1n��KnEP�g��/kׅ���ӯ��3uʭ�d�Ӵl9�k�n���;m��u��R�㧝Ւvs�.C`�q�(�j)/@��g �m�΁V�|��{�?\ti;������I5q�.M�hRu�y��@|�G �wD���A"b��;�����ot&�0ɽ��@;������*j.��4��I�`�{��|�sqe�>��Xa���o3 \���<�9�<�{�~�#�rʪù����x���&�[I�仇h�çY�!�=�κ�x94\R��Fv`�p���i����zZu�y��@\�F ��US�d�699���\�ff~�2g�d$+�o�����3�ݫ��M���G����x��p_���>/�3 \���Rs�?@��
���J��{=��l%;���=�V�1���{�?n:4���ӈc�r}��4Ԝ�i��+f ��UQ.�a6�����͵�l���pͽ��3[mm����rE��"br	9��'�B���/���=�7v�1��W!��ZXq�����Li�$��{��ށ}�������\o�V$��o"���@|�F�k���Em��Np���l�9"8����p?��3������?Ӏw�{�>O# s�r�Dݗ@U�a�>�� �&�@|�F��yN�e�V�LQ��ԉ�a�s�3l;����B;Gj4u�񮞱u�m�ο��~>:�RJLr4O�Ĕ��o���z�p޻�t�j�����4!��E'z��0sX��Np�ow����W���44�&����ן�@����BS9�ݻs{���x�zs�g�37$��s�� �6�@\���c�����ϳ��ￎ����$��$�ye���m�0汚:Np��ϳ�K��<�4��5�fIifL�f��#R*mf�E��緱���Û\\%�u{2UE�]���5��F��3@�I������x��L��&&9�]�^����7�f��n����PrOkex�&LX�Np��j��m�@�[����S�~���%#$H�&
n� �6�@\�F��3@�I���˛^'��G;�7��8�w��<��h|ۻ�>�P�
�C�&���I� �mb]��j��+'=M��Is���)�. ��Cx[c�ۜ�t�h�ڋ[#V�{0��1ֆ��U%+�-�d�i�y�rѸԾUbF�3J��y��`(��%Pu��B�ɧ��5s5UE!��c�d����g������f��n��]׬����u�EI�&&�<��r0Lۧcg��/\&�ҶH5�:�9�%tn9�����㾿6��?��x�{%ӫ
�]%ۋ4�l=ՙ�6���Mø3s��m[�� �&F���� �X��'8y��}�.o# ��PN�CfEJ!N���j���fL��ݻ��*�<�X�'0C�x��Ĝ�G��.��oz��g��{vS �I� �B�*�*ff������F��3@�I���� Ӫ�WDV\MWIc4�I������g �~��+PQ��qɐ0m4B��^�����n��
U�md��	��������ASw�h�9�56�@\�G��3:�m��:���5Ĥ�#D�1%$��{�>o# �3@�I�@�!Bu%YvW�sw���0Ic4�j��oz��F��sOj� �3@j��Sot��`�n$�8��$�ħxt�j��oz������:�Xݍ9��`��n�a�I��]�|=a����\��n3��^x����"fG�85&}$��wm����`��hRs�7Цe���UWz�������U�!L�ۭ,|{4�n�TD(�R�9�.s���Ӫxs�T6�KϘ扄��BMyDUyӻ��o3��ڞV�Bdō�Rs�@j��Sot��`��h`�.$�8ȧ͉) �ݽ���8���t�j��H�: j73C�gP�Pb3��'v8��5̑��]����LM�<q��@M����y�n�S�]{W �m�@����w#CNci��:���/R�2k�٠7^���ҭP�B�=S<�ήw���fg�g�E���f�o���Tx�N`�cĜq}$��[���_[���Xj�!(�W[�{4�(k�GRm�0�����8���^��;n��e-�8"2LA�5U:whG�m����͉5��H�M�ic�D�:�#������c����po���^��54�@|�F w�SP�B츸�����NpM=�7��r����g�f|����q'��E>lIH�����~n��(��q�,|{4��skC���������8﷔�9�h5BQ
~�{��湧&y�{3��UT�U� �,f��'8�����ʿ���*��_����VoY��4o{��� �j�YyW.]kY����.k��;\����U��2ѹ�^p]��dZDb�{;8�gc�6xn3����\0<�΍��t��-���ś6Ɏ�G&����{vp����^�� ��ƛY*DRr��a������Od��f�.��m�[�t���U8�n8�
�d1;MY๧I��7mٕv��[�I�������Z+�[a�*�x��N_6�p�n����rn,)��x�����W9�g�O}G��湠-�w`?7J���S�j�0v<MĜQI�.�S��y\��T��	�B���dM7&�s���g ����ڸm�ހn�a����c����p�c4�9�5��@|�F /��XEɋ���ڸm�ށ}o3�n�yN��ڐ(Ռ�Hd�6��1��n�m��<!��a�y2Sճ�a��Z�����I�")�bJE�;n���iP��f�$����h����$�N���7�������� x �7�-�f��I�����S��������E@U\`	r�hRs������8���N�� �Ģ��u�[Ot��`	r�h
R �u��'>rE�;�oz�������ڸ���c��r� �j#�K�͎����!p�K�'���Lb䰦c������3̈ȚnL1��:�������ڸݷ� ݮ�s��	������/a)Rk�٠>�{v�t���X`�����.���m���/������!�,
HI���4�Y��WDU��qTM!"�"ld���f�	F9��K� ��	��� �"�
���	f�J��($�dD���q1`0��&
���W�0<�QaT��(?��Q�UR�>��S,�c9D���:W�D�����@|�F �x���p���	�c�';�/��P/^�O��ǳ@^<w`b�|�#���f5�y��[�]b�m�sۮ;hL�:�ͮ��݇Y"�dP�C�����ܹc4�9�M����0��˃��Ǌ���.���[���_[����:`j�0v<M���9�� m7���0��hRs�'�C�14ܘdi������-��yW~���W,�8H�D��!�M)�w���*�w��Z��i���(���O�5I� �ot�Ҡ5%�4�����)��bQ3�R���s&ӭ�y���k�v�y�ek�F؂���B~����_$Ǐ������.n�ށ}o3�[����mI�?�R,4�� ���4�T���)khP�K���@����6��:�j�v��n:�Qci�1�:��O�5M� �ot����7�q+1�i��S�:��p�
z�~��iP��,�I-�G��	eM��  �4���De�N�9:�1�M� ;;]Gg��cp�mGZ�5����kU�L5�e{3�آ�N	��x��;2�'k�K65��2�xq�3d�]�ZlӍ��k7bZ��N4<n��3�	tc�ub���*��s�G;# +�ks���;t���-�u���-33���mz�jCg�Vq�;^�۱��x'�����w��j��7%�e�A�t:{=O����4sٛc�I,�6ݧ���������������xR��(������t���O�s�W ۞���LCM'&�s�v�g ǎ�`y�1�w{	L%!��ޜ��<�73�_����]v��m�@�o3��jj��Ȧ����#�j��4��7��&�3@���L��?�N.�m�@���8ݼ�@��\sַ\��F�*�=t�Ў�;-������=[Χ��t�N�u1���(H%���Nw�]���6��:�j�v��k�!�6��UET�\`	����}�z���s�?&��]���7�q+��RD��Q
w�@j��4���} �yi�4-��ĜM�1� ۶��]���6��:g�e�j�sٸ�Ɉi���sW�M�`����� m7ށ�h�X�YqLN�n �H�qa`��.���֭���=u���4-en_ns	������:�j���Ͼ�m�p�ښ�29����'8t�nh�7J�o2�I�6��)2cX�lI8��oz�y�;�%n�t�]��w�����M^�4�F �x��np6���ZC�7�n|�6���7v����m݀�T�(���7NqO�����ݺ6`�͘�n��g��׏:��rׅ��;��_p}�t�eql_}����n��6��x�*َ�`d��pmH��� ����ϰ.���ݼ�@��\n{7�1190�G7@i���x�>��� �m�/Wr6�7������yN�uڨ�n�<��A�Y	vQnx���ښ)��@x����uڸ�}m��o# I<f�C��n���X�&�=%kc�.Mm�m�u��$��;v2��$�;3��K &8b�cX�lI8�������7J���L�H��|�n�����q��!��i����8��S�]u�������	D�,	s2��)$'��\�3@J�`j�@M��&�U��)"X��>��]��~�oz�y��ϰ�m�:�i����ԋ����<�{�6�F �<f��79$w~?_���&�%�H  6�Gl3yY�	���"�y��m�\�ݍ���A���k��W 4v{b�T�lan�xzt�;+uvݹ'�%a1<%����n��5;[�g#����gz��M��[p'���aP۴5PrF���^���v9V]�D�utqv6�ɨlp�qۮ��ݑ��*�:4HN=�����%�s� 8��N��>u&�j6����������I�e���4�F�1�=Z��8B�(��9��q��;�9A���ϻ���wܟ2bӒb�)9�?z�g �m�:���?]�� �W�#&)����P�t��74����R���jh���ư�'8t]��~��ٰ�L�ݥ@<{ZX0�Wz.����\\�3=��l%P�O��݁��J��m�:׵p�[j5&	O���@|�F �<f��'8�ot?v��7�<Yo�٨F��uѡd���0]]��=n����\���wwO�!��y�_�QU3W��T���{�7���.ۉ\�b�%��<��k�5�ƥ*8�v���T�:e���0R67#�L��_m����p�@��\n{7�1jI1�{v���1�����2o֖g1�}������Ɋ|c� ���}��`jP��7׳@n=۰>mҠ/�V��q��a�i�% �mu��.v�Lh�j�\=�4���O����O�֡����PE]�T���{�so# |�S�~��rC�1�li$���oz}@so# |�3@J��}������7;�=m�p�Ng���gsR1U�W@C"�҆*���d1��G�M�0�F�sSj2���?�������߿���~�F��7�n32f�0��4�9�&�@�o# �ڒ�s�,i�!>���j�ء)������ۻJ�c�X�}�?m�㦍�,X:�j�nXՓ��N��\]�2���{yظ�M3n�&Zy����c���*���
"���9�6�q;�6��!9ށ������e���s@|��̃�O�'T��ހ�:�絥���sA�$|����� n�SIX���dXc��:g1���w`|ۥA�
"���P�y��}�M�/)�7Ci���ěI]� ����y4�T������쿡���v�u�i�8r�&N�z2r��Km[qV=ewn:�k3)vs*H���9۰>mҠ<��,�c��ID�v��~TIZ�x�q�����=v�g1��m݁�n�B�J ��3-G1Iƚ"���������~��8��S�Um0�47�2L#�@g�w`|ۥ@y�X
"Fg1��=��܌��$������g ��L�39�h�n�ދW�P���%5I"C,j+p��&����e$ 	$�e�")5S�J�-kI@� J� �M:� �
lR �p,�!0B�X� �B���</	5$w�o��<ЬℲ�$+�A
��Œ�H�1)eH%]�݁�*��6x��<��X(8B7���z���    � 	-�< ְ   �         ⫎y�p���sۮ,�b������'�	-�	�北]�Vs55R�[�H �%�d+��4�[�Id���\v�ʹ�i��������m�G:�����6� �#GZ���2���q��҆��\�ף
ǤȒ�q��"<�u�&ӵ/��,F�B�E��GM��;M��r�J�+��"��@uS�յt���Uvl���8�'�͆j���cJ��#HJ��"�@D����ڒ^a,�����
�q�.�T��bPH�Qf"!l	>�s�J��įnFꪭ����+�Bi�E;Ŷ��m5�n�D���M��6��K�� uT,�0/#�v9e���k���I��ּ%&e�����mv�t�v�U���0��N�*�9�Z��-�m�lSUu��Zw�\�Z���`��A�yV���ؽ���ݕjv�Gh��e��s�J�;'FұvĽeL���kTZ���ִ+�e	�ݫQ�jڒ%^3H��U욒�X2֦]����YC�li��򎖵����BG��B�.�/�U��j�0�` !RTӵ�:lm�h�3�5k�z�O[��X�z:���P�'��QV=��ycy�9��:�ݩ��g`*���6�P�G�(D j�ۧsI���\�UV�vcbՌt�@�ېS<\�UU��N,��Q-+*�W��(1�<+�K-�pBޚI-��X��N2��5� 4#���t3/Ums��j�ZU���^an'��U[8�S�ʪ����ؘ�0m�l�kkź&�D�]u6�m�lH��  m۶�Vmɵ�bLQX.��F�����Jk[E,�jj4=��q5<�&�{M'�C��¬�A�Q��ت�P `1�ݕh�
3m��p��˱�톧��(��b=g���	����5� ��,�n٪��i{f�kY�Z��@HP�(��
?�S��� P���T�P�辊��>
 �.�}���Y�f�d� 7%im��N`٪�l��rF�뛮0��c5q�c�u��c��Wtݵ�p���[uf�q���ŝ�� ��gɵ���׳�י۲�>�\�Fl�����4�n��\Ao�h�T�8=v�P7;-;v�$nT!��::���y��m��s�T�w�6WX�m�tn�爁+�81̈́J�(C	��#��qJh��st�s�R9�wy�.�Ì�F����;�Ny��A�|sb];��{.�X�t򾠈PȖ651O�p��3��^S�fs������t���>rEb�3�`����������[o3�z��:}�g��o�LMLI�����sot���9����� ���|�'��t&{����~)�ݵ@f��,���(Q�6���Y3-�y�F<x��p]��@�ڸ��ށm�����v	HE&D!&Hܵ�Y�\N_6��S��n�`�m�n����v��������\��% cO�àZ�\}m�@m�Z��3^֖�wDw���N�w��Z��}�{�<>F�bH�"���T��e����Hז.>���Ԓc�7;�-���.��:���/���՛��Q��B Ng ���`7��~m݁
mҠxX�B�a#Ƥ��k�p�oz��8ݼ�@��@�V0j52���V��P�.l9�+u$��K&k�9t�]�>g�>9�!�Q	�����_[{�o# i<f��78�'USu57�|U^����4�3@n���m�L�����F�1�bx!�������sB����I$+Q	Gy�g���o3�n�ĬƜ��'��74٘��m�T(��������29191��p$��~��ށn�g ���:�j�h�̓ƛ�Xa�\n͂�֎�'�a-m�\��sF�䰦c�����s���Bdy$��'9�-�N��L��9Ԕ\��{v �V�橞ĩ��
��0I�4�9�<�{�7�����.��c�E�I��Np$�����jO�s�j���ĚI8��ݽ�� �ٵt?}�����꤫�~�mm��	��AUw�jـjv���s�rI���#�E!!�O����aɯ=X����\v��̓��Cr���+������G��5D�Wf��s�7I��'�F�ںp۸���N��qt^��P�Lm����P��͐��m�w�b�|�H��v��[��?���~{�ٰ7x�hيx>�����qL�a�%;���>{�ٰ�9��{3/z�e��%>X��ݲ��5DD$��^́�����(	�DBS!�1\E*T0�C�������	��  ��i{n�	�	Ҳ�vJgR_������lZ��ιú�����#���8A;(t�'b�Fۃ��h��gz�
�!%�(���LܶlfƷa�5=v��v�c9Cu�C���v{�(Uu)'c��k�x�q�Y	ƛ�FFcE�n��,����n���˘�Gٞ&F]����mu��
�����w��l�:�B�n#���ou%�T9��^;p�ܺtVc�5�ؠG�Y����˰=[K�i�����c��wg��������rI�ڶd} jv���o�I#��CI' ����vS�wl�t]��w�i���R!邪�tݳ ���>��� ��@����bo��!�p햮��78$��}�nـ'�%�WD���/�6|nh�Q����7v�e��}F�Y��(dh�.�U�]N���s��{x�l���;s���e�kC�$�$�	&B<j�pn��@�e8v�V}�׵pi���O�k$�qL�`7�elB�D@�B�K�>{�ٰ7y�4�1݀c���ĩ���n�S��@n���>9$�@m[8�_+�Y"I�ȲG98��j��{�6���m΁�ɫ����CI' ������/�� ��j�^��.m���H���}#����M�Y�Jr��޺�K�5��p�F�<���X�r`<c����p햮�u�\ۻ{�<���bo��&�8��sz�DD�I��f���݀���o��q��"y>�.�u�\߾��yxpC����H �G�5��� ������v�I�� ��	"����I=�;f��s�5I�m7w'�5�I����)�.�j�vS�]���yQh�X�YqE��⠩�胄���;'f���K�lq�u�99cF�Ͼ��9ɍ�>X�@9v�V�Ҷ`6�@|��'.IsWi<�$s���]�N{��ϐ[o8����us���>č�o�72	��L�9Ҁ{��`?>��x���3���UJ�m�&1���C���31}�$�nmi@k��̀�:�x��	@����s{�;�ʾ�٘}��2D��&�8�-]��p�����P	B�_='T�N�zs��!vwaqp�.��հGVݝ�s�׶<x��'�<O����{�>�1�g1r18a���������v�ށ}e8�-]�p�$�ɐpjs8�oz���l�t�y����30i��W&B7�I���;f Ӷ�@i[0�{�	�\N�S�@'3�]���/�S�6ۻ�	B�~�J�21�L˞t9ʚ�������'��6���y�Z��}�o$�B���)$�I$��K5��K[%]���#�x��B8�#�/)�ܪ���l�Ʋv��d\�]��gZ^�%q��mѲ.W�uV��}�c��]c���8��ݱqT%���\� kY<n�����`��rCU=t�(.�������v��#�W�9���09W1�зrb�z���,�&z�!�n	fu���s����87�=h��g������	>���;tq&���[NRP-��)���v���gWZ�:se������X�"��Ѷ�HNL������@�����j���>���y��ʩ[cRITQQ3W���0ݷ:��0m���YlM�$InC�[es`?7J�!(�6ۻ�:TcMM��N#���/��8�����m����v�I�� �J�U �n��BP$�%�����ݛ��g ���n� pLY#ƾ�$��śE�n�F�2d.����ǌ��P�x��<�D�4�$�s���g ��W@����-���Vn'r&�A �»���7��LQ�BU0
�B��BaR`�E誦�< -o��ʽ��T�*�2��:qw��]���ڛsv� �n���P��60�r��HdM���8�}�����y��-]��g ﲪV��r`Lc�5{�4�F ۶�@|�F �ot?v��7�<Yn�]ڵ0�+77м�7�m�mv;M���m�mX�c������м�	��M9��-]��m�����r�q��<�g@�m*����@6���
}/d�$�(59��oz�y�9�0��RI	���t�R������8ɛBthH@��a&d`�5��p�m e�1�p���4�� ma&1��Q��Q�~M� l�4
��~A\A=ϯ��O~]�����yq�"mG	����o# m�s�4�F��@7kˑ�� �m���-]��P���m�T������{�L�Y�lB�+8�뮱��v']��e^�.�ۮ�|��"��d��q�D��,��_�����Tm��7J� ��s`c�WV)�#i4�$�m����m���v�g ﲪV�Ԓb1�Nw�4�F ۶�@i������L�o��.GT�L�y�A�
��ń����oz]���6�qX8��J�������0�{�4�F�۫�hkn��I"�|dQ�3���']���&ӹX�+��4���uu�4�c3��(�*l&�0�{�4�F��s�]���6��o.<dL�LhNw�]��l���wf�׻J���w`����S�L1��p�-]����{�.����.�a^%o��'�qt���I��y�m΀�6S�Ȉ%1�Ф��7woz�}��}��wmXn�vl�Ҡ21(�(H"AM
Ã ��@PSD� ��J�,��3]����*[d�  ݮ��m��k9՛�ת�ܵ���[n�#lA6F�H=\�k��s��$  ֨19.���m��8�Bт��2�b��uv<͵����� ���[�p��{y��ˬl�J�n�F�R�I%�γ ,�jY��N��ѶY]=9�xy}�]un��Nw��L���8����l<�֤��E�ǝ�t�#CWY��b������owy�ww���=���zc��t7;����q���\<�8��&�x����;����-��䤓�'&������;l�t��8���@����bm��`�&����s�4�F �Ot����q.18a��!�qt�y�wv������e��~Wn$��LJ"��$�����5�nt���)��\xȘ䘐��@�o3�v�l�'��$�������J��'���t�r���A����,�ya��,[��}X�!7�#�X �i�p�-]��0�{�>v� h���I73�;Ѽ�9����xsB�	a�Q��@�@�	_�����I'�'l�5�nt��v7ESLRL�������g�DB�s�n�vlz�P����g��T�T�]��Nـkv��7��$���~TIe�&�2 x�R��ՠ4�F �Ot�� p��vL�ŕьF	��Yv���=��"��Wcgn{!��lr\nSG~{���>�8mۦ���`<n� �1݀����\��{�6����$�$�Ģ '3�]ݽ��S�_�Z��y�� ���yq��;��'����(��s`�BT��A�f
��m�� ݯ.G0�ĂL"�����s�4�F �Ot�� .�u���XG�qt��8 ���1Հ�������5�2\���e���`�K08V)Ǣ����D����wk�/7Bդ	Ֆ: .A�]����݀�������7J��,�KlJI1�rw�]���>�0��W@����.���*�2؛�}<J�����:I�`$�@|��pV1<���b}�]�32��g*��}�<���}�^�����Z@D���T}�^y������K����;'By�@<�w`lBIDnmi`o��f�y���2Z9<�����d4��l�f�֎���ls��qh�p�fqrXS1����w���r���B�Ɇ��a�`�ӝ��0�{�	�:VO�	0��C�m�j�v�8�m�@��� �e�4V��5��G�ɰc�@cx��Q	$Ϭ�1�t�n,�$�1�93�m�{�;f �x���0�)d������<m	9ށ}e8��}�fݲ���g ۶��<ϳ�/�m�Q��� � 4�dn�0��i;UPyu�x���h��&�O=�p�B*���Ӹ�ZDr��t#P�����d�G]nZL�m+�3�T�У;���2q�:��A�ʆZ���϶vu'Q�nT�F�H���t۫���s�6���k��1���6�ۭ��wOb7N�iw݁��nT]=���=��zP�i�=��]s#:�V�v�SFl�TD��+���{�߾�^��~_�M�b0s�<��vi�#�&�ӶԧVsu�RI�!42� ��74<Fn�vߛ�ZX1Ҡ1�w`?7J��cS/�;�y�󤩞]�t�""�1�w`>o# M<f��YawT�qaUq�&���yi�4���-4�n�q&)#����y�n�e��*	%Ǎ݀c��q>�����$���O�4�F �ot�y��գ��w�'��jD��&�'����=�����/mh��4���j�s�RIuS��w�h'��&���|�}��}��ݼ�@�:��ȢK&2����M'���O�4�G ���ES�<C�Г����8<t���@<�J�Ǎ݁�&�3<��OW9��U∈J%������� ۶��_[�����O�py3[���yi��O# M<f�e��f7���	,��d����"P�	����Omێ��Þ��yz��ﻻ��w�v��$�5����v��v�8ݼ���.ِM7�7�R!Ȝ�@�gW@�{+:T<n섢!G~S5+�cD�`�s8ۼ�@��w�/AaBEe$�S`����}�{goz�y� ��m ����j�:T<n�x�PD%�v�ި�|�#"cNL�	��@M<�4�i�`
9��ق�[���=\��ܭ�6� ��U�<M�.4p��)�ls�܎!�C�x@*�@M<�4�i�`	��@�ؓ��6673�m��tϳ>�>���My��e�WD���Փ5�h	���&��4�0��;yW���k��[��al�k[9B"�7v<t�x��(���{����.?��$�Nw�m���	���O# M7�J%U1DL~����c��Z�Έ8�����!ck�W���=t/$LOI�q'�73�m��Xx�P�IB��<�* ���dm}Np��y�n�ށ����6��:����,�$�!��ު7vy�T	DBI��,<���٪��%"hǉ�����y�4�4�0�{�t�������*�j� M<f��<�4��_{���_/s�|�'�a���Ƃ���M�ps[4o���J=Y�r᷆l 8;�䍂���L$d��E��Յ_ �O�0$��lp�.1,IT5	�4
bANYijC1Yr0#`��%�X3$�M�=�zk�'[�\8����2�����B6�!{���S�6�$ă �,�T|��f{�i�� )@ � "�m$x�``      �   ��,Z#�L[4��f�`!���hon���4�%ږ� �Y��y�[�첳U[@P
������C�F݇��u5Ӵj$�F���u^�'bCEyǭ��%�����ƒd����ۮ؎Љ�N[�,�
k*�U/ �U*gv�r��W���p'C����m�PsZ��I��.��^Ku�vW��I�+�vof�Q#g�ܲ��@umP'���J�j�%Z�����W��[{km��؞�T�rL�S�t49V���=f��/K8
���G��tcK��k�AjX�F�F�0v�V��Q���q�y��4��������*[��I�^Y�D�jH�mp�l]UK����[�r-AK,n)Rۮ6tU�d�m9��d��[Q�᫊�c�\���[nV�v�^�e����X��u��\k����7�ǙvP��d��
�WLW+��7* @�Z���3.�Ke�Ef��&�N�aWZ�n+oIb7�^ �Ʒj"{<i�,� ��T�5Nf�n�8���4a���Y; ��e1�ya���V�	�]����ݎr�pl)�*K�I��m� ���7hV���(t�I�:�3kJK\�P;�غ��� ��J\@,��d8`7=5�>�n�`�,��z���<r���&#nlgvۆ�8G-T�뛗k9a�mE�9Ƕt���UU�ȓ�R;$[Umr�1�#�^W�m��K��8�^U-�jes�S�+.P&���)����YqIV�U�Z�Re��C�Y��jyZ��McS�^"���9d�hK��հ.��Ojv�O���8��
�  m�[�k&��mUT#�q;�xM��__m�;G�f)eX
�U�eBn�U枪}S��Z�[�.��(Z䕥@�.pݷ�h���\���*�rkl��+����/^����s/;$b�b��\R�9V�v��ލ�Y����o�=��<��QqD�/ ?�����WB�����t������I� ��\띹Y+q]�հ/b��)�F����۠ܽ��v��u���Ä�8㭓���pv�8�P�*�̬���3Ƅ�r@P��ݞ!0x�e�C�=��gC*eݸ�8F����5:�l��w8�ͷ���R��lsR��c��:�����S�0Ul������Lש��t.���q�O^=pmڷ��[;~�{������c�?V];�����|�,t.�pq��]�pn�.��-�O����w�������qS__�VLL�`����# M7���8ݼ�@�v�>dd�""`�� ����HJ"&G���������J�/����M�`7I"��9ށ���@?��,؈������݁��Z�}�"j����f�� ~O�4�F �'vD(J��@�NK�+�Ɏ��j��:T�J7߾u�*����_%�8!F9�#�#@� ݻM�\ɱ�����ۥ�phn�;�������F\��\7EU]Ɓ�7�t�����h��p��%"x��������U���P�'�
.���i`k{J��ݽ��}���$j?���m���llo���=�,�Ҡ���@<x�_Nw��;�IS<�,5DJP�^ڠ?&�n��y�x�Ͳ
Ⱥ.���fª� |����0��j�8���n�"��ci0k1�55�l��(�V���%�s`Ǳ��U�.(�Ƴ�l�Yww0UW�i�`��4��ϳ>�v��mx�<�!�ɉ��6�p��i�`�{�6�F 4CRT���.��໼�@m<��Ot�̣z�!��BP�D�����;�o)�=��Ȳ9�Q����U��PB�;����iP�t΁n�g ��)jbR'�x��rw�6�F ��3@m<��OtK �g�Y��Vҵ��Vc�Y^{b�J1g�.��9�6��	��}�;o��g�e˖� ~O�6�F �'�i�`�L�����w�&&ytX�[2n7�`n��@?��,�b9K�;��d���*�0�=�O#��<f��y����n�E�bs��������kK�t�9
I��Q�ُ��<�!�ɉ��6�p�o)�>�ݼ��m�@�o3�w��eJ6�K ��&�bw9��'m����䩭�ۍsG��1���9Ŝ� ��ЊI�ݼ��[���0��h�GEe�]\7EU]� �ot���O�6�g>� ��)�0r6�x��s�ݔ�O�6�F �otU.`)�MU�T�Q5Wf �x���0�{�[���?z�V�O��p_$�à[�� %���t�x�DBJo���k��l� f�,�S�!��x�^eW������q�E!��ㄳnn��A츈�r�����iE�q�����׮���;�]��Iv��ǥ����wpe'��.�.��K�zs��9h��#U�pg�l�vMca����۴{���<��~�{Zك5��&y� ��\m���ѻ>a ����l�����lݽ۵Ue������k*8;ve<A�)�\�n�X�f�$Þ-�v��p��Qn�Ӫ�h'�s�^��۰�J�ǎ�`7�� ��q��p��,���v�9�&�3@m<�4��	�K��qdU]�SUWi�4���M���g 7�Y�D�ư�2��:��0�{�6�F �x���謹�&$�����m�@�o3�m��tv�8n�
��I�"saGN���'q�M�-p�:�����Eg4N�;lr6�x�hNw�m���v�n�g ۶��{Z��4�ā��Ϊ:e�BJ�Q���J�z�n�۷��?]�bO���'�n��4��	���&�3@�l��.�'�
!��6��v�8ݼ�@۷��-4�n��!$�"s�4�0��h	���&�������{���mв�b��zC�[px�Z#�Z��v"�<)��+��竭�FNyZ��O�&�F �o~�4�0}�TIA�1L�E$���o3�mMyi�4�#�.ț������U��:Te�%	@�CK��Y �H�y���������s8�����!�	���O# ^i�h	���s��@�R���"�cm�����t�y���{�6��p�n�`�����Q��kk<�ָ�9����t`.0��N�m�q�K߲8%�c�O��y�9��v�8���4�0�Ɓ��d]w��r]L�\`�=�O# ^i�h	���=|Pn�NrE��9ށ�o3�/4�4�"4�0|��	�K��e��T�EUU� ����O# ����$R"�G*`?�=���9Q�VmQ%�S!�Ng@���p_c��n��<v�J!(�s!5��ʘ��$��9]z˄:"d����p�25�k$�gt%���yC������v�Le����n���F ����9'��/@�N������B�j�@�o# ^i�hݼ�����Z�;�X�6Uq�/4�4I�`G��=�<���/�%n8���G�}�΁�����Ot&�0�Ɓ�L��.�����f�f�� �����F ����9'�ʺw�?�قR�P�K��_{�=�{��?��q4�v�L 
��v�`4�\�4��9�x䍨
ݳȞ�3�Ƃ"�8��<� �qE�`�a8U�:��"W"q�vt`��`��ZG�6[�mr�q�m�;�g�r�]��mv��Հ��9�{�}$;�� f9���x�3��u�ܼ�n2�р�h�n<�]�q�8�n�tk����]�򼻓+si��v[I��y&�v�<q)lC�:���� s�'�u�կj޷ٙOk΂��Y-�a�x���Z.���c�<�k(uge�i��D�(����p�v�:�o3�z�oz׊�,��cX�m̠3���B�1��@o�v���U� ��Z�J)�Ɖ'3�{v�8�7��y�Oc@|�te�V]MMI%U�`���M�`�=����m��p�?��͎F�<NN�x�PQ��J�ǎ� ��w`Z���W�M�bطX|����0#�c����K��^�d�5:�N�y�w ӆ;UUWry.Y�,�9r��/2I�<d�;���g��`c�J���2�B'�"���|�|�}��9W}�os�ٟ}�~�L21��q%M�����	���>��4���9�©�O$NH�lNw�m�������v�8��{�6�U�gЎǍ�3�?{�!B��*����o* ��Z6�15a4���28�x��.�7�\&q"��`���V����g�������4������O# }��:�QY�r, �!�3�_޷��t��:e��:U
��C>1��!���ށn�g ���?�|����t?~�_
��,X�$��$����XNA�L4��?���,HL D(��v$�$Bׂ	����\����fA#��2<ǘ$h^j���4�Ș���$2��D1LO�R�L2���b4J@@H��`9@CEDA1�I� DE~�Ƥ� �!�,I
*v�AВ��K-ŲX�H�V��J(4l�k
�"p��2�� �=9��BS��%l�!�2��4(�0ƙ1��LgXcp� RcHdb���J@��Ʒ�?�z�pS�� ��N&	�� �દ~AQ�"������RC� ��%�r""�""ߝ��*>����q��<}�<:�p�s�T��ޖ��T���@�o3�wuh��dG�tX�@	BI?f:��J�c�:��o�pII�(��J7$R�/.&ru�;]g�廜��9��<׵��n�t澎$�I��n�ށn�g ۷����p�h7q��G$�9���@c�L��J�Ǎ��
F�����>�x�7�6�p�������p_m�@�o3�j��mQ%�#!��iX�@{3��Ҡ��4�DwW������?��N�InL���v(J��@^6�X1Ҡ<�����X�u�%��=v����s�^]��l+jM�V�4Ŕ�69�n��\��6v���7��jm�h'��rI���'c�ě��;���O���c�@{3��ҭQ
&MnIzs�M}qeE�Y7{��d`�{�>o3�wm�΁v�Q̌r}�&�pfc���T�nՆ�DLDB��������cl�9$�Ȝ�@����;��V�t�fc�R��Fn�{�A���  �F���N�Y;:Zt���q�q����%�u�s�q�(�����������38:v��*��0Fw�@�Rr]v��=����;�h�Z����M�vP�gvx^6j�����ԑ\�{H����gk!�r�q�T�Ob��v2xk�vVl<���6���H˴��ˮ�a��1��
�[�qٷQΩݸ����c��q�s���(�,������pm,<���)���hr�F��ILm��A�yēs<����t���9$�@|�F ���9���I	��*n�0�O#">6�����6�{�}QY�Nx�!�3�km݀��*?B�S/wvՁ��*��2��#x��';�/��p���@�����>6�{�=���v12¨����m�h'��&���p���x����!�D`����\���ɻ[�b���۱��;Zi�>ևDb��6�eE��U�h'��&���`	�{��2���B8%M��m������	� ����Àm��΁wo3�m�n;�$r87u{�>v��Oc@i<�Sot�1�}���i9�ݽ΁Ry����� �}P��D��H]eM��F��y�jm���0n��t/��AF9�� 0m�F��T�&ќ]��`��h�4W��g_�ܿ}�ї4�8F��ɝ�����@���ۻ{���g ﰦZؤo�4�z��0I=���0M��3N�&A Ong ����@����(R$�3xۻ��T���k��<]*.������0m��7��wz�8�L�s#�GQ����m����;��`�d`��T��ή\u;'s�4k;=:�ֻ�YיuK8K��R��J��Tmny�����)�?67��ws��r��5��@I�UPY����,�73�{޼����8m����g3�<��0PB#k �o#@i<�[ot��`��0�X�'��!�3�v�{�/��p�}��9_���HH��=�㿳�z��6�)�4Bs���*�!LBm���:T�n����{��,�n�N�aκ���r�s�c�֌qg6��ܭ�z�y��E�ɇ�����# ]�# m����0����y���@����-���>o# I,�#�ȅ&E�Ud]%�g��m݀��*5)�ۥ@<�K�m�`�$M̀�Nw�[���33)P��T�N���`7�\�{�����\�U� �Y}�\�0�{�[���>��a�n'd�B���)$ �ޛl��Kuת���m�Ov�j�]�d�A�a�y,�vca뱣v6��	UnX�۶�����Ӓ���g6�;m,��^r�H�շ���w<f�2��'I�1v0��v;U���/f��t�
����O8Ķ��8n`�i�k��nB�H9U���[�3�ŗ�ؑu%F�jN`�����$�;]`�.�r��������{�����wقRC�&ئ���9՝���C=�uC���5�>�����"����&
DmdM�<�{J���w`7��∅r�iP󒱾,qƁ�Crg �n�w�[���o# K�F}��o�D7TM�TIR#����@<n��%-�@=����jb�9&��M��m�`	r��$�@m<�R�[��&�!w���ڰ�J����u`7���]���7����9�H�B��וl�uZ�n�=���':u��ms��m(	s���L�o!M����ށn�g ��-��\�x�P��szs�;�Ozt7�5�<����9�P� �*D�}��]�=�����$�@I�UPY�$�1,i�3�]���7}��g���ށn�g ��.�
Dmdc����0�=�O# i���H�����46nL���ށn�g �o3�n�y����ӭ4����ݭQŮu\���pn&�\ؘ�,χp�BV�~ϱsg8ؤo�':�y���0�d`�{�t�4IN�j
�j�0���呀.I�ڼ���-��Ӏ�Nw:�y���~��yo��!eEm2���5	t�ۥ@o۴��A��xs��xvK����r_�@m<��l����� ������$i�a ��@�o3 i�0�d`��@]�E�[n9�j�|�Z�[9�n�L�qï9Ӷ�.�	+��48�}�{�nWo�Y��9���� K�F �ot�����1�,�N�rzJ��WK�t�b�7^���?��h�=�"��ʂ�株
9��P�w`7���(�x���t��-|\�������v�6"%(Ku���(�e*��M(J#�������*��'��'��73�o�# K�F �ot���rUNɚ����#c��[�:]p��Sv2�6읭vw��/�m�a�!]������m��Ҡ���o*J@g��P���F7��	@ng �m�@�o3�.V�.Y�>�d��C��YuE��]�U��������.K# K�F �ot�1�}	&LKm��g�����g ��R����R�/^ڠ�΄�&)�(,L�t�y�[����2U��w�ʿ��H���EU\��������C�8���s��l@p��*���`���_����������@��3���������������{���~���ُ�����տ����DJ�������_�:�����������������U
D@���������G��UX���T����������'ʑ�����K?�?����_�j��_�O��Ź�@@�TaEI@��HT�	% 	�H@��!BQ"DQ"B�1%�

TJh@��)F�(B$
@�P���`%		FI�%�B �"A�BB��!	�$�I@a �!A�!dR�!�	@BY�T�adFE�P� D�d� VQ�$P��f�@��F!$!%	FF ��d$Q�!a�e�!Td@A�	F@$�D$AHF�RQ�IP�`HF�`��F�bA�Q�P �B� �aE B �`E	FA�	 Q�U%@ BA�TeAP$FA�	PV�P@�P	FAT�aD�D�e@�`BD�a!Q�P!!F��%$ B �	$a!TeY@�VP! B @!QH��@�H��@��I!@�$�	I@��	@��Q%@�%T!U�I@�	@%AYG?�l��{�d�*��������?���s�������������g�*������齿�������?��#_���"��}�=�ng����������?�����UU�a�<?�QU�����=�lT(����-�����jx�L���r���g��ߩg��UVo�����?�UU�?���������C��?��o��UW��w�@"���7����������"��\+��bS]\�,�W�-%
!Uv~,��O���x<���w<�}��UU��|�Ʒ����UWW�o�#�����0���������)�ژ'& Ol�8( ���0�7�    }         P       �  >@P
 D  �(    ���*�� ��     �T)
   �  0 �� ** �4��ͼ����^�r�[�w*�� �*Y>��&���zV�Ԧ|��2҆!� j�{��V("t!�" � �=Ň����֜���t�� �(  R (f�O�+� �=)̀)�&�Q� �L@���v ���� ,�8�DJP =4� i� 	� 3���viE@�(�@)���S�bhҔ�� bR�i���  p`P
  �  ̀ ���n�@.���ɪ����{��}Jd>�-�[ru�qwMo��z\w}j\���=��z�n��C���w��q�N�,�r��_p �M��r�ϲ�����&���|>(	P J a5T�}�žl�&�7�}�MQ��� s���һ�����Ҿ��ܥ�P nRž�:y�xӓBŕ;�;�X��˓�^��ݶg']/�O�_d�>�5����g]m�wm�� �|R�@ E  ̀ ��1�t��wo����D�ݩ}� 9�ӓ��=�/��_.��S���G�}�\�������Ϸ_m��{u��ʠ��9>�S�^������{Ү���=R���맽�a{����r�ּ  4�Sm%J�  ?�M�*R�  O���J�2 Ob�Hڢ�2�E?Б���   ����)�L�hx�B���~~��~����8Ҧ���|�(�J!_����
���QU<�DW�PT_�"���QU<D=����R*DS��.��!P ��`��<1e004�g�|��[ּ�(�0�b1`T�B�H0�0h��!$6��(F��)�H0��n.k�H0�F����&�3�Ԑ�O1޳zߞcE2 F�RA 2��ro�C@Œr_	�̖6�a	��L�YHVVV�Ȱ�!Iג G@0�p4���S�8�捡G�����Ӳ4Ța1ލ��_�jivq��2�]�IS5Ji�x�܏^s�K
E�X�����C��0�4pNJ��� � � A�
���J.��h��#�C70����5`Q�V�f�xxl!LB �lU�Gh@�������7�4��W�R�� �4�&��n�}�<�$HS3[���c\��ߞ��D�F�a����k��F���[e��y<���!H@�R5�R<)���@@*�A]�p�4�q����,X4p��!ͬiT��!�ev�3E��B�4��B�kE7ĂE(`4#Z�(
�w�o�<H�7%Ց�!�3&I�����B��)�Z�]�{�y�!�`���ES�5�E7p#H�0�A"WlJat@�H��D�t@��Wz��l��f��d�,c�^��=�g=��ozx��ssɛ9�Zw(T����˾Г��\�U:�9�w#�xl�L�-ެ����s�6|�����75��ך�4p5�K��B�,���K�����"OX����F �@#d�B�����0)�B$p�;�$�B�(A�������Dj�7�nj�%��t�m�&�k4B�f�s|7s|���6lC�CA
�ѨW$(¤X�c���b�#B+ "D4��&xރiǌ��I&i D�&���CS�Y��hi��t.��N�B�a�D<���f�7Cf���h�8��.�+�1�7�����nc�^8
�l<.c��Ј�H���DX�}<Uy��Ϥ�1��1 Q`�,)X��QQ�Hca"kz����ߛ�.xl���	���*B�B���
bB4ל�0��
h%�%����a���H���sF�KL%�y�L�㬛֎�
� �y�̺��A��nzK����rz�g�=�����d��p�YR]{�>@�4����G���w~��!�_5����6�ЂF#.Ӂ��x�.
b��j�����D�d��X���!+�U�4~4�ؑ�2{�����CF��2�Mx;�oz"]����D�����I 61i�߷iJ}��ᇡ����hĨ1�R	��@(�H&EH�AD�J���7���#g�&�Q�5$0HC	��H�\�L��.�Gd�0��CF��Y���f6���B�拏 %0.��PH��x�W;(�c�ޮ�n��� �HHF,!�[&�Ƒ�����V,��	���y�>���F�0�c$ �zĎ��9��L��R�HGx!@������RYNxa��Maw��9yi�|39gy��M^a�ˣ|*!!0����$a2���4:p�x�i
c�]ɜ9�����%�X�<��H]4É�!ta�6d>Sk����LR����8j0�04�"ŤR;H����$����M4�^/�Ʊ���
(HA( B �h$"T ���рT �&�,bBh����1�m8	��`�`P#t�8ǉ��kf�D�@�7��l2%�7���$Bp4l�9iHD�h�Ð�nH�7���m�
�F�i��ɢ�Ќ$$�e�����aI@�B�`b�A�J q7���#S5�^n��H��#�sp�ᢾ$Z@.��0Z�@�0&�p��+�ME�n�\�N}H���1��y�{ѧ��6�B�i��9��h��Kp����4��,��p5+"�
��y� �bz��`H�B$(,�VԮ�BH�����!	m������,���/7�����Pb6����ǀe�j�{�~(P��td��^T��]P	�.�����
�j�M�����5w5#���]��k^h� q��ͩ����i�x�+LАC� ��2�.����@��BI+)H1$��,CIH �"B���m�i�2`I-�s����\�$�.��I�-p
�Ѣ��Y��ْ"$��i)��I�j�8B��$jZ��C5!��˒		(cp����ˣl��0�&	�@�Z�HIc�=Pg��N�j��=��'�Ow�<�מ{���t�"M'�2B�����H�V�(AwlV����!
@�H�� ��D�$ vz0(a���&h�%�9�1�b@HŁQ���� �X5Rt��1��Wr:T� U P0@�;h���F�8$$�&�h14lÃ�nhf�	+�<i"��0Ѽ8D�I��� S3�)��k##�sz�z�F�n�\�8��S<},d+���p8�0淜��%2k|6�!�ּ��v�1�Ԏ�:]�Hh�`�"� H�0��q(�$t$�)���~��쇀�E04/)`�CJP=����с�!h��@�b@�$ 5"D�'�!���i��D�@�*H�t��B��ŖIX0��2HY�� 4HID�xR�����7&�D��xЁ=	ՊI20#BB1b� 24b�
mh��$ ]��i��%3G5�9���JH��x�Ͷ�|�4CcA�F�F��f�6�*�����@.@������IJ��P�H�d5Sp!$#
�*�+IurO%�h�.\�����4/�b���
]n�����.;6'���0���l�S+��N1��6�ar����o7ɾ@,�B����h�� �%�1����[�7&ə#�t0�9�#��¸B0$�t��2�)5�`��d���G+,Y�a!h����:cd U����2�&@���d���"aA�ă,c�7M�C�#`�5�k��0`�MoP&:�\�4!H�J�X�<M��   x.�j`�B�)s�߳{�s�1�G'�h���SdZ�
0
#ȴP��Ɖ�Sc@��]�s�#��[ֵ� h              [@      �                                  	 @                           ����s�m��m�	]6! � �a���5� dQ��m��8���  �[uY#�6���Uc���mn��vZ�p  m    ���m�ŶM*�ֵ&���	���	�U� &-઀�`6�M����Y%��p8 ��BݦZ������Ӡ[� 	eݶ  �v8�  	  6�Z��-Ǥ6�[F�N��m� �mء����-�  ti$��\z��5i2�F��I@$'M��@�UC�VC�kg)[�]v��l6�fդŠZ�nl $9��cv�ՓXL   ѭŷZ�B�V�@R��l�*��(����ᢁm۴�m�   ᬗ�r�0�`�\�o�$�h������[hhm������ m��m�ӗ�� 6����Am� 8Hp �S]�!�'+m�m�PUÇ�e�Wj����h ky�2qÃR�^��N�gZ]j�].�4P,�Y&��7[��m Tٸ	 5��a6�R��w-6JB-�hٶHr�m�]ʸ�f�	 6��6���h ��6�I&� � �I�[Am��.�i0&ײ��[�B����mB(SU�ʪ�U��S�9v��meɧ�:��d�mC�y-H$�D�����.����]�vΊm�  kZ� �۳l��� ���l �L�-��� ���   浀-����|  �` �I��  ��'  �ۥ��kS� �m�mH�	-�"�m�  �($mp�9mh�@��e�I� �J� �l�@	�v	6��@��4���i6-�LImְh��� ���Ӷ��m��Ͱ!�moQĉ$:�$I�6��,��,��	 [@��zݻ[p���m�m�M�v�d����  p�$�۶�M�%�#Ed�S �mUU]T���O(�  ���e�`��['��m&6�mHBK�v�H-��M�$ ʗd 	��[&�nN� �7����۶�$�C����X [A��٦��"M��!6�.�m$-�  :�) ��M[[�@�R�J�
��  	  � j�& @���qm�>=$�   	]7l�6�mf�6�@mzD�� �` H       ������@ �M��`I�  6ٶ�-�  �I�-�γ` h  �m�E��  88      ��    nط[�]��O���-� �-�mI@p� H       �   p��߾� �<��t��@$ ��&�$ I8v[],��p    9�X�u�  8	     �6�L�XА -� 4�������   �9���yl���HV�Cm�A,���6ͱ��m�^��� m-���I$  =6��P�ٖ\ �XI�ۑzΠp �湝��}��  �  �w��χ    �l�]6m[,   [@8����m�v٤�Iit
i9� A��1���ê�"Z�e`�Wl�(�6� �(!�t��U���:*�Zp0�i0ڥ\N�Y[�m��v�[�@8��}��|��\�v��m� 5ӵ�%	gP�"��d�v��I��j�&շ8�"A"@�uV��l8�5� p^��6����&�l�����YV&�i-�Y   8k5 �`�"Ӵ���4NSS�Mt�JR�@   �lGD�A���	�l-�>}>�v�X���&�K4ܭU<��
�nB�����y�f�p�ɇf��)�� 5UJ�U;k�p]+bB�][k���
��ԵTpY��ۂŜ����`d[B� t�]�jͰ �J�q�۸V���؄��R�*�R9ڤ��)6�ܔ m�ie �� �ʴ�آ�y�  p���6� �-r �E��y���hu+ʴ���,��ێ�Cm� �	^�N۶ V�-���x +��
�N«\ګzst`�`'@��e�6׻I��  �4��cu���N�[��l�-�  �lt  i[mm�I�J�<�
,0   �M�  5�̑�jMp�l  ��I���[� l 6ٶ�5��x` 6� �z:��6�� �e�6� [v�6��m�2���ěI�	 vհHJp���m�&���@  l� VӠ p  ��@Hm�mm��BC���8mt�	 �N�l � �l��,���AB[U[*ʡ�-P�`#i��� t�6ؐ���v  m�$� -�  �ۤ�d���axt��l �p-6 �8��0�k*RC�!tԞ�YZ���[� �NX	:L*r/I��trv�r�-\S^�5�J;^ͦ�6����`݂��U��A���wD�UUS���x�Ǝ�>UHN�m/-vh Xa����6�nYL�kf�ۤ�[E�<�Բ�~���m�۵l��������<���}�� �HŧkV�vs� � 7m�m��  l� $���8� �i�m�U��ֻ��,��6ێ� ��    ��n�-�� 6�D���p�j�F�M�*I��&���h  	I�[y��6�-�   �   �>�          8m�K([d[[l-�  q�߶��M���'8$���[x�[qm�6ݦۛy��@  Xd��}�} Ҷt�m�� �m��     	 8       V��ĀH�`l����� [@�    ��    8[@q �M�[�,�q��         n��08s��M����k����WX��*v��I-� H 6�Yg$� @�g��z�    m� 	 ��-��U�&՝���`��l�	�}���ր5��9m��� ���ݰ M�f��Ԇ� mm�r�   ;m�l  � �0    �n6��m�-�@m��@GWUK;e���F�        ��B�:�j� ��m&Ä���H�$���� -� �n�v�Y%  :M,���l��� ��M���ko`  �m��h����u�ں��A��m���nlְ�  H[@ ʾOUJ�T������Z*�@��|���uK�,�\�ʵT�HrҔU[@A�b����	���A.��v�;   �4P 6�6ƓM��:� 	 8��t�B8١˵(h{�J�k��6�E�U��m���3)��Q��+n���Z��LpPb̓i@�J�ʚ��w/�x)iʃU�6ڝ�[�m��8�kk'9��vYM ��ACU*c��j�ٶۀ���H������i�`�n�X�[m�NL  �`�� ۢ��ݰ�V.�s` m�0 	���f�*��z�H�V�RZR��dUj��n�kj@��� Y�i�`�iY����2D��   [d-� �K��:F� +�Z��
l�^��Ā ���  [xp�H�[@ ,\@  �`������h�`$�-�[d[E� $ A�o��%�  � �m 8r@ m��m Hm��6� ���� �mm� t#�> �  ���` 6�   ٶ8�Lq  	e-� m�@   h-�$v�.I($��E��	6����ll   'Nz�n��� 6�m�A��[p[%$��v���m�   �������e�fͰ ��ki�mm�  [l�d�����m m�6J�M�d�`m�m����t[h��M��r[` t�������oP趏d�k�Q��  Hm��Kmd��m�n�����G�!4�4�U�+<����� �p��0.� ��{��������{����a 	d���v�?�W�/@�v���Aڬ ����E9�!��@�"hҢ�OOpQ|��(o�NFM�L#�

�t(�x��DChb��J�o�%A4�#ϑ@�@N �� ���W�_�� {�=T�TJ?#Tg�z(<M)��y
�FԠ�[@�8���@ iU<G��@� 	"$�ABE��H1`��U�EH*��| &T�/��Q0給�PB�z��:=C���T(��
, �+�=�E�� ��F��H �$H�$�#+�>N��(�OC�`H� >����E�(��	�k� �+���Ep�D>X�l�pQC�\<D]�APLO�](�<"����AUڏ�A��*� ����6�  H        8     �	W5�$�%��4�۰�2�U\��b�]�՝����<�:
�^���0����dS�1���+m��q��x��s����R�A��l��'ct�m�At�S���e:s6�Ai���mu;:�^��weNw1�:�6��Ɬs�i������R疀��j�e�RT�UL��M�˚f�B���۝��;d ��]R��ʼ�e퀮6wb��n�,1kgc&��ţ7(��n͛Sp�{k86l�Gg�	��l픪�R�@H�Ckn�n*��j�VY^��8�v��F�	6���g-�����+UUVʻ]�Q�`-�PH��UT!��U��U;̥���^��=��\���\��u\	�f�V��wg��*��@��"�M��p�G��#r],�73���@�k\�m���1���UZִ��#�}�m�m�X�"skS�9��r+��X[��h��.8�-x��� 
�{v�n��mu��K�l��.0���j�S�j�()�*�!@cR��vu'�+n�۱��mv
U������ڠ�8l`,5<��YP����UW�u��xݧ�Pm&+P�n�nZM��|n�ImlnSXr�ۙj��24����.�T��\�FBY液@ ������Rc&���&@�ivm��$�XѣSa���K�e�SKj�7Y'*dZ��)A��v�8ڐڕ���ɂ6�7J�m9����l�:M6��>"�G �j{r���K*�<����J�=��=��h�aU	�j�A�on���U��<�ꍷCri@0�����'5�mD�ʪdp�F��%8Xy�U�V��i��@ �<�֧ecTB ��u	�0Ầ��s�)ej�b��/.��^���E�<p2�Ay�[��(�<�̓"��9����v����-3ڨƎ�k3Z55�f���4���}z��
�U4�*� 
��y�w�Ā�iY�&,��ח-���(�r©Wnk��`�y:��8���g���6m1�hQ��LS��z\=�:2ۮk�"�;.��8��)�:�^5p�<۴�m\Gm��\�`�Z�z���$�K �ȝW�x�\�*�݌��)=[�݀���vs��!;��u%Ƒ���)��*㋎��������Or��ݬ2� �� �Q�����&�s�M�����q�r�۱� �c�;m�v{r!����+�C���3�;]�}U}U\A�����a����)(���ǚ�a(J��'�,��Ձ��u`|�hRA*�#i�`w+&���7]���U���5���t�(D˫��& =nL@7�Z���=��sql���IIR4�q�Y����@s��@z䘀u��n�e^f��d�qL�=/gq��&�qn���2��w7N�!$�9TԈ���"S�Jt����y���O`���1�rb�J�f�]�3N����j�I秺�o OH���� 1H
�<H����mN��s㖀#�p�2�3h�.���D�I�[�㖀�Ot�;��z�'�%D1��ś��o�:{�I���Kͼ�)(���ǚ���+&���7]���oiҔ�u(h�P��U���om��d�N�y��t
�ص�
�`�%��ٺ�H%R�m8��d�����`qf�3j�3���Н"J�����1�rb�r��������m�H4�q�]�vc�[�Ы	
.��E	b�^z{4�1n���H��NQ)�R;�r����& =nL@t�W���)9Pm�����VM,-�vӍՁ�X��؈P�o���(\R��;�@�qW=m�nR�v<J��1Z��˱ӭg47*H((HS����H�!�:��;���x�9�� ʙ.��6�Cv��2�q�rb�r���[�����dn4(���ǒ����& =nL@zS�*��) �J���;��K�w]�ś�ru�hb�UM �@���V�֣I�IB#T�,-��& �-ΜT��Orf��[n��i,�֞��np��y��nWkn�fp��v��Q�Y5�ij�[�ճ ����q��3+�Ŏ֨��#���Հn�ȑ�1��S��vc�Vr�T���1�rb�J�f�]Yy��f^^���8��b���x����r�hH��X[��[�㖀�N*@I6�%�����R� Ԏ����`{ﾪ�vo� ͭ���9~��ܓ`� �R�a$����wwN�}���?	 l�k��>v4K�s$�ޙ�N�y��g\�;]�������rކ�;���u��ގ���n�`6n1�p�ݫ�8��|>{�`�Uj�f�;mAyB�2�̆C�K08�^�f,@^s�{�&�75����\��5��%��A�����K�9dIB�f��_P�ݖ]v��\��]a�nw]6�i��c���A�1J>������@���mŕ��Y{m��9y��O�ú��Ǩ����Bn˛��O�ΜT��b����f��
E$�R6�Vr�n���}��^���վ�3�3����'Lݢ�˫ݤ\��& �- �f�Xw6H�nP�@q������@7�Z�qR�I��,�ͳ6�h�ʽ��y%���@u�1Ż����mzR�=J�A�NEf:�\u�c��ш_m�ʼq��Q�Mr��8�R��jH��l�`un�8�u��5X��B�JB&��S��������K��$����ÓN���y��̬�X�)�U)8��R����$��r��� =q�@7�f���8أ�D��UW�-ɾV�7��b�$�JpZi{����J���3+&�����|�}�`g^j�1Wq��Q(�6�S��պ^�{=��]��]�c:�N;6sy�6n��JI�d�Ј�'�s]�ś��μ�`w+&��͒8�U 8�rG`zܘ��UvG7� �M�@z㘀�8�"S�Jt��������VM,�"���&�ݺ�ٹ'�Ͼ��9��Z8�R�m��,�d�����`qf�3�5X�I
q)��{����Ɉ�`��O`�������@p���dע$mp�{m�%Z� �+у���)*P�1�e�x՗,tfF�w4����Ɉ�`��O`��Ǯ��tf��Ĝ�Q�"q�ܚ_�dm>i`vu�XKn�R�P�L���AH���J���`n����7]��ɥ��ն��Bt��U��RS�׵`v^�X��,'�I/��g�UU\%Ni`���H�R�w���[���͛�9�m���#oގ�	ذP�jG:��㺲m�2�ǵ���8��W������sLjc8Ӷ�k*�w��͛�9�_n�����:H��D�m)����b��b�� �p�+6�ʉ�!w]����`w�4�;�M,ףz�!Ɯ�F�����였�{6l���+r�ě�(����&�s	�����`qwu�}\;�I$�I$�IWg����c:�:�+��\n���3i뙺��eҹ'X��hWe�4�ay�~�'���n��Y"�%�Y-�v'\\gTi%���Ӷ.9�E�/6ݶۖӻHv���E��; Q�	"U�\��2��l����:��P��a�t»�z�`�N |����[v��g[7g%����;�<�|k�����m���E���p]�����Z0�9��׳���>z��ލ��,�t�pF�S�ɘ�;v�۱u��Z�(H�%N�m�t����8���.��y�����q4�N��"4���������6l��G���Jq�ێ����9ך��}�U}If�<XY�v��D�!���BR;�y���a4�8���.���:Mʉ6ڎ+�����^o� ��y���V���E	ŷ=�V�&��}���&�s��+�q������I"HPID$)Ĥ"i$�!`qw7���r�ٰ@I��!�di��H�.�����W��g:�U���i`qw5��FmF�"j1L�33q��-͛������6�K�$r��R6�Vs	�����`qwu���n�IguoM:�(�Rp�K�&��Iz������}�ޤ�7�n�Iw+/Nq$�U��_f���@���w[�l���֧���
�M�b����z�Y
*�fqճ �Iu��Ē�y��I.�e��$�VM��Y�������IH�Ē�y�߫������I,[<;I%Ǜ��I%�)i#����m��v�K0��s����_Lݾ�*<"��E1@O�`AH��b�D�z\C�$�mA�����z#��_ph�n B#B�(�@�F$`�d��@"I@�a4�5���FH�! A�BH$�j�)T���jH�@d� � B		BA� @��bBD��B)!$	
K �����U"�@�#
ҲEa*#(ȃLX�P��EI!0�@���F�!�D8]�л  �6<#Rd�D��H�%F!GzގpPW�E8(�~:`� z�:S��	�*h�4��Q;]k9�{�e�̶�3��o��@�����[�+B0������߇i$���~�������v�>����s�����rfF��5g���^q$��kv�K0��s�%ՓGi$�W�?���}�=�F��`�'��{>�@�4+��n�vryp���ݣcb�Z�] �7,\6��RK�7i$��W8�]Y4v�K�7_8�Y�4�ABG��m���Y�o+����}�6�-�����y�%��[�Sm-�/.A�	����$�-�������$�[�n�If��q$��܍�F�R�&�������[o�����m��=���m�5�)�Cﾾ��i$�7��B	ʌt���I.�����ϳ7��$�^Mj�Iq�+�m����9f����I��ms���������!"�ۉ�{����7��iG��[�o+�I.��դ�����/�USo�'i!-���!N%$I���W�&9uޤ�-�������^�ϜI,y�s:���o�O�Ü����֎�̷5���v�K�}��{�m�o|ݤ���}�o�]�Ib��ߩ���}Q�"N6��F��K��o��I-�}�����g�i$���|�If�U�
8�N�m8ݤ�M���8�X�x~�6���y�%�g���]�ꪪ�}��m�zHI$�Z�z��$���۳��&���z7498�7d����e�#�Vv�qt]�c��Gj�Y��B>�;<kg�p��ɴ%u��b�vM[<#U�*���GoI]pù:^�7e���;��l����vM�X@X�:�aڔ3���:��OhY�{N��v�	�@����9�e��	��⺇�r��u�/2\��p#^N�&�5����~�߳���W���J��r[z�7DZ�7B�2�4�Χ~�ϵ�2I/"r��{�Cr8P��C�������>i$���~�ZK�5i.7�o�\�I�\m�b�Ɠn�M����|�Ic��\m%�o�\�K����v�In�Ʀ"ܕ�<�~}�T����� ~���W��Ib���K�UM�o��Ē^{KĎ�RnSi���_������I,[<;I%Ǜ��I.��դ�Y�F��RD�HB��K�&��Iq���K�&�i$��9Ē+i�T5KiR�;F�as��N)�k��aƳ̱���.{ ��G���X��K�iFgM��� �����K�&�i$��?�W����Ib���I-�F��Iē�����Ē�ɭY�z�UE�@�����6�s�%ճô�\{���U_�U$[�z�PP��*umƭ$�4���$�VM������$�^Mj�B�ĵ>SLM��D���$�^Mj�Iq���K�&��Iw�9Ē]ݹ�4�RQ�Չ%ǻ��I.��դ���ֹĒ�ɣ��\���$�I��(4*QJT���i{s��9�q�<[�c��ٞ��!�^}��lQ���%e�?����~����z�8�]Y4v�K�s_8�K^R�GB)7)��JF�$�d�o�I.��;I%׹��I.��դ�]ݣI
q)"M��q�q$��h�$�^�q*����U�!G�� m@z���}�v�|�^�����߯?��Λ5g����7ٷ��I.��դ�̙��%ՓGi$���ڍ'N&��D��K�&�i$�����RK��Iu�k�K��d�dz���hz;	��I���>�rq����:6nx��i�^g��u1b��9�Uƭ$�d�o�I.��;I%׹��I.��դ���5>SLM��N7�$�VM��m�׷��I.��դ�̙��$wuڊ(�E9CQ�;I%׹��I.��դ�̙��%ՓGi$�3M�QB��m�G8�]y5�I%�3[�K�&��^�����P����$��KI�ܦ�bR5i$�&k|�I?�����|I%׹��I.��դ��mz���n��Xñ�4��U�[`�sX;%b�Z9�8{f�rƹn���sXP	���%�g�i$��5�%דZ��Y�5�q$���O[IƜq���i$��5�%דZ��Y�5�q$��h�$�2Q�Q��I��r��|�Iu�֭$�d�o�O�m�d��I.��|�If�U�
8�'Q6�j�IfL��Ē�ɣ��]{��Ē�ɭZI-�#S�4ćDED�q�q$��h�$�^�q$��kV�K2f��$�V���$�I"JI%�خ�Ά�&^�<�I������8d.��k��[�[���H�^�c�l���m��y]�t�۵.*�뢺�� ��]��L���d��)��X��۶�9ݰnr<��7��! U;�Ź%�G����byx����z�pƃ4�.p���.:^��l��6����V�!�q�F����������i�i�_}����/_���т�m]:�e�8Põ'���[v�X�A�r\Ŵrk�ұEt��QCn�$��|�Ē�ɹwm��u�ٟ�R�皶�~�fn�m���$qE
jTm!G8�]y5�I%�3[�K�&��Iu�k�Ik�ZH�E	�M�5#V�K2f��$�VM������$�^Mj�I.�Ѥ��16�Q��Ē�ɣ��]{��Ē�ɭZ;K�n����O[�qFG$,�Ɉ_9��̴���3%f�]�ͳ�(���{v�Zrr9��	���M7�%���k��ٺAљB��~m�㘀m��@{����L�4�H�T�m�`fd֯�p�We}ꪪ_U}%@og�Vo�����}��ȍN�j�J"�m�Ձ�������`qw5��5���v��:O�(�Cne���:�33���R�J"{���）QF�J� Q�`qw5���hs� :㘀�IW�J�3K�+�Iˋב�^s�'Lu�NÞ�kk�C����҄R��ڶ�+$`�% �ljG�3��-�{\s�sID7O�16�JF�w&�ꪤ�^�;�7���ɭX�����pn(��䅁�x���{���(��(I	DD%UY&�`s�4�9��ڍ&D8�RR��@z��@6�e�=�`��b��P�ĩ�&ێ��ɭX�M,��vs]��]ǮЪR�5����/m���Y�wo��K�Ļi�7:g��Ӕ�'J"�m�Ձ�������`qw5��5���v��:O�����ŕvz��@>{2�簰f�)QF�J�R�vs]��ٖ��=��9�GW��/%&����5��ɥ�չ�¨��w�I��`ݣI�i���X�@z�&L@z��@6�e�q��@p�cn�k������m�S��N�����8��m���Z^e'M��q�@z��@6�e�U���Xs��`w]�&D8�$�����k�TB���ͩ�;��X����X>&8�6D�q��5��ɥ���K������7��N�*N��D�r�����X�������aB�m�����#QR8�m�����`qwX��S`}��,
T!%�)JZ"��#r���Dhı� $U��H�=+n
kj @�+�b�mIjI#,c)-�,��!�4�R�fr @D"��.BBC¦#ZT�C0��%�HD>C1�� ��!��a�HE�͂ŉ��FH:0c���1Hb&��H1P��c�j�& Z�$$A*���(,4<H D�B!0�B,RA# '3Sh0�#���`D"�q	 ��L@�	�4�p`d�B$�	 x�]h���0B�B);��;�>m�kX  p �`      ���    �PtE^^6��iΦj�9�"Ʀ�6��z ,��f]��b��є���D�I:wk�m��[/j2�p�E�����ٗ��Î�,t�+Eӵ��u�plC����6-5�kZGZ�V�(��t�����l���]]��9��=���l�c��	|�����&�( �����h��+��b�5jB��<��,����=��}�#t�Vk�k����,�!��/n��l&Hy0?����H�Z6��X��M���]�����YI�Uኪ]ɶ�I�U��ct�ꩥ�.�V��r�V�KU��9,�d�M�`�Y-�b��5��� ��' ^�OP]V�2�L%�u��F0sl�F�AՊj���UVʲ�aĭۢ�2c�-v��ckX�
1��z���a[���e�n.���c��6j�ƺ6+��+T�d4��ǟ�`��D۳�wu�h�ĝ�Ɲ�Y�Jհg9����r�YB^�۬��-�@���dBN����5)��@n�e�YUiK�b�q==%��ے6s=���yUU@��ٳ)���2�I��ʀ�&R��!����;WXwG\�'W[�]����i�gE��f\�"��6��ZT�76�<�f�H����PՃ��+v趘��� J�ؓ��iu���6�R��T�U	�l�.U��`��\�����d䓾�g�}n�[&��5C�Hx����V�*�G����vf�A�UjP�/=�5UU�aI�%8Z44��R���݄k|���Vҡ�e���IW�%��U"7.�.�:�b�:Ĵ�/-�T���^!�U��j-��(�j��%�C�f�q�<�fțK�ۨ�.�T�avyn��Dm�<�-4���'kכ�F��G*�VMi��U`���V���nӉ^�]*��� L�4"�G�nʥ�i��Xf*��K�;Rᙩ�kYn[4hz��wC�T� q3���@��������ww~����$ m��0Wn.��)<��6��nN�Z�z��m��ƺ��Mu�P��
�-�>q��vm��}���!�t��(e�5Yb�����bw\�j-���<�m�2$pn{]a����)	ݶ�^1l�Y6�Npۣh�h��A��z��3Od�R^���.ѱҭX�#`���9�c;b�-b��p�*�C�(���ہ�f�m+l�U�
�y��	�d��%�˩�3Pƥ]��Gs;����n���s���]�����9�51E)QJT�����y��5��ɥ�չ��7r��:)$���cR;3&���m�͞,^�;����;�F�Ȝi���X�M,��v{ꪤ��|�ݞj�Օ��6ۉ��#��V������ɭX�M,c�t�&D8�N;�����=�hs� :㘀7�+M���X�J=uΚ7o\v݆:N������yN���n{p]`�Uk�y����6�e�=�`��b��b?���Y���M�9y��
�|�~oq���<���m9�a! ��!?E(�P4ț�b}���6��bX�'s�{�ND�,K��r�9�&TȖ'�~����]R㚓SVff�ӑ,K��?w�m9ı,O3߻�ND��"}��ܻND�,K�~�fӑ,Kľ}�e֮���K�WE.�Y��Kı<�~�m9ı,O��}˴�Kı<���m9İ?"̉��w�m9ı,K��K�kXB�sF�3&]k6��bX�'�}���r%�bX�{��6��bX�'�߻�ND�,K����ӑ,Kľ}�uN��g�����M=qk�w�у�#�q���ѣ�h��i-Ƶn�{Z�:g�M�r%�bX�{��6��bX�'�߻�ND�,K�������}���%��w��9ı,O�����d�L�̚�Lֵ6��bX�'�߻�ND�,K����ӑ,K���ܻND�,JB�;��|B�T¢��x�'���+��f���fӑ,K��>���r%�bX�}���iȖ5��D��H���w���ND�,K���smp���#�G՞���$p���%%�\�bXX�}���iȖ%�by����r%�bX���m9İ"����}V}T}^�#��F�SJTM�rlI�9�i7�}#�g�fӱ,K��߻ͧ"X�%������r%��ow�����Q��\�C��l\Xn������\&�
��T(��"%$"Wv�ڑ��\sRjh˚�ND�,K���ͧ"X�%��w�ND�,Kߏ�ٴ�Kı<���m9ı,K��v]j���d�5tR�k6��bX�'���m9ı,O~>�fӑ,K��߷ٴ�Kı<ϻ��r%�bX���������j�I��ӑ,K�����m9ı,O=�}�ND���DȞ���r%�bX�{�y��Kı/��;$)�8�%JB��R>�}H���~-9ı,O3��6��bX�'���m9İ=SDTW,K��;6���{��7����^�g9������ı,O3��6��bX�'���ͧ"X�%������r%�bX�{��6��bX�%���wV�I�Vj��th���1M��Xˮp9��i�E��\���zmsٵ�E�Fa	g��{��7��������ND�,Kߏ�ٴ�Kı<���l>	�L�bX����r%�bX���A2G:pm�����#�Gԏ�ߏ�ٴ�?ș������r%�bX��~ͧ"X�%��{��ӑ,K�ｳ�8Lֳn�\�3SiȖ%�b{����r%�bX�g��m9ı,O3߻�ND�,Kߍ}۴�Kı=����j٨\sRkVe�M�"X�%��}��ӑ,K��=�siȖ%�b{�v��bX�'���ͧ"#�Gԏ�n�"�(1J$�������ı,O3��6��bX�#���v��bX�'���ͧ"X�%��}��ӑ,K��P"�O�����  ��s��m�ڻ�n��ǳ�t��L���]c�toc��8n�(&�5c;��'t[�^���M�R�%;�[R��k����skOb�.Ûq��5I0W; ��hnvn�k���RW/+i��pmֺv"��v�n;@bs  ���(�#�lj���c�5��$�����1�ۗ��Ex-�C�qF7/\�u�vC��繃vh�;�w��j��)�qڲ��R뫥��8��k�p�=���Y�YD�v�_Cũ��R.F�S�%�bw���&ӑ,K��߷ٴ�Kı<ϻ��r%�bX�g��m9ı,K�zN�j5sRfL��Z�ND�,K�~�fӐ�
���,O��]�"X�%��}��m9ı,O=;�ͧ"X�%����v]Yfjf��Zњ֦ӑ,K���}۴�Kı<�{��r%��ș��fӑ,K��߷ٴ�Kı>�Rw���&��\�us5�]�"X�%��{��ӑ,K��ӻ��r%�bX����6��bX�'���ݧ"X�%��u>�$pC�܎��R>�}H�����iȖ%�b{����r%�bX����v��bX�'��{�ND�,K�wy3�m҃s������<��#���7�������n9�m-φ:N�Cviz�.�358�D�,K﻿�iȖ%�b{���r%�bX�g��l=Y�L�bX����6��bX�'��ܼ֭��d3Rjh˚�ND�,K�u�nӐ����MD�5�����Kı<���6��bX�'���ͧ"ʙ������∋8�Vȱ������ŉ�}��m9ı,O=;�ͧ"X�%��o�iȖ%�by�w���Kı/{�{��!���\ɗ5�ND�,Kߏ�ٴ�Kı=���m9ı,O3��6��bX�D�_~��ND�,K���~��2j�2e����r%�bX����6��bX��@����ٴ�%�bX�����ND�,Kߏ�ٴ�Kı=:jó%�JkRjM.��5���[F�Yfw�Щʮ�{r���8���b7�����w���oq�����ͧ"X�%��{�siȖ%�b{���6��bX�'���ͧ"X�%���m��XtfUd�~{�7���{������Ӑ��$r&D�>����ND�,K߻��iȖ%�by�w���J}H���g���$pC�)�㿫�ԢX�'�o�iȖ%�by����r%�G�E��j'����ND�,K���ͧ"X�%�߻gnp���4j���f�ӑ,K��߷ٴ�Kı<ϻ��r%�bX�g�w6��bX�@�����Kı>����Z�jd�I�Y�56��bX�'��{�ND�,K����ӑ,K�����m9ı,O=�}�ND�,Kߏ���Re��ɃZ�$��������w#�GnLY�t���.Iw'ju*�i]�Y�ND�,K����ӑ,K�����m9ı,O=�}�ND�,K���ͧ"X�%�{ߋ�]a��ֲ�L��m9ı,O�>�fӑ,K��߷ٴ�Kı<����r%�bX�g��m9ı,K�zN�j5pљ2�]jm9ı,O}�}�ND�,K���ͧ"X�%��{��ӑ,K�����m9ı,N�s����ոkZ3Z��r%�g�@�~���r%�bX��߿fӑ,K�����m9İ<���Puȝ��|�ND�)�#����B	������R>���=�siȖ%�b}���6��bX�'���ͧ"X�%��w��ӑ,K�� �k�����VL��L��]M\5�����v�ԮC;�q�ϛs1�6�a���]m�Veɭf��kFfkY��%�bX����M�"X�%��o�iȖ%�by�����Kı<�{��r%�bX�Ͼ���5��F]�a����Kı=���m9ı,O3�w6��bX�'��{�ND�,K�O�ٴ�Kı<�������i���R>�}H����ͧ"X�%��{��ӑ,K�����m9ı,O}�}�ND�,K��ߦ�"�.�ة�����{��7�����ӑ,K�����m9ı,O}�}�ND�,K���ͧ"X�%�{߬�XC-�5ur̹��r%�bX�z}�ͧ"X�%��o�iȖ%�by�����Kı<�{��r%�bX����������q m��gT\H'j�~W]�Cb�c�%�b2�/V3��ۣˣO0�B;N7/9.X�n^zWNYk���#v�a�te�\>�� �ggk�Y>ɴ؄�{i��d�{t7��u�ӫ�C���m	Ys���Z�e�r燞+�z�y�:N��#��+���-�YM��w�>wC�+Ս�����N5���Ɛ����7�w�y��6��M�g�a�ι�S���v �o,]�5���Mڻ ��9wD'h����iu���Kı<���M�"X�%��{��ӑ,K��=�siȖ%�b{���6��bX�'sӹ�uasR��5��jm9ı,O3��6��bX�'��{�ND�,K�O�ٴ�K�����K��
HRB�|�8M��33Y��f�iȖ%�by�����Kı=��}�ND�,K�~�fӑ,K��=�siȖ%�b{�O����ֵ��5�35��r%�bX��}�ͧ"X�%��o�iȖ%�by�����Kı<�{��r%�bX������.j��ֳ�M�"X�%��o�iȖ%�by�����Kı<�{��r%�bX��}�ͧ"X�%����s�j;O6�Q���Mun��np��z��܏klFtX���u�ml�����N�m��ۉ�Kı=Ͽ~ͧ"X�%��{��ӑ,K�����m9ı,O}�}�=ߛ�oq�����~���8�#a��ND�,K���ͧ!��FA��.�;�bX�l��M�"X�%������Kı<�{��r%�bX�����5�2[�W.Y�5�ND�,K�O�ٴ�Kı=���m9ı,O3�w6��bX�'��{�ND�,K�ޓ�Z�M\4fL��Z�ND�,K�~�fӑ,K��=�siȖ%�by����r%�bX��}����7���{�������#sF�깫m9ı,O3��6��bX�'��{�ND�,K�O�ٴ�Kı=���m9ı,O���u3Y%���Lrf�qfm]2�ݓ�1y�ms�l"��kQ��Qq�6kYzJM������7���{����ͧ"X�%�����r%�bX����6�g�2%�b{�~��ND�,C{��}�,��\g�����{��7������m9ı,O}�}�ND�,K���ͧ"X�%��{�siȖ%������p���u/-�{�7���%��o�iȖ%�by�����K��*���G��H�#$b�ؠ������h��-,v#�	!�FR $Bb�"�+��-���(}�#�0`EA��a�
��,H�
�A� �Hu�
�F�	 AX� �\] @!��H�\�=Uu�(�}6OAAb��iQ]��E"���@��1T��@~En�]6z�;"o>繴�Kı=��}�ND�,K���$6�c�"p���ԏ�R���ͧ"X�%��{�siȖ%�b{���6��bX�'���ͧ"X�%������51qt\?=ߛ�oq��'���ͧ"X�%������r%�bX�{��6��bX�'��{�ND�,x���}���}��8]�y-�=�Z�u�n� &���r�5��<s��-®��x�{s��W,�.��ND�,K�O�ٴ�Kı<���m9ı,O3�w6��bX�'���ͧ"X�%�|�I٭C5n5�e�֦ӑ,K��߷ٴ�Kı<����r%�bX�g�w6��bX�'ޟo�iȖ%�bw>;��Vf��un�kFkZ�ND�,K���ͧ"X�%��{�siȖ%�b}���6��bX�'���ͧ"X�%��ړ��jf�f�]]M]k6��bX�'���ͧ"X�%������r%�bX�{��6��bX"x�Ow���ND�,K܆�B
IHu%6�w�p���#�B}�۽�ND�,K�~�fӑ,K��;��ӑ,K��=����KĻ��{���ml/\]����s���a�������M��И�u����*t�OAu������Kı<���m9ı,O3��m9ı,O3߻�ND�,KϾ�v�9ı,O}��9��nS0�I�Y�56��bX�'���6��bX�'���ͧ"X�%���o;v��bX�'���ͧ"X�%�|����j��d�&�K�k6��bX�'���ͧ"X�%���o;v��bX�'���ͧ"X�%��{��ӑ,KĽ��I���2�Y��K��"w��~�ND�,K߻��iȖ%�by�����Kı<�~�m9ı,K�zN�j�pѬ&�5v��bX�'���ͧ"X�%������ٴ�%�bX�����ND�,K߾�v�9ı,L@?���kj��V���+��[��Rݵ��ml��OYcׯH���м�9��bvL�n-�u����f펲����G�v{v�ۃb�)v
��M��t:M��Z٭ٳ� {��l��S�a��ϾcuŃt���X1H[��ZB�x�K���\c�M��+ɪ�,/v��r0mƢ����n��a��K����V�Ǝz��[[���Y�/���{��|���@�����v����vݰɇ^�����8��Lq���kC�b3JAu]�֧��Kı>���6��bX�'���ͧ"X�%���o;v��bX�'so��\>�}H���f�7�cpN�iG���fӑ,K��=����Kı>�_gsiȖ%�by����r%�bX�g��m9ı,O{���ֵ��5�33Y��Kı>�_gsiȖ%�by����r%�bX�g��m9ı,O3߻�ND�,K��rw5�sWXj��˙��r%�bX�{��6��bX�'��{�ND�,K����ӑ,K���}�ͧ"X�%��vg55m�\��3V��M�"X�%��{��ӑ,K��=����Kı>>�ݻND�,K�~�fӑ,K��߻��0�2�v$[6�ċ�6�����C�y�uss��ɺ��zw�Rjb,��]������,K����ӑ,K���_v�9ı,O=�}�^D�,K��{�ND�,K�����-ѫ..��ND�,K��}۴�(� ꂲ(+�6Mı,N���6��bX�'�����r%�bX�g�w6��bX�%��'fh�[��a1�5��Kı<���m9ı,O3��m9ı,O3߻�ND�,K��ͧ"X�%�����q� �\M�{�7���n��X�w��n	 �_~�lI�==��&��'by����r%�bX��D���fj]�K���f�iȖ%�by�����Kı>>���r%�bX����6��bX�'���6��bX�%�����ܝqhn5����N���q[��Eֻ[N�y���J�l�-�n��J�v�������bX�'N��6��bX�'���ͧ"X�%��w�ͧ"X�%��{��ӛ�oq���}�]��1=�r��w�Kı=���m9ı,O3��m9ı,O3��6��bX�'��w�Noq�����������#0#o��D�,K��{�ND�,K���ͧ"X�� �P�x;TCg"n'ƾ�fӑ,K����iȖ!���Ͽ�SSgj���~oq�X�'��{�ND�,K��ٴ�Kı=���m9ı,O3��m9ı,K��^��d�F��L���r%�bX�}�ͧ"X�%��o�iȖ%�by��siȖ%�by�����C{��7��~���:y;y�)#=t�^�;nG��1���"�7�;v�n�A�p�ڻZ�jh�F��	u���Kı=���m9ı,O3��m9ı,O3��6��bX�'�o�iȖ%�bw=;��Vf��un�kFkZ�ND�,K���ͧ"X�%��{��ӑ,K�����m9ı,O}�}�ND�,K�O����t�M������7���{������r%�bX��}�ͧ"X�%��o�iȖ%�by�w���Kı=���Q=Tnz�Z~{�7������w���y�m9ı,O���M�"X�%��w��ӑ,K��b��KϷ���{��7����뾵�'����SiȖ%�b{����r%�bX�g~�m9ı,O3��6��bX�'ޟo�iȖ%�b{�w�55��.Ytd��s;�aal�]�rp��:۪6{�v��1-Z
�րN�0#o����7���x�;�siȖ%�by�����Kı>��}�ND�,K�~�fӑ,K�q����b,��^�O�w���oq����ͧ"X�%������r%�bX����6��bX�'�߻�ND�,K���Z�%��՗	�5�ND�,K�O�ٴ�Kı=���m9ı,O3�w6��bX�'��{�ND�,K�ޓ�Z���4k�.�6��bX�'���ͧ"X�%��{��ӑ,K��=�siȖ%�b{���6��b]�7�����FiH.����w���bX�g��m9ı,O3��6��bX�'��o�iȖ%�b{����r%�Y�����继������?���� T�{]�P�<��u�M=���e��r9͓6���9��n��F�U�aP�GQ��x�bcf���K�Z�����UĲ�-tZ��{F�����퓱��[���Cv�<l��ңq�\.���1����]��@
�Ʉ6�q�z%�B���>	y�^BX����/bv����F��Y퀺)���ǰ��W
un�c*�����=��|�O�Pg�Jۛ���9��JgG�u�9Ӧ�X۶]�]�^ y���i�l�U���6j~����7��b~����Kı<��}�ND�,K�~�fӑ,K��=����K��{��m�}�'���W*��w��ŉby���6���RDȖ'�w�ӑ,K��>���r%�bX�g�w6����oq��_�]��1=Լ����bX�'���ͧ"X�%��{�siȖ%�by����r%�bX�z}����}H���#�����&�MDH�NM�"X�-��{�siȖ%�by����r%�bX�z}�ͧ"X�	by����r%�bX��{l�殮�K�kL��ͧ"X�%��{�siȖ%�by���6��bX�'���ͧ"X�%��{�siȖ%�b~C��?kZ��%3Z;v��I�WK�ݏ�le�A�8{I]��YT8.���������ll] ���7�ı=���M�"X�%��o�iȖ%�by����"X�%��{�si��Gԏ�R�m$�GMQJB�9ı,O=�}�NC�5�I?�]<�Ȗ'3���ND�,K����iȖ%�by���6���%�bw>>�t����f�=ߛ�oq�����ͧ"X�%��{�siȖ%�by���6��bX�'���ͧ"X�%������e`�b?=ߛ�oq���y����r%�bX�z}�ͧ"X�%��o�iȖ%��'���ͧ"X�!�߿�~o�D�Q���Y�����{�������m9ı,? �}���6�D�,K����iȖ%�by����r{��7����߿�᭺���tA�{Y,��4j�9ǞM�C$�[)�ݩ��F�I������;�Xbz�ym�������ow�߷ٴ�Kı<�~�m9ı,O3߻�ND�,K�O�ٴ�Kı37��"I�騉i���R>�}H��=����DBı,K�w[ND�,K�O�ٴ�Kı<���m9@�,K��m������]Z%��m9ı,O3߻�ND�,K�O�ٴ�KDW�T�h����o���r%�bX�g�w6��bX�%�~��Z�%��շ˭kiȖ%�#by���6��bX�'���ͧ"X�%��{�siȖ%��A�3߻�[ND�,K����5��4\2����r%�bX�{��6��bX���{�ND�,K����ӑ,K�����m9ı,ON����0���D˖�Δ;Qv�л���g&�ygq�z��7,qs������O� ��&.�o����7���{����6��bX�%���[ND�,Kٴ�Kı=���m9ı,O�~���i`�i?=ߛ�oq���|���Ӑ��1Dr&D�;ӻ�6��bX�'�w�ӑ,K��;��ӛ�oq���~����څ�s�����Ȗ%�b}���6��bX�'���ͧ"X��%��w�ͧ"X�%�|��o����7���{����}kOAu/9���K�,O}�}�ND�,K��{�ND�,K��{��"X��k�
m�:<ș�~�m9�Gԏ�s|>B$�m5PM8_���Gŉby��siȖ%�b*�{�m9ı,O�>�fӑ,K��߷ٴ���oq�������h��;D`�nb�[����W8vn3�y�GnLY������f#b�z�8���J$�G�\>�}H���.罭�"X�%������r%�bX����6"��bX�'��{�ND�,K��Yۭd��tj[�˚�ӑ,K�����m9�r&D�>���6��bX�'��߳iȖ%�b_=�u��O�M}L���/~�G�A�G:h!W�,K﻿�iȖ%�by�w���KRı/����r%�bX�}>�g�w���oq��_�}~�SX�M6��bY� dOu�߳iȖ%�b_~��[ND�,K����r%�b"؞���6��bX�'~ԝ��f�Ѭֲ��k6��bX�%���[ND�,K����r%�bX����6��bX�'��{�ND�,K���B`�\E> �͘�H) Ȣl}$	4K,�%$%#cH�
�ZQw�h��"A�5�3[�R�$	!$ @|&q� t�������CUK�@�`�BsF�R�$��	���Y���#!1��x̷Jm��P�A$�)�X����r<��F�g�`�G<��	�� ��"ʌ�4)!b�T
2�DВBlSLc��1x:[�����}����;���l   l      6�    �j	�e�T���9�c�z���vX`�����ݸ���\�G
��6H+`D݈ػ<�ҵf�ms���[-t)��f��ې�F�W���P�j6�m[���3�y�,�k�#�Lfu������F9W�ېh�dɕ$��v�
���z�.��8�/-�Z�[IӁ1��6��:)�/B�EOGPb�䗶�"��������QK`���ku�3��R�YL�$��jNm��׎��9�,8Xmj��v�e$`+���_]��J�L�UV�x��6Q]�m��2-[)-U���U�� �Z��
��	.��w>���Bh8���tU9��m6U���c7+c]�:
�y#j���Ҷͫl�9֬4��:�\l���Mk����:�<��nQ�t����g��[��f�bM�t�+�X��q�	��@�3��u��]����p�[m� �x8���۩�]�n�x�y��2�6�u�����)��.ٔ�V�u�sל��n��vʙ����D�����'��[k�ʩ�*lV�^�Q��#�:��R�(��ɴC˯I���10/`����P]�Q�)�����4#[Ug�|� �M��*����*e3]�b��g"v�mPn�S� 8��ؓ�s��7$�����p�b@eX
��-�m�E�Zt�*�UUL�N�.�>��8v9��T�v�0�IĪ�+V�d�Q[J��Q�l��!NC�MUUrm*1Y ���[^2���icv�%���@Ȩon��ڥk��f�+lL�:��<�mڻ:�v�zx�<ƥuD�Ǟ��Y+k���Tr�3ڸؔ�mR$T��*�2df��r�T��y倭��nwF�]��:C���$�+�P���D���s9�v�v�)V��ûN&���%c(*[����]
�ְ[Ś#�VĻe��\��k2�fR�� �"#@�PC�ڨiD/�:A|M��?^�ww����k_� m����F�+"�,v�{3�F�h�rn�������]g�,�g��n�x7f܋9壃0\1!F���EŶ��dmm=]��j�9�R��]��d�P�p:9ݎr8�V�Ŏ+��y�=�����s�[v�l�$���-gnN^��ń���[S�[k�x����:H�)⵶힥χ���gJLk<
tl�h�۳t�$��Zɭ��n�f!�ӝ��	=�����y������t��t2�t3�������m�T��a�3Z���%�by���6��bX�'���ͧ"X�%��}����,K��=�siȖ%�bw=�N�\��4[�Z�356��bX�'���ͧ"X�%��}��ӑ,Kľ{��iȖ%�b}��}�NAVı,O=��9� ���"������{��7��������bX�%���[ND�,Kߧ���r%�bX����6��bX�%���2�ST��Mh�u��r%�b�b_=�u��Kı>�}�ͧ"X�%��o�iȖ%�'���6��bX�<}��o�;c�����{��7������m9ı,O=�}�ND�,K��{�ND�,K����ӑ,K�W諾_���?R�QR��10C%9P�u��[������\��bٻ^�oG2���l��t�:}I&�R\2�.�6�D�,K߻��iȖ%�by��siȖ%�b_=���r%�bX��>�fӑ,K��|w;$����|�~oq�����~���NC�؉�biD�K���[ND�,K�g���r%�bX�{��6���2�D�?wD��Vff�ѭkY��n��ND�,K��kiȖ%�b{��}�ND�K��߷ٴ�Kı<�����Kı>����֭ɭkVkE��kiȖ%����>��?M�"X�%������Kı<�����Kű/���m9ı,N�d�h��\�E�5��3SiȖ%�by����r%�bX�g{��r%�bX��~�bX�'�O�ٴ�Kı>�߳�G`Bz#,k�t;m�@�=�+�ۀ����ГvMwZ�\�:ȭ�x�Kı<�����KĲ����$������a�����ʓ?B*PJ�f�� �9�c� =�`���1 n�-$`!)�C�Ԓ��4�9��,�
�P�!(��
��mՀf7� ��H�Q������r/�_�}���9�`� �d7dRt�'!`qn�w6X�&�;�Kk�8�&����q��Qծ�e�wk�+�8���l"��\�@F��8�{4Cn%*GPJG`�l�;�M,w&��3`l�7RH�u%&����s� =rL@�5}_�~���,�yʉ��JJT�����l�`z䘏��~�9ϵ �7���v�m��T�n� �se��2lܝ7M���<�;����Rg�
�8�w6X�&�;�K�w]��ݥ�t�Q5ڹ-�7`�Q�G�Oʙ��#���z�r86��p���꫎�Y#	O�&��4�] =�`���1 {���Qܺ8	�@'*��ri~�H�������pͺ�2��N% �M�r�۫ ���f�IL�ڰ;��X�8)R8ڂR; �se��Y�V;�KW�������@��&I"++v�37Pӊ��@z䘀=�krL_���BEV��|5� �:���k�in��H��&�'G�G&�X��v$:��K�qmZ4mm�m���4&:�C<�i�Wr7�z�g�����+�^AB�3�Ɲ����v��u��L����-��uE$u�;<v�^�4m�vx'��.�6#C�.�<��6���v��hv���hxi�p�:E��x�vN������8CV��ݶ1u�I�2�f��2�/Q@? o}�����㋵a:�X:�Η�����8��;F�s&��l�t�v󵸝L�t0�p]M*��n��XKn�����%	v�ޯ~��7}���#ciG4ۅ�ź���{��ŎՁ�s��P����l��B(:	(q�`uf����ug~�.��Ż��3�V2��6���D(�ŏ�`w_4�>��XOqՀwv�$j�'�j�NU���������y���;2�n���a*2����[Wm�n]vݱ����l/F;n�����ٜnB@���F�"�*m�r�����̬ۯqsg�����i8'QH҂R;����W�W���u`w�4�8�uߩ#wҏH�qIR��ۍ%O� =�`���1��1��u⎥%*F��V;�K�7]����`w+6���sGr$6�Ҏ*k34@zܘ���ϳ�9S�Hs� ߟ�������8%[n�ɨm����]��z���b�z�ٺ��kնZyT�բ�b��{�����N*@{���r; ��U�*>H��6�vr�n���	L���,�{V��u{	B�*��j?5A��5E'*����XY���$�E��B��Q}3��`wv�����ӉH�Jn���8�u�]�vqc�a興S�w�����ɩ��4�<ܻ��w�st������Vc�P���ԥ�"k�*��>S�u�<V1��]c�];)�%ԥ��h�s�d�T�uDT�)�����]X�M,,�� ���=�%��:����%X�q�Ә���{���c��!B�U���D���Q�M��`b��;����N*@w=� �K��hiz]�n���V�����;V{�e���]���;yn��$)�B�g�qR���@yӊ�7ǀ�}�_I��������t�v��\��.��I�8�I�y6^�v���x�юg�*XƯlujN�e2��ͤs� =m�@z�L���:T�R ��^���*�`�,,�v[���ڰ;��/СD$�L�=�jS�tIPQ�`ug���f�Yﾪ��������y��(�rT�*Jy����V�O�H�� =nL@z�L@n�[u"N(�RR�n��`w�4�=�{���ݫ��ڰ<�A�7��pm��Yi$�"M��u���/q�{Z��]�ې�^y5��Eӧ@��6����� �Pm�����Ͱu�*I���z���s�w$Kg;���i�G2򮊌���)�e� �]�jL�͹6K�:��h � y�u/��lڅɩ]�Yv��pvb��m�Tr��3]n9�J�T�����n��pn�S�-����jɗ�s;Ѯ�+TX��[q�>yY9:��4[���ц��1�ciG6ۇ@���8����f�~� ����3�I��T����"��V����	DL�����,,�w� �j�QHJ}�JG`n��s� =nL@z�L@Ԇ�U���m�����u`qf�8�u�z���X��:�m8��Tcr�[��& T���*\��`N�6�m�vn�N��Ok��뵅:��n�vrr�(@��zh�o�������X��<�W�v^�X�;Vs�(QHvw�v��G�i�RDT�)��3�7J�Q_�t��vo����<�w��,�w�#�Խu"N(�%*D�%X�ڰ>�n��%�{/v�Ƕ��4w"��J8����7]�ś���3���J�n��֦��s�H���T�`}8�X�	�ޟ��Ձś���ɲI�Q�����u��{;�p kc�u�����hWɵ������. w
)	O���R>�l�`w2i`qf�8�u�en�:_D�6���p�;��_�DD/D(��2wޫ'}�`f4�2����"�T�Ɯ������q���P�S1
JB���T"SL��$B(bcCbI�q� PbA$$�3F$�#BP���`A��̗8[��  D�$`Q������H(���%� B��@��0	T� `�Y��@�	�z��HHx��==]#�0TQ�U8�/�|
> �����97���}��,�3tM7aCt����_}_R�}�		�o`���1$�&�\��h�%6�vpɥ���������:��;�7]���f�9��N*���'�ٗ[���V�wMg42������>ۧ�B�Ŷ�Q)*D�Q�JS��Àf��`}-��>�n��!%�1�K1�W�JM����M�����`qf�;�M,�M/�UUU$�=F�9IJ/sq�>�ǰ@s{�I���BR���JGaﾯ��m��1�i`}-��IDDZ��� P�~@ED�0*���ڌJ�s;��`�n�4���R7�@z䘀��1�{ߪ��W���o�n~���Z;[p��S�����y��KE� rpٸ7O:�s���������O� �B*�cR�ߝ�ś���4�;�4�:���4�I�q�R;���JS&1�K��۫�(��4J$�ێ��4�;�4��W�}Iu{�v������M$I�JJS��������`u{�v�ݖ���Y�ߋ3|;�t鴣 �n\�����=��� ?���=����p  ev�,-Jr��Փ[��bãI������5�8��3r��t�,4�e�n���
�D��kjS&�S����$����6�,�^rb�.t��n��<��.g�ͨƵt��k���	2gc�nv�̀ 6�۪�؄�.�ۗq^aJ�ݥ��6.Tg����w�eSs����Ks=���g�,�RL��Y��%��B&�]��Q���L����/np��k���۝��bm�F���%�j.�����v>|ß��v���w}��j�{7�@z㘀;���S��4Ф�0ɥ���2��^:��/Д(�DB����^�#��NhN�HX�OŁŹ��9����4�5v��L��41�p��JD���X�����2��3�XTf�n$�8��'�ř����u�����,��'>.�׵�CۮQקI�m�R�{����sn�`��KR��X�I=Pk�p���~1�o`���1�nbs��n��P�N&'��K�U_}�_z��$;S�@O��=��኷n��mF��p�8�5�Y������R]�g���ŀw�&=�D�'�IVӘ����,�8��P����X{i3Т���)�$�9�M,(�w��vu�XNc��9#S�Yñ�uXru���tr��W":���ф�a.�M�����m��V�����fXK�VӘ�Т#���Kg֑��$QSC��8�5�Y���d���d����RF*7�MĘIyWy����@>��AG�� =q�@n�dj:�$J$�܎��_Rܩ�VuŹ�����`oq)��8��(���9�5X[��,�vv�j�?U}_W��u�� &�*��Ӝ�z�C��ˍ��M��ױ�����3!�ɮ���|��p�7N�Q��qt_���Y���<�`sj��Dǵ$����ř��_$nS�+�������`�C[
)�JR�t������V1�<�W������en�:_D�6�h��9�5X[��,�vOW�X��X	�P=D0Uk��Y~VWk_��e(��qX�� =m�@>�r�x���L��+�<�����tK�lp���rXw\
o��{r�לvE��P/?6߇�������V1��A���=�J=#Qԑ"Q%&�vv�j�9�5X[��,�w�|���Jm&7C��$������
�� 'V9h7-n�Rm�bqX[��,�v0y���<�`i�Ɯ��
H�[sf9h<r��� W���w{�~�w��q m�ݐ���T�O%˝��0�]�CYγ:��I�b��Menzg
 !���R)���]�NYuG���<�і���b0�ð��Ǝ�с����s�V}��=��y�nu��h����i��u Y��J��$���=��<OT�#�pvc����D�'�>,5Y�v�w��fnb�z���9]���v����G	�6	�z�{P�}���{�?8�7�tJv�KrZ��I�tz���e5%v=`99;u��S��Ld�n�MqSlIǠg��+��U�Ź�����`��$t��4�t��9�5X�� =m�@y��%�L���n���qX[��,�v~����+�����3i4�mҒ	�i�a��'؀�d��x�=q�@I6���I%E(nG`s��fM,-�vn����\%	��*2&�T&�;���h��c�ܛk�q}�vӕľt�	��o�B�r�Jq1��n���7]��j�;���PCiFF�����Uvu���c����۔�������)#�8�u���?RY�����`���%)I������|���ՁŹ�����`��$t��4�t��;��V��7]��j�潄�$����;W��Iں��VM�
���`z�&�x� �:n��$QSCr�-�v[�f9hr*@u�ܫ���̫���+/7nL@y��9ȩ幮���F�҄�R�$�v0y�ܓ�~�f��M��z�
�XQ��H$E��h� r�S	aB!)P�S�P���>��`d��X�34�'r��N&'Գ}�U����:�5��&�35\jhmF8�s���^:�7�!�w��3M��{u`s���:%5D`�MԍB�	M�Cl�v��v�m؜o>�wl�oN��A�L��%
H���v0ɥ��ݺ��\A����kУ�JRm$�9�� <�T���1�������_|n�/��M$�!HX��ՁŹ���UIb�y���+^�����1��`}/X�n���sa�Jyr!!��P? ����'����r�k3���+/7rL@y��{�f� ��z�D�j��TQH"D?䫪��[��a]h��vAݥ��Nv�pQ��v�'�%8�ӏ�wG�Vf�Ձ�����︃��`{<��"N(�%R�n�� �9h_I�\���_~��vn�Ơ1�j1�؜V�{�����`op�X�5X7Ri�5MJ��'��X~BP����Xe=�;X���UR����g�kС��*mI��c��}�Z���I���~��@=a�~H)�SJ���J� � (BHK�Ѡ�� �1!P� A��D�E2�*Q�,)��a0�A��T��b�4P�-"@���Jb��*a($�Q�i�";���#DR	�aHHP6�X�P�:{�wN�����#��6�  H        9��    ���w6�[����:T�������ɵ���eی�v'�u��J���%�&������]"{4v�E e�b���U��;'j��^Z9����Q��t;n�d��FB�ͥJ�K����l�F���ض�6���c�ʗmh֍=�J� 4�)�l1���qWN:�>j;k`�ry�Jn�.T90]&hw1�AEA%:.�T��cv�N������ZsX�@�;`7c�6$4�͸nFj���
'6wKZ��	U����<p�'M���FK)�-4��$l	�E�tI�� �OZ�ʻc̵]!6�d��c�в[�K��.��$,�n��wf��y��U\�X%���ܹ��[��z��6b\k3��<���g:��i��ȇI���<��[ϳ�MV��ͳ\E"-]��F���s�f�V\�	[kЌ�s�R�]�^gqB��ڦ�n�$(8`-��\����6�(�/06�R9���h]�	���wd ��&۴]��j�����	�V�ڷ5�j�[]:�*��ܚ���Pq�zۑ8-�i�Ks�=tEղ�H9�'1u��Q�v�����U�ȭ�p�
#��e
U]ס��=��M�gc'�L�S� 8^�[l���ڧJi{D�d�M��[\��m���� ]:��HʵUVwBC�l�(l�b�U���jb��Y�yv�����A���٧�]$ͣ0�V�ƳM�۔��ۆ�r��ԡ/+p5lx�:�Iv+�9��d�[�[l��;kr��]sՖ�65W�a�N�8ŋrN�����A��G;��Uc��f�-��GoNQ�U��֪���^���G֍���]5�a:Y%� *ݪ�U�;	mv�R��wn<��70��<�ʬ�YV݉���8A��M��ֺ��P��氶��P�Lն�M�p�"�� @V��f��1���Ѡ����OS�Q�A9�h�x"����~�ֵ֤�kZҭU96+��g�N莧;��j���]g��]�>zN[$�ۛ:�Z$�t��9�Ű�����Y�8M��nǭ�&̷S��*lv�):�v��)�n=lV܋%�� �IU4xuܕavl���c���[���q܅e�uUX�/Jbр�;2	���`-z��)L\��<k�i;6J���v�l�X�G.�7��8*L��U1��rv�mpθz��{'���ێv9�����q��e�= 0��=Z�>�bM��.�ν�`qnk�8�u�^��A�V�lO�W��r��D������1�����Z�$���H��D��RA7M8�[�v�3e��{�����`n�dj:�$Jq���s�`s�uX[��=T�����Jx�'r��N	�K��-�b��b ��srV��3������F�\Z������˸�dCH]�lm���1S�}�Kg<��J�~��� s��<�5��- wD�{MF��FJ��;�/�}ڪ��!�Db�Y �T�E�$! RU�� bEb�S��~�b���Z���.��2�%JrX0͖:�U�Ź��;��`��$t��`��S���d����1 w9�>�wO���?3�4F�c�+�s]�w���3��,u� �մ���"M�:�YqS��*qu�/:�{m* <dP�/�v��o�r��C���⦜|o��gk6X��V�w%#QԑR���7w�sP�r��� =|�_�#٩O$�	T���`w�\���~�Ŋ�",$		 �ʩ~�}�U5՛�`��,w5\q��JS#m8�-�v�͖���a�ꪪ��=�+ ���O�5��J��75 >�5�Z���f��rԛ�LY�ڼsn�t��l����=�8kɃi�]��o}����n���]��| �=��Ss`}/y$������^�#�Pp$܎��1��s]�ՙ��3��/��Y��q�Ƙ��X^�;�3]��Hܭ��;��VPfj �m��tӎ���u`Տ��M͂�DBP��9��`o�Q��T��%7#��f���K�s]�ՙ���v3`�#u$���Ԑp��[���]�Od���	M%�e��`BHG*EC���\�y�ͷ����|�Ź����������K��Wt6��c��,-�w���1n���o���٥���|�g�&�A���J"P�9V��U�gV>Y�Jg�y���׵`�@�"�%JI8�=�%�[�`u�4�>���7����U�f�x�)O����Ԏ��3f���3]�gV>X�Z���JIm����9� t�Ztʭ&�v�����{4�̩"�g%���<�ܽu���z�ZX��6����;h��n�:G��Y�/X�:��8�M�b�Sv޶��Yxc�,U�ϱy.ðnm7>�Cs䞒LZ�p��n9�wl�O��[�d6�m���.!�ю�uh"���|�� �*Y��׷��9��1�|��n^�Q��a�۪2�tc��!����qѭ����z�kc;-�;Z��k>sv�7ih��Y�n^��&��"�I���F|GMRE�y{ߝ�ՙ��3��?�}\A�~�1Q��1�ۥ$����_9��9�vIh\s�(��0R����3��,u�=�}_%���1n���Ji"R)(Jpn��1��s]����a諭�-��K��Wt��m(��V��Ձ���Iv����{��s`w+#�"")DM	F� �Sr��=�������yQ�6�������'[��I��@����k��f��y��U}�^�; �j�P�H�Jm���9�?VW[����� =m�@u4�Ҩ9D�6�t�9�5X[���UU�]Y�v�[�`j�c�Q�,/sm�b��b }Njݎ+�35n$�H&�����`l(J^'���=��x����T�'��Y��=���s/m���@�����j;Q�PKV׷7nE���vk+�a��G��=��=q�@z��@F��n�"������`s�5_ﾯ��#���`uf��w6X�j��t6�n����Ձ��Ykn�6!BX���y�偹���9�3`�hjR$7w�s�5��-�b �=������n; ����y�����`qw5�Z�b6����;p�P�J��qn3��y���-���ф�ӵ������Ҩ9D�6�nK�y���ܘ���9�	}O*^�A�����V��$�p;�,u�=UT����7u���q�Y�v �M@{��@u�1$�&�^��n!J�9#���UIn{���=�:�5ܞ���O��� (o7�9����&�%"��P�X��VV���:��|�5D(Q����$:c
�)�=[��og���oev���h7n��3'��II&��Ir����}���_9�����=� �<&�ze5) ����k���9ך���v��5����2�&�q�vM@{��������R�WPq�1�#�X�M,��vs]�gwe�����DQ��%!`uG1��1 >�P�@����\K����sgK��IN�۝��-�ؗ�Nz=-���'nUӞDٔ�2���WO0)�s����a"V��o!6�9�ơ;t�և��7����=�����.:�����=�HwUՁ�튶w[%r�*"v��y�'i�V�O �m���kN��V]�&0�a�1!�tv��s�π�6��)�z�v�qY������rPj�x *m��[M��K�m�����J~Y��ny�/=u��e�qղr����z8ܖڮ�w]d��^q�Ʋ��V���w��@����H�� $�F�Ӓ��R����3����sn���vf�{�M$I�%�87��7 :㘀��1 >�P�5���q���`unk�8���;�,w6��;�=Q5MJD�f����b }&�=�*@u�1��~��Ϛڸ$⍣PqG]q�uθ���.�C�3m�p�bnA2V��:w\f^f� }&�=�*@u�1��1 s4�#�
q�1�#�X�mժ��V@��,BO S@�&^:�;9��:�/�2l�t�y""p"���������k���9�۫�35n$�J��i�`qu�@����H�� �$7/6SdD�����3����sn���vs]��]Ǯ��q��}"Q������lm��8�N�N=c�����u�ۆ�b
�nѺQ�fn���\s�swvX�S\lMD���\���� �M@{�T�:m�e��H�$vf� ���?����`�1B*���W5�@�K�P�	��CdBhU�kE\B4 e!RQ�P"� Tb0�02Xk����	P�i������vs����?D ��!��!�C@���U��M�+�tE ����P'�k�8�� x�5���A���=�{7$�n��!���Q�)6���3����qR�9�[ssnfnU�N1F6�rK��u`unk�8�5�wvX���w�Ј��>u%���]v1ܰ]�EvW�ぷ�+ۭ���S��/EDNR����1{|�,�v�ݞ�ﾪ�������"ĘIQ;���@zۘ�I�7 :㘀�tn��%6DJ�Sr; �����u`unk�8�5��Ji"N)(����%�����]��*����8�5�r�����vX����'C�&�ؤ�\svI�x?������g�<['b1
�%��x(m��V�vwg��1�khNɶ�v�]����5D�O-ƭ�wm�nb �&�<�T���ۈka��S�(m'�owe��H�ﮬk�+�3]��ص��B�dm7{���7 #�-�nb �&�5wG���'(�Iʰ7j�8�& 	�j��HX7,�3o2����ʹ���t���qR<r�$@|A�U_�=ύjMkZֵ�[@�D�v��6Γ-D�S��J�ε����a�sć^��1���'v�/Kہ����944��v���܌#��y5^��w]x���K�9��w*�/mV��x�-t'nn!,٦Q��\����z5�n�2r���ϗ���vTfp�yFz��� :����W;�s�O���@#f�%���]��R:N"���n��6�7o7m3Vd-�|"!�:(�nꜚ�\��"�+��w��x>K��`Œ��WPv���i5r������0�iˣ]25~����@y��9h��@>w{۷�HP�ܒ��f�X�5X36X�vX����'D�6�RU�9h��@�����Gswq�:jR$���9���7����f�X�5Xw��ᔧ�PƜ�9�@y��;�����9����NޮӚ@���{8���q���,��2v�1�1�0p�v.�Ig�s:QJj���n*@G�Z���9�@K�d3p�'(�Iʰ7�5\����uU��AvIh�M@F�X7,�3n�7W&�*�6�76 ���zJg[�V���ͨ�pr����z�#qRv9h	�%��e�y��F�Fi����T������vX�G��m!Ԏ&%MJ�v��)���=U�O&�Y�Ս[�rX���?��_�N�m�I\����޽�`������� �ﮬ=��F�GM�D���96�77�	$�d77y`k{j��y��W�{Pס��R�)9��;�{��>�߶nz
)�*� 8���vՁ�~�9�V�(S���ԎI`F�x�'d��'I�r	��hBNU���U���d�� 77y`<�j��Jղ�Q�J��a�K�=r�:���]�z������&L���Bx�ݖJQ)��n$�J��n.�~�	�j7 #�- �P�n^f��w<\�"��`����Dɭ�]=�z�U��1Mjȥ)Pn9V�EH��@zܘ��"��{2�,�Er�5$�y�a�����;�U��ݫ%
;
BH3� ��u�T�Pr�"�+�7]��������r�n����y��μ�$t&��N�*qL�z�^���m���\q'��A�"���7������ w�R�9CiH��޺�;��V��Vn���jqҨ9N5y�������x�=nL@N�U��4�R5DR�BNU���U�����%��DEW��j�{��`}!��q&TMqXY����Ձ�ͺ�7j�3�n�D����ݫbQ����5�ٰ>�n�'������?���$ m�k-;"�u�N���&���|v���y빶Ԣ�[q!m�\]d�ִ��ݍ��Lk+��Va1<]��[�V'��n��P8�Մ��<t2�E�մ�={(Y��G�7�tji��I�����2K��ɖ���85]�od;hm����#��Ş~-$6��W=rJm�k3tNGT�N������5��y���G4ݸ�g�ճ�DS�i���U%�d͗Y.��XfܝY��n[��[��Ong��Sd���Ց4@!$$*�4��h��ٖn����?ߔ����Ɉ	�*@>��/r��$q�(Ғ�ǚ��W�URGV����{�Vs6��;���ӥ�"@�H��& 'H���H��@�M?U���3.�q:EHn*@F�U�����]{�;�g�8�T�M�^f����㖀��1:EH��F��n���P!�pI�P�v�&�7A��h�����u��E��N���;Em�I$�qX+�N7V�v�%����]XA��A���)�J#���rbu��[���*@zO� #�- �Q�Q���DJ#M����Ձ�ͺ��}�UR^׾VV�����Z��JS諕\�+(���{�5�ٰ>�n���Ձ��5�Н8�iIV��h[��T����=ɛ��k��&	�e�[��=�/��vMו�k�M;V�7W���{��|�c]�.tU�/�uϾ�� 9����ܽ ��=��)O����vw%@9��Ձ��U�ś��_W�}I�=��J��N�������Հ�͒�]R�P���v�v��Օ�Hڢ)���`<�s`}8�X�ڰ�JS�����w�cq'RS��G�ś����@sqR<r��̕�����^��lK��k=s/m���|�;����f�e�U�;W^T*���Q�i���ݺ�;��V��Vn�:dz���O�W*�\Vs�؄�)�]=���j����X�SZ�	�㉡F��`n<����1:EHn*@���ʸ'(�")"��}�}_.���������;VX�DB�J]��f�\�oŕ{Xm^e�� 'H���H�˰8�u�Z�b6�I&�ӁJ&�A�����X�(m]��u���>�ae����5f:U)Ɠi��X�۫q���BP�}!��j��kkNUJ9<�p��6�㖀��1:EHn*@qf�ĝTD���,�v�]�5(P�g�V�{6e#
*�f�{��y����"�7 #�-ś��Ι�p�����U��͵`<�s`}-��[�`|��!B�����ݘ�ȼPG�F��|Qb���!��ܦA��3 4Q'�@��O)�B� @�H�I��2 Q���V�K�UW�A�š� �24!_kX#q�( s�S{��b� `�.�0�����F衁�Q�D�4�� A�b!)�# ��,���^<�B"E`���wwy���������6�  H        8     m�GL�j�ڮ�uI�m�T����:�8�]�-�rzGv�9h��-����o�|�V�{7�臓��4t2NSkl�n��{T��f�0��Mh�l�Ȉ�mc7S�t�qĚ�4-��WL�}�b�R�T��7[�Ĵ�1�2n���y�Es��j����-kkm�
Curl燫!�Y���9	z|�X5�>��l��"$vQ�S���M�cvg��k-�љpA�k�SYcgmC���g�"b��@�R�φ���ṚےrY%5�� m�ɲp�N�$�lK)�-4k�#EI�J�L�� 	m�ݗm�h[f�$"t �V�[�=�#T��giG,��l�u��.�AKP�T�n��T�;���ٝ5�iwaR�B���FgE�N���r�J	�3���7h1cfj��X�d3.���+���4X���A)c�\��|������흞'�;"�ꀴq�';��O��cvFd6� �µ��"Wm4�UF�;h�]th	Ӳ���i~|_�>:�p5���'��kK^$��My���lڶ��`(mVrb}�>J�iw���c����k��[l�������	m� �]���^��n �]5F�
������	��R��/��(絶�Ԇ��uUUUWU�C�+/<�YMU��RN��ț ����u�P n�K�ʻ-�4��(YI%dL�ʵR�U$m�*Z�Z�ו�����ٶ��q.�� H�k����g���[k�OR�7�Ԫ�+�6���ʮ����Z@Z�q)AQ��˒�g��۸ڹ�X�Ź�.����x���nӌ�]C���X yK�
ԦJ�9��[i�ڀU�rYvU�ñ=���P��*e�P�䔲����dUv�����
�df�.����:꽕N�aa
W�2(�Q^|�b�Q�\U��ۄ�%vR.:��kZ�2 /@���| �(MtD�j+C_w~�������   etݝE��ud�z�O3��-ШNs=g7!�PYغێӞf�)')"�=:*��Cq�2���mJd�c����I,����^�Y�^�lN�vxRݷ�rGVE�F,��:U�7kf]㗈��yhӍ.��Ѱ7僭��BF	ӭ�$����z��*��n��2�aǋ<�㝎'�/L�4qk��d��Q���Xx>�{��y��Ϗ�m9:5¦��<�n�m��N\���^��b���I[���$o_绽���#�ĐN�(Ғ�~{�X[���۫36��7qk��J
@���XKn��$�������u�oaz!DD*�~�
�$S�G�O+�`o�֬�v�򈈉���l��Ձ󡲸�T�)��mʰ33n�ך�,n�<�!(R�����kkNUJ9<��R$��+c�ݧ�_ ����՛����<-�r^.�.�闶ےB���uw/�z�:��ǜv�X9��2�ʹ�ɈT�����3�����:�6�3sn��Uj�Q��!B���}j��}6ӍՁ�2lN%"����$�U��ͺ�3^j�8�u���VwT֣Bt5 �<��qXz"!(^�����;�U��6���f�X�-r7N:r�(�����1 ㊐�T�s������>Rs��HD�f���ݫc�w#�]�.u9��\����p��M�����\(\�;Vs�c�z��d�V~g�Ď���i6�X�۫5�h[�8�-�!��n��D�5�`c�s`}8�YP�ET(Qԅ`	T���B#""��K� %��� f��wVs6��⣻�bpT�J�t7����g7ޫ}��`w1ڰ1�5`f0ǵ�ܨ�Q��vnmՁ�7}���Vn����]B!?�ՙ��/K�o'n	��N9I��a_X������mئ�~��j�)�ID�S�G+�fﮬ1�@zܘ�q�H��e�yA��'*g�V:�7�
&N�ݫ�۫��u`�����R4��+����ǎ՞�3���=� ��
| �OSU3�U��$�^��X�ڰ1�9�����Dv!(N��.��������i6�X�۫�Uo��p������u`�{���
���Ѫ�z���2]�DTtp=a4���'l��OZ(�	HE	9Vk�Vn�� 9�����36�M�Uɰ>�n��L�^ڰ1��`c����H�a���r�ێ��o�X�v��%2��́�{�`grx�2%"����$�U��ͺ�3^j�8�u���VwT���:	I�%X����=���mX�v�D.�������߯��B@��U��e� �)�I��Wc[P����6�GNzN�Z�nyy�p�lK(�G[0�ףj�{D���p���Е��cb1N����;Ygln$s�`�]�3��w]��/8ɂ��q�1q�8��qљ�u���j�����[ϓ�3Sr����v�\����ۀ�(�6���j�˓��]���9�˓���l��7'a@��su{0��������q����^�b�Kv-��Զ���ɷ��B����;v5m�[��DM/$I#J)"�5g����ͺ�;��Vk�V��a���ܦ�JG`f�ڿ�
d��Հ��́��u`|�l�*��J�	��r��mՁ��U�ś���ͺ�5f�IHE	9V��=nL@8�~�nO�H�yn%N��`qf�3sn��mՁ��U�mj�ZD�����I�_��� �/kn�������_Fx����ao\�	!�ܩIĆ�|}���;��Vk�Vn�;�]ԉH��}*I9�+����D8K�G8W�}6N��`cͺ�3���'I�:��F��`f�Ԁ��1 ㊐�T�$w3w/+r��H��H�=_.���������f�X�5X{����EJnSM%#�3^���H1�@zܘ�+���Y����V�J z��{8ۑ�83�e�;ysŕtm>yN�"]���7D��.��O���v�u�l��I} ��Ke�^aHE	9Vk�Vn�7&�s6����ĩ��c��6ӍՁ�8��z8��(H�`@�Q��@M���T�z���?j�3)�l �����a�/^��omX��N7Vw�u"����$�U��ͺ�3^j�8�u��4�9���FEQ:M�d代����'��m����!�.���-�r݊i��S���&�Hu%�)+�o��X�& {7 	���ʽ/v�ۻ���@zܘ�q��T�z�U�w�*{�D��4�R;7&�s�6��{6e�Ձ󡳜�pd���I�*��f�X�5XY��&��������Ձ�t�N0��"����@9�Z����*@sqR����ߧ��>�㫣	y�G�\h���]�k�wSm��c>;p����;m�8��=ݝ�|�k-��i�e�|����@8�7 y��̧X���M�
D���ۤ7 �-�rb�s1V��{(�J�I%X�۫5�=�|�V����{�VwT���t��RDiIV:nl��v�<�ߕ�n��s��PRQ"J)"�8�u���Vs�c��cn!$�8lޮp9�UR�U;�v6x]"�a��b��58�:w޺��N�㖔
VѨlk��Ķ�ŏ�k�Śޭ9�������V��N��d�5.��͍��l`��c�O�l\��&�<��g�]��+&kQ�;t�OW�v�Q��//2�zn�pk�4���c�,먅������쯮��Ʒs)�*ޞ]6om��[���Z4�L�@����G<�m\�t�c���d������:v�D�hy8�v�Vt\7tX混�\��G�?��7 �-�rb����!ȕF�M�Vs6���RF��f��ڰ1�j��)�e�\�O�{E��m '��ր��1 䊐��XA��A�&�*!��Vn�v��;VR���`6�:��k�U��Uʰ1�j��B��7�/�~~�8�u�
�ܶ=��&�@:�SCѰ�ܓ�v�sv����웋������|,�Qu;���(� �RQ>�$�J��� �<�`qw��u`{4�8�N�D�!hܓ߳���Qآ:CGe�����j��c�~I%
d7\�9ʧJ
J$IEVV����ݺ�;��Vk�V���>)��N���H���H2K@zܘ�鄆nR��S��I�*��f�X�������\�}�`f��X����A�$;�`�����|�rv<KE�0֭�]�/.*��u#DU �BI9Vk�Vn�� ;�T��]t�{y�Y�m�Fn���b� ;�T�s$�������3iֿT��BPێ��{�7$��~ٹ�";��,��t�aZ���LTb� EM}�~����FhV	%<@0B��c����|C2W�	!�9 !Si��SH��"�X�5@E4�OAGf
?" b��S�<DOh
J+�����RD"��@� �T�I ��(�_�J� Wj�:�5���� �RQ>�$��V�
"'ߕ���f��q��1�j��i4q��!Ԕ"1IVk�V��J#����wmX�;V�O�뜘�Lt�sZ痞��N��n��v�9fm{c�u$����jn�N��Y~�����1�j��q���A�ǹ<�i��JA'IH��۫�ͺ�1�s`}=n�W�J%T?Q��R���Ene��f�O���d������rmՀnV��H	!9Vk�V�����ݫ%	-s��� �$������rOJyޗW3R�˫�1�M�����<�����/��{j��{����ojF*R*P'�6ܨӮ{m���>;���!ك�P���pjz�m�-����h����*@w8� �Ih.�3���ID�I$���j���BIDU�����~�X۵`s4�8�N��J��5�����*@w8� H�n�fU�{�o&g����O[�v���%��DBU��zl_��� TqO8Lҙ�) 䊐�*@9�Z��b�U3����  t�/2�v�bcW6�l݄Ku>ԁvuǫ�띞�\C�=u��۩���Pvk�6gF�E���W���7(�A�nf�/���M���$zn�\M��^`^Z+�3Y�k6[�rǐN��ݵ�8�L���3�n_��!�7>�l�=�`�=:e��u��h��cc�Z��\R����[!m����CtOҠ��p�Us�nRs���_�w{�q��8�aB��m�3�6:뎓v��06�n���`S�Q���j���3�P�����R̒���H� GR�ҨH	!9Vk�W���ꪤ����������6���*��(��hp䔊�&��z�X۵g�
g1�|��`w)�=�'r������j��qڰ1�sa�P�'���`u�f�D�RQ>�$�J�;�۫5������ݺ�1Wq�@�DJM��ď=[�����v�k�Χv����V�6;!s�s�q��!Ԕ"1IVk�Vw]���u`w��V��쉴D��D�Q��I���f����"b"���U��{D��H�ʐd��B�~���{��U�� �R��H2K@qwu��n�:T�q�#I7!`w�T�s$�����*@ԸnbH	!9Vk�V�����=��7ޞ,�mՁ��{	$����k��td��۳5��2�8:����H'�^�x�5���(��hp�t9�ś���٥��ͺ�3^�3)�=�'rP�(���&���d����1}U_����WR%"����$�n�:nl�	R�P�(J�(���V<�X�&�6'@�J��`f�Ԁ��1 �� 9�� 	�ݼ�5)(�%qXY��W��վ�����Ł��U����?�Q�B�R(ش�Q���ճd�r*����×r�v��]�Q�5���I�R;7f�r�i`f��`qf�:��G*M�ʑ����;�8�76ӍՁ�񗰢���^^#h! 8$�)|��`zܘ�rl��fS�W���xe��f�=nL@96t�� ��Z Px ��<�s�+��Z���M�B��7���K�D$��DBOV��o�ޛ�������^���t�{U/<^���M�����������xo.I'n����"�)N�874@s��@9�Z����`�}�4q�:RP��'5��5Ձ��qg~��򈈅T��{�����QG��߿;7f�~��kg�|��`�C[�T� ���v7�XŜe�����
"{Ov�^�xq�CiO�i&�,�d���ID$��v~��j��ݫ�J9
;��W����nvΗU�V״��1�۫n�Yu��\
i��λm�z��8���%�u�ѤS�)x"�lG7n	X6�mV�S�klR��skOb��&J�z�)77m��m�["I��q���6Œ���ڱ�`�X�؊���tj�'0ɺYvI�vⶻ/5��[jN6,����v��Y2���/93����kk�K�J/72���Mf�f䦵Y�:��)����o���I�;7K'�Ü�û�'�
p,�v.�t�x�ݖ�����KK�Z���T�,uś���ݺ�U}��Uqml�`wG[�J&�n��!�I�>�n�mڰ;�8�77��ԑ�N�Ђq7%
��v�g������"�3�[�`v^�Xb�_)�O�H�p�;��Kz�U�ś���ɥ���5�����J��`>�s`y$��=��o�XŜe���cPI0Q
&�H�(R���Km��Twka�d�W]�rn8�}�	q�DU.z
�v���6��& #{:{纬��z�/�9D�IH�̚\�(,��		@�秺�XǺ�,�vV��㤆�j�iT�8XŜe��M͚�B��{/v�n��Z�������T�,��h[����=����w[�#t���C�XY��̚X�ɥ��{��6�j�"t؅*F��ϗ|,�.�m�x��)�;v4Y��L�$��P�ə��*;Uuw'rP�(���?y��;��Kz�U�ś���Vip��I�V�ff�t�	�%�=nL@G�Z;�kR�:lD�"5I��޽�`r��ٹ���F0XH(`!$"��BH(@"��$�Q�`�(�E<�����<��]��Nn-�6�����+�7]���K�����ID)����{�y���1������@G�Z�=�vIh,�v�͒T�!�*(r��"I]ut��Ǒ�@ǅ��e��q��ϳv�D����=��f�&�eH�iHp����޽�`qf�7j��դm$��!`>�s~�'e�Ձ��́�Y�X�Y��F�P$��C�XY��ǎl؄���Ɵ4�7+vl�K\���n����f�������ܓ�����	]�	$���u`}�V�L�H%R�m8��d��޽�`qf�7j�9��
2*�����jWkkn�E�n%�oaL1N��[v:��ݚyT�N��IB#T�,��Vn��c�%P�;@�o<X{g��*�y33�QEqXY���Wԑ�{�`f������_|�n�ȑ��"S�Jt������9�� 'd����1�*h�I���4��+�UT�koŁ�{�`}8�Xy$��|{6�l�ʩDR�IR��7�uXݛ�>��~$��kٹ'�EAU��
����EAU��
��PT_�"����W�H*
��EU�
��X*@��
���  �B�*�* *�� *
���ET��@ �D *@`*U��B"� F� 
�EB� P��DE��X
�H
� X
�*�EH
�A`*@����A"*`*`*��
�AA��
���qW��*�APUj
���EAU��*
��PU�����T_�"���B*
��*
���PVI��y����	�` �����Z��            }4       �  �*DA�%P(R�ET�� P��@ *�
� 
( ��H H  ���  QTU��( $3`���C�-�ʸ���er���}7ǾE=�����c�ׯO"�2z�� �w>�������W�{�C��Ҁ`�v�x����7p �=oy���Os�f�=�/x�U\ �� QTQU@P
R�l�窦6����=���E8�U� W>����&�qe�O>�>��Pt�q��S����M�>�� >�K;_y�ɯ�94����}� �)�޼��}�_Y|����n��> @UU ( c` }�ڗ���� ��QI�  �ٚ 3`�� �)F�� �( 6 ҉�@  &Ɣ�1 
l  H @ M� b ��� 8�JR Q�;  0� (H  (1��� �� M� c�O�>�J�w�{ʧ-��kٽ�:^���0 ��ɗ���׀�>��j��
)�ϥ1we9|�z�7C׼��������5���|��}y�w��ޕ� x> 	H�*�l
��V>�Z����s�MN�}�K8 �������)�ٽ�������PzK'v}o>��� �|�s��o}��` =�S'ݟO!�&�ox�:W O��[ϹO=�-95s9����   "~���)P  "~��{*�)�@���R��� �@��T��)S@  "���J�ڥJT @E4SeJH� �O�?����Y��o������]��{���]�� Uz��� ����� ���`EW� X� *�D?��I�������
�b��Qk��]$� �A�� 4��ԥ5
B(@`"P��V'�1�
�4�̖�!�1������ԳG1%�,�BP�cM2�\0�X�$$V2"B#b@˭�ϧai�oL+z�7�)�x������eeg��0�}�t� љ�*�Y.�#��]��4�4M3h�������d3Z��{9���D��5L#V���r�Sl���M�5d��l�X��M�eI��4i6Ji2f�C.p�7$&�V�3F$g�*���y���3{z�w4l�b� 
:Z&��d������f�XT��aR2��#ă!���V$H�P�b]��&��IB�`B25jĂTb�t�"�J�5^�è�@��!sz�W��>�|)\ }"�� ��8d��A.�u�[�]n;�ٶ�V,*����A4�(D(hǱ�@�.�h]K�&kSF�4��I��wx�!JD��ٙthx�h1�*���8;&$J2,CN�3��!R�CJ|���D!F!,k��(lCCF"�xi!F�
A'�!Щ)b� F��6��hcB�7.�B�!SH˟����>ڐ)l���4g�aCZ5˩�q t�o|�7��h���(A�@4D�"�9����l!�4B��Ea, �#�K�k�kSR�bjbHMj�MXZ`i� ��DB�{ψ� C����Z���, �� �X���.�>1j0(0a�# D H����-!P�3����PѲHd�A��N��p����i!�H����8�8��
i���	������7XW�2H~�]1!��~ܡ��[t�78~D�h0���a!�֨�� ����XkC�l��F1�P5��~d��M�F����š�&�~%��	]c>�@���H�B$jk_��k?�� �1)$d��A��M
° @�B0J��@p�$���8���Ҕc@���E��@�~HA`B$��WG��� �"`��"At	� �6	��~8�&�o5�&!���@��"�@��*��؄�qv;���6]�������?�u�@!��'���ӎ��~SFvp�~6h��n�?�G⤥ӎ�g?~6l�6a�?�ji%���4V4jB��IB�?Hr�Mc
B������j˩0v�h@�L$6�xf�sF�ns�%���
��?a�q��x��bB2��C
@�+�*B�b�I���g�ɸ_����~"IGIB"HF#�0��ٝ�>�Ȭ?g'g'�~	�g[���u��w#6K�0���#�#��f�r�#(A�M&ǃ� BF!Mk��x� ��yIk6��nPp>r$�Xaa�#I&�d��0H1`@#: ��$i>��wO��W���W9Î�d�XƄ(ā 	2(A������!+�ALH
EL�7F����h��F,3YB[�!�����]fkg��Ɩ4"W�����u��Y����~?m���B�6�ݼ��Y�~�	���aMq�X�i$p�я�!@�o?���Û'B�����S��DY�}��W���a�D-ֵ��]ϫF�����D����5�6u�f�kFJkԆ�, Ō� H F�p`B�-4a���@�Q4�`����*�D�#��]I���?�����d�4B8���$Z0�!�c],hD+@�i�3��j�����O߫3a��9��K�?�����\���f�Ys]:t�~B6D���H�Qћ�yyj�0M�	M+ �`�*¬h�hE��F�F�+��oL���Z��� ���d"�!c[)R������U���Hk�X�J	;�~��&�&7��\��
�g䌬�+aO�h����t�J�z�T�Z�����$��f����R3S��#�
2��$I�\��$&1d'��m`����}��g��l�t�u3��H��v���,"$
�*1(�+�!	fmi���*��������u�Q�.�e/�Mf��G6O���vs'��uY�ĺ��a��&������MB�9���p0�H1av�o�Zټ���8H@bB��|��d��B50��֤$��,.�]1/�K�Յ*Ț���uu�# �j0
� @&��}��D�v[�V5�'߹tA�!HAd�n1*�_��� F"Qt���Al�0bV]����?�8���o{�C9��|C��pņ���p���l��bB�,�7��Ya18ƚ�5�M��̉FSl���2D6l��4a��o''����+�����*K1��
&}�;�x���{���.�駁��8�'��R"�Hb;�#�3�!#�GG-oœ���ᐚB<��>G�0)�8*i"X��Q��N �C��o��nS9�J,�#��H�XD����L��S�!�XY0�P��dbF�h�dn;$"HJ�Đ!���v��Dѣ�\�o�E�Mf�dx��x�h�fc���RM�B�8vl�`�ӎ;0XSN���M�:!�B�6o�q���n�3Y���m3��p\f���l��;�������qػF5�`�����fv]�*��1��I\v�LF5ӎ�n;1+�6K�`�6i��k�6����
�C��d�.�6l�r0�5
H9�͘H�ц��m# �h�a�#�4c�d� F��7�SHG�H�2�y�'da:q�SXD�@ A��,
#shn�nϦc0����0�X�)]EJ�[)��v�(�Ąƒ�$J�H#�m������v�.���p�6ʹ����c���l��kk��̦���@ R*�,��C�D� ؁�$��"V�����u�6IHYw�[p�#dH�a ����đ`@*@B&��F�IBY��@�0,(��	�	�`EF�ɽg#u���F ��b�L	$i�3��i
�6m2�WpjL6m�5��, �$�uћ]�����&vjYF�&��e���
��pht� D�E�!�bW��F�#0��j��I�c!A�B�1bA�,H1��l����c<�	'B�(GX�FAcdM!�d�		m�F��&��6n5�t%u�4jJkGi$5����o�"]:0�ȗXѐ�XB�HWI�E��>�����a��֊t6~���[?=��"�	�����4&.�cGL�G�>               ��                                    � �                    � �            �0�                            m�    �              -�l  �Za�۰]�L8 �,�*� h  I�v�mH  $  ����4� ml�,�U�� +*�����l�m�����   h ֭��m�H["I��	A�-�,����,kx�C��*�|�*��UPY �z�m�]5�Z!6�UJ��mʰ
�pUl���^��`'�����-���/ZV�h��ckmU����H�b@$�kz�඀ ����X�b�nNX�)V�.ہ9�i�iQ�۪ev�-<����U]�����LևH�` c� m�m��Z���-��0`  ���{ﾀ p -���5��ie� m�#��u�ܼ���`A2j��v��mPquUŐca]� 8ٕm'����1h$`  �7-����#���md�mU\�O�%��Mr�l2ӤͳE$  n٬�'d�);7pM@� L!�l!��ղb�	�$�'ju�������b�K�r6�媪U�3R�@ ����V�y��EH$�m��۱`@M�.S   ����TJ��\��-mJ�UC��9�� 	�Վ�n���`���S���k�m��֊ 6ر��$�4U�6��ށ����nܩ��m��P�m�F�D��l�nݗ��P-�
�-��m��H -� ��#� <��庫vU��cZ��^j@h-��!�l m �`$ ڛ����Oc݁ -� Zi3��qE�	X
����@[Du�sm�hݶ �H qm:Y[[�{YfG=+��pV�UR�Kh�˼�&��![`�����+�۞$�4��`2�؄�s��mSmu]�N�am�H�t�n�
m�l\�`�½9亸
�6N�]#$�ۥ���g�X`"mqn�[[l5�    ��F�` It�؄�p႖�
�d܎I�m�6�@6ؐ	lM� ��� � l m���s2� ���UU              �`�  -��  6ݸ�m6�[M����nm�pq�kp��K� 6��V��� �Z��t�m��s��ۉ�7*�A��Z��$H]6�pc��m����Ih*m��pm���`�n�d�[-��l�nm&�m  m���ז�9�*˱��M��k����E�V� �u���8��nC��{b��u[T[t^Zv�n��6̆�`� -�y`%Z����1�F�9�� �bŴ#�zԌ�l[y�m�� Rxe���WN.f�{\;d H 	�Ud!���j�d����`  %�۫b�6��Ԅ�*�Ö��'PA ��l	��h���մ���vM�� �{Mv�lhm�ݛc����Mz�d8 nI,�am�p-�$m�/U�m�,����h$�t�-�[&��}T�}嵐�-Pl�[���k7"�Hq�@@�h �����UP9�Z�8��[d�  7Eݶ  	�8����m�I�mI� m&Z��`	  �[vض�5� 5�!P�ڪ�y�UeZ��W�2�p�  	 �6��$��lڶp  ���˘ր���M�6�` m�     o��zmm�$o-n @       iXI���W��5�@    ���$�H�J�o6�� $ Hl m� p��  �z#�Z5�U]��Qq���@m���jG6��     �m-� p$    ��ۛI����|8  n��St�20���;�6��r/[mg-��%-�;^� ��	�
��Yrt��	d�� �.�   p 9,�[A!%�m�m%��Hm�$�     ɷm&� [�^l       #����,�B���W�]Vxk)eI��m� .�m�Kz��'8��N�&m��  e���*����Ьl$� �  m��t�6�n�]]p sj�  �k��b�1K=�ק�ܻ�c 5@     �۴�l����n^��ݼ��>���L�    �`-� -�I  9m7m����j��ݤ��y�ӡ�.�~�_:���j�MtP�&��m��
P  �Ŵ	         �`��  86�` �f�� ��� j��@�k�m�+5��'N2I$�m����$  H�v�   8  M���<[@�H -��wR�p �f�m� gZ�m�l����9��2C��m�L�l	�� m�I$��l�k�������� -�M�m������ar�.�Xɥ�S�$�h��үT���T������� ���b� 8�@IK�l�׶˪\ 9U@�U�Y\nej�   �$��	�,�p��Kz�p���{	h[WV���В�9��l� [@�  8 -�m���`  m�%�\�<v�.�U@pW1�d�gN�5�i&Z����̝���qۜb�������jY4��[�['���tݨH۶):�-��6� �ۀ�@�v��  @Y��(�V�o6ͱ p 
���:K�.�� �6�-��� M�` l����]�i2@ �u�r[o8I��e۪VV���)Y�-��m�    �4�iu���]��    z�=�ݶ��YŴ$m%l�[�$)@ -��9�݇   �l m���Ӌ��l-�[� �I�H  �f    ��  ٴӭ�I�      mo\  ݤͰ U�UUJ��3�
�PKh gYxp�	w%Ͷqz��`i3m��$kX�����U+++r��@s(�u  qm�nհmoY���oVB,��HM���"�c�v�볫m�m�$sm�l�m�l���ً���ְ�  [Cn� $�����-��6�wNZ88  �p[[l,�:�ٖ����)E�  �6� q'6���?�!J��uWUp���@���6[EUUHl��F��VU���I��K6�3 N�
�MU~]&�|V���V���-�0 ^�mYv�Z�)��*�����{-R��*���m� [^.�m2\��Iҗ`�p    kC`ͷ^�-6ۋ�Z ����&�[\  �V��63=T����䁔�5�� q�ȷ�"@<$��
��@2�.ܽ���n3 ղ�Ut [.�p�H6�4rܜ���m�$ �֛` m[   � l�   �=�9n�    �[v�I�  m��� m���R֮�  ��p	�[Kh8-� �hE��f���.�t�v$9m t-����@�m�t *(N�����&�vÖ�!�V˪��p�B�ҭ�À    �+v�j���   &�Kn-��,6�ҹ&ҭ�t�����[@  �l��i!ƶF��    m�  s���� -���,5����~q�p*�j�P'XNC2�no6݅���͛�Fh��z!�+f�e��  햁�m  -��������� H���}�-��m&�m�� ��       H�HՆ�  ��  	$�޸ H�q�`     r@  �6�V   �PHi3l  8 6� ��  �  m�    �6@h�U��m8m������mI�l��6ͻ]������ �3�� $-��ӳd�ƙ���Y,�r��܀9IіH��6�"�*z���&[I��m���[@e����	 N��m�k��L��n݀mf��Y!�p�m� ����]�U��R�R��f���`�-�m�  ۵-@n��6�mm�� �m�s�l���Z55Pq����������ɫ�33Z֤�?� S`"�
�U_�Q� ��Q�I�� l��@��Lb��? ?Ȣ�MbAE�	��AS_��"�W�U�� 8E0���R ��D�u≱�"?� 8
/��(~�v��G�P 8@A�l]�E_�
������%"*E`��!��!�U�*	���]������@�@ Œ'PP�R ��>A�PMA�uP!�T>�O�)�L�! �Y �V1Q"ȡE1R���"�w� t4
hQ0���C�G`���E�!��~Aڠ � �*����QSG1�)�
p�"0HDX		E!ńU����t
&	�V��*��_���(�@E���Q1T|��T0� tP* iTLDR�MP�1Cj ��^���G�H�D��pEW�?� ��B$@�� Q?�	5�߳3330 m�      �m��  l� m�    �$  �5Y'[�M:��;m�Y��E�d��͵�.k�+r�`Ψ�nXb��uR�Ł8e������Id�u��:K����Y��)#�����(j�LH�NGLs«�����Ŋ�>�H�X�F׵�7Q(ݙ%�I�n��M�RΈ뭡�X��rR�]ɉ��F݌x��1�֩:P#F
ay��X�D��޵U�le�F�I� @ +c�U�  ;m��4�V�is6Ջ�Q�Z:;'A5Ҽ��&�J����#�{@�BA)q1����u�2�9�s��T��Gs T�"�vG����P�M��VA㲩VV�ͩ���S[$������*���G*6R��6�4�Tm�m�9oCc�j���i�R.{�����#3T�p�����̋I�=J��
���y[���W$#[URv|��b���mb�m�v���v��9��ke�L����J�r��t��;�/m��qm ��A��z��kY9B�Cmu��f�7G/N���9��@e��IS�����n:ۮ#EUQHd�Nm�M�4���A�<�������[ZM�Vnv�N�ԩN3L��0(�fM-�h��� �,���&�v�PCnl�[TiUiv^��pu�㋋B݆�ɽv��w�����[��P��yv`�'��N;�wR�Z4걀�t�kڕ���vh����s�F0
�vugUm�`��YV���/`ݽv�q�M�.gv-�[iVU��6�[j�LFtl�D���-ɔ��N�q^k{U��u5fRx �n.	�*���x�gI��T�%���'6C/idm�� �n�M�Ha�hG��`jU�m���IH.�B���3�;h��c��L���Zl�	_7ڕ[r��xv��v8��5b����h����>UW��b� S��D�8� mT�^�����<�=��`0�Rn���*�J����y7/CXŴ��=#����CF��%�3�1N�&�x"��@Ԫ��Wk�=lۢ5�ۋg�
R�n���I����֓�2dl��C�����u�;Og�M�qX���X�YDw���3]�<\��k9�"(qgG$��ioG'<jS��y����l`,q�$*�5����w�����8�\}���]�˃�&�s�c9��7l;3ݎx�'�enG���^���(���������o�@�aa����I#�܏@o*Z��G9���Dɏj� �{V����oR��#$q�#qh�e4׬�<����uh�َD�qI�5��z�����ގ������^�hm���rH�H�sP|� ${��t� �j �ݼ����B'\�9�7<T�g�CTz
.SNM.�aw,N)���e��w=�h�lG5��b�8uƜȘ��i8��?z�k���> ���� 	� �TJ���K����xgڀ��1#ܖ��u"��O���Cp�^�@��W�[�ՠ~���=�\�eD�)�4fnn�:��@H�%�>�@��a��J�y$H�r=ގ�����s�D��@u���3.���7rR#�#�<i;[��=n��T����nw\9c]E`�͜�\ΝL�,|�}�`�:9��s=�hnM��H)Rd�E!��f���@���@��)�3���:۱�8D��y&�f�7$�}�nI�������(�Q��g��S@:�4�i;�lq�����uh�e4׬�<����î4�D�F�I����S@=z���^�oGV��b�D?�m����v��o6N1X�K��R�{&t&�9�n*1mO������բ����m� �Oڀ��1#ܖ�����&�ʢ��Dln94/uz�Z�YM ��4�á���H�&���rZ�_�ꪻ:9��sx�z�dd��4�n-����?w��䟯ﻭ���W�? .�V��ڠ��f�w$����Y32\�E&H�R��h^��z:�߻���yUo�Im���Ra�Hk	0��K=;�#mt�����2���'/�>|����3����w6�֋�`]��|����'Ǖ-X�}�s�׵`vR��f�c�7��@���@��)��f���@�yc�1�#H����-���@u󘀑�K@s2�5I�����Cp�Y�٘��Y�w>�@���@�l���/䲨�dl����3'�6""9��utn֖���ܓH��C𳭨`D�D����V&�����QO�*؃�i!�mjk@���f`l �aۧi��Tu#"ۭ��Wt���l�2cuw`�v;qez�^�rZ������F�����0�6��G����W:��9&���j�v�[��sR�U��ݗ���n.��%-��K֬,c�y}jT�^*5n�ܗ92��m��Β'Ul���Xҥi���q[ҝp��l����	#�/�wϑ�ٶ�Z�!�����v��<f!P�;F���gI�&x���ymm9�	m{��E���5֫���w��z��h���~���������~�����ʴ�Q�J2ITUMJUS4��L����q �{V���z:�+l�	 �qI�5� tsP㖀��K@}&� ��I�"�ɠw>�@���@�l���K׬��+`�m�87$MŠ[�ՠ~�S@=z���_6�}��߽����r�fwU�Ӻۀ��>��Q�����)�D�^%���4�#H����/�{�ƀz��s�z:��ΤRbp269�4�~�o��<��T4;��׷w$�����?[)��#�TX����#cq��-#ܖ��M� ��>�(�L�U$T��U+�""!n��V��|h�Y�w>�@��cz��!#�)�@�l���g���_�����@���@�h$��e��&LmLK1]=@sҮ:�jU��F[
\�Nn���E�Us��RH���C@=z���Z�Z�e4��dJL	$O$�GU`fN5{���$n��V�� ��4�$��q�8�ܑ7�oGV�;�w�sB	AE�AO�G[��nh��@�yc�1�#H����-L��G5&Ih	�fS�Rbp2691��z���ՠ[�ՠZ�Z�`ڢN	%&�@�5t=�N��숱Ola&��˛�Ӯ�a
�QbGB����&�k�h�uh�V�z�����J�y$H�I�oGV�k�h�Y�Z�[��������ח�N�L�,|�}���h�Y�Z�Z�Z��c��RH��#�C�K��M��-ޏ�rT���@ϻ���'��u�\�3I�"�ɠw>�@���@�l��z���`�T��ɎA��7������x֎�����;�v� �@L�4�7Nn�P+��lq��"n/�}���~�S@=z���Z+���doM�V[�_��f���z���K�����D7 ��4��h�uh���=�E�Y\Q
267�s�z:���h�Y�~�(����I#DRE�[�ՠ~�`�:9���@:�����?n���� ���"���r4��M���h݋�퇚��r\1)�@���D�����: ��I5��+���cn)'���]e:���p���8�l�y0�rW#���%-�:��u`T9��6��[���]�yv�����n�]���S��Q�;q�Q0X��������(�3A����;�,���v��f��gBt��8gR:���|����O�����غBt���������]�R�i�6�h�&�^�d�2��aG��X�ѫS"����w���<�Ձ�8Հ�T�`y[f8I$�Lq��4׬�;�U�[�ՠ~�SRG[^��I�U*���3'�ʖ�������guh}~���V�rF��&��-���-v� ��4]�@�yc�1̍�"i��@�ڴ�?��}v�����j�np�NRT�5A㬝���r&"h�|�8,ENN��.i!3�%��#�4�"�����ƤZ��h�V�oGV�k�h��,v˚��Mk5��'{���E�b�+����T�`7-� ��V��\I�y$H�I�oGV�k�h�Y�Z�Z�^7��&HH�JF��-v� ��4]�@���@��p�
I��qh�Y�}����}>��7]N��mX��{vɔ�*hX�<�{\˵v^��u�� ��\m�V^9���+��MK�fk�.�L}I?vwU��T�`7-� ��V�I7C��8�ܑ7�oGV�����|��h}~��ՠr����F�4��sm&Ih�MGT��U�ʯQ�B(�~�6�UB�A�� Sʍ��tK4�a(���U�6&UMhNhD���U^�ڄ*�$f^��*$9n�<��> � ��H�@HA�!d�
FH��TlH���@�;~AE��4x��:"�E��A����ʦ���PC���P}�k�� ',��s^�����^��L��Y���Mf��rqT~�}��{�����O{�:��G9�KvwU����(���*��J��z��$����*��{5��@��׽w$�}�g��O�kг�)?�&�-�]�%�kkS�M��4���l���K�m��:
ŰIa�I�������?+��������%�;�ð���yHթ�e��o�_�O���w�A�����V�T�{	�v�h����I�8G�w_��k�h�Z|���wvnjQUUT�*�R��̒����%��~��]�W�ξ�ƕJ� �(��{�srI����I�ǉ9qh�Z��M ����� ���K�;&G��G�\p�N����7j���v�GC'M�i�2�,H4��9#��"&�n8��j�{��-v��GV�W���FF�&5"�z٠Z�Z�j�=èŖE��$nM�j�eKV��n��fn��#���U.%�1S)(�UJ��G9�ή��;���Dq#3v���[�Pk{13j��EQU5)ULҰ�"!n����؎�ݝա�}n���fg�g��I?�l�)#m�UU*�Z��v�p����<�Ov@y��<���t�A�2�Quճ�Z��J����k�c�S	�)lҲr��L:�6:����Mf���]t ,�h�h��l����4$�y:���g 4��	E"Wa�׍���wYs�;�/Zr'5Cv�ݑ�t�S/N���E#�rL^��\�3�5�v+��lA<d7���}��_2���Is��\�L���X:��l۳Y�X��i3Ŗ3ut�95$���$Rc���{�Z�Z�j�:��Ɖ0$�<�(���ՠ^���-v� �����V�HŎ87$MŠ^���-v� ����ՠy^X�s#x��lqŠZ�Z�[4]�@��ՠU��D�7��ɍH�޶h�V�{��@�ڴ]1#�|q-t*7�[��:�r������D�>��a4�Pe݇cq�JS�Z����[V̩j�n[_���s��ڰ1��x�0̗5f\̻�w�]��h�$b+",��\��k޻�N��rN�j߳���>��ꉨ�	i8�Z�� ��Հܶ����n�ƤjI��qh��h�V�o]��k�h�^��&�'�B)���$��-d��>�j ��ݼ�����.�X��Ǌ�)�]���η��z{W78.�aS��+@U�C3e�MŠ[�a�Z�Z����ՠy^X�sx6�nC@�ڴ��4]�@���@��ԉ�nb&a����h��$�-��V:ڪ����c�ĭ������P�5R2Hܚ�ՠ[�a�Z�Z�z��T_�e��d��I�o;����9���]�^̀ܶ���C��3wfЯ�Q����RnN�۹�WLN+s��ȱ�������$j��'$4]�@��W�Z�Z�v��c�HԐ�b�Š~W��-v�޻�j�;�]r"L	$O�)�k�h��h�V��^�@?rJ�9C��qh�L��\s?{ޯVW�^���RZ�yc�1̍�"m�I��k�h���]�@�t�h�D:&��Ls	��A�q���kd��r��y�wnT^�Tb�,���m��(���?����V���p�-v��5��,�5R28�z�ՠw�\4]�@��W�{�k�Yq<� �DRE�w�\4]�@��W�Z�Z��S�n48��ՠ~W��-v����yZ��R5$�G��>�� $�- ��&Ih�9��  �a�.E�8�N�������rv��NGz��O��ƹٖ�pn��nv�ʺ�i�S�T�a�tm���6��t���z�h�m���F��J��;;��YڻH6�X�ٵ�dscM���Վd�6�v�{s�֊�ܷ���'��-�u�A��ç^Hd�"JԔ�]�����8��w�k�q�oe�+���G8������"~{�����������ٻu��Gh*I��];d#�^ܕ���e'gVN_��㯙]#ur4f�U5T�T����V{)�`u�g�vC�o�@>�/���G䉸��K��"#�������׳`fN5`y<Q.���"&ؔ�h���׬�;�U�w�\4
�]H���dlr!� ���o�粅�}��ft�|}�$��L�E��$nRIwN��I,ʧ	ZI.�l�RH�U���p��,��u���,P\��W<��`�u����I�)�qѣ]j��)�tg��I��w�%�T�+I%���Itʴ�Y��~��U�xި���#q��1-I%���g9����<nr��zf���w���IwIq-�g��6�n�G�� ��5���$z�MI%�:�ߗ�ۮϱ�I%�ߏߒK�+�D8�'�B)
��Y��w�%���U���v��%���y?�~}�� ��߶bv��X��I,���$�[�w�$y�*�IfV5����v3�ͦ��^Z�V�����֌+�f�l��DuZ�KĴ��~ww�ﷷ���"&�)1��$�n���=e&���W��%ϥƵ$�|�R)1���$�%3Gz�G�2�b9�L�M��ޤ�v}�jI/��?~I/sSe�F�jFff��7m����r�~���Wv��A`�p��gz�G�2�$�}�+������T��U.�%Q�Neۄ�$���w�$z�MI%�:�ߒJ���)��n4UMD�I%���Itʴ�Y��w�%ϥƵ$��A%���X'L�ژ�=Vyѵ�	�ҶGJu����-ӛ�R`+�Y�l�����>���}�|�m��~?�RK')īI%���Id�w5H�I��E!5$�t�~�٘�\�\kRIzݧ��$z�MI$�$���0�LNH�������Z�K��OߒH����K�u_�$�W�;#�<dQ�Rd�I%���Itʴ�Y��w�'�@bVc(U�B#�2F	h-*�X�&��Hȣ����w5��]�m����E&7����p��$�YI�$�df\�ޤ�NS�V�K��;Ԓ�&S������01l=����ȋ]���!�&�����Y��E�Q$�:��ZI,�ƻԒ��q*�Iu�gz�G�2jI/��k�YP�db�I��%ϥ�W��9�L�^ݽ;Ԓ3kJ��Y��w�%_W��)�8�#�֤��n��RH�U���U7W��I'.�%ZI/NQ��ȣ�Ra	$?~I#�RjI.�ƻԒ��q*�[>���I9kmȇ �D�HMI%�:�ߒK�K�$�[�w�$y�*Ē�{�g��b	P%IT�B�B��*�"l��/��DЙ��Ut��K�$��kL���Ҏ���`D$$�$!$@�TC*��4:�ܤ���1�-VBؐ`ht�#����N�.��2b���A*B��`A L5�4-A ��� �(@dH1#�MB���!BF	`ԄRF2��`��+O@�W��b� 1�HЉ� �X��H-]G� �`у$X�X�4���F"H�� ���*@Q�p�� �#�>�"��`@"F,��a�Ӟ������          ��l�z   �I�       	 -� !MV�.2US���Zεkn�����Ste �˗d�ss�܃���z�j�f��ڊ*�pݘ�8���6<�1[Wi��(�
-�	n�M3+s,�-�c6�=W/T`۵hع]�m�FT�Gt�k8��	Լ��sB:6Bz��W$@܋��e�5�#�;n�Nʃ���ӄ)R�v�2Y�	�r��Y-��I�ooPZ\ft�Qf
��˵�$���$�O4�� U@�V��'[)QV��׶<9�Ӷ����T��Bn�a����2�(���j�mĞ:�bN��G$ZtV�#'�����]'[��LJR:]����K�+M�b�9�Zt']���T�ԏY�R�muUn�嗶r�ԭ��`�k�tT^�k+f�4Ѷ����i��Nv�3AlUtjj�ľn( ͠���\KjU��{2�]5[C�2A i#�^s�Ϗ�o�����<��v��&OQ�rnMU�H�-�Y&���q�A�ڧ�����ِZL 6�6�Kki6dlӡ�
��v	�4�DԷn�Ÿ�V�,4Qr��`dݍ`�N+�ݜ��U�D��U)Ү��XA��<���7ntJ��B�s�I�X��"�n�)���;��J�T�iL��XI���i��l���$��tপ�\�J�e����ܧ֪�N7.�i�sJٞ���n"wtvQ�Gn��l�t;��ڬ8�ؚ�\j��kmȆ]�mv�F�6z�kS��v �ejt�s��UP>Hnp�[8���,�;[m�:T�f�6������ll�	l���tF�n�;gdJ�e�Z�F�3abZ�#��0.œ�Ĥ˄��R-���pj�S��e�2�%g�e������TCb��k�����T�J�mT��mPG<b����c�m��n�_>s��>/'@C�.����Q�iJ
���AJ�Yq�J]j�  � %�A�t�b;A���<������w~|��` ���'x��=�I����[�k�����in{Y�	���k��k�/T4rŔl]6R��u��G�fj���	f�Z��F+^Ĺ�k��;mѪU�tAQ����u���[��q*��۲ð�����ݛ��z��ӄ-'V�v���>|�a�B�ʹ�7e��gXR�c�a�n�d`��z[�}Gkqs���^��.��g�pq��u�H��x'��ȕv�r��|������|jݓ��î��؉��Z@����Y��Y��SÒ&��U}>��I/��?~I%�,Z�K�u_�$��,uƜ���F�I���]n�ޤ��J�IfV5ޤ�,�ԒU�]H���267n�$������̬k�_DG&e�[�I/nޝ�I{��,�5R2H܋RIwN���Ŕ��I%���I/:t�$�}K8(�y21F��H�~I.].RI~�i��I/YbԒ]Ӫ��$�q�QXǃ�]!8�#�N:�i�v��e��v�F{Um�h�2��0���5jd�ݟ����I%�N���̬k�I,YN	��^�����G ��H~��K�X��a�DHȐ�e��wל��׹�kRI~�i����͵[���C�I"x܊����n���$�e8&�Iu�gz�K�X�$����(�A9"n/ߒK�S�m$�[�w�$��Ҵ��9șnޯ��}�9��ҹ�.�v~ ���ޡ#ΙV�K2���$�r�J��M��)��n�=��턹��1C��g�խ����!��Y,�n�i�$�M�L�ޤ��L�I%�X�z�Y9N%lr:�>���~~ R��D���դ�̬k�I,���$�[�w�$y�3~SZտ���S�h�5.j�.f^r�{��]�m�{��r�j�S.L�vf�Iw�U��IW��f��mncZ�K��;Ԓ<�i$�+�RO���"I/>�T��Q�)0���$�χI$���+�Ib�pM���v��$�tJ�Q��;>�s.��tvۭ�a�#�����<soj%r�y��[1Ud�b�i$�+�RH��j�$�[�w�$�)ũ$�䕰qF8'$M���Iv�I%���I,�t�$�ec]�I	��^$�ldQ�RdSRI~�i��I.�bԒ]Ӫ��$�;�MI%_�E"������$�t�jI.��~��G��Ui(��DB]n�ޤ�:U ��*�R2H܋RIwN��䒫��jI/��?~I%�,Z�K��"��	(��˱D�=�٭�Wn�m	��m�˸+�.���
ӱ�����Ӊ5�G�������	.�l�RIfS�i$�+�RI�L�/ȉ	��8MI%�ݧ��g�cm+g�jI+e�~��Ur���KϭS$�I�I!��I.�bԒ]Ӫ��$��)5$��v��$�n�\�(�I�5J����̬k�I&�����]n�ޤ��-I$�ح��<$��&���$�ʖ��Iu�gz�K2�+I%�X�{m����y:y��y;��� 6�m
��W�؎v%{n�I�s�2\I9��h�m�v��]���gF��6湹q�v��yneɧ�z�<[����m�.�p���sϭ�\�f���.��i�&�nud3eX]<� �l�n�zܧQ�\�6ӷC���k/\t�� pWc<�o�v��x�C;W��e1�����$�m��\d�k<�$4,W>a7Z��8y�w{�=��8���4�e*#�\rM��āc�[�R:9�pV�.răH�5rԹ�+��� ����� fS�i$�+��ȏzRZ�N���[,G��E�S�b�����߱�����I�z�Ԓ��v��L�<ڨ�SQ�#$��@�}V���٠~�S@�t����w����&)"�9z���l�� �9h���U�DHH�FH���e4wJhϪ�;�Z�]�iY�&8��l�1�Z.���(���ͷ���s����2�p��]=&,p�)$JL!$����M��Zy�^���M��"� �D�� �9jW�^��W��#�و�� =�L��"9ăGv��S��T��MZ<�߱��7�@7�Z ��vLnH�ȣm�#�?[)�{�S@̜j�y	�-ٰ51J�����dJ��=�L�7����%ńܲ�z�����̙���P�H�2������={���}\a4�P�n�Ė�5��R2H�4s��V��YM�Қ�k���&F(�1I��jٽ�#��絥��֖�q� �`�)��	���@��S@�t��3�?���k��\���Z�8I�%&���=�)�uv��կC����W���@�_��ȤiH�7"��:d��}�& �-��p]�7���Cr��tkW8�7��.e���]n����M��T�nL��kQ=�Ha���1 �Iho`�s$� �d�㍈�6�R=��h��:�V��jנU�:�9�Ddlm�ho`�s$�7�- �Ih�T
%�R�eUIUS4Xo#���{[��>�r��I�u���芄Q? hAC6��3eo���P�QP��X̤Ձ�[V|�9mXȈ�t�G�K��٠\͋(��.��X�ss�@�حknwF�h�:V�iw:�8��,�K�=��`wΙ`c�Ձ��MX�SǤ�I ��)�@��)�uv���U�uv�����N1H�<ݽ� �onZ�Z���[	x)���@�tUh��h�e4]���5rL�8�Ej-�v�����˺������?>o�   5&�6�	N�][�=e�t�WIt[˞�v��4q����tX��X�$Ʉ�`��l�E�uJ�z�M �A4of�琶�t���4I��،X�כ(����l�*��K<�T0�TՎ,�֍��\�]a�����(����mL�K�.xǩ����]���@p�gm�v�՞+Sz�M�*K6\�mc���Gќ��w�{���_���	���j�rN�㒅7��/�ʚ�y�.y�]�ӎ� 2�cV�r��bh�.�e4]���ڴw(�j6�d��hs�����'d������.x��<��(�2G����/��@��)�U�^�~�ˊa2BF��@��Z��� 9��h�^Vi$RH)0����?z�hwW�{��V����9��=�	+��T�7mvSARON��َѺ�GQ#(\����|���WH�*�hgqR<�V�m��߿�����U�z�����S@/![	xG��]eˬ�䟾�/n��|�@P��TU{ك�P���}& 	�*L�8�Ej-�ڴ޲�]���ս�"�G� ؘ)t� ����f :=����"�6܌�7��z��@��M������6��I1L�,P\�١	:��I��Y���܅"�Ĳ9�ͷRZM?�dCɊb�$q��սץ,y�>�G#�@�ǹy�Ll*������I�=zS@�����ֽ����w�O�BI&NHh����}w��ٴG�}� u�D�e���X���"Q�cd�M�Hlp?0_�� �F�Db�&f�1�Hȉ?�TKaqx������Xb�@�a!, �B���@a�2p�AV �I𫠿
��C��@`��T���D�!QW���] �j�=@֕ m\@?"�V����k?k�5��>��ٹ'�|�$N3���Ȥ4^���ʽץ4޲�y
�H��q8�q��ʽץ4޲�/Z�m����w߿~v3��M�P#=j��m�]h¾�w�`r*�n�,Վ�f�]Y"q��64�����?Wj�9zנuv��UDZH�d!�}2K@;�1 �I���������Ԍ�'��ֽ���ץ4�ڴ�k���&)�4L��@9�f :=��Z���/{��ez�8O.)��	"$���)�~�ՠr��@��o@����I�nU�����U��qtn�k��i��;N��9fqe��QWvL@��	��V��ֽ���ץ4��Y"q���<m�Šr��@��o@��M�v� ��l$Q�9$R(�z�&b�� >�%����>�2�"q���r7��b��h����9zנuv��UDZ8��b�UE��-�b!�n�@{;�6�Wf�A>A��
Ab�$"�`E��`T��빙�����35� ��]��k�ˤF�'6[u�Ol�úO!ҷfC�܋�PI�b��$�I���h/N�#gk��ѽ�[:yKc�����o��c��� n�R��;`�0ƶyq==�ul����u)�d۵O*^b2��79G��6����ٻv꽦�nk��ӭ�F��en�n:�)���^Ew,R"5�U���*�(�FΧ�7n��E��������{���̥�����k�������&��s�lDueն�Y@Y�+)lsu,�:A��o�����	m��G�@wd����ߋ�fV��Q�d�=��f��Қ��Z/Z��(�\S	�4L��4^�@wd��w�b[y5 �2���AI�&�{�ՠr��@��٠z���y�Y�1Ix��@w�b[y5���%�$�Fe���Og��uwߗ�r8��w=��������E-\b����s���YD+E�Jپ��rg�@t{vIh}& ����!��٫c�'����뿻�?{�;͎s�vn�ڰ<�vl�%Հ`�ɧ�26�B��=�j�9zנU���=zS@�,B�rF�jFF��A��I���j��}�7h�.x��y1LQ�d�=��f��Қ��Z/Z�\b*�0x��ĦH=t"�d�x]�R�'V�5H=��suk.Pn\r<�pȉ	&Hܚ�Jh�h�k�*�vh��y�Ȥ�R`���$�x�%��PI�@^u��H�)#OcqhϪ�*��w7CJi"D ���e4�l��V�E�E"rE�Ko&�>�`�;��x��̹&H��8�r(���e4�l�;�U�Uˬ�-|6��LN@DC��K��	�>������k\Cs�괛n y�D��bSi�Hhz٠w>�@��Y�~�S@�T��5R3k/7P㖀���@}&� >�P�w�2���1F��Z\�����޶hϪ�\�tȉ	%Jj�6�oK y�Vd�V�F۝��3�1ݪl�;=J���RH)(�� >�P㖀�-�@}&��'���6����7%��t��u��|��%�{@�lsI	sr\�Wd�7P���NM��Z溽���޶h�B��2'$�	���uz�e4�l�;�U��7rL����I#�8���hz٠w>�@��W�U�:�9�Ddm��!�w��@�}V�y��@�l��֨+�!FF��qhϪ�*��h�n�~�{w$�� �����33333 l  ���b���*'a7H���F�-��<R��ܚ1l�f79���V�w=�R��Rnm۵������o��֧��$�8��)�[�]�!��1�1��.�izv�k��Ӹ��UR6�ù�����	Ϟ.5j�z@��GA�0uIh˄4�Z��l�m�WD����luq�͑7Vb{(6۰�&��X+�.��-�:��aG�߽��|�o� |0\���+�Y�v�G9{u�ó�]v�p����v�]��n�cY��3�j�Gͷ��}Vrڰ3�ڰ�Հy��UEQU(�����:�2��q#2wU�ۿ-��f�ԑ�~>x�r)$�	�����h�V���^�k�hϱ��H�Ix��C�����~{�6rڰ��/mn� �4%�T��RF���@��o@�ڴ�ڴ]�@�b�ėُ�#�PrLC@�rс�.9&�d�ɶխ�(GF�p^�vs�$�wt���j���������$���|��7-���u�ճ`jb�SP�"*gWD�dܓ�u���4QW,�u����8���e�G9	ڠQ;EH���4�Z�?�ZWUz�S@��)�{��P�b�	�Zg�b�Ml��ZX�Xls��kuXE�'�)�$$a"�@��h��̈�m��7guX��3`b�&RtR�]î���P��hnۋ\k�h���K�7D�;8��_���v��ݽ��)�\������$�<s1$� c�����4���k�o�ٙ��[ٛwkK�t��s��$���b�N89$PMŠuw��l��3�?���(� h�M_����;~��ܒw�k]$���qȣ����?����h�M,��}��qc��6�H7I��J�3*I�,y�,���se����ߛ�/���wp�!����c�x�U-k��cr�{p��b�aI��\��VWq���wfcش=�b���F���|�s�ށm��=�)�{��P�)��UMM��No�Dr#興��>WŁ��?ƁWuz�w�2d��"%*���,��,�r""��́�Z����x�r)$�	����?�/ｿM�={�krO�k��nJ"� ��������h]�G!#D�'�ȥY�l�s���Ml�ͭ,��4���p�G1cO�c�����zL�l<�5�M/Gg�7�*s7&[�i�d�ܽ2�q��@N��6�����+~z�տ�L�H�RG"n(��L����"9�1�_�w�=��f����Z�n�SP�B*fT�TX�ZXf9��G!,r�f������b�K��U%L�U3E���s�e�����<��X}Ȉ��������ET
��t77���G ;�� ��nI���H�� $R6I�Q�(�Z�a��lO�9��(��2)e�/�Tt��!�
hȲP_�Ij���Ytb�~A����Q ��b~�	1VBD'xH�O���aXX!"FƱG)CJD�����g�
�m:) t0��U���&�"��"����#e!��j�?��WHH�cH�0"�?"���������          -��`  ۰       ��  [T�u���q�[�n�����t�LS��1�,g�N����q[v�Ԫ���ؐ�=�]�M��10r�J�WAǚ/�ۮm��X�9n�{Rl����а�N���6�VfR�����U�F�`}�k*c�"T�"S]c�tV�;�jkes�Q���59M����A㚬n�f^�DmY"湶�q����+ɳ��(C�-HQɚ	V�F��l��M$�  *յ��#�%U����sM̅�ë����v�����v{i�ۋNGx�`��7r�I�;;8-�pA����×Iiv-]��.5q��[��;�.$ōa���A�L��EC�� c�ۈ��<�O+P��r�ivY8��UU� ���i���ݭ�lUA75����][l�'V�Iu!�I�J�Z��Qܠ���0�$�x�eX�:�o"�Z����d���]�p�2F�;L����A1�U�u�4"��m� �UUU*�*��K��d��#U�����974��5�=�^3<�v��ŉK�]�rlT�U�i�[�U�K�
��IW@l�T���f�F�Ƅ	�h2��嶩��Ҟ�`��f0ݔ8#<����V5V�1N)54qud�'m)p'C����E^��2��ڊd�+]E<�Y&{b��e��r:1\s(��73N�!���+���&��:Wr2
�1�'��sp�V�`wB�c��q4t� ���S��ѱҪ�z��Ob�h+�YV�j%[�

jXݸ�H:�<�KÙ�P��ڷ=[��KW)�KN�c1��	'Rյ8©���l���@�.�T��앫�55UEY�)htW�Z�̹����@����-�B��T�d�g�MB��3���{%��n$�������)����l�Tt�
�l��v���UX /
 �AC�D�PТ?
 ��`���g��������ne�0 m�[-^�е�wM�Set�=��0jV���]n��KZS��N���&S��9���i/b���l����0��:�n�m�*�bD^|֌=	R���-��m����t;��[�..ۦcJNYÒ�i�[Wn���㇗`�*��q��ݺʆK���nW����.��5�ZG��<�f֭��w�v�B�)K��ڴ��VQ�eѶknj=B��gC�Ⱥ��[�s���w�|�'��L���D����}���YM���9��r�̀�\l��5J��UT�� >�@;�1���@tqV���������$h�DۑHhw�47�-��H�@C,���mƤ�A�����������nh�����?�}��@>���I	#J(�I�����t� �����e�?���q��y犌P���b ��%�`�zc��(�J/k5c����{Hm��f�����o����z��k@�빠~����&5$��4^���B?�GJ� �js5�kp��Ł����9�r!#�>��B��8�����=z�i��J�>4
���'AL�!#	�7��3?�k�ŀۭ,^nl>��vl���Ȥ�R`4ԙ�wt���W�|�W|���]���%̬�@�:�]�bр���c��y�z3F��Y9mset�TRE1�H�$��"��9zנ}�_�׳iȖ%�b}�����?�j%�b{����r%�bX����Vk.j�Y����5s5��Kı;���fӑ,K�����"X�%����6��bX�'u���� ؖ%�}��^3�̶fk33.kY�ND�,K�w�6��bX�'{�p�r%�ʈASS
v�ț��}�kiȖ%�bw]���ND�,K��ۢ{SWF\,�kF��6��bY�)Q=�~6��bX�'����m9ı,N��kٴ�Kı>�}�iȖ%�b}��ja��f�3�a��Kı;���m9ı,N��kٴ�Kı>�}�iȖ%�bw���"X�%����֬��˚,.��F��7h�՛�c����E�ɹ
EI�$�h�g�ض=��]��5m3������X�'u����r%�bX�{���Kı;���ӑ,K������Kı?jw��<\0̙�&ff�6��bX�'��m9ı,N����Kı;���m9ı,K���m9�T�Kݟ��Mrk2�fK�I.��"X�%��{��ӑ,K������Kı/�{ٴ�Kı>�}���{��7��￿~}.gRj�Z+m9ı,N��{[ND�,K����ND�,K�w�6��bXA�D��W������Kı/��r}�d�,���~oq����=�fӑ,K�����"X�%���~�ND�,K����ӑ,K��;��������3e�T�3\�dhǳ��W�p��vy����Mz&e����-���p-����2�f��Kı;���ND�,K���6��bX�'u����"X�%�{�ͧ"X�%��x��=���.f��Z�ND�,K���6���E5Q,Ok����r%�bX������r%�bX�{���Kı>��x�j᫖f�5�5��ND�,K����ӑ,KĿ��fӑ,E�,O��p�r%�bX��w��Kı?}:͞.a5�kRfI��m9ı,K���m9ı,O��p�r%�bX��w��K�A�;���m9ı,Oڝ�.�3&f����ͧ"X�%����ND�,K���6��bX�'u����"X�%�{�ͧ"X�%�t�<��y����;Ο�?@ �  l9��v�k���)e�ekc��� �p�#>ܔV!^��h뮮vg9�dZv܍��WJY�W>dj-��m�t�έ��a��6�h�N��,Z��Ed�!�6�놡�Ev����t,��d$�<՝��VFp�v3ϴ��
�a6ڦ��ے�n���@�t����m�7[m���%�Ϫ��:7�9�q%h�8�1�M6Yn��@ ��3�˳\�.�u���)6�,1"<h��9$ɜa���EƲ�k��Ԙ
�x^�l�U���|�7���%����6��bX�'u����"X�%�{�͇� P?D�K�����m>��g�g�g�����!���.{�}D�,K����Ӑ�D#���b_����iȖ%�bw���6��bX�'{�si� �bX�������̺�j�f�M\�m9ı,K���m9ı,O��p�r%�-���؛�H�o�����H��צ�kZճZֵ5u��$���}���ӑ,K���{�ND�,K����ӑ,K��_{��r%�bX�׎�ښ�2�fkZ5�a��Kı>���ӑ,K���{[ND�,K�}�kiȖ%�b}���ӑ,��ow����>�z0�Xkp�������cc�9�t�뮢^ERi�]b��8��噭M�ͧ"X�%��}�kiȖ%�b}���m9ı,O��p��_�5ı;���m9ı,O�<͟�̓XfjL�3Y��"X�%�������*ı>�}�iȖ%�b}����Kı;���m9ı,O�e�tx�a�34e��kiȖ%�b}���ӑ,K������Kı;���m9ı,O��}��"X�%���/��5�s3%�$��d�r%�`؟���6��bX�'���[ND�,K�}�kiȖ%�b{�o�iȖ%�b~��_��I��n��=ߛ�oq���{]ﵴ�Kİ~������bX�'���6��bX�'ｿM�"X�%�����e�b����)���\�>n���Od�e�nS��蓞�1wl[�9�k5c��rj�k��%�bX��}���"X�%�ｿM�"X�%���o�iȖ%�b{]ﵴ�Kı/��k�a�����f��k3[ND�,K�{~�NC�B:���'�����r%�bX�������Kı>��������j%��������z.4���{�7���{������M�"X�%��w��ӑ,����
9"o[�涜�bX�'���6��bX�'ݘΞ�\5r�֦�\ɴ�Kı=����r%�bX�k��[ND�,K�{~�ND�,������6��bX�'}?���\0���2L�kiȖ%�b}���m9ı,}��m9ı,O�{~�ND�,K��}��"X�%�������<[�f�:AG��]�֧��tK�6N�v�(�M۪�a�9���B������S?=ߛ�oq���ߦӑ,K������Kı=����r%�bX�k��[ND�,K��S�乗32\�K��M�"X�%���o�i��MD�?��kiȖ%�bw]�����bX�'���6�������w������)Ԛ�V譴�Kı?��kiȖ%�b}���m9ı,O}��m9ı,O�{~�=ߛ�oq����r}i�d�,���"X����ﵴ�Kı=����Kı?}��m9İ'� _;Sr'�?����"X�%�~����Tl�o|��Y�Y�Y�~�~��=ND�,K��ߦӑ,K����kiȖ%�b}���m9ı,O}����j��p�l%�\��/�.�V��b;6n{\�K���Dz{/��Ҫ�M�"X�%���o�iȖ%�b{]ﵴ�Kı>������bX�'���6��bX�'���)���W,�jkW2m9ı,Ok�����bX�'����ӑ,K���ߦӑ,K������O�D����'}?����a�35&d���ӑ,K����m9ı,O}��m9��!������6��bX�'����m9ı,O�e�tx�a�34e��kiȖ%�b{�o�iȖ%�b~����r%�bX��{�m9İ?�P���￵��Kı<x���.e�̗0��5�iȖ%�b~����r%�bXG�=��m?D�,K�￵��Kı=����Kı;��y�O'�wyӿ}����`�`�W;���n��z��e3�GbӶnK-��v���i�ͼ�p�κ���%e-��I����ٙ�4G�g�۶f�3҃'n�ֺn9M��$YβbNHq�����
��V��v�N���R�o]B��Lq��l�kS��Z�t���f����-Ė\��6l�QHf�X��=��ζ+�z�d����ǃ$>��_�{��C�E��^,۳sN��tv��F��%����`7��X�W%�x�.�s'��Kı?��kiȖ%�b}���m9ı,O}��m9ı,O�{~�ND�,K��M_ff�W5�����W3[ND�,K�}�ki�
�Q5������ӑ,K������ND�,K��}��"ؖ%�}��^3�̷.fkYffkiȖ%�b{�o�iȖ%�b~����r%�bX��{�m9ı,O��}��"X�%��x��}���.f��Z�ND�,K��ߦӑ,K������Kı>������bX%����ND�,K��$�����Y��ѫ�6��bX�'u����"X�%���ﵴ�Kı>�}�iȖ%�b~����r%�bX�k�Y��}���ԃŜ��n[�^�q<��Wn灺]���s�+���::_|��O{ޮvq�$f�r%�bX�k��[ND�,K�w�6��bX�'ｿM��3�MD�,Ok����r%�bX�w/����a�34fe�fӑ,K�����!W���������bk�ߦӑ,K������r%�bX��}��r%�bX��J{\�2�f[��ə�m9ı,O���m9ı,N��{[ND�Vı/��ٴ�Kı>�}�iȖ<oq��~��ѝOMagEo����7�������Kı/��ٴ�Kı>�}�iȖ%�)b}���i�����~�����+`���%�bX��}��r%�bX"1����O�,K�ｿ��Kı;���m9ı,K�ŷ��50����j\r�h����
m��{h�vJ���״�y�|���cox�Z�g����u�u�'��m9ı,O���m9ı,N��{[ND�,K�｛ND�,x���߯\�Eƕ�n�����{��'���6���@�MD�=��kiȖ%�b_����ND�,K�w�6��bX�'}0��&fYfkSF�d�r%�bX�������bX�%��{6��cE�qH�#`�X����d!(��XlCF)7u�DP�R)]�W�8���Ut���&����@�7�сF	a%�%"�X�0%�)!�Q�`F� @�R� DX�#u
��
��k®U� �� @�4CP���H��c� %A����uN�"A#IUaE4k��>آ�8:EC����P��t|�E�D?��W�C����br'����ӑ,K���ߦӑ,K����6x�a�35&d���ӑ,KP�/��ٴ�Kı>�}�iȖ%�b}���iȖ%�bw_{��r%�bX����B��p�2fh�ˬͧ"X�%����ND�,K� }�M��%�b{]���ӑ,KĿ��f����{��7������ֹ��MY3:%��I�@uv�q$ۙ�e�j���m�ss����K�s3-��d��6��bX�'���6��bX�'u����"X�%�w�͈	Ȗ%�b}���ӑ,K�����3��<Ί�=ߛ�oq���w_{��r%�bX��}��r%�bX�{���Kı>�w��Uı�{�߿v�3*�DX)�����{��������r%�bX�{���Kı>�w��Kı;���m9ı�<����o�8�b3{�}O:�:��>�}�iȖ%�b}���iȖ%�bw_{��r%�``��ڔ~xi7bk�����Kı=��/�5u�ᩚ֍kXm9ı,O���m9ı,N��{[ND�,K���kiȖ%�b}���ӑ,K��T����<g�&�㞭شXX���/S%�`Rs�n��b)��;aߝ����|�=���,�jkW2m?D�,K�������bX�'�w��ӑ,K�����"X�%��{�M�"X�%����vz�0��5&jL�kiȖ%�b~�}�m9ı>�}�iȖ%�b}���iȖ%�bw_{��r%�bX����B��p�2fh�e�kiȖ%�b}���ӑ,K���ߦӑ,lK����ӑ,K������r%�bX��H{\�2�%��d��6��bY�Q;�s�m9ı,Ok����r%�bX���{[ND�,K�w�6��bX�=��~����gEo����7���'u����"X�%�����������X�%���p�r%�bX�w���K<�<�<��<�;�?}�� �-�*�W��v5��9��Yz�]��ܖ��kgy���RΉ�j�
��jjA��NB/qjsW)�`��dQ�݈��<��۝&�Ѱ�D�.�88�=��#��ٖ*˹�v�n����,���r��O[t��6�Q��;�������s�ZF�����\V0����5vܵǆxɪ'ӇT3�zryۭ�����{����m��k�]��l;WX���5<�.�1�]�����u�a�s���w{������kZ&ff�Ks5��%�bX������Kı>�}�iȖ%�b}���ӑ,K������Kı/��{&�ffe�s3Z̙��ӑ,K�����"X�%��{�ND�,K����ӑ,K���w�iȟ��E�MOq���������عҼ��=ߛ�oq������Kı;���m9�����w=�v��bX�'���iȖ%�b}鄞�30��3Z�5u�ӑ,K�;���m9ı,O�g}v��bX�'��m9ı,O�w�6��bX�'�]��3$��5%�f�[ND�,K���]�"X�%��}���ӑ,K���ߦӑ,K������Kı>�ޚ��kEцZ\ɚ��"�[�]q�cu���P��g3��Mqu���,.�.fL���Yv��bX�'��m9ı,O���m9ı,N��{[ND�,K��v��bX�%��C�2�]k2\̶ffND�,K��~�NB(�� �MD�;���m9ı,O��z�9ı,O���m9ı,Ow/�u��)��n�f�k2m9ı,N��{[ND�,K��v��b*�%����M�"X�%��}�M�"X�%�{�I��k5�h����-��ӑ,K����]�"X�%����M�"X�%��}�M�"X�(�bw_{��r%�bX����d�L�fK�35��\˴�Kı=�{�iȖ%�a�￹�6��X�%���{�[ND�,K��v��bX�%�},��u�\U��L��qY��%���\�pvTuH��i�]I�x��Nu*�]�"X�%��}�M�"X�%��w��ӑ,K����]�"X�%��޻ND�,K�L$����,�jkWY�iȖ%�b{]ﵴ�Kı>�{�iȖ%�b{���ӑ,K���ߦӐBı,O�<��˙&��Ԛ�f�[ND�,K��v��bX�'��z�9��j&�k�ߦӑ,K����kiȖ%�b}���Ip�2fh�̺˴�K��g�v��bX�'���6��bX�'���[ND�,騝����ӑ,KĿ��!��.eֳ%��s.e�r%�bX�w���r%�bX��{�m9ı,O����r%�bX��=��Kı?�S��`?��Vѝq6�)�F��G@uͷ`W']3o����t�F�/�w��{sCp[�Y��̛O�X�%��k����ӑ,K����]�"X�%��޻ND�,K��~�ND�,K��I��k5�h����-��ӑ,K����]� ��bX��=��Kı>���Kı=����r'����b_����ə��r�f����v��bX�'�s���9ı,O���m9�K����kiȖ%�b}���ӑ,K���N����\���ֵ�̻ND�,K��~�ND�,K��}��"X�%��s޻ND�,/�V<C���(~�O�����r%�bX��a'����,ˣZ�̛ND�,K�ﹴ�Kı~�w�iȖ%�b{���ӑ,K���o�iȖ%�b}��o�y�0�ᮻBL�nѳ����,��]&�;:9/k�GMٌ�V�l��]5�������ow���]�"X�%��޻ND�,K�｛��j%�b{���r%�bX��������d�љ�s.ӑ,K����]�"X�%�w�ͧ"X�%�����r%�bX�w;��H,P�I��h�՗D֦��bn	 ��}�ؒ	"wﻉ�$��w;��Kı=�{�iȖ%�b{���jfh�̷F�Z˙�ND�,K�ﹴ�Kı>�w�iȖ%�b{���ӑ,K,K���m9ı,K�'�Y�ֵ�ffj䙙��Kı>�{�iȖ%�b{���ӑ,KĿw�ͧ"X�%�����r%�bX�P�;�;����� A� i�nʁ�+�MW;am��>q�Ek�c�]���e;���:��q�\I'd�Ur��6s���"=b9J�l�W�I������p��x疥�)x�4�\��i��Ua&s]O*:�\B��� 7N��D=vl�1uu�c�kzҜ��ɬ�g��Y�4빺3�َ�^��%�j�1�I<͗ �8�m��e��+����3�9�Gbf�N�;*���ى�t�؅V�3ś/l��;��}ޠ�Ҩؙ����%�b{��]�"X�%�{���ND�,K��}��"X�%�����#�!�r�����%M*�J���f]�"X�%�{���ND�,K��}��"X�%����kiȖ%�b{���ӐD�,K���%���]e�tf��6��bX�'���[ND�,K�{��ӑ,�@!��������ND�,K���ٴ�Kı>��7�.d��3Rk	��m9ĳ�*��w;����"X�%������ND�,K����ND�,K��}��"X�%��g�.�%�ə�Y�Z�m9ı,O}���r%�bX����r%�bX��{�m9ı,O�����"X�%���q����=���az�-��2��ژ�${X��ʫv���P�'�w{�]���Bk	���\˴�Kı/�{ٴ�Kı=����r%�bX�k�{[ND�,K�g�v��bX�'�����L�����kYs3iȖ%�b{]ﵴ�:5Q,N�涜�bX�'��z�9ı,K���m9ı,K��u~��j�K?=ߛ�oq���_�߮ӑ,K����]�"X��MD����m9ı,O�{���r%�bX���_��L�*Z�?=ߛ�oq����{ &�w��iȖ%�b^���6��bX�'���[ND�,K�}�kiȖ{��7�������#b�������KĿ}�fӑ,K��b��ki�%�bX������Kı>�w鷿7���{����oܧ�F�0̽xi{>^��\�����Cs�zcb�]�mW@�M_=ߛ�oq���~�߿u��Kı>������bX�'���6��bX�%��{6��bX�'�Y��̓Y�5%�f�[ND�,K�}�kiȍ�bX�{���r%�bX����r%�bX�������bX�'ݞ����3&f�f]k5��Kı>�w��Kı/�{ٴ�K+�$X(D��R(2*B ���H�"����LFQ?�DȞ׿��ӑ,K��������bX�%��C�2�]]a32ٙ��ND�,K�޻ND�,K����ӑ,K��_{��r%�bX�{���~oq������?~���Vf�<r%�bX�������bX��G����m?D�,K�����r%�bX�}���r%�bX���Mj��˙	JLN��Ȅv�3�_(�:�s���ζ懖��t�-��W��%������7���x�_{��r%�bX�{���r%�bX�}���Ȗ%�bw_{��r%�b�>�\��HEK]�~{�7���x�>�w��Kı>�=��Kı;���m9ı,O�����"X�<ow��o׏�Gj�yk|�~oq��K�޻ND�,K����ӑ,@��_{��r%�bX�{���r%�bX�za'�&f��eѭ\̻ND�,K��{6��bX�'����ӑ,K���ߦӑ,K���88��������ND�,K�O�l�u��d�IrL�fӑ,K��_{��r%�bX�{���r%�bX�}���r%�bX��{ٴ�Kı;����)��D&�J�u�V���ҝ�A䛵�C�����j[:���!�f�9ı,O���m9ı,O��z�9ı,K߽�ڨ�%�bX�k�{[ND�,K���2��	��噬�ND�,K�޻ND�,K��{6��bX�'����ӑ,K���ߦӑlK��r��Y���5�n�f�fe�r%�bX��{ٴ�Kı>�w�iȖ%�b}���iȖ%�b~�{�iȖ%�b_vN�^�[�5�˚�36��bY��5�߿�ӑ,K�����6��bX�'��v��bX�%�{���ND�,K�����e���������{��7��������"X�%����]�"X�%�{���ND�,K��}v��bX�&�H>�! ���?M�d�E���CZ৘�b&�G�H��KJ�G :�"F.4(@ДK(>M��Є�B��HB5�B0�%cV�B4+D�F:��$�����H ��9��ڼ�ffffffff        [A��  ��        H� UA\��:��U��U�M�x�v��T�T��Λ��3D��IzY����&0��!\v��Rqv�ʽ;Z�l::�{;V�!uz;]s1s��Ӹ�m�!ض�*'N�>͕����yؓ���9$���6R4��ť�#=qš�Gq$����QD�7U�gk�Ύ��m�y���a6SDz��Ɖ��Ɖ�؝q�N��l3���Y����N�t ��nn���ki]�[i��6  �]7\�P�T�������vgt��f2'n�*fI�:���*4�v�[ ��y&ݞ���'���盫�#�IH���6W\�Uv�vQ�!0�<q4���m���,��05�j���ԦT1%-�n��
9�(������[lcb����#E��P����I��l�����m�f��VtdȰ�Ѝd�m�^� 
�
��[U@����n����dwe��[���ə+��@<��[�Di�Hi�Rn	g���3�*@j���S#��k���{�H+!5 !���m���zy5[*�I��a����M��Μm�[��+aC:�I�y3Q���&�*�$���0W6Qa���h�e��(q)n9���6\̹x��#`j�VV�W����-�U|ӳ��$9��l�B�pӍ�!'�F�2�����D\[=qu�c��g���K7OQ�sS�Nt��Eu�d�3�eʆ����ܒ���k��Uy`��6i�f���.ђ)�uۄݺJ�QH�U�3�Zږ�U���Qԫq�IP�;5�J��l�MK��j��^e�j�g���t�$�S��F���UԄ�]�^y6Ԓ��'U��G#Yt��۶�n�حPS�i��ɷ9���ZvV���i�x� m�'V�1�r���Ɇ۷
s.����`uDg����,�&����`[m��m������?%DM��J'���m� ��B �)�#���m*������  �߽�� ` m�mt]H�+��T�N���n��󪙹ݴ�à&�MǇS^��Ս$3�s��5����7V�n\\7�Ƚ#�Α*�xx�ջc��RY5��.f�+&5��J%+/c������C���!g���:�ܝ=���l�W��q���:�-ɒ�,M����,���/r�����V�}e�"ym�*��l��;Z���)m�ڣu�p�1r<b��ǎM˸��t-#�n{7BI���G����s�mM���bX�'����9ı,K߽��r%�bX�w;��"�'蚉bX�����ӑ,K���a'������jeѭ\̻ND�,K��{6��bX�'����9ı,O���m9ı,O��z�9@lK����<\�k2kR\�5���Kı>�w�iȖ%�b}���iȖ%�b~�{�iȖ%�b^��fӑ,K����g���sE��f]�"X�%����M�"X�%����]�"X�%�{���ND�,@V����]�"X�%�{���2�]]a32ܳ5�iȖ%�b~�{�iȖ%�b_���iȖ%�b}��ӑ,K���ߦӑ,K����z..���m��N��tv��m��]ƺݵ��n�jgL��#l?;��{�|��әn�f���v��bX�%��{6��bX�'����9ı,O���l?�~���%������9ı,K����?�!�B*�����{��7���}�m9?�O��a��O�,O}�M�"X�%�����ӑ,KĿ��f��w���7���{������,�T�əv��bX�'���6��bX�'��z�9ı,K���m9ı,O����r%�bX�׎��j��Y��f��3Y6��bX�'��z�9ı,K���m9ı,O����r%�b*�'���6��bX�'ޘI�I�����[���e�r%�bX��}��r%�bX�w=��Kı>�w��Kı>�{�iȖ%�b=����K�5%�j���w=x�wۮ'���^�n\i��s�+�t+���󻻯��{�鉴���q,K�����9ı,O���m9ı,O����r%�bX��}��r%�bX�vz�z�.fe�35��ND�,K��~�ND�,K��v��bX�%��{6��bX�'��z�9ı/}�Ohˬ���fe�3Y6��bX�'��z�9ı,K���m9����HQJE"@dd��CB��]��ȝ�}��Kı?w���r%�bX���n����32]�a32�9ı,O��}��"X�%��s޻ND�,K��ߦӑ,K�D!������ӑ,KĿzj�Z��[��u��e�f���bX�'��z�9ı,O�{~�ND�,K��v��bX�'����ӑ,KĿ|[|��u��g\t���E�*r2�n���p��Q�r��o���9�e����*W���G!������;����9�9��g�_�-�Ϟ}i��7	4d��/c��-��t��"!#4x��dq"'��"�9u���j�?z�h�j�?x�苊L�`�[��y%�>�@s�-{�C~����R��@�|���ɒE)#qh�e4s�h^��+��^J�ػuo$B�@��M�1�]�[K�.��e�!���'LK�s��c'�L���/c��㝎s��ͭ,FT�qG�H'�9��h^������;ٵ������s�DL�}����hU5S5��jl�ߦ��2Ϣ9I���_��~�\v���Ʉq�l/fޖ��V��͆��DK���*�����Q��F�#���v��������'����$���f䏕H) +1���XDX@��}���  6���K#m��z�k�b�l�����l�:CVr��6xzӫeI���N�N�)�9���]=�j�>'�7lI^�lf�s�a���m{n�`�Un[%��
�{Y��$���͹2��1�H�p،Z9j����z�`�;��u�^<]#�����f��eYf8ϲ�4$k��6Fx�v���s�`�B[�=Y��z4{�5/;T���]-���<�1NS]v[cC�l��e��E������H�;Y�Z��K�GHH���rO���<�9�<�������z��g؜ �$9��z��ڴ�h�נ{���ɒE)u6������؈��I��6-{:�ì�71I��@�;V�y�����r!<��`j1�٤��<��#�@=z��g�?���l��;�ՠ�$�c.)��bS >�ɵu�3��A��*qQ�l��+n�:[����pQȜ�ҊI�y^�@�;V����܈�r:��{V�Kbv��S%MVk0����~�{w ?�S�PP�����@/��@�^����\Q�$���SE���Հw�>�r9�-{6���@�<BIm�LmI�z��\s�K@>�-�Y�jU�TMQ2
&����x����9ȇ������@=z�޴mj��!HD�E�U�0���۝��^y��g\�:�Mqu��ݧ�D�2d�G�D�z��4�h�hW����N(��$JdUJ��Kj��Dr>�G92����ߦ��XU�T{��%�I�aZ��w7$�{�u���? �O	��#����Vs�X����sB��SQR�*�����Y:�l�F�=-� ��4�J�mF��a$zz�- �$���@u�1 G2i��cU���$��VC&��0B�o`��<s��Վ�Oa������K?��vҵFE��z�������ZQ�Z8�l���"�^�g�����ș1n��Ѫ���
���DG=�&\O&9�c�M���zz­��Z��h�/�E�2d�F�I�a�G#��N��|�s���<�Շy�_�@+����L5��z|X)nb�%2FE�w�� tsPq�@>�K@UU� ]��r}���R�0���� �����h�\]�t��|�|>)#T�w����������� o�ߕ`y<s`g�X�mh��M:���s$J)&��z�<�j��Kj�<���G#�H=�؝����0�=���h�j�^�@�^�ʮd�LD��#"�3�ڰ<u`y<sa��q<�5X��}�Hԍ5#RE��f��z��aV��v��g�{$�I$�UUT�����-�;����\[Y�0%ـ�H��:Ӵ��]n��ݮ���<q�e
B[��n-c�{N����u�k��uط�;���_5���9��>V�4�ݫu����ʲ�6&�O<� �����"3�U�j�lv�����ڹ:�<�<oc#[���!���<]�r!u�랞��8hg���*P�&�q�&J��d���'"��Z���n���l��t��$�^F�T��{[x��<�����.��Fn4"^GLa���\=sYv9��m�O�f��:�3���9�:��{V8�r#�S&HH�8���Zyڴ׬�<�W��gX)nb�%2FR�3�ڰ<ug�܈�"&Z�~�_���Q�N�(I"O$�#�@=z���zz­��Z�p�N�&�f�̷.fnI����rO��_w���W��- ��4��J��ƜR$��g��=�\����b������u�Z��x�Q�I�	#�;��Zyڴ׬�<�W�r��Y#�)��Nf\2�I��w�t�2�T�"#�¨sb(��!���s��'׽��$��V����"�<�	���ԑh�?j�9��*Z�Ihr�R�D� �jj�>��8�u��'cU��v� ��4vTD\S&HH�㙺�}���d��:9�������.B�b���:��Ÿ�Ӱ��h"�IŎ�q#·t�������wϖ(�1I�ȿy���^�@=z���U�T{����r	�qh���:9��*Z�Ik�z����4���MB9�")&�w��w�ʴ���u {�:$ �������\ Њ�!��r���!CH��A�!�ʨ�H� �A�l�`T�"VT%ւ�*�E��kJ�m���"�a�"� E(��4$M1�ЅHRQe`ѕ"�!pփIhM	=4�
���e֗߿��!�/ L#E]�;x�
�������T�T�z�_�ՠ$��w��p̸ؤ�L�I�w�ʴ�h�Y�����K��M��̑Ɣ�HܑL� �$���@��-���O�����х����M�i���Y���{�-�\���$��k6�,��:BC\�2��UK��j�<�Ձ��o""9G=!�~�X~G
��LT�B�Q55V��@>�R��K@�:�{l��L�����yܫ@�;V�$w����h��
E���L�e+���G��V����X8�r�����2�����H�9�I�8��X5�t�����Kj��vP���[�%�u����G7n��Oayܦy�;����&u�4<փ�t�=�"3Ж��I? w��w�ʴ�h�Y��'rF1ƅ$nI4�V��/?�Z�_��z��*�u�8�c$nH�E�w��@=z� ��4�V��a���8��$�h�X�9���*Z�Z�*��y���H(��� �c�y��<��]�׽w$���srN�/E���舟����   m�tWN�Ux2�J�N�/h����#Y�d���s=Z6��R���6�N�]d��)z�|�|���z)�DGIsg�H���͓It�jj�24'eVN�������M�C��:eH6����ZԜ̓Z�����R�1�L���m&M�s��CWM���D��]�3�yX�:��tn.��Y�e��Ǔ�e�Pr���|��E@��Y�JN�ˢ�Lֵ�mJX�z��]�@XWN�q�4��6�k��TV���DLS&HH��N�eZ�v� ��4��h��
E���L�V��Z ��nj�J������$y�y$�qh�Y��@�;�h�ڴ�e�n<�(G1�nn� ��d�h�Ih���?w'rF1��r'	$�yܫ@��ՠ�f�{����mPd�$G����\���-���>M�n�����Vu��&rď.���d/45Gͷ����>l�f�{����U�ue�#N=L�də�w$���sqA4�GC�����h�Ihd�6昤�94��h�r�?ٙ���z��Z�_����ɒ<x�@}���>y%��j ��	�S�R(��$JdS"�?s�h�Y�Uֽ��U�Uxm+&52&f�✗�f�av�3�L6�lƙ����ĉD�$y�y$�qh�Y�U�́��o"9��s��q�D���*TT�MEMUXcs{Ȉ�D$<��V���@=z� �ܝ���Ȝ�I��>�����w�w�s@~@_�{����>]��@�W�GS#rE2$y%��j[��T�3:��8��$�h�Y�Uֽ=.�<�`o9�G7kHF�(�BDա�l�&��q���\Og�<��@g魃=��'B�"E388�L�O�U~���T�L��G5Υ��%^���G�G�w�ʴWj�^�@�ֽ ��:�H�s�)�L�@�v� ��4]k�;��ZV�'Y#���&H���.��4
��=��U�$"l 
 �x���wwrI����(�G2L�I�Uֽ�����Ǖ���k��`x��=�IdD�*&�B'\����m��S��E���iz"6z�ka�ܵiv&�8�L�Q����?>�����ՠ�f�WZ�Up�$q�1�7$S"�=]�@=z��Z��V��hΡ#MF����h�:�1csf�"8����`f��=��`��q&	�&�˭zyܫ@�v� ��4vTD\S&HH��M���X����] �{V,nl'�y<����� A�m�mW=�B��+�8�WM�"{lܖJ�8�V�)����ns&�/ms��d�J*z3���`�;��
�6�L�ᵘ�1v��F[����٤V)�qf�՛�ۓn�dV惧���-vђ�X⻠<�&�K�X6�ݳ��cS�m�ݢZ҈�J�\tOG:�sr�Ū����u�ݖs���mlW�m����v8˗sH�w�?�����޷5�s2\!�f�"���&���Z���:ڕ��7qvrƺ��\�a�ABF�)"S"������Z��h�נw�ʴ�.V�A<����V环��$4�f�y;�Wj��`�$jD�(��.���r��ڴ׬�ד�#Q�I�I��w*�=]�@=z��331W~��|��d�`�m����Ih���v���- ��g�<g�']����={	���%��U�Ʉ���H�;qQ���j7V՗I5��UJ�<�Ձ��=.��9Ȏ���-�_f�O#�$�8��9u����o%+@t�- tsP�Y�b�$$x��zyܫ@�v�>�����H��@�����3�$jbn)�TR���s�6�U�f��76z\5�uk����r	�$qh�Y�;rb�J���Z ����mѽH`�rd��h��)��źy^2�n4�ã�DnK�f�۟��w�����ݚC:d1������j��Kk���� ��a#Q�I��M�}�ߟr��u`x����$5���UMA5S9�]w$������~�nm��EH�h	�E֧��srN}����>�-	��rb�- ��4׬�3���"��V9[-1SJ�(���@��- �$���D�>M����K:���J6��T=x�n7K�Ʌ��	�:�覷X��e��9g�s��#x��&��w*�;�ՠ�f�z��}�u������L�dZyگy��$�j�3^Ձ��XҖ'��'�L�Š�f�z��yܫ@�;V�^������K���%��������Kj��G#���}�{�߭����Ͽ����K��ͻ��*Z�Ih���:9�q��6�իg�����:�e�Bc�J�{ ݅�˭5�Kķ��t��#l�U�����X�:���9@���-�џ|�(�$�$Z��PG5 �%K@>�-�.U�#�$�8��^�@�;�i�fbW��- ��@�eG�2�	�<qȀ}���d��:9����'Q�`��&)"S"�����@=z�$�����'ߵӷrN;������% �X�YP�P�jB��*A�(լBBc��TT#B@h@�H�,1MUH�V��R�B% H�� YBF���*M��b"�VP�!e�,U,�E �M��p���Z:ٶ
H	x�D�@1�,+�%�AM&m�q �cŅ!P�Q�B)b�������ĉ`l�iP�HH&�����������     ?�=  [v�m�  m         ��  Ӭ-Y5����9P��Q{m��Zڋz����7��\�]	Z.�x��ƀy^<��[r����n6[pW]��ό���鲜�� ���z�W|Ny���D�=n�9�m��Gl��	H5�s�r�0$�<�.�݄L��e��:��]q���t�S�uK����v[�EC�v�%��gg�s�ѥBm�&g�V�� j��A�2R�m�l�Ul  ���7i�f@�5^���Z&j�m����G�
!y��gt��<�e�;Gx�.�;�)��Q�R����,d�k�KK;$���C��u:{D���l�s֦��S�\�G�Έ��76�5]����2Ÿ!nA�+�^J���^�4ֶ���ۥ��pe6�6�(��lv���j�B35U��f��<X�F�2[��ک]���,�\�5�T�X�m�\jm�.�%��2�֋6vv�/C�.V�'�.]�$��M���E��u���kvZ �`�m� �I-���%�q�
,��m�d�D�����읕:K���I�0I@x�eu�5T�^�C�\Չl�M�KQ�K����.�34�`P��M�^�����C��wY ��1B!ɶm���UT�ތ�H4SJ��G;e�u5V�f��vP0SW2����l[ f�S �@�b��u{I���g��k��If�}�]�썥�o:�Z���3r7%����;\6��CO�$�j�B�m3�)�zQkd:��dWpa��v5-R��U)A*��Q�q�u�[U��.�J�H�)��]�r\Zö�8�WT��&��5m/-\�:0�M�lv� ��(�n�^[� �uu�Al��ej��j�� ���}ݶ���kFIm�H��A۵$�7'G\ϳ�۷!�H$hr���<�n���M�v	���fZ�V�q@�)��J���A0
"&������
hz��@(*�G���ky������� m�{_4�D�v��ìZ�Z�/|������ɺ�W���N�d���ݶ[�5��Bj�S]9Q�B��Mh�8��=U��P����p�[s�m��[鉍K=!�ݠ�c��s�X�K#Y-��W&�ܓMӛ�����HFm�s���n-�&��77�;mF���ֈ�p��v톃sa�0���k��nIx7D!���{����̀�w?��]g1�5h��D�q�t�ڻ:ѦB������>d��_��{������Z��]�� =��f:�3���-� y�55&
)���7�fg�$<��V�� ��W������f꟢F6�b�7$��������Z��3?��#��M �~�+��H�51��E*�Vr[V玬َ�>�"��|���}�H'�(�$D�h�:�>�D,ok�<��Vr[V��?hj�'F����n�\D��q��O�1�[:2hՍu�t�����;�����}���>y%��j�4p�
�*�������3���s��Gb�"�����.������'��o�c��$nAlTMIRMM%QJ����;��:9����}���%��V�L�
b��
�V�}�L�����X�r��;V�^����j ��d�h�Ih��������i���5�s�]����;������lP�n�9i9�R�]R�VR\L�j����j��Kj�<���u��X}[��9�LDmɑL�@��ՠ�� �u��V���-	�E/tݳwm F�nj%W���w��H��
O�7�o]7w$���n��\BL�M"���MU�܈��&^��`|���X�mX�u`y�G
`�+$$x��&�|�U�~�j��f�{��ׄ)�dbx)��2F�K$-E��;m�)�����:�i_K"�YL�
��Gn���Pjdc�%2)�~�����f�{���ܫ@��+���'�I�qX�uDr9ăڰ7'cU�ܖՀ^����M �u���jϢ��`�Հw2e�U*�ESS4MUU�܎s�[������`>�nH��Q�?��a���y�'/~ֻ%T�J�EL�TR��`w%�`}�qk{_�:ߦ�|�U�w���dB�#�&�,�"4�>)��S�s��	�M\�ɵH�1�y�BLRE��� ��4�r���Z���*	�qHMT�X�:���������`y������$fƣ�h*����bbjj����`w%�g���F��`�Ձ��:����JdS"�?s�h�@=�f�|�U�U����X܂y%T4��:�>�,ok�nNƫ�/��I��;N��;Ϗ�� l kY<�v�IzK�/R/I8v����������n�����]+�tv�؏�؟����U�OB�n�G�|X�$:���:��8؀[�Qs˚M����e]F������4�U{b�vvu���6��ǱXs՛Gk��kj�0<�`rv�ؑ�Y3���v�C��n�����vl��1{#Z{v؂Y��:���ٳ��T�? �P���w5�vjM�I�u�������y�V�/)ʥ���
�v}X�5��[��r'5&
'���@�w*�?s�h�@?rW�q�953R����\5�H��`�Հ{����u�Ȧ"6�dZ�vZ ��@���- �U��F���E�r�� �u�Wr��zϾZQ�����G��ssPd�h�IhrL@KeX���	��pY����S�{n�hD/����o�Ȧ���[i�+�Cv� �R��K@;�b ��:QX�TMIRMM%QJ��������s������(���M�?��1ˆ���qSQcr	�qh��@=z���V��v� ��)$a&G�z�kڰ�ƫ=-�nl�'����q��$�Wr���Z+k�^�@��m_�$����ۄ��+�n���l�7���%5$V{N�d�X�갭�H�51�&E2-��Z+k�<u����?G��ߦ��*Jb�T�b�-����Y�uw*�;�ՠ{�sˉ�q0���Y�wuӷs���! B��6�Q2"""=Ȉ�<��`5����D�8&
�������������ƫ��nl׬�=pκ(8��JdS"�d��w$���@9���>��˿�I�^ݛ�1v(��P�]�۟LA��A�Җٳk,�$�~��}���%�5.�=ݫ ��V9pՁ��Հ<��0�#�9&�z��Wr���Z�٠�W�q�8�q�����.�3�ڳa!��Xkڰ9un�G�27$��E�w��@�PG5R{��UU�(Q W>�:v�I�賽�r����x��@:�4]k�:��hrڰ>��s���#B*y0�SUE)�S^�jmӷ�¸��x�u��9�U `���cc�����-���Ԓx�����:��h�ՠm������	�Ɉ2T�L��rjۓQ�tPjdc�%2)�h�ՠ��7�4�f�͝�V&�qSE5B��s���f�˭z��V���Z{�RH�$�I&�˭z��j��Հf7VG����8�p�B
�#>�{�33333&c  l;#M�u�q)V�W�i�p���v_u7c��/.�����:ᝣ���4��[�Ѯ��T|9�մw-�]ˏe뭉�n'F��
�������U��=�&�X[��� �c'�.�]��M��׮u�S�u<=��m�,���V���n5�޺�bcL��7�<g�ի���U��Yx������1�|��������rZ�x��M������\��rkT\g������(j�q�r�:]��u��bp�������d�_�o�������v� �h�Y�yuv5#�SrdS"�;�տ�~�hkڰ<��W�""�#t�&QAUEN)"�~�h�Y�z��h�j�=�\�PN0�9&�z����Ձ��Շ܈����Ձ�'d��EQS13SU`c�Xr"9+ut��M ��4���dQ��q��|R9���I��Y�s]�˨����nw\9c]EѮ[88522G�ȿ�� =��@=�����@�u�dp�r�3Yw$�w���b�1Ut ;P�EPy��.�3�ڽ�9�H��Ƣ�E#�<�$��_���ܫ@�;V�u�h�+���q�ѻ��s%K@>�- 9&��j���H��Fӊ)�h�j�>��Dq=ݮ�f���j�1������O�z����^89���g�����8��Tj֬��Y�V�;R�$��$���@9���d���*�����M ��4��Zyڬu{��r8��'d��EQS13SU`=��Vz[Vd�DD	B�8E� �b�F!!�}sjD���R$�H�V�,L�Fi��а���(JDa�� �
��"ư(B�!
�D�H`��\0���b��O�H�@�
B��	u4��s4'�D����� �R"݇YpGb8� m�sf�DgD�c�]��+��$�"`0`@�U��(R � P"cAا",H��#"Hb�HH� ����u ڪ���P�Tv��
��CAS��+"�"@! �#"�	�
lE�,���
Y����'����]�#�L�dZ�����O+uX�ڰ<u`c�X�Ƥ�B<��8���@�fg����@{;�������(**�����9�JF�Ÿ	���(���C����3�:b�T���{$�?>=��.�3���:�����-��&U6(�q�I4�r���Z{��^��ٙ������#q�c#i��h���@����������-"�5B85"��f�z��I���۹?������� �Ȣ|�'��u�߮����/�u�.�Y�UMU�y���#�����<��`��޸�*�D�"2A��$Ox1�����4�fU�),�z���P�6�w�a<�!��@�w*�;�ՠ�� ��4�]�#�L�dZz[W���A��Xkڰ��W�9�G�$|���9�BL��#�@>���f�|�U�w��@�n���E#ȞHӎM ��4�r���Zw���������_6�������,��T�L��njۓǫ�<�?>~�  � 6�:�f�p��B�j׋��@��[r^s�u�Z��\��5�鍨{�۪.����ǆ����ώ���t&Tm���m��W��Thm��\6�z�qՉ���>X݉��ϫ1���<����z�Z^;����s]��,$Ѭ��M\e�1A�%C6x�m��L�
�V�0h#:ػKЅ�5�����;cX��nӿ���|���l�/7j��k#��2�!���]����֨�f�ubzR3��\�F"������V �X�����V�yԊ$�A$�ԋ@/u��?��"��6��j�<�`{%8�8Jh�$M�G&�˭z�V���Z{��=��?�A<�!���|�U�y�j�c��N^�� f�4J���ƦE2-�ڴ�Y�r�^�|�U�~���l��sncjbM)���cq֮^�m��]6�N�����|�	5��ȔRd����~�.����Z��h���Q(�y�qɹ'���[�?�S�#��+� ��v����3guX�u`bq.I�q�Ĥz�V���Z{��9u�@��u�ۘ�26�QL�@�Z ��@;rbvJ���e8E�H�LjE���������ϖ���Z�`ڸ6B%Ĳ2����C���q����m�6�s҅Ƅ��sX6�`�$�A�lr94]k�/�ʴWj��f��Ʈ`�'�$#x7#�/�ʴWj�^�@�ֽ��#�h����jdS"�;���BO������j����������?s�@�����J)	2G��G5 tsP�T�7�@G"�ܽJ)D�F�rh^����O���w��@=z��0m*��@nc��g���5��l�ӽ���[��#����.�b3�mF�n1)��w*�?z�h�Y�y{��9^N���SN(�m�>�@�_9��*Z�볨��E"$�n�_����@�;�h�e4sW0W�Bxfnn�:��@>�R�t� u�W���: :Ef�A�
�w�����v`�'�$#x7#�;��Z�9r1�ߏ ?��<��lfU��=��.g0ui��j燶�Wa���얌�U�KKVS��6K�S%�t >�@�_9��*Z۹S��(�$��C@=z���^��w*�?z�o��_���࢑�O$j�j�X�l��jϢ9	{6��������6�b�7��@�;�h�e4׬��1s���*����ܡLIS*I��V|��ŭ�tX�z�V�ٙ�������I$�I#m�UUUJ�ݤ�t���J�sRk\�u��ď�1en KClQ9A�
�\�Fʔ���gk�y��7j��m�Խ��^��\�f��.��eЕ-ڵ�׆���h�&�Ge��r���Sj)�6���{X�1��������ax���ˣm��v��9�\^n�,�K��Qd�[7�㝪�y��Q�ܻ��ں֋��\�P�<�U�}�Mj�ɣm��v�)k�1C�Á�GE�b�[smfvԎ,�bލ��K�h&,�0{6�/c��\5���P{6��:��`��<�&(��rh^���q��t� y���H�D�-1QTT�5S`nNƫ�t�>�"5���_���8�R��#$q��L�@��)�����^�|�U�r�jpr%��#QHh�@�g�s�����ϖ���S@�lJ�i)!�0Q%u�>6��^�vۭr��r��I�$���Z�y�7f�V' �࢑�O$i�'�9u����V|韜�GP�Հ=Z��&UL����j[���;�];w� ��"(h`I �XP�Rp�z�W�)�@$�_9�	pfL�NA�dm1ɑh�e4�Y����K�_���?��{��H�N$��4@���s�T��6m\�e��c��C�ɠy{��/�ʴ޲�{��<�b*�b��Q�;�;elkkS�{n�m9�l��j�����Nt�q���+�W+1QTT�5S�7'cU���S@/u�����(ޥ1���8ԊdZ�YM ��h^���r��+S��(�$��C@/u��?_�w[�"&Ł��P��T<��DM
��n����rN��?���Z��4��8��<������t��ĵ�� {���*�q�Ĥz�V���S@/u������ڹ2"(�G�C�&���e�2�7k���u��C�U������w����4��F���=�O� ��h^���r��<�E"y�A�"f� y���q#=�rv5X�h�`��1F�#�@��W�?K����q/f֖��X��	0�0̗4]k3[����������'����$��w7%��D| n�޷$��|7�Lq��8ԊdZ�YM ��h^���r���iY	�����`�F-�1�K'V�ힶk<� P�/V,����5�[K��N5R{$�??>=���s`?K���Ϲ��G=!����7ﾸ��rF�F�rh^������s�5Xͭ,�:���r! {���*��8�bR=�g�@��)�����^�U8uƜ��"6��ȴ?ٜ�r�oK ���/c������VQ���LO'�lr!�h�Y�/����_�����I7ϳ�'� (��� (��� 
*�� Uj ���@����
*���
*������
���*��F"� ��@
� 
�E*�T@��DU��D���A�*�"�"",��H�� *""���"���A
�H
�U�����DU��DT *D
�X", ��`*��D��D�"���@T *H�,UV� U��ADb��U��D`*","� *X","*� ��
�@�"�B�B�X��H",
��,� ��"�",`*"��D`*`��DH�,��E@",�T�"�T`��H
�@�, ��� $�� QU�� ��� ���Z�(�� U� QU��EW� _� U� QU�`EW� �����
�2�ȌG��&(������9�>�n|I@�      ���@  ��  4 t� �	
�*��REP� � (�  � 
* � P�TU*@��JQT�    5H � ��   >��\[�ܯyeɥ��Ot���
�}����Y���w���ŻOo}o�����͗7}����� ������0 �`<�|���뼝.�&�������y:����n�r�	��� �Ą���� �'P��}�����n{�׋+��e.� �����q���w�� � /Y�:!�X��'�����}��������}��˖��ԯs�
9ײ�t������{ow� ���(  ( �̀ ��\��\^w�<^������|�ռ�N��:�ŹU�@*��+���G�s� 6��=�}�Tx }7�jq�����һ�:��w�� �����=�|��|�/^�oR���
  �P���������>�N��__]��1�P�@0�����3� ��)Nt  ���ܥ Jb4 14��� 4N��b n�:P;�: ���݈:P3���ΔPwX�AF&�P qĊ �� Q���
 �Q�)�w)@���q��x �o��/t���};�YU}���_|� ���e��sy�v<  ���������B�o'���o'��O{��{o�y�� _O��J�۾�]_;۫Ϸ޾�������  z�)�R� �р����j��@ 4 ���R�*�hL�"{RM�A���hb)�������  �M�)$&@4<S��(�����?���:_��5A���Q����% ��3/�\ES���
��Q_�U`��*����'cg�$k5I���K!$��_�GpH��m�SFK/�'��l�� @��	�����H�հ!  J�P�w�U�r>�2���$a�y�95���e?(b��$R���# �R$+���B��16�'�q��l�E�h|��I@��!���H��FC�f�5�Z֢X)���U� �30L���}A�ɫ$3�%5 ��2˘e�R�5
������!�����+�͍E@��W�����y�T�N��M+AcVLd�p�5��9�M��P�	��a��PӉ#
s�o��+�M���ǐ�J��s_`��ٜ�h�g
�P�Y x$�1���B��I��b4O�?2$k�i �Jq�m1�	%�ю.͐,ii�۷�M�k��6�1>B0�@�$ aF����&P|]R�s����� �/�'.��K7���N:���ɳ��Ȱ���bh��I���j	M���)��xG!��~�@��1ౡ��̈́�1+�S1۷�D5����!F�N6a��28�l�d����v���l`���!IWD�P�6���Ě��4��	7CFI��v�4d6KBW�ީe�ݥ6F���0ܺ��Ի1ٴ�D
�3{bXMa6RM�iz	���	�A���BB�~tb�0��	iH Đ�!#�A�20�]BHR� @�Y%�2]3%$	`�4�Z���fH��̬`ȹJI	Yml)k�b� ��;�0	"#���j<ͧ!		m�Y	eM0D4���F+����
�f��y��]�aN;6L���#��ܒ�hqv$1`�g��Nr�۽:�a hbT�R�ۭe�,�����+Ł~#tb�h�D�U5��n�M����B��N��/�����6�:D�ֲ�������}�������cX`Q��f���G�O�220�X1cf�փL$��CC��	k��H�5�Ó�H��7��޹9��-�s��ѷ��%�������؄i����}w�R��N-�XaB#H�R�R:H��O�B�����8N0�!�2�	���!�(EEl�`�F$ h�x����T����Yђ�hCh�
C�(B��bƚ'�P"B:`m�+���	��X艁��"Zh1��q9���A6��)���7&�C��MD�I��ĉ��G�F���$lL���!a	Np9�)@�����qێ͘~�l��:��&9��l8�BkSh���i����0�6�y�5�a�d�ЅH�2M�rH�p8M�ȗD�$��pX�8Gp���#0L7ŃRH��$�!ty&��#yd6��<p?(�aCI+���!a?~�NkY�9��A$-B���"�?�cM�C�$(CDL6�He� NI
�B��,)�������d#];���Lk	`U��E�So*��7/
JD���
P��ۖ�C�[#5l��.��i�
���ėU֌b�@���b��.�ת{��*U������#�#P�2$��%H��cF`A�H@#$$"� �"�$HWD��6p�(h!��V��BSFr����n/˶JA$U"@�B%M.(AH�]����㳇�f��5���M�3z��xq��HNi���a)��\J.�8�i��8�a��ta��04с���k��1y�+��
�u��|*h���_!Rt���)�/�	u�����(j�RaHR#��at�.��.����m�9,��]/��HT���@�Q�`P4T0"��i���,cWJ�LM���(l�bX�M
D��1� P���ؐ)�.�F0`�E0�	)�iq`�!!M+����A�:nfcl�[��?j~��� Ąj@���0
ƚ4�h��18�#
i]��h�c����*<���}sjR���m��8_�
�����VB,u
i�T�E "Ađ"$v�BE((V!Z2ۛ�,?�aͤ�?$HP�D��1�$)(D��D4aϹ�M�j��|.��ߋ�*E[�۬��Xj%`@4���H���&w_�x~9��i�B��X����BP���8�]�X�)�w0�T���xp!!�(i�;!ͤ*J2聁f��ld�9��lvm����� s�ȅtMË�	u��!XY�p��rnht+ #��B3�M���Gd?<bR�5,���5
&� 8Gd	���iJB�u�������#�
�H��"�1ѦcA �tHq�e*���֡��"ɣF��%4i���Rt��	@Ө�5�.~�Ѩ�.�z��ф�hHj�@�@#4M]0��޻���ѣZ��K;�r� ������������фXФ+I�	YuYR�
X|�G<挚�0(�Y0�Y�X0t�����G��#]&!�"P�$hh4kI.����eϴ\�	�#��^hF���@#�]]�H�SF4�'�5�g �Fwm����$(��AMkY8p�NW��JwF�eщ�r]k%60�PBS^��MU�_"�ǅ�Rs��0`m���x��@(�$��/�*�����R�\�h��Iۺh��K���[�Y�C�)���_�4�:���WL�%����"@$H�Y��+��8pFta����tl�#��4�1����ȒB����p �!�
D�
A�.&;�y.�]Ͼ?)I���.$)q�É�aXSi	M�!hE����
���~�CF8~Bю�?�LH?�PҘ6p�~HWN.Ï�_��.��vR5ӎ��K���i�pӴbPӉ.�!�h�Me�]�B��f�p��"�H�8��)�K�xC/c)������Y5�CgƳ��~4 :(>�Xhֹ�l�r:4�i��Jl�4�цr��k�¤o�Y:�w�/½M������ ԟ�5�y�xe���2���]m$$�d)�4"04L]� �d6�:74˺ƗZ��K�4��6h9�P�oAw#%�Yɬ��Y�H-[�-y!�aY��ƑW�Z�a$�<��T9T�z��
B��"XŊWY��V�| �
0&��h� ��@bT�B-.�o_a�}��d.��7�o�n9/��Б�;"�B���1
��0 b�v
k}��_֤�>��w�i��!ѐ�e�.�9�����N�H����h���Ӑ���%4ozeҒ�2� 4��$`H���%'���1�mkT�%&@��m�%}UU��C�B�_�~4�B�!F�B�%4�A��H8$���B�H~�q@�Tu�Z5/78f�5�$�>9��_��&��1�J����dCj�!R~��9�
�IMJm6�����]o[� �F�&��ڒ�3a/�;81�����рI�LHƑ
K�	�f��k��h͛aN�5�G�XFmO�F-)��E����0��OOs�:�6�u�u���ߏ��� m�  �       ��       � m     �               �                           hq"۶�r�Y`[uuN��V[�6ٲ��I-N�� 6�`9`ٵ�m&�q����,����[A [\���o[�^�� ���G6�6ıwl��
�UUP�t  U���
�-E�'�����KZL  c�ۗ��m'��m�&�V��8;e��p��-�6�M�Cm�M�lmk7Z�X��F�Z5怪U�UW��M������2	����;5W6��g7n�j�L�UR����U�e$�N�x	m���!r�+���iU�\  貑\I�l     @� h f�      �� ���V A�Z�k�ݶ mmff�^n��jV"�M&�0�@3��-�e�i]��\���k�c"d��T�Ie�`�s[Pz�Q�s�v���vT+E�ԵR��W.Y]��j��P-�[%y5���m�\���E ���nC HA� 5�i0 ��m#m5i���9mm;mfБ����v�hr@@��jҔ.ܭQ��z �V�[N $�4��@���Q��j����V2��m��p�gj�.VF�d���4]J�&���(F#V�̖�[�%���U��5R��-�:u����. m�մ-� !#    h ��  �h   @                     ��g��ݢ�`	�V��>|����A+�K���������1�)�0 �u*��tʵP�못h
��@h�uUUՕ� h����Wg9nH ��-�8�[p%�\6�X4�e] t���UN���EI��n�l�M�$ �a �u�����WR�A�Uj�&:�-6 �/H���U��۴��m���m� �`  ��m����vÂ��ݶ)Im�*@pm�:�m�ړ��8��sk�ɛ6��A�Wl�+��ᶍv�m�K:��$�[C��u��6 �nٴ���6�ժe@���m���������y�V�V5*�Q�:i7<5�܎���\�]T[]d�I��p����[�:�.#9�g%�����8 	!�f�Ÿ    p   m��P�m��`h�-  H� �H�Ğ-�  �m��lm��R �` M��     �	'I $$X���  [WM�t-�݀�P H �R 6� <�� �m������f�\ ]�[U�`N@ kjIY��˕�� [@ ��}m}�$T��W���0=U@:����m�6��   ��[@ H �vV�yM��ɹ���&t��� 6�` ��P��ְm�Mz��\ގ�$�&���f	��,���V���� �  �� ��ݢWl�A'��6�'�` �-�N�H �����>}� 5��0mpp i 6Z  [@��e�mU�Z��:NN���J����p$ @ �  �m�YL[@��( ��-�$ඎZr�-/YX鱭�:g������9x�   ,�6�Ӥ�-����m�`�ۭ� -���l���Z#m�ۡ���V�ZccU���k �����$�P �F�x��U[@`����6�y` ��k��g\��[봁���۶��K� ���m;|���m�� 	e-����Z  6�^��H�׮�㭯���a����Ӣ<� -�n֪̭�[�mu(�$t m��  k2 qʖ�6�v��H8�&�Hm7K��u�D�@�I���m��z��.�*��U),������7U[� �n :A�� 5� �8��p�-�,7l�[l  mm�6ݎ$-�mt�6m�i�����{ͳma�N��`N�i&�-�m�6���m�:�x�A��l�/K�� m���k� H$8�`�ޠi�  
�j j�m� ����@m�v�   ���m [Lh́#m��� �j�v��� �d����������ۭ� m���$m�-�   ͗���[q�Am2p�����n� ����         �a�  ڴ�  �J����l@����    p�m�8m�m   Hj�ll�@��~�m��6u��M�$ $��H6���  p6� ��s�o�m  ЖU��W6-�oP ����l�K\���� tZV�:�6���\����ZfMvD���� ���i���6�i\�.��/(�� �`���2�H[@ 6���8���f�~w���K��  v�<��UU�5�T��� ��[ �B��v�j]��a�ZU���cr��kU�Q��3��+(M�m]Z��e�V�hp ݤ��� �   %���m�m�Y��H�nxH6݁:  �3�lP��e��V^��(�ڴ�n� �	H���[��m΂@    6Z �oZ���� ����` l�  ��   ����l�zc��`�d��  h m��6�  {u��e+j i3�� [m� �d�@	�l��n�I ���m��  $��i6-���m۰�e��t^�i V͗bW��6j8A�� '8���]�Km�mg.� �[:\�� �-��vE��l�0�;N[� �		]�랗j�Z�U�
 6Z���d�]��1 [$� ���m��m]�j��Ʃl��C 8�UR����Omu��j6��-X�e[E�@�8�כ[��)�y��L�W]R9��ll�@n���PZf�kj�M�$� -��bF\�Yx�m���`������l,�&����6�C�tm����H}���P���ط[��`,5�-���E�d� m�T����!a��   m��ykk(�Y�eC�U*���%���YS�%���)Y^����Ij���]��+`Hm��p/-UU]T�J�R�:�@��\S���8�RNm�lH-+eZ���e%�V����!m @lp A��K�����	/Mv �c�[%����% 
B��]mv�
�c� ��n�  ��`� p6���m���ۭ`���&�Kh��Hm��▪�
S(�yV�@[v탚Ȧ�i���b�  �-6    H�� ��c#m� �����m䅜[p@�m�6�-`   h[@Xu�-����� [A��;M�m �ض��չr}��>t�������q�j��R)3l8� B퍶n۰I�Up ��t���FꪩЀ��HS��<�U@��0���i88[-����m�i�Ca`�@����	h�>|��\�8��8-��h�N[��������NT�l�ge��6�I�U����] nzZ^�z�  �h �Fv��F� ��f�(���ki
^YR�y�mv�I�  �j�ne�$ 6� �[�m�n�,��8�cl�WI��J��U�P�'�d���ڠ�WG ���8�5�iVj�[n�9m  �ު���u�Ҭ��䊀
H���Π6ۭ�p[vۆ�>�ﾶK��aoYy`���@T�Vԫ�T ���nm��d�l�6��-��JH�[��H ٷa'$UPA���Sh��ƥX�yd�'�m��[�[-�S R�q+�MMUT�[%� ��i5�q�]W�I���V�&ĵUR�	�UNR�u�H� �	�jݭ�mi���     l � ����0          �        m��  Sl�v��/ �� 
�mf�6�,�f�6�A�  6� @ P�Sjڀ   	 a@    I��X��0 u���P 
���A�s�u�Gt��r�.1UT�[C���p���m\&�Ǭ��ݰ �$�mfv�u�[ [BAmRK#� ���6� -���ul�,�t�	 ۴���3^�Hm&�H	�	� �ށ�m�m�*�� ��G��V˶ųe��$[On�H�\�U�   ���n5�՛m��vH��w��F�md����%LΪ�y�����w��J�/�|����P?�+���Wm(@j4U�Sb~D�H����(|��D'�Ue��t��Q�j���c2B
BB�D������+ �@?�"��B�tڿ4EM
 *pG���| ��C�Wj�E ��D��X�;�Dz�H��@:�Q���P� �(p��@"��M���}A��*�Sb� ?!�/ �� �@"������� �D�)�D"��  }�|訯[ g>?"��E:y!�`3 ���"���z�%�G���
� ~�~���)�&��:�:CA(@�������b��A�X� ��DD�� W���uHbŃϐؠ|'PW�?	�""A��(l@�҂?(� ����⢟�G�
l�=@@�R ��A�E��@�mT� ��&`@���?��**?<:,<���^���� 'D"�Oʿcm�6���   m�\    �kxF��ʵ�gl�=tn����g���uĪ���]V�!e�-���e|JA�8]�s�� �`m� t��m]�v�a%E�z�k�eu��L�r�*�n�pBTFP@��3� ���v^w2��g��M�7����*�C����"hV)n55T���UUP���wOjR��:��msi�"a�\ݷ[������'��%@9���$��<��:\`��n.���s���t�w]r��=
0WZE�U��@�j��/Mʽ��F�.H����9y�ZͺT��G[m��2l��Nɕ��ȝ�6_:�V�pt���v�rsױ)����vѱq\��"�r˷ �m\�i{r%��m	�= (���&��{"�u�cQp#\r��x��1���	�6���;�m�2lٱnMІ�+���-ۍ
��jc7mP��;��r^k�1S]SÚ�i�\� �գOtKUnk�Mh m��\�,��cN�s2���CΛF ��{��v�F�J�
��f	�H���& �O\c�C7*��[;����0A��.�V�x��[ra���N˴�웳�9��4��h,��-�`O]�	%�6��omV��cm��筶\Bф
�3ma�^	��T�ɧv7^.{v�-��Y�٪4:�jv�HҾ���K�E��+r�q��r�m��.���Y��h!9��:nlM�j,�6Y�2�N+#6A�� �m�a�URMن�»��iv�����l\�7:GT=K��TjD��(��1��^��,�$cY�;ؖ�;���)��rX��F��Uum�*ݹ*�6ډ�m��N<�mճ-D:2�,�MSY:v�I�8Wu��E�����d� m�H   �mݍ��Sik��7� 6�2���׍�Ć�m�	؈5�9A��摎D3�]�5;=r:ぐ��[�j�5. ���D��"�����C@+�SU�����ww�w�~?[��j���X7Y��񭄻]]30�PIQ��Ö�5�9eت��`˶�]��7'֦�wI�,v�㣲��X��T�z9�ƪ]���\� 6�]����nSp�[qe�L�uq��E��) �l�v7VE��ctO[��;a��-��8�0C���	��q�j6���ce�۫���:S��t���ŹC3҇g����w���{��s��ۗ)�D9x�69�er��l���ܹ^_�h��i�����s=빠s��ݬ��4�/�=�֬{��T��e-�%L�VޭپJQ�
!*�������ۚ�[��s����G#qd�G�:��F�t�0=�%0h��_�p�d�17����h=n�λV�~�3>�S�h혲�"�,,�ʼL�F�ے��J`n�k�����M�.�Ֆ�ss�m8��(O���<��5���,�#�,�V䀍���YY���)�:��F�u����1��X�&AF��h�ս*��X���	"H���P�
!{�{}j�չ���[�`�Y`AFE�H	H��;�]��i��)�:�I.�ϋł����^b`E�4��ܔ��rSw�L/�ʌ�A�H��6�h�h���.J`n�i�H��"E���3�e�z��۳\��c�R�iooU�/,v[�\/*��`����],uT�͉�%07z4���i��)�n������Y�f,Uw�����.���ڴ�jٙ�}���ً�)�L�k2��:w��ܓ������� �Պ(~D0��]�ܓ��wf䟻=1XcQ%$�L�L�9�j�/����Ѧ]#Ln�]ϲ������̦뒘�`E�4��ܔ����?�����аr`�&Q��K���b��6�R�5�J@;Q��c{��մ(ȲI)]��ۚ�[��s�ՠ_;V��kY��CI��4�F�ے��J`n�i�)ҔH��d�E6�h�h�դ���.��s@�m��9���~#��ȲG�yL	�%07z4���4�����*_SH"T�����]�'�g�H܊)�qh��s��h�l�ݛ�Jug7Jf%�:Nj�K�܉�K�6���<�=8�����;����F�ھ��5*��2��sM�5�9vu��V����<�_HfoZ�3��y���ˢ�V,����ܔ��rSw�L	��s@3��7~�C�(�r-��Lލ0"�`{nJ`�J�2�,�W��Uf^SIV�O&S�Lmڴ�j�=mk6|��b� �rf��7mX��>�����͵`u �H	F,�F %ꄣ*�WD� !�XDa#�(�!�P�w����~۶�@����m����;7a��EͬHJu�m�[8����ct6�)�	��:0Nq�H���kTls���I���ŋJ��/ϟ0a�����>���<����C�NqئweR�g7��^��4��/N*U����h��-�FR5�4���6�s�7�s�z��^#n1�x8���q��m�6�6�Z��o[W8Gh�4�un�k�sy����=7��p�U�e:H��k��'R��,�l�z��]Q��u��L	�%07z5�|���L�09|�xO��dn,���|�[����L��֬[�j��ջ6�"rM��W�YX�˼��F��F�ے��ՠw�b�~�D��$ND�h�Z��rSe�LI%[�<��XcQ%�ĦE&h�h�ՠw������h��Z��d�$9ڶ"s �%�Ocn-�`�1����,m��;F���0P��Ac���E�=������L]#Lm�L�)\+/*�f�5��eܓ�ﻳ~(�����������}��.Jm%Tt��<���ŒA�������9�j�;]�@�}w4ޫ."(�y#�I2I3C�""}��l���͵`b��V(��|G#qdLr-�ڴ�s1,��/˳�Xz�f�32j�*�ކ��u�c��M)Pu��F#i�j"ꅻY[�f��#�X�!�e�I����m09t�0=�%06\��ݘ�\�2�(m74��V,ݵ|�$����=������s@��XcQ(�rbS%�7$��w�rO��{w<��S�	�
���B���֬]�j�����<���Yy���rSw�L]#Luڴ��(�Y#Ɍ�C@�}`jލ0=�%06\��6B�enڣ������;2V�v˻6sj��Hz_l5\s���m�~���Y;���nz��]�"�`{nJ`{fA��Ѧ�՗Q��Hܙ#��s�ՠs�S@��mX^͵|�$�d�t�hp:t�s.�U�e07�gၻѦ����{�`�'$�r�S�ƛr�a�\B���+V�Z�>�ǹ�%��#�>&��M�>��S]s5��0̫̫��ս`{nJ`{fA��ѧ��?z羼�vB� g�W3�г]/L�Qi'h�$z�C$[��9�Z�� ���u�+10=�%0=� ����V��hw�e�E�!��)���K�Qq	U�֬[�j��ջ6��S��%�<���4��s@�w�s@�]�@�l���y,��̆<��L[Ѧ���dg�V�O&�ye�DH�E$nL���9�j�9���=��V��mX�":"t�ΕU]UU=�g�����Y�4+�0�#	бغ��h���t��[��]�߾����]��T��{n�����*3J����l�!�:=�eu ks���a9�Ee��J�c�^mu��j�Kphj��Z\��9�mwF\�ZzYwhu��-Yp�Ws. ��t���:,�$4��G�/K4��d��n]1Vܝ�nѨ��H��z��������Zz&�5mۏ�liӇ�MMڝ��A�NY�:u��"NL'�q�R7�7"�����;�`jލ0=�%0�WQ>�̫�0Řf`������i��)��٥�Jd���Z��2P�ni���1fm��ٳ�BQ3��Ł��j��
�l1��i�1��I�<�Z/�4�09oF�킹��W�Z«++2���`~_.�������뒘�3+n���̐i�M�,m�D�v�n'l4�P�$�<����t{��'6�N^Z�ef`������i��)������ݩVঘ�6ʙm���70��4�����n���ٰ;�]� �|��"$k"�7&H�h뒘�Jf}�U[�`E:4��ʖa>#��dMȴ�j�;�]����9�j���_��9S&7Nl{6ՁСr�����`nV��	(���ҩU&��S.��h���3��Ὡ�f�6�e�.���a8���C�ֺ�đ,$��9��_߷4��h���ϳPw�����1��i�1��F��n��
d��37�X�v�@3���,� ��$��h�}ݛ��8��� �7@\~a$�	�6Q!I*1��{�l��jՁD���2�� MJPE��x�A�TSAt���ѥp� � �	�QiCA��(�@�v�	�$���b:"�T�E���Q�id��CZ@0M�J� �4�h�w@(|�D(����!�T��*+�M��N=Q?
b?�Pc�E4��o��(r�=�{7�-���W!��S��Kt���Q
s7�[�xｳ��r�?}�f��"��t�=��74�I�r����k�9ou��!��v}=��6f��I}!��������r���%���.P��!uɴ⪱����]s�]�5�1�NX��9m�R�m}脔L�o����$��}���֬��-�a�IO�}�p:tܴ�j[vmwM�Q�B�Tn��V}	%3�w�֬���!}�5(P�Et���sM˖US�D%;���`}	r�����g$�{k�l�jWCcs(m75�	]ӵ�����BS!��vСv�y&�(t ��yHEO��������B���k�_욹nji���rڰ>JO���(Q��<��PwO�0�ITR5�MW_W\��)a���Z�qn؍��C!$񞽡�9�\Z)t���^�N���rV�?���������l�#3{����՝
���v��U�d�d��5]�U۹���VrP�g��Z�gs脾����$��>�*��&�9����W�	)��]�f$�ϔ%�t�f���J"d=�ҩH�lM�ꪩ�`}�/c�鳔$��f�����(����܇�AM�N����舉�}�`foZ�����a�>��6�#"#M�t���۪`�s�//n�u���U�juR��2;�&�]󤺩�3�8��»Zl�&��w�l����]ڵ�!��UW�X�6�n+]F]d�k�P�m��������*�ԜO]��A �zq���h�r�sE��R�Oh)����x\�3�j� �k�l�.đ����\BX��n��l�;Z�܃ۣ��Vu��tι���œ����T��T���Q?;A�M0�&
�箢 �d5>�3�5L:z��t�5�9g4݌6ێ�k�CD[\�}���������;{�r�􇲻�B�O(�o�l�jWCcs(m74��W�d��`{+�z���6BS���3��y��̺�m���j��=��6�wOB��37�X|���,�(�')�)2]K���!L���6f��IG��֬.">P��}�`�*���L��&�[�6�S���7��t(�C�]�`oWt�D};O�O��ۚ�SئU5;+qp�ϩ��\�]�W\��4u%\�g*s{7[��L���>�Jw��V���΄���wO�!$����ֿ(I} g��*��F�S�޵5��rN��=����Fc�%h�
 WS������ ����$7��_�B��$�1~�ߑP:tܴ�nl�_�M�D(S&f��{��D$��ewM�؊�:)�&��`Ӫs`n�i��F�ے�.J`n�T��%��"r'3@��s@�]�@�v�����8��m��Y ܍F78vԑ��6�����7QgVTȢ�R9���s���ƢQ�$��I3@�]�@笃w�L�0�s��(�e�^e0=� ����{�Lm�LZ�X,#�y1�ㆁ���h��ٹ��S���A*s��s�rO�w:X9�+X�i��n�]SVJI��0=[%�=� ����jI���Jr۪*�Vޭٰ?$�{z������w޻�;kHZ�b27&'�]\[s7%v����0������g��K�xWm�zY���1����Z=e4��s@�w4uڴ��~q�9�$�{��U�`{nJ`{�A��ً.B)�L�9��w޻�:�Z=e4��s@�Ea�D�NI�k310=�%0=� �����|�Z�!(�(Q	������7%1K��̦�d�Kw����ti��V�v��Y~�B��,q�dd&.Ύ�Lg��\�ۅ[\+K��dv�-f�����H�ci��Y��;�]��v���h^�Ya��l�����z4��ܔ����d�#A$q�ɚ:�Z-��}�f%��S@�w4ev��$�d��ȴI�`n�A��Ѧ�����_�pnE&�!�w���=�]��v���h�c�ܑ��O�j���N�{PuX��$Vau��3�iXv�SU\���n�ո�tDU��u���m���S�Զvʁ]!��-��e�sέ�����\��[;]v��FH]P�;�Nڮ��5,͌���8�J*��=l������ڶlM�٤�v�e8�FV�t�]�5����N絓��v:ψ�q��n������E�`�s3Z��*��D��y����4j�.��i#V���7[O�R�6���Hε���c�#�I�%u�[�D�'�I���?u���vl�^��j��35�`f���(�R�i���m��V��(J�=���35�`ffڰ�iF�9Lj��.��)��2��0;�4��l��9j�`�8"(Ldr{�M�Ѧ�d�����A���t��P��Q�h�����^��e4�Қ�~��,��dn6�N7�<=v��Ϟ����{t-Y�����8[j�}:�	#�nL�9�j�9l����S@��w4ev��$�d��ȴ[)}
X��4+��|X��Vޭٽ���1#�~x_�pnD�G����R��͵gD%3��=���=�jV�E �Ƞ�R�빠s�ՠr�K�S��Ł�+��Q.��ӦU&�Lm�LI�`n�A��Ѧu��@�θ��b'0����mƎ����N����l΀[������8~g|�GZ��V]e�W�ݙ�d�`{nՠ�c�#�	�G!�w��ބ�ɻ�j��Wt���6NeJ�`�C$iG!�[n�λV��>Ͼ�DD$%U�N�����`fl��Cu!$q�ɚ�}���j�9]�@�})�[n�̮�Đl�̍�E�[rSv�SI`{nJ`:�R���=�z��9И���,t�4ʱ���8B�D�:ݚ���]�=�6)Л/��ҘH��rSK���(�#��A�Z��n���$s�ՠr�V�޿U�w��A��i��fb`{nJ`IrSv�SI`��,2,��Q��Z�ՠw��nI���7'�41~�P�
$�A�Ā@bD�@���(F!D���HF2m����b�ʬF��}�|����������D���E1�Zz�V�~���h�h�V������2H�7
5��I��.��d����bW#�z{h����%��cd�)$Z��h�X��<�_HfV���zUC���mӢ��`}�ݛ�J"&N��2�������]�?� ��#�@��́�Vl��.P����X��嵋*1��N�qh��Z��hz�fÔ$��>�39�U��9���H��-�s@�]�@�ڴ����h��(���%d&��N�@u.|��%�\$@���AҠ`@� ;S-Bk&�хǡ匁v�$BBHP�VA�<H�,XŃ �C_�������_٨ ��(�0��0k�H ��U�͈�X�ef��bM4@� ����`��@*���Z@�,
�#�8�b]�C�(��#�!�dHkR�0cm��0!��K9�@�!Jf
@�J��"�␰�t�07 ċ0,�)HԔ`�B����X2P� k�����D�" ~s�UX�m��m�m�   �����  &�v����m ڣg)�6vz�tKӞg؋�!+\���֪_i�Y�9jA�7n��גe��;,�h  �������p��Gn�6 ����2�;���]�X����ڑ�[=�=J�jV5�i�yi���nݎ��
�nn�.-��m m��5� ����ݭ%�*[]zzđ՗�m���z]�XRt�-��Ofݣ\<�[	5H@�;`;b���5Y9ݝ����n���ŷG@O9ӵp]s��@V�����`�K88M����-PZ�
�j�y�g-̌�䙇h���cٻ*��^RY����](�e��]d���dx���ec`���q`v���v�BT���W�x�q�	z:vנ�,�=mj��pK��<ŵ�:6�%��A)q����/'[��i��v���p��� 7Sv��M��Z�z�C�]��Md�3�:��N�]S�2Z�� d%b�;rݷ),��M�Ē�@m�[�'s�H�.R;u5�6Wgm��j(6*��U+��1�z�]��=�y�5��n���=C�q��Wl�Һ*`+�\�<��y��!-J��٪�;���褉2-N��<��enڃ�
Il�%�&���D��d�)�9[m.\V�V�'��q�����p��:vI��c�L�{
01آ�=�@������K'7?��|�C+���jY1��u�d��'p��tl�T<NΆ%����g��N�Dx,嗶,��Xj%�!Yې'7��jd�;X�'<��֕j���(۶��n�@�ˮ��֭���,�p e��Cc��6�#�⥨
�K�f�����:��Z��^R6ض��N���D�]͖�,���ĭ������y$vʫ��N�X�(iK�����z�   H,\�:[��l��c� 2BF�ޝb���]9\ 3ҹu�@�~>o�	+)���j��5s�8
��S!��2hժ�x@M��E�!� �M�����T�s�"��C��&���3�̓0]/9���}��ä���8��۬t�n��ZR��[c��n�5��trN-��1��9�=���ll�ٻ+���DHs�m�G<KkJv�t�(��F:��G�H"r3��u�����-��9"XӴēE�͕�t����B���Cu=`�Z�˕�g[�e.�u���:�N�,���Ɛ�Ye�Kz�)�D��Nܻ��{��u������,�<�k���7��6��^�ʆ��mӞ[`��

d�F�po$�:���IrSv�SI`vLR�1K�t����7�芣2������X�h=V;�Ƞ���q��޼ٰ7wmY�BQ3��;��l�ʜ��̆6HҒE�[n��mz�ՠ{�ՠ����d�a$��ɚ����.J`n�J`I#L����N��k�6�74l��IӇ��7jv���x�c�'-�:��v��gڬ<�ї�L	.J`n�J`I#Lm�Lx����dp"n=�~�}���b�"�D!��֬�wU�n��	)�wZ�]ӕ*��Sn���֘RKd_U$�u�L������8��I&hVנ�4yڬ:����X��br��1K�.��$�)��rSI`mI-�ڋ��}��udn1���D�{n'm����q�˕5��n)�Z^�M/+8���;V�m��U��������h���X��̆6HډŠz۹�u[�`f�����7�2l�s�P�lT�n��Ձ���`f��٫���$�"Q�����`vgZ�>�YP6ɪ��̦K����`t���nE �*Ȍq��GF��;�����i��rS��L��]KUVb�{q�\�ţZ��Q��N�6�e��� ���.�k�����f��6߿~���ے�.J`n�A�:���MH��$��v��ڴ�Қ�����a�Bc�(�r-�vSw�ߒ�����rS�)dWH�"��di����S@�w4u����l@X�#���}���[ZǦd1��J7����9�j�9�j�;�Jh�yV���XH���M��\�{Y�7d�a*�ĕ�R�'7k-�cD�G>�[�������~�>m��%07�!�%�
�0=�Ɉ����ȣ�h�o��#��Ɓ�nh�h�R���d�܋@� �����rS�rSvb�s��,r(8I����9�j�9�j�;�]��tYr��5"o$�4u�L	��f\��F��`O�/��� Y��B��;���hֵ�������u�2���wAB��u�W���;L6)q�.��r�Vዩe'���:ضu��iع8��+]Z#��*��n�d�c��8h��m��[r@n�0j
Tx݊�ۮ�m�.z�je�����ϫ9@�v��Z�yzԛ�Ml;ns���2�-��m��K<Tݘ�.'+��B��d�vb��-n�i�r���.���{�]�C'7H�%��{��;����:Օ�f����n7�;a�wP�I<g�@����];����r��B1F��~����Z}빠{3m!D}!��=�)��r�n�SR����WД(S&n���]ήRK���q$���z`�C�4��5$�}���Iy��s1��6�q$�n�jI.�lX�����ɜ�I/;cԒ\��s�%�]�Ԓ]��3�I%���ĐOs"�H�$�=-\�I{�t5$�}���Iu�����!71���+����mu>I�i٪a��%�6�I�r�mra���n���+G�����I%�z�9Ē]v�~�8�K�m\�I{� ��X�Ƞ�N���y��� �	��rߵ�f�m���z���۰����*���|J��L�SR��)$�q$�����I.zZ�Ē���jI.�י�$��te�E	��Q���祫�I/z��y��K�}�7���z�Iv�X�cJ'����'"�K޻��$�g�������$�����I.zZ�ĒG�����lm�c��3Nf%���D��Vι�,i�q��Ƣe��:�<�V��n]KnGRIw޼�q$�]��I.zZ�Ē���jI.�lX�����ɜ�I.�c�ٙ�6�퟿.q$����K���s�$��W���	�G$z�K���r�~��ܛ�� ����޻�p�IW���I.z��"2G�I0mȹ�m���rn�o��r�o�w���|��}����J�~�H�ŎE"p5$�}���Iu����ӜI/z����ߦ��'VZI�r��܁�6��:� �n��s9Q�U���J㮻6dT���L�Iu����ӜI/z��y��I�Z� �D8b�G$�UU^���bI]�wF��UW����UU]vǩ$�=V;�(�G# ��8�^��I%�z�9Ē]vǩ$���Jܩf郙O$m�I~�����o��9m��{٭�m���g9m�tM,,�P�]o_��fgk��UC��Sm�)ɜ�I.�cԒW���m9Ē���jJgٛ��陞����੟���$��uT���L38����3lЍ�k=���ubr
�0Vݗ��ϳ@�V��� ?��?�����t5$�}���Iu����z�Xђ8�y$܋�I/z��y��I.�cԒ\��s�%m�A>�(�c�B8�jI.�י�$��=I%�KW8�^��I%��,�0pq��M�g8���|��jI*�k�K޻��$�m�s�$g]k,)�4��jI/;k�K޻��$�m�s�$�m�RI~���}����v�HW��z[����)uuLj��8TYx��(4$�$�B�E��*�ͼ}�p��]�5��$�E����J��Q�C��s!Y��9�����76x<�s��J�7YCr�k&�-Y���g����+Q�Msn�+���g��scmÐ��������[q�+�v�m�Mxx�m�4&�;M�䛟�>���\�5�\��2��R[�Zߏ�?�s��~K?H��Ľ3�Ѣ:��:���U˝q�V�4v�*�e��a�#�R�4��rT��n�������$�]�MI$�m��I[�,���C�nGRIz���9�ٍ��m�RI+�g8�^��I%��b��d�9$�nL�I.�&��^��q$���K��g8�K�W��r$���9#ԒK���$��wCRIz���Iu����[��FH����
99Ē���jI/[y��I.�cԒK���$��fg�߲�����8�&���mˋ�י��ms�'@΢۲F�p�:��n�~��\�!#�9#�RI~����q$�]��I%�l�K޻��$���c�LjD܊L�Iu������X�DBL�Z���r�{�orn�o�[��Hκ�XR!�j9#Ԓ]v��$��wCRI{��9Ē]vǩ$�/�.6�dpr2I|�K��f?z�$���s�$��RIu�_8�U�36|9���F�r�����s�$��RIu�_8�^��I$�ەbOY!̔+r�//f��;/n[�*��w=��s�PvϑDnY�c�N��B�ߟ����=I%�m|�I{�t?}��}��V����I{���D�9!G$z�K���Ē���jI/z�g8�K�����|�K��f4d�	<�M��$��wCRI{���/��	IF4"V$H�I
$�K){�(�\_́ �Fi���H4�N�A4�F"���1D&�@@B1����3X0���&���'��O���@bA �`�17
H�XČ"�R!!�R��-Ma �	�%���;�N*uH"mPC�#� ���|���!�M��O����l��v�_��ݶߵ߻�r�{ۺ�d�8�d�B8�jI/z�g8�K���$�]��%�]�Ԓ^��߇�5"nE&s�$��RIu�_8�^��ܛ�����r�|*'{�ެ�\-6�6��N ]�ne\l{X��
��*Z�Б���:n�h�Iմj�I5?������$��wCRI{��ffg8�K���$�o��Q�89#��I/z����s�$��RIu�_8�U�36|HC�Q��K޷��$��=I%�-\�I{�t5$���qc�c�Q�nL�Iu���햮q$��m�H���w�9m��s�&���t9!G$z�K�Z�Ē���jI/z�f��l�ya���T�'Fɏ����Gj�0�娞Bg[���-�خ#]]+=�yFH����F�Z{e4z�� �m�k�h���qb�"�q�@�&06\��ݙu�I߇�5"nE&h{l�;]�M���K������3���a"$1J�M����6g>,��V�n���Q����D��;�)�~ȍ������������BJU�F)�"���A���	DH� ��c���[UT\f��sr\H��u�7i��D����<Cs;�Ѷ�fi��U�)#�7[u����A��e'�����s�$��������m�l�Fq�Oe����]*Z���Ss����4]���e��ۤ�<�7[\�m�Z�kCv��GF�9����m�%�d�8v��h
���v�k��m��0N�'v�j��l��s�d���7����y�|v�vۦ:�\Ӳ�T�d9wf�f��!�@v��W��j�U:l��z4���2��?~��0�1����0=�k����H�rf�w����fgʍ��`ñw�LgKE�^eU����Yy���̃vd�`����+ƌq����rHh��7z4�7d��d;%�3/)R���//�F����̃{e4��2Ǎ���1Eq�FG�l\�v�m�F�nt��62;z���9�j����D�r)3@;�f���M���{빠s:�X�)��E�@�k��~P��BIDTB���M���=�ִ��h��ҭ��djG�2ލ0�1����J?�6���#��qw�r w���~ 种�~�,Lr	I"�ɚݓِ`ñw�Lu��WfiW�c���Z�%$,�&�q9��ONSF�H'#t�`���3��k%�W�ِ`ñw�LvL`yl�i���)��;�)�w�����4v�h���8�ō�	#��?~��7$��w���WR��p$I%*#�%\�>,�^��ZJ�"�ƤMȤ� �m�;e4��h����c�D�C�%RM����07di�nɌ	Ȳ]Y9�Ӻ�7pp��A�=�p]��qP	�7�r�k���&5vhT���Jm���07di�vɌِ`J��Jω6���$4��� �m�{e4�Jh�ŏ�A)$Q�3@;d���L��`n�� ���pSdҩ�.��݇Nc�;_��j�|�%
���`b�{J�T�4�2��̦��07z4�;d�������2cģ�9�&Fǋ�s*�.�9�'�gnt�r�N����ݮV6y�Щe�a���w�LvL`{nJ`ol��޺,��'�H��I��یm�Lِ`n�i��.��eT�s䢊I�s�ՠw�S@�}w4��h�Y(2'�H��R-��ލ0�1��)�+��L�� �RF���;�]� �m�:�Z��K�$�������~�J���P���<{>���d�ohWg8�q<&�&�ce�S1@"t�納휉'^G5�{v��S]�{a6���c`�.�!Ѷ�^����vwv-�a �0\Z9d��C��귳R��rz�멎���uw[���l���D��=b� �q��s��sZ��vhnL�Ѧ�ͳ�qm����F��v�"���v������lb�E"�U������w��	�3X;Q	��]�������[�mVV�r=X��]��Ö�0ERG��ɐjInL����s�ՠw�S@�}w4�����lNMRt۰>�n����39�`foZ�{l�9���hƤM�H��@�l���Ѧ�&06�����+Wu�-Jt7-�e���w��`������Xr�9�|X����)Ժ�:t:m� ݓRK`ñ�F���ֺ�K���٘Iv^�w:S�0���Y�=zuj�k�.ӿ۫���}޺d��h(���[xO�����ץ���k�G�gs�;�����8��nǠw�Sϳ옘��K�$����Հn��ӻ���2t�.p62�e�R����`�@궽���]�,FL��mӪmXtD)���`d�uX��,9(Jw{�V��H�)���i�Rt۰=;�V興Y�||�u� �n���߽��np�L��]DɊ<���̖j��N���kOm�#��m�������nJ�����Y��=�w4ݶhVנv�\X�<y"�8h����!B���`d�uX��/�D%2ws䉐q���q�3@=�ߦ��mz|��(�o��f�}��ܓ��wT�C��M8�r�a�D%9]�Vg>,��V�"L�w;ݲ�he1�*��Ձ�k����Dn�|� ��vU���#�`�9�<R�F�!㜹۫M��>E5�b�:e�h�������{��h���!Ғ5� ���� �m�U����*�c�L�����V�n���B_�"!U?�~�w��X������ �I��G$�:�ڰ=�zY�3��j�3;������R*�檉nG5N�9DBJs:��7{�nI?~�srEU
��|q�������.,x��<��I4��V%
s;��d�uX��,�?vʇ��ue���.�)q��.�� Ap�%gV9�T�ʸ�9'��]l��u���`�cjIlِ���%�	?~��;��?�j	ϒ�)&��m{�%�DBUF����;�~�`��Тd�l��C��nJ�:u`fs���ݵg�Q
&L��`d�uX��
��MHۙuL���S�����`zwv�?DDD�u�`t�s�Q-4ʚmӪm0�1��$���0;�i�>�������$I��X��$��lMf�
��n�h�)����o��1$�"A�FV$HȢYj	����B�[@�@���]!�j�N�����/#��@0��aRS�H���.(R��'b��ʠ2��	 ��c�X� �y�@��Q�^
X`B����B �`@�w�X¶�Ic(�H�,��)C�������q��      [z�     �uMwDk�i-��<���R���a�(��7+�Ŝ�Mu�������6�Yw7,s�N��Y:\�ie�A�%Z�J��^:��m<����}*wio,�/D��GE��U�6n��m�b�{g��<>;v뭩;]�	}`�Xݎu;[f�m��]p����� ���v�ڷM����ٌ)��+�9�qm������X�v���c�ZiV���&��^,1	��e�H6Qnɛv�+k	i��P��ڽaY�RZ�
C��ĹJ+n���]v�m�dJ)�W��2r�����]/l�6m�Ca5X��vU��Z"�Rq��6�OUm� �\��&̈l�6ݲ�aؚ4�	�u���p�*��6���j�C<�E�:�9n�4�	���q-�F�3�<�Wl!l�L�;G�q^� b0M����55�U���rQ�X��=/H킳O6�RI��F �H5�f^y������%�]�$�� ��P�j����72�ػ��}����-���cU�Z=b�w�IY�@yʺY{���B���l����J�Sv��I�s;��w2T�N�[�N�K4JQ��f̘ƅ��9I�7Nv�8��g�� ��v�k�:tLge�;'1���:s�Eg3�y�M;u�'AE���/
gP��\�8M�-����u�;9��y
3�#]]T� �
ֲ���R,�$�ɐ��ۑ�h�C��Y�,��x�4�1�����SjuΖF��E@�$��esvי[C�xIUj�)��õ`x9^.Ŏ��f�,����D�';r�.��&��[>8��]��v�2vf�1J���l%�ۮ:0,���3bzst��� ��Bf�;x�VT$�CyP�ޅ���t�]=l�	�t�`ld ��AV��I�=�a�z�7m�����*�A��,��Ҡ�\�:B�8�d�<�۱�m��yR�Ɗ�ҷ{���ꆅ_΄	�^��>PzQL  ���1v	���ߟ{���ֿM�`Yf��)�n���Bڦ��-Ӻgr�ݤ�4%�]U�l��iE�+i��p�e:�`wiݶ��:��8۶��]��x�n�a�݊Z�����T�Ӻn��`����Fҧ`����/=]�x�t5��Bc����ک�SJ�mf����;i:�p����v�j�Y6lIs���&Wp=q�&���6���-��&�{�ܭg�����hY�w��3�1�s+���L3d�c�g�7f�n�Y�`s��7OF@�\��&��wk�Ϗ&��6�q7��<U�����M޷WD(_H�����}J�U-�U܎j��� ��&06���|��3��J��t�KM�n�`n�Z�l���̃vdݐ���Yv�mSn���9����s�����a�s7�V�WW)�4�e˖݁����ݙ�F����_|���~�����c�p:u�5��8㒛r�\xU��KVڵ�kq/:S��I���6�O����ލ0�1����Ů�UL�t:l�=��W�Id(�JTB��:���0��݁���`{�����M��t�2��nj�V�����K?L�s���޵`���DSeULӚ��a�!BS������Ł�fڰ�9�����}J�U-�Uܔ�0`ñw�LvL`{fA�w��>�JzWi��ۋ��יbm��z����!Z�j@����t�s�fy�Y��w�LvL`{nJ�_z���~�~<�R���$s4��h�h��;�]��H�y������.[v����K?D/�%j"!�x�~������'߻�ܓ��OJ�朦�rUK��á(�ξ,����&0=�%0%w)��tfe�^`���� ݓے��!�m�~�{���KGRZ�&�mC���b�W��C��y��{e07�9�f5����̼LvL`{nJ`ñw�� ��Xу�m���LrM�v���39�`foZ�/n���Q
d��}I��6��N9��~�������F,�v�������*�6S�R62���`�L`{nJa�/����<P�w��7q�*���4�mSn�`�L`{nJ`ñw�L����߿N��PR�6�m��&.�2��k�E��9[@�.0<����g7hk��˖������ץ��fڰ/[4��ȜY&H�I"�;�)�
Q�DU��Հj�ߝ���vl�^k,���iG�����hs��9(J&}��6v�,̙[b(i�N�n����]���vln=,:!DB��woJ�M�UUL�MSn��ܔ����F�-����%�w��������?��jBj���u�{Q2Ɲtv�"�8�[
0g�Cjb��vZ��:ku�5�V�+D�Ln6G;i���Ԇq;J�k�nq&4�g(.��yTѳ��\��zM��э�VL�3���ͺt3!�/�f@���ݝq�u���s,��6[��R��!�=��oc���V���-�Itckg$�;����\�Y֒�nNx-����t�~����g뙣.�FkR�ۇsa3��'a�鬖��4$Ύ�:֫s�͂��F5"m�Ĝr.�Y�hﮫ ����J}!��;+��]C�ӑ���2���m_�J"d1gs�=�ܴ��o�}��G�����"����LL�~��ے��}U��n���Ԥ�j��TҚ�	)������`n�� ղc �ԮK*�b̢�ۛ�ץ��#3���,�vӶ��`ő8�)�����f]��rB٬Q�9hI��n��J쵨:N�j�y�Yy���LVɌT���I/���-��Ɓ����i�&A���&h�����=RK`{fA��ѧ��?K�cF�m�ƞLrM����@�l���z�hs����+ƌjD��\�:��>��6��� ř���wv��K��q91�B���z�h.�T���%0;��jZ�X��� ga����t���&y�H&��ay�7ף<��}Q�a����~���ف�[��wF��_E�*�%&۰>�ݛ��Jd�Wt��֬f��	B��\T��t���N����36՜�����>I$����}n��Wl�8��k���Ғ8��@��w4��Y�r�V��Ģ}Ϻl�]b)�SR���j�9wL`z\����)��Ѧ�"�WѦy-\���"�#�svsMԦ������r��cK�c�27�G�l���L�L`wti�r��ݒ�hƤM�H�$�h-�f|�m���\�����[������banLR61:����j�ř����f�>���ʐ��(�ĜnE&h~W-��`{��l��v��
����}��=�~�$��$�G3@�v� ���`r�0'"�R��gZ�7pp����q�qv���Aˬ7�UMZy稘�٣�9�@�7Q����ߟ~���`r�0=.J`N���ό��$n7&��z�h�z�h�ՠn�IB�;�eu�M1�-�T�`j��V�[�gBI)���wzՀv՗Ә��72)3C�1w���h9�Vfm��%�o|��}J�MH�b�I"�*�@���o�g ��zՁ�����%����*��6ۡY�c\㧭�݂�d�uĬ��4�qk�5���R�;t��F�x�J�;s�^f����L�u�n��q��z/kʱ�2�h�^v�q�bL��քxp��\��h�D�d;r��	�ssm�^;&�1]�t	��X*Ʀ��»nJ�v'�z�\Y0Ѱ�i�ݮevz!Mc]&)Ș�1��n�"�0���Us��i�ڷg=�c��'̯]a����ݜ�[z�t�:�9�n�+s���ds'On.�h[����c�8�����v���{e?�︃����@���C�H�oq�j������$�L�|X9�V��j�(�:6���dӥ-�f�tՁ�ϋ�d��05N�0:�JW��U^]��(WW��d��05N�0�������jW8U2ۥN�X�`j�`z\����-��.��N�C�K�v�;���AV�G9��Dm�:ʀ�M���w_>|N~m��8�,�^������L�����$�A$�����g�CNbln4�Ȥ������9SA��^�� �����������}w4����7�H��76O�j���mY�D(S8�zՁ�?ߖ���q���<Hp�F��;۶�Y�j���vl:!%
g����}2T6��R��Tܶ�Y�j���3t���v��j��W��l�Л���Ѥx��� ]٦9�f�I�7m#��qQt�ڷ�sw������x���:�������W����l�����V�i�q�Rq�N&L���s���3����3?~����\���4+k�/���	72۪m�`ffڰ<��j�Dy/BQB�w��qbB@"ň���� D�1 A���] :U HHd`@0&�8)T��|U�DF�"21 �!���e!F��3D���4o`R�$d!�R �w�(0"�p$�J�0Go1c$�0`0$Il�$�H4���L"��� �F������G�"� 8�P٠4�J� |�TAO����	��滭���l�=mk�9�lRH��4?�BJ'o|�OwU����`ffڰv�������i��I�����fB����ǀ��֬/fڰ=��s#����&�J�箢�4i����s���S�vSZ��\e\�6��<����SS�m��ץ���j���m�I(�􇧻�����8�Ě�G����;��ܰ>�ݫ�k��B�
d���%CceR���̬�����LT��ِ`wfڰ�Ӆ��r��S4���:I)�wuX�|X���?$�*@D(�0F(�x �6>�k�M�!��X�2'&H�I"�9�)�w��h���h�h�ϕ����H�S�J�F����e�Z:�v���rnI3M	4���	*v]J��ʢ[m�6x���05oF��%0=� ��%Ҷ"�eQ-�-��/fھ�J�3+�t���h��՗��167n'-�ޭٰ>��,舅3��j����s@���1�xԈ��@�l���nڰ<��jâ"!)�}�`fs�T��jf��t��ݵ`~���{����6�ץ�Т5VN�UM�Z����a�u���ŵ
a2WC����N#i�ԴV���7XW\��nt���š�n�N��d�����<s�N�z��n�۰88�:0q��{n�n�zn�qAp�ob�v�;v|��`�t�5�m�s��S[v�l���3mJ��;n��Y�5�b�{2�N|�]�ע�h�#�(HL&�¥n6�UY6,�P\�eN�\NJj�PM��	f�wuLɭfh��ܩΎ��ր�.���J��t�M6��I�!DBJ���J��dҚ�Rܶ�V��Lے�ِ`n�� ��\Y⬥y���f^&��Ll�07di����vo�A�PCZ�����5��SYs����O���4��]?4���7(ʕZ!��D�۪l���(U�����O�07nJ`{fA��K�V"�e*���m��ٶ��P�f>��g>,{vՀ{4ZK��%1SG�ŷ3vk�e���Q�k=�S�<񮭀^�䭹��N�9�\�-�]�m��?~� �̃vF���L���Ћ̽h��[�k2�I������ ;𠗼I��0?.��`nܔ�����]e��j\�����j���m�:!$�s+�lg>,f=�*m�Jj�Kr�`jލ07nJ`{fA�����~�`�ʌ��b��y#��w�ՠs� �ݑ���� ����~�(�]��iK�]�6M�9)�.���6�����5�9�#��E�)1�8������=��V��m~���C2����jUp�6)$��h�s���z��k��"d��Ub)�R�n��ڰ9t��vd����07di�{�+bh����u5M9mXtNg_����j��8�{�`gk�U")��UW�fffS�2�05oF��6l�
w6��KU��9�M����]{nf�Dg i�q�58m/R;+E����}6v���rbQE��?~����w;빠r�V���M�ʐ�H�����`y{6���]�`{��l��W�L�������C��G3@�����9]ٳ�DL��Z�5n�� Xf�j�*�f+u�0=.J`n���ti����F��P��S���rO�g����B�I"�-��s@���ʷ{�����>�ݛ �-[% �.Sf���m[�8B�n��p����Ǝ�J��v�`�
�4�C	<jG�f������٥������В�Pn��j�;�J�E5T�q��E&h��9]�@�m��1fm��GBQGmt��S33D�U��Sw�`�y��ۊ�U8���QA��Z{n������ץ�$��s�7_�1�d�[���L]Ѧ��0=.J`n��=��ww�~�>�O+6���&0��Kksy�����\��N"c�ˮ&���ki�c+Ļh+�9�>�j�=�ec�6���nI�;f6��6θx�ց���dq��`-��l�9�!Ծ�KeBB1�=Y�l<Wb���r^��v �^)8I6���<�='/]�v��؎��]%�����t������ȉZ�h:gi��'��ظ0��ww�{��|�;����h3pu:�.u�lNv�z5Z�8��X�c�tan�=w�����ֳq�A�<��}�~4Wj�7di�˺4�%+�fR���`����L�`r�07fA��}'mR��62���r�́��j�ř���	%3�ϋ�]�`f�Ԫ���Sr�ՇBJ?DBJ�w~�7?�@�v���s@=����6�q�x���$���L�09wF��~���������\�q�Hr���v��E��	���:z6�#]]��{���M�j)US%�M��{��l{vՁ�3mX�h��tNI&5#PR9���ڿGBJ����X���ٰ3ww<�R4�r2E&h�z�hVנz\����� ߺ��EyF^Z*�tՇ�Q�*׿�U�����=��V,͵`ݕMP�S���۰>�ݛ�_������r��j�7ۮ���F7�{n��Fr�L��q�eܐ�5�5�*�ɞ�]
��M���N�M�����09wF��1��rS=�R��4��)�r�j�ř���D�vw;�]�`nfڰ͕�4SUEU75M�ڰ��>�ݛ?D(3�Q��l�.��  0D�ARB*�E�TO�������n�/���Ҭh�9��N
'$�:��0;��06�K`v�Up�m��[�d�Ḿ�ݵ`~���
9ww:��?��ڴwхx�Li nx����v��u�L�ћd����<�������bǐ�F�5"$Rf������ǥ�����BK���V���+���x'�9�k�Z+�h�Y�j�L��{�ST�U9�nlg>,��?BQ
goZ�3�zl^�5��HA�R9��=�w4�}vnI����r*�*	� ������4����za2D�r(��4�}u06_J`{fA��#LT9B�e]�hZ��\TEH�d	�7R�7Kѥ�{q8��`��鎼9�r�-�]�m��S�2���_/�A˧����0�cx܈���@�l���۹`y{6Ձ��ھP�%2vW)�&�m��j
�@���s@�w�s@꾯@����33mJ��-�QR܍�j��BJ���[�`}�zX~P��;��+ ��U���"q��H�h��h��,���ٶ�KbP��Ҕ�J�E-՗D��I]1�@"K�],K�mN��]�~%*Q�9�`1����.��u�?khP�PD#�qm"ͨ8�l@� �L2�BR��^la�	,$��I(O^�޾���ޝ===��>q��      �6�    Hm��;l���s��[I��c(�m����UvQ��<\�gl���2GeNiDڂYi6�UJL�a D�dj�m��l�m�n)jHN�ø���΍���k��]�"<5���:ۍն��knD��X����j�i�ܽ �2�%�Ij�v�@j��Pw.�\��a,n�^H�l<xf4���q�+�b�p�U��R.�6B���R/A��kVFeL��u�+�I8��T������.i�:T�e����bt>V����,B9z�T����	МJ��;�-yƥۗ&͹M�z$�� ��%�R�⤞�N�S���b:�K:	q+)�d�b��3��W+�k����<c.zo5��.ga�=d)v*��m�9�Z�8*B��t�'x'c�=F��=���:�
�I�On��J��C����գV6�e���=&�\��-��D�����n�Wl��v
%
�;(�i
��0)UJ��c�8z�wi��\��q,��B�,��]8��,mF�{�����d�&����%i���=q:�L��[r�@�"���FtɌε-N��n;R��Yݬ�-�e��P�MUE�p�1�=�b5��K�آ6�h�=�'St-[]��ƹzި=�v��	�Q��L:ipۗ��ؕ��<���-']���,[F�&rvZ2�ӥs��HӜ�ٵC��R�DH���vt��i�F٢�cvͽ ��r�)��v����UU��56�.�T;VxZە	�.�/�&�uY ���n�fv��`�����5�ǯu�� ��p�A�C����""g6�oC�6�]um� �u>�jބ	��J�u���ⶎ�@m�kh � 	��ݨ�/L����*�Vr.���+�U�JK�c�'Z�(6�&뫛��Qt��A[s[�Gl�fK�fR���ٯ�ੵ�P(�� @J'6 UJ5~Ah�x�'UE� lD*�Q(��9Q���Mpx
}��ֻKs35nk33#x�N��8mN��m�flCd�i횅$�m�j��B�-b��&u �Z8y�db$�c8��\c:{8�z���6m��H5�nH��B�.�� �u���N�j}J�S6v'gsnSa����ͻ8y͐Kf�:/:�����퍻�t�;RY�r�ltݵ�a�kq��5�>sm�花���arn��u�\�is���Ё�峓��dѓ2j��AD��m��ض��5k:�c7�)+�g���٥�$�dHq9���/�zS@�mܰ<��k�P�%	%����`~�]R����̬˼���#L[Ѧ��X{^��	(�3��UX���E7.[�L]?4����d�4�7�e�1�lMȣ���v�S@�l���ݵa�%
qf�����Ҋ��UJ�2�W���2ލ05oF���@�m�4��2%0Q���̉;m���d���@�����۴bԮG^��S�=�{���븚�ڙn���L���V��mX{^��%􇳟n��T�岩Slf�ܓ����߁�J��~؂B6��X���=��W�(S!��ڕ��A�<O#s4���h��;�]���]� ��c������"�>��,��V��mXtDNWwU�Ӫ���E&E#r�n�����mz;e4.��58��d�pZ[�zcM$�t��Nr=A:�����n*z;wR��4��)�r���zՁ�$��d�4�7e)�Y�]�w�Yx��jIll�0;�i��sm_B��ݯ�T�t�R�nF�V���'�w�74 ��$H�*�Q�!,I(j!%e,{j��ջ6��	��'��p�=�w4�}w4{^��(P�(QY���X��ԪLr�V�33/V�i���d�]��;��#�L��2"4сԞ�=m��Fm���7m#��uSr%�7O���_7��sM̲�t�D���^ξ.�)!I
������Kı>����PI�&�X�'N���ӑ,Kħ����5��e�:5s2�9ı,O�{~�ND�,K���m9ı,O���ND�,K�g�v���%�b{];�y�s,hm�uM�����$-���Ȗ%�b|}�p�r%�bX�{=��Kı?{=��Kı=���k��f]Y�.k0�r%�bX�;�p�r%�bX����6��bX�'�g�v��bXE������m9�RB����b�7TMSs-�M���
ı,O�{~�ND�,K��޻ND�,K��ND�,K�{�NG��7�������߇J%�I%p��Q��5^qH!�FooT��������)��L�ɐ骤�`���|B�����}�p�ı,N����Kı:w���,K����]�"X�%����L��h�YnK��˴�Kı;�{�Ӑ���j%������Kı>����ӑ,K�����ӑ?�j&�)!ow�)1�eR��6髅�
HS���p�r%�bX����6��c��CQ5�����ND�,K����"X�%�~;{�x̷&��E�&��ӑ,K?�����6��bX�'����v��bX�'�w�6��bX"؝;�p�r%�bX���ަ��K5�Y�CW2m9ı,O��z�9ı,?�#�����ı,O���"X�%���޻ND�,K�l!'���������������ؽ=��y��Onە4+���n��P�WF�3)C�'#;�`)v��#e��l�Y�����:�m�M'�յ&��ͣ�3�z�n9��K�stu&:HنG�U�P�ź1k�֦�@k��nq�t��{ Ѹ��Kn^a����ϒ9�aN]ۣ�Z畝m���S'n���o���\p�3�6��$�zL���"L�gI-n��w����1����X�<:u[\����S�g=s�R�&�eW\і���9����B���w�{��7������?�ND�,K�{�ND�,K��ߦ��,K�����ӑ,K���S\��2�̹sY�ӑ,K�����ӑ,K������Kı?{=��Kı>����Kı/{�y�d˭[�f[�f��"X�%���o�iȖ%�b~�{�iȖ*�b}�}�iȖ%�bt�}�iȖB����e���6����|B�,K��޻ND�,K��ND�,K�{�ND�,@lO�{~�ND�,K��ߋ�kY�Mf\�3Y�iȖ%�b}�}�iȖ%�a� Gǽ���~�bX�'�����r%�bX�����r%�bX����&L��uLɭe���oN)$6qs:|%�Pm��!xz-	�Ll����7j��{�7���{�����m9ı,O�{~�ND�,K��޻Uyı,O��m9ı,�9�WR�)�S��%�p�!I
HS��ߦӐ�C��*���K�����ND�,K�{�ӑ,K��Ӿ��Kı)����2Y���B��iȖ%�b~�w�iȖ%�b}�}�iȖ ��b~��p�r%�bX����6��bX�'|v�~&e�2L̺�j�.ӑ,K�����ӑ,K��Ӿ��Kı?}��m9ı,O����9ı,N���5�L3.��˗5�m9ı,O�;�ND�,K@�����Kı?w;��Kı>����Kı/~�����285��ŷ3�4g����L6ݬ��Nl��Jݸ�aDc�����hPZ]��ӑ,K������Kı?w;��Kı>����Kı?uo|��)!I
H^ǲ���UHm�l˙6��bX�'��}v���1MD�K����"X�%���p�r%�bX����6��bX�'�w~.��f�5�r\�f]�"X�%�����"X�%���}�iȖ0�@����P_�?��?�ı=���m9ı,O}�޻ND�,K��ܲhɗ2kF�XL��ND�,TB��Ӿ�ӑ,K������Kı?w;��Kı>����Kı/ޞץT��u*�&5-�/�RB����|\�bX�'��}v��bX�'�w�6��bX�'��6��bX�%���=?�
��f�k�"s3Չg t���Nn(�pqh�];l��t�~;��ޜ����Y�5	���i�%�bX�{=�v��bX�'{�p�r%�bX��w��r%�bX�{=��Kı;��o�ɗ&I�˫�˙v��bX�'{�p�r���H��w؛�H'�׽v��H����n'��?�5�������&�Rk2�Z��ND�,K���ӑ,K����]�"X�%����]�"X�%����6��bX�%�}O72�Z�e�0�ͧ"X�
QD�����ӑ,K�����iȖ%�bw���"X�[�D��0/�sq5���m9ı,O����3XkF\��d�˴�Kı?{���r%�bX���iȖ%�bw�}�iȖ%�b}���ӑ,K���{��u��^�OC�v���񛳧+6�E�ۥ�#K�I�d�Uf����9ߎ�w{����w��zb�L�M��%�b{���6��bX�'zw�6��bX�'�����"X�%�����_��$)!ow}!I�[&�tљ��iȖ%�bw�}�iȖ%�b}�{��r%�bX����m9ı,N�����,K���5��Mf��ѓ�m9ı,O��{[ND�,K���M�"X�%����6��bX�'����"X�%�N��������M����$)!I������"X�'{�p�r%�bX�w�6��bX�-����kiȖ%�b{��߁61�754��.�)!I
H[��+��,K������Kı?}���r%�bX����6��bX�'âx���V���lvtA���x�[L�:4�:�,/j'&�j��9�y��F�k��9؝``�7y�OnK�u�NPg��Rv7���@���)\�9U�uH�gzK˺6��Ob�n�'=��6ݩ6�W���_�^�������W������Z5�Q�)��5\v]��8���K�c�絖�nV�ؗj��=9;Wm�Tw���������&�պ�غ�y#��%�&:jZ�x9ۥ3��)�m��c��ͻ]C�BM���%�bX�>���"X�%�����ӑ,K�����Uyı,O��m9ı,K�ާ��r�V�Y����iȖ%�b}���ӑ,K������Kı;�{�ӑ,K������Kı?}���3XkD�d�fL̻ND�,K��ߦӑ,K��}�ND�T������Kı>�{�iȖ%�b|{���n����e�rf�m9ı,N����Kı>>�m9ı,O����r%�bX����6��bX�'}�rɣ&\�u5��ff��r%�bX�w�6��bX��E {�����ı,O�����Kı;�{�ӑ,K�w��Ӿ?�v5�g�U���r�ڲ���ko�^Ç���xх�p�e�e�f�sFa.a��Kı>�{�iȖ%�b~����r%�bX���iȖ%�b|}�p�r%�bX���C^3%�ˬ�%ֳYv��bX�'ｿM�!ͪ�Ė�`�2
06�iO�PG����K\��m9ı,N��m9ı,O�{~�ND�WU5�~�~�
c()���.�p�!I
HRA����ӑ,K������Kı>�{�iȖ%�b~����r%�bX����9�̙5&�.�k0�r%�b�؟w�6��bX�'ｿM�"X�%���o�iȖ%�b}�}�iȖ%�bS�O72�֮���᫬6��bX�'ｿM�"X�%���o�iȖ%�b}�}�iȖ%�b|}�p�r%���b��G�8�6F ��9[���fQ�Mڹ44�إ����muhF���z/�k��UHt�ln��/�RB����|Zr%�bX�}�p�r%�bX�w�6��bX�'�޻ND�,K��ߤ���R��,�2�|B��������r%�bX�w�6��bX�'�޻ND�,K��ߦӑı,O���B��M�m�p�!I
HRB��}�iȖ%�b~�=��K����	��!�@��3Q�RP��zq�Q�0<f�p`IhP��˲%b$H�$���� ��
�j�
�H�
2����`8�ߘ[2�P ,Ё.*�b���`D�q�����(�*B���%Ԯ�Ћ5k*���[I�7��h�X��BV,SC*$5���
����L��M��Ne4$�.u?�H���]�AV�à ��>D�������4�'��ŉȝ���6��bX�%����r%�bX��\U:L��!�Sj�|B��������ӑ,K������Kı/�wٴ�K��>>�m9ı,T�¦�2S�t!S�7����$���6��bX�%���6��bX�'����"X�%�����ӑ,K�w�����?���N�#	��*��ۋ��E�xAP�i$�Er7U��ٵ��.��.e�~�bX�%�}��ND�,K�{�ND�,K���]��@�Q,K�����ND�,K����������۸_��$)!j����Kı?}���r%�bX�����r%�bX����r%�bX��}O72�֭�fK�WXm9ı,O�g�v��bX�'�g�v��bX�%���6��bX�'N��6��bX�'ﳴ�fkhˬ�2fk.ӑ,K?�������ӑ,KĽ￳iȖ%�bt�}�iȖ%��x�u���9��Kı:}���7Z�S3Yr]f�.ӑ,K�����ӑ,K�����ӑ,K���{�iȖ%�b~�{�iȖ%�b}�w�{VS.���G3��<�mu�G�g&��"�6<���[qs�{T=h�Fn�7|�~oq������}�iȖ%�b~�=��Kı?{=��Kı>����Kı'8��Н9�R��Sj�|B���O��{[NC�:���'����v��bX�'����iȖ%�bt�}�iȖ%����s�NiЉ������$) �?{=��Kı;�{�ӑ,K�����ӑ,K���{�iȖ%�b{�����!s2j�2�]�"X�%�����"X�%�ӽ��"X�%�����ӑ,K�����ӑ,JB��̫�Hm���j�|B��bt�}�iȖ%�a� !�����ı,O�����9ı,O��m9ı,O�4��"����w��;����_�l5��-΍��7;[�u���3	�W�xd��2��j&ؙ$�9�ٱ:HMlk����`�ݮԛ��ud�ЌD���]�r�":�V�j�6�`����w͹�n��!s�֍۠�س6�n�0\r�v�IXî8+s��sF9:�qˬ��و9�ܘ������{C�b�=��CK76�k�[��<Im1��[����L֋�-Ѐ���͜�2kN��B�$F��*p�Ȩ\�D�M��ic<���F�t�^(��<���w"X�%����=v��bX�'�g�v��bX�'�w�6��bX�'N��6��RB����e�E'T�ln���bX�'�g�v��bX�'�w�6��bX�'N��6��bX�'�����"X�%�����i��j��˒�5�v��bX�'{�p�r%�bX�;�p�r%�bX�k�����bX�'�g�n�)!I
H]��H4�-��Ӧ��3iȖ%�bt�}�iȖ%�b~�=��Kı?{=��Kı>���\/�RB���8�⩪9�R��k0�r%�bX���z�9ı,O��z�9ı,O��m9ı,N��m9ı,O|eou�Jd̚��\�.N�M�m�bڸ�mb̘��s�m�2E��ںݗsZ�;�������7���{�����ӑ,K�����ӑ,K�����ӑ,K���{�iȖ%�b{����fB�d��e̻ND�,K��NB�:�W��u"X�;�p�r%�bX�������bX�'�g�v��bX�'���Nc5�MI��W5�m9ı,N��m9ı,O��{[ND�� V���g���r%�bX�����"X�%�N���s.[�5�����ND�,K�{��ӑ,K�����ӑ,K��}�ND�,K�{�ND�,K���O#�E'T�m�n��)!I
H^��7�,K��}�ND�,K�{�ND�,K�{��ӑ,K���{��.K�\p�uʹ#N�i-rO.ξm��$�t���#n��F|,�LXf�ӑ,K��}�ND�,K�{�ND�,K�{����U	�&�X�'����v��bX�'����,���uu��ff��r%�bX�;�p�r�MD�;����m9ı,O�����9ı,N����Kı/ޞצ��9�R��Sj�|B�������iȖ%�b~�{�iȖ?�| r'"k���6��bX�'����O�RB���wxM�̔�l���r%�bX�����r%�bX���iȖ%�bt�}�iȖ%�b}�{��r%�bX���=�d�!s2j�2�]�"X�%����6��bX�N��6��bX�'�޻ND�,K��޻ND�,K�_����S��KI���$,��z�4����dw#G5ՏK<�s:��r!���gj������oq���<{��6��bX�'�޻ND�,K��޻ND�,K��ND�,K����\�WW3%�WXm9ı,O�g�v��bX�'�g�v��bX�'�w�6��bX�'N��6��bY
H^ǲ��Ӣ��e67Nn�)!H�'�g�v��bX�'�w�6��bX�'N��6��bX�'�޻ND�,K��߬�u��35�%�k2�9ĳ�"��w���m9ı,O���"X�%�}�fӑ,K��qU b �n'��}v��bX�'��p�9�2�]k2���ND�,K�{�ND�,K������m?D�,K�����ND�,K��ND�,K=�ǿ{�����^����"�ť�ٷn&�J�ꎞ�ݷk�n��?ӛ����p����ε���&a5�m?D�,K�{���r%�bX�����r%�bX���p�r%�bX�;�p�r%�bX���-�ˬ�&I��m9ı,O��z�9ı,O��m9ı,N��m9ı,O��}��"X�%�����fL23&��.e�r%�bX���p�r%�bX�;�p�r%��� CQ5�{���r%�bX�g���r%�bX�͙W�SL�Srꛦ��)!I
H];�p�r%�bX����[ND�,K��޻ND�,K�{�ND�,K����\�WW3%�WXm9ı,O��}��"X�%�����]�"X�%�����"X�%�ӽ��"X��$/Т.I�u~t����۩�J�x��t݊��v�&�����\�톥��<-G:�6K�tv.
�΃��P�Y��k '\�'�;��I��8C=gmN`�,�B#�rN�$0�S��������Z�^��u�6��\�{%��歬�m^y�Q̦%�aM�ch������u�������[lhv�M����:�A������e�od54c�S�"lޮ�l�Mi��i$�z� ;p�{j�N&�ooU��a\%�2����H�k�g<M�����X�%���g˴�Kı?w���Kı:w���Kı?k�����bX�'ϻ�LֳT����f�.ӑ,K�����ӑD,K�����ӑ,K������r%�bX�����/�RB���7�R�66MM�ۦ�9ı,N��m9ı,O��}��"X�%����]�"X�%������
HRB�q��6P�̱�h��ӑ,K������r%�bX�����r%�bX���p�r%�`�bt�}�iȖ%�b_��5�l�]f�.Ys5��Kı?{=��Kı?w���Kı:w���Kı?k�����bX�%����k�2Қ̇RaӪ�!��y��t��*��i�֪�v�-f�i�����D��{��g��'���6��bX�'N��6��bX�'�w���D�,K��޻ND�RB�f̫�)�PSsUM�W���K�{�NB!�!�^;���'���6��bX�'��޻ND�,K�{�ND�,K�����e�us2\5u�ӑ,K�����ND�,K��޻ND�Q,K�{�ND�,K�{�ND�,K���O35���5��.��ND�,�������ӑ,K������Kı:w���Kı?}�siȖ%�b|����ֳT����ɬ˴�Kı>����Kı:w���Kı?}�siȖ%�b~�{�iȖ%�b{_{ԙ���ue���ʇ
�\���n�\�k	qonz�J��eU�_w��}���u��g}��Kı:w���Kı?}�siȖ%�b~�{�a� �$����&�
qϊiԺn�9�mڵ)���M��K�����ӑ,K�����ӑ,K�����Ӑ�,�$)��W1̔��-�p�!I
H,O��z�9ı,O��m9��"�M��D� �C���'�w�6��bX�%���m9ıRB�6U��4�-������|B��b}�}�iȖ%�bt�}�iȖ%�b_�{ٴ�K�[��޻ND�,K����a�D�e�k3Xm9ı,N��m9ı,K��{6��bX�'�g�v��bX�'�w�6��c���}�����j����mڥE�It�u$��t�6y�!u��*�c����ܺ��.��iȖ%�b_�{ٴ�Kı?{=��Kı>����Kı:w���Kı?}����#�:t:n�|B�����}�pr"�%�b}�}�iȖ%�bt�}�iȖ%�b_�{ٴ�Kı>~͓�j��m�6�nn�)!I
HY��ND�,K�{�ND�,K���ͧ"X�%����]�"X�%����O8ff���f�̺�iȖ%��'N��6��bX�%����ND�,K��޻ND�,��E�n&���W����$-�~�*�S�UI�h�a��Kı/���r%�bX�����r%�bX�}�p�r%�bX�;�p�r%�bX�u쾓Z�%�fe�V�\�a3q,���z����7<ݱ��@Mų�Ź�a��qU�������ow�g�v��bX�'�w�6��bX�'N��6#Ȗ%�b_�{ٴ�KĤ.���\!�1Kl�tۛ��
HRB�>����Kı:w���Kı/���r%�bX�����r%�bX��m7�k�&�.kY��iȖ%�bt�}�iȖ%�b_�{ٴ�Kı?{=��Kı>����Kı)���.\�[3S3%�WXm9ı,K��{6��bX�'�g�v��bX�'�w�6��bX�'N��6��$)!I��Q�:tT����黅�
ı,O��z�9ı,O��m9ı,N��m9ı,K��{6��bX�'N��H�#`@�U�|��£7>�ݤB�iX`XQ�RQ�X�R��@`�#�p����ߔ�u�6�5�.�:�!©�4 <1e+4J�0q�R�-�a*�i�H�+4�P��j[�)(A2��4i�"�!Q�@���H��4%�ZQH�yEpWY�`J���wN�v������      �6�    ۲	rR[5����ͭ�{c��n��.Em���1�l��@"t�9��t T�wi�۲���m[�HH�6��'m�{4��/DI�WE��6zmRݩ��.��-g��q� �2�G���f����N�+R^��1m�1��4��ZeV�Vΰ�+����UU�9�՘� �61��%�qu1Plq��n]t�͎p�I�KW��r��QP1-g m�H���J�vƯ�mp+mt�:�]�!s���3�H�+=��@V
��I��Z�]�[R9z�+h�:Y
�S�R�Ɋ�ɕ�8� ��Z��* lps��ۡ]b�Ռ(݌sJQu*ɵ�qձM)t۳��ss�Ji�e�4)�Z�P���mc����V��6ݚ��=<%.�2kr����i%sӦ��-��.Y���ѻ��[�n\�v]�L��R�Q�m��V��p�v$�ݑ���Ɗ$�	�=a�N�=yp=BS��g�%*��\C�F� UR��mU���x�5��]�EQ	� �Wx6�x�dݭ�n���p�V���
��S�q�"bEV`���l�=�7�-eUiUdrTWR��R�(����+T�;>v�3[Q��T�
W(�6w3t�k�:	]�;a�V��'�\�mڗV�%7�6յ�
Ӌv�$�g��m�l�1��pq�e�ln�n��]<6��-��3Z�T��\�F+�\�mSѳ�\��ٷ]M�Q��9&��J���	���4�Htp�.n����d^��U$�c�\Uv�74ʡ�>W$H���Ċ�B����Ƅ�]+4j�{i�6�L=$�]�G���p�i�(vұ��6p�[M\F��#�,��"1'�p��kH}�������m%���J9�����9�۶�ӵi���H� m�v� � ��l���i��ۤ������n�-�{S��:�yƑ�Z�3j�aJk�ԕ�Ǒ]��n�N؀y9
��}�{�{���QR�iP�+��W���8��`��G���F��T;�  USA��5w�hֵ�fffff&z+��	�<���/*���pL�6��KEj����+t^f��v�W���8W[g���]����ù�4�4����b��'/��{w��zt1P\E����ڎC#���5F��� 4��9�1g�l�l};�`�Yn��Jvs���ܕĈ�fG���2�W�z�퀇\�q�Lc[	�l����� &�T�4X�n��nt��|��ky�sY�a�e�їF�	�1�yK�+6�X�6!4����R*��fͥq��w���}W%�R�&�E74��.!I
HRB����ӑ,K�����ӑ,KĿ���iȖ%�b~�{�iȖ%�b}��S�I����Y��2��"X�%�ӽ��!� !D�K�����r%�bX�g���r%�bX�}�p�r'��*!Q
H[�����]Rr��Sj�r%�bX���fӑ,K�����ӑ,���j'{��ND�,Kǽ��iȖ%�bS�k�Jk.�P�����Kı?{=��Kı>����Kı:w���K�,K��{6��bX�'���k��a���5sY�v��bX�'�w�6��bX��|{�ߍ��%�b_����ND�,K��޻ND�,K��I=ugd�������L��Qvzjg,n9�3��)�Ьa��s{7Y��-7|�~D�,K�{�ND�,K���ͧ"X�%����]�"X�%��������oq���}��:�&J����9ı,K��{6���Pࡊ��]�"j%���o�m9ı,O���ND�,K��{�ӑ?��MHRB�}(��E)tʧC���)!H�'{����Kı>����Kı>>��m9ı,K��{6��bR��1�J��e�i�����D���￿ND�,K���m9ı,K��{6��bX�'�{~�NEI
HRB��R�0m���n�ni���%�b|}�p�r%�bX����m9ı,O���6��bX�'��m8}���#춬����D"C�"Ts�T+�5��*��%m���m{�m��p٧�\��5Tڸ_��$)!O���r%�bX�}��m9ı,O��p��%�bX�{�6��bX�%;�����T������)!I
HY�}6��bX�'��m9ı,O���ND�,K�｛ND�,Kݝ�|!�1Kl���e���$)!I7}�iȖ%�b|}�p�r%����J�@�(~�"~�{��ͧ"X�%����M�"X�%��{ڧ1��&��˖�a��K��j'N�~6��bX�%���ٴ�Kı?{=��Kı>�}�iȖ%�b_ӽ�0�sYnY�̚.��ӑ,KĿ��fӑ,K��c�������Kı;�p�r%�bX�;�p�r%�bX�������OC=.��p�ȗ��2��n�����F*rf��um�_�v��0�4ֳS5���Kı?{=��Kı>�}�iȖ%�bt�}�iȖ%�b_���iȖ%�b|���ε���ɭ\�k2�9ı,O��p�r� GQ5���p�r%�bX��fӑ,K�����ӑ,K���l���35unfjk&k�"X�%�ӽ��"X�%�w�ͧ"X�%����]�"X�%��{�ND�,K�Oo�Z�Y��S5��k0�r%�g��Q5����iȖ%�b}����iȖ%�b}���ӑ,K�P��������?����r%�bX����ֿ���]f�.33iȖ%�b~�{�iȖ*HRDf�|��S&�޵`��`nT�߼�o����sr@�'k�h�0uW�b#��C/mF�QT�s���M�D�2��`r�0t����)��v�[��e752�V,͵���C���uwM��͵��x��NFKd�)�R��������f��	L��^h-���s���M�I���L�09wF��L`o�}D��E�A�#r-����?�忹� ��;�ץ��\BQ�6{ΕU6�m�Y"]2��Cv�j�b�l��:LH���]%�Np�V�u�Wc�X�ol'/]��nը�j���O��l�8wl�ݎ�s�c�ۓN]�=T�V����ʤ�V��J�E �a�Լ��ϟ>o��0ݬ��R�<=v�ۋ98�Y��#m۷.m��#
<ڤ����k������t끠靦2�u��d3Y��e�� �E6��k5&��z��\��ɞ&y�벙�ܖf��"ݎ�A�N��d��k#�u�L������L�&0=.J`oti���F��5#p&7&h=l��#����@�?4���`�
�,)^U刬U�����)��Ѧ.�� �I�̙[h*Zb��SM�s`{3mX�6Հ{ٮç�����ީVঙ@�.�3�ti�n����Ll�=������2����b6�ʭ�ҊP9�����] :�;.c(�Dh��:5��WY�b��Lw�0=.J`{di��޻�<��������$�9]�����$�6o~�Ձ˻�� ��]�ߺ���l�$�jF�Z;n�����w��@�v��� IiIxe�a����� ��rS�#L��7>j(��1�3@;�Y�r\������ti�5]P��ς�������8�c���X�!к�����mRάq��C"���0RM�ڴ��j�ř��~^�7{�?wL�֊�kW�]^efS�#L]Ѧ��mń�ͩVঙHm�e��Y�ٹ$������ H	��(uM��""�"=[��M��oZ����FKd���-T�V�s7����>����]��~X_��h��H���9\������ti�{����
�n��LM��u͡j�QI�]f�މ���sE��/<��g��=Q�y]�%-�'���L�&0=.J`n̠��I�$c�s4g�w4��h�ՠw޻�ie�5l���܉�{����L��WI��S���i��"���1I&���Z}����4��	$�z�I/�_�٠[R˸4�C��8��զ.���.J`/��/��/�/Al�hMƆ:��i6�.9����Nȱ��m��p�k�Fv�������k�=3�t0ʬ�Z������.J`otk@3ޫ* �$��� 筚˒��`r�`yu�"|e�]���t݁�ٰ=����έ�`��M�u���JD�jF�Z}���H� �I��%07fPLT�1I ����w4��h�չ'����?���A �N�����!5S�k��V��ma`
�z�X����[977j��')�������u����4]ֺ�,��.w�m���mv .�
��gF�I�1���t= <�7b�i��6I6-N�6yٞwM3Rb�OM\��{qV�L���~|�\\�ݵ��q׵�`��nwDFVp�(���X#����<7F���n�\V���9�u�E.�֤%Թ�ֲ[���C�>���w^����~w�?3w(�YYӫ"��ru��8�FV����ݱ�u�"f��S���;�Ϝj&F�LrL� �����k�h�`r�`�
�)^Ve��+v��f��d�޵`j��V�n��(H�,��4�8�6ȜZ����{:F��L`l�)��K����ah��*�109t�0t���rS�����h[�g�AH"2H)����Z��Fs�޵`b��V_f�T��1��J�箢��ײ2�&�M��6�x��;��E��yS��0�%���K���i��� =���۔u�˙�V�f]f]�?}�vo�+��$�RJ>Q��7֬75��ݛ�d��!�N[��[l�:j�ս�0t���rS{�L��]��X�dn�$� 筚k�h���������1�dX⑘F)$�;��6DD%����[�j�>��`�ߪހ٬s;�[s8�c�M��-�c\yT��N��dó�lj����.#��\ʼ��F��F��L`l�)���R��M2���mX�vՀ}���������W�%27zS�9l��m�L�V��v��fϷ�	�44��հ��H��bH� FO�� �n�V�V	�B��{�� b��Cql���bD @��@�BF! �H�U��R
�
X(�D(F�!��$X¬*�c
�*B,"�K$���4h�t+	*�����jƱ�������L�
A$t���PRA����D�P��������� �T�5Q�����J�5��(�"ji�Eg?	'��e#� V�cH��bBXb�(�t�Ь e?&�
, ��JA �`�14j��tBִ)Ј��1"�c�F ���O��ܵŐ?Jd��?}tp��g9�1�a���+���Aꁴ ���b���A^1X� �"H��D^(#W� iM "���Q�=�j�ջ���VJ6N��R��n��$�%9Ϻl��V/[����@��~E�7�4�"r-ٛj���ow��os�=��6���ӵ��ZK���;e��d�lI�6B�N��i�ix,DDu0���qU�2�09t�0t���rS{�L��7>j(��1�3@9�f���f��nڰ1f���?B�T���X�|F)$�/���Z}n������[4����,r@q���ݵ`b��V��v�BHJ�  LN��M��߮����7��)���j�ś���%9���3��t��� �iD�4�Ci�H�,�����8�h�LVݬ���mVܥ���W#pr���2)6I	�9��[4�j�;�w4g���;�~X_��b�BE#������DB�3{�X��Հ{7]�Q�L�����f�SsS%74���֬]#LzL`l�)��2���Y�LRH8)3@�z�� ﭚk�h~�
#�U����������R����4��`�ce�L�`r�`/�"7��������m�E&�$�C��G�;l�.�$]^��3�i���fR�i#m�^KG��m��Eȗ��I����n�q����h�]��9�=��5�q��n��p��cq])� 7���q��Ҡ;J���U٢AГ�[�I,�@�2	�e�׮[tWc-����v�ě�Ǟ��A�Y�㶝�ÃuX���R�1���̘��[UU�g:""��κ�������w�������3�����j���1r��ĳ�ۧ�`�yF��G��)7=nŹ���R�tKm��W���nڰ1f� �[4v���(����@�����H�~��=_��@�v��ֳgÉ���i�`b��V��f��(Jg:�����`�)��l�������%06\��ޑ����Ɂ�:���l���H��;]�@���=��s@@=�'f"d��G�<uٺ��'!r3d���8��m3D\��,.�e���Ȣ&!9�Ɖ"r-��s@�z���v��ڴ����1I35����w�7�P:TN�PGd%҄��	.Q_����ܮ�>�m��������j7̊L�9���%0=�`r�`w�s��++>2�/2�.J`{z4���4���U��X�4��$qh������g ����j���*���-�7/-9�Ɏy����X�8&�|�u��R�2�^��v�!W|�~�H��rSe�L�0ҖQ ��!1'3@睫@�v�����=��sbGr����l���H�ܓ�k޻�~�����ڨ�DC��P��9Ӿ���=�}۹'��Ζiȣ�$I�h�������<�Zk�h��)b�dp�f��7mX�������ٛj���O����<����G�m�;q'X�:=/���1Ń�m5��H$������)��$��F��F��i�܂���5�@궽����1f��پS!��\әsR�6�Vf^[����H��rS�rS�ֳgÙA�$���]���{w$��w�rb'x+����F �G���?k�ύ�'�߻L.% ��H<I��9�j�?�?�����ˠow�V,ݵ`�1�e7I�6�Q[v63dV@�0ܫ�ݫ�,\0�F�R9�^m�n�H�Qa>#���IZ;e4�զ����rS��O��+3/.�ŕx07�4�ս`{�J`{fA�39�WC��h�Lt�ڰ1f���ٳ�P�}���3w�X/V�[.Tj90s"�4yڴv�h���N,��X��Urd�rS�u.�����.�������Lu�LIo�������?g����`�N��vغ{g�[L�k��3��Ц�ʗQZ�n��[&�a/S�y;��N�tq�7U��l��$mț�SKz��c{�IӺ�`��m�NJV�~q�|�#�׶ϗu�m֨���p���`����H�k 1��u��N����J�N֎�Y�����ZЌ�G�-�ZtlŗŻ&�v	�V�$<rb�b[�lg������{��8 ��~�p��4��P̚��55rt=��{`��Nf���.�ݗ�N^��و��n��IȚ�$��@�o����]����%􇳟�uR�4��SY����Lu�Ll�07�4�ϗؐg�V~��QH7���k��hِg�U]'��~i���ԉ�f]�ffe�0=� ����V�i��;V�Θ?"�ㄑƉ"p�;�F��/�t���6_����̃w��S��8�&
���L�fE�����ܖf��#u�����3��]�����NR�+"�05oF�뒘�J��/��I�������5�)&
dRf��;V�P�R"'@,
 U*��$	d(_BJ��=oK76Ձ�ٶ�=�cw ��Hb�G"�/��@�fڳ��֬mwM�}항̧5YJ�0.�/)��Ѧ]#Lu�L��f�R�4��S-�`b�F�뒘��`oti��R�W�������`�F�Br��UI��.����`z�F�1�}��;�V#Ue�����Su�L�0"�`{<������	$�-�ڴ��s@��w4yڴt���$�0������V�ݵd�%�!%�DE�$�yU���@@�A2���-����@�lAa�H�r'�L�F�뒘�Ja�����������5�)&
dRf��;V�:��F�t�0&���Y�R�YY�n'r�g;���:\Ht^����Ţ�t���{��ԝ�ܗ��%j��I?K����`E�4��\��7`�T�M�-ӛٛj�)���Z�;_��@�v��ֳgÙA�$�Vnڰ>�ݛ:"�mwM���j��~�:\�2f��̚ѭk��T��οߦ��������V�$(Ē������Wu��J:N�uCmӦ뒘�`E�4��\������mr�b����5�n��8yى$"Q��%�ۦَ�n����{rn�k�ڭ]p�L�0"�`{�J����$�����-����1F���h=n��Q'������=�����S&qZO�cQ%$�L�L�;_��@�v�w�L�F�݂��
W�b²�-���	(J{_t��֬Y�j��(�c� �t�`�U.Sm��t����mX�r��/�\03ՙ6�(J�_��_�UW�`AV�*�� ��� �����_�UQA?�TF*A`	E�0Ab#E�!E�P��Q�DX��DX(Q
�E�A`1*(#E�DX�)E��b��DX" E���`��bE��dQ0IE�DX�B
 Q
P�Q"�DX �B
�DX�A`�AP�$ ��E�� T  1DX�DXB0DXD@DYT!E�����
�*�� ��AU�
�W��_�U�AU��AW�A_�PU(*������)��
]�f,�4( ���0���          �        �   @ T�
U)J�ER�T�����  �U!H��(�  P R�  @ %
�8  1@(�( +l(�i �@�� P@��@�_[qg*㻟g^����{�^x �-�����ξ  �7��}㷍_< ��^}�/z���^�����P���[���MQ����W��<�   �̀Q;�Rx��-�NM:q;�*�;ϡ�ҬM]94���H�����r�=���N6U_{� ��J����3_Z��U1���(�UU�U^�v�����uB�(� � ��  P 3`�{�7ۋ\m�nW���-�烛t�'2go���U}�P����U2k� ��}��}�ż����<��\��{O-����ټ�S� ==�&M*�}�_7v����O]��|���(  *E c0 ;�V��w����ק������J��
+��i�5K=�>�>L��=����[���ϻ)͓�W�i�e;�|(>���v�N�zy4������y�@�o=}m�����{랾�������K���TP�(	H�6 �U.���nyoos�����}� � i�@@�@ "P �� � �      �(` � Rl�8� �� D aT4� D�6 iH� D�  z��iR�=L� �"������J�  �=U*M�T4  ��R��ET�F�"���Jm����hL��M�)Tڞ�4�SaB�������������L�̧N�8�nޯ�"���,������QU?�EAU��EAU�aV"��DB�����Jj;����+3���������"��CH8�����DM$�!�K�L
@"|ũ�CB?��ҡ�x�#	"BMn���l����.B�6�Hؒ P�Q�`A�U"1��$4@�hu�6�,Ґ��1"n ��D��
���Iu�63���T�w��R!��$�6��2�4@��$��jņ�9��,��A�ad��$#�$ӣ �du��h�bId�H2o���m5p-��|X�P��i$l&��@���j��~��>6�.�{8M��G�~���$�8�M_���āe��c����EbF�1�Sgƣj���d��CP��Y)
�H����s��S��M��?!� �����}���?r��p���@��Ɲ4����>D�@��"V)~2��4fM���~#I��'�k���kT�k&���ąt|���|$(�{�ֿ}5���bE��B���Z.�)RZ�]���ɲ���$	��#���M: ��u����� \'5�Mi�~����k!O�,.0�}�5�!Oàb5ѭk6_�����"��	X�$��	C��#dIB`P��8�v���J:l��*&�ǀ1��;!�
F����M�xE���ț!��HS��cjqHtC�x?���M8�q8bD3a�a���]^�p�0�M$T�����4CR�>�ы
l"�Y�LM�3]2Xc��.�l��8�BHXP�Xl�A5q,)�%%3f�l�M
��͆ؑX�`:2�f�cV%!�j٥�{�SF*�Lau�7�	tfM�]����1���� ��H@�pc(�` �b�@����G�!iH�64��D�%t�0*�0�BB%���p60)�0�SfĒ5��rIR@��H��B�I)��X,et�D�	
l)72J����{5��ZM�4M��h�2) h"4�"I1t�1$m��D� 2I��ٳ#m�!!�mzA��bq�-�j�0�R�%���
�i,�n�50��@��������$:CCn��7HĲ `�5�d+�Ò�����A܀ƚ�q*����bHB���+
D(:@��!�D�@�����[g�t�K]����?d4�$J���7F�"h�@�D�$��*2�c!CD0,0�E��	��`E��D�	��[I,i���FH�	؄!5e�O�?�.�l�ͧ��c)`��� D��q���+J�	�@���?m��6b@��	�"�D�H�C�H@!����L� B�-���"~��~@�~�� � H�TӉ��r���B}hF��V$ H�!���0P��J� a�{��Lx]B	���� �5ֹO���LO���`�hi$$H4tB A�hd�XGR�� ���F@�XF+a %r UsW��~ia#�7?-P�Ԁ��e�R�hpp�F�1��hi0vH%d4a�dR����1�2 j&���$H�I���� �`��2M��HSF��n�Y4f�' �ču����i�!%u��o�"F�ip6qwI��܈lx��e��|��k��?rk#���@�9�]����ߕ��w�+�P׊�
��D+RY5���"A��ɸ�p�4�9#����Y��J����\7���&)���-Y�k�Ʀ���f�D?( �?k{�}��G��s��p(O����8�Rũ`' ]f��3��nl�Ӄ&���I*�� �Y�(op�A�B��������a�~8c�)�b6���HF*�`A�X$S�ƺ1����`B%�!�g���6pbE�M;�M�C��C��CHn�	�~����CN�	���5m	a��tM���8[�k��+��my��F�SQ��Zn�����tᲁ�L:w��ܿMk� HSF���FY�B�?K�Gz�.���9���)#��C55�t���i *ILۣ.��)�ōt�
�&�0���E�o�(p0�с.me4�ƛq�H1�k6J᳐$*�͒���ԦH����i�0���oY�%�q���T6)�@���@���JE�
�*:p����aR�A4�1�4a� H�� j��	$�p�#4�nBHT4�(m0ٵ �F;ܑ��B�hLh�(i��JÎ�7�𓖑�,�[$	d7]?�:�t}&�q.�D�
P��HB����R[s�4�F͢`��be��B���P*���O���%#�p�F��� 0X�a"p'�3F�a��N�`��ӆ�B��>�A�#A�`Aj�Y"D�`��A��#�Üif��u�0ٹCP���26Jc���(6d�ȶXR����4h7�@�SQ
����$�XFB�i�tH���6m0��L�{�D��WA�Iu��I�?h�7�������f�,al�akter!��G8J� @"h)Q4~Ц�6��7�7��ԂP��;)E�	 �E��`�`x8�m\?H}n<�g����000>@�HA����O���?���ڒ"Ă�)!J���RR!Q��m@�E�	 Q�XA9,! @�	(��)��;
! D����@���b�th�l�$����C�$
!$ijU� WXB�0*FHA��Jo
�F$4����qA �5�H�0��h�N k����U�)�"Z$hK&j[�Ӿ$Hr0�H�HЊ�b�bR
V,H�����.�L!�AHX��`�с�@��C[��$#t`m��U�f�f�'8�`J�3g	ČaH0�
h\�%�5f�B�1���R�ܒHN2��l!t`�
�i~�޸O��6,B	�bD�b�`R	
1	���[��tX�j
F���kCA{�u\!#6sx�̫��l��?���(i�)ŋ
q"�b34�b�1��-���FےI$�   �|                      $                                                [@H                 ��                                                            ��         �j�m*)V�.�j���fmk �m'\ְ -�H9l �f�mt�    ����n�A�� 6� l[f�F$�p���mm�8�� ��m�h �m   � �  m�n�ۭ�$���` ���8 �t�Mt����8 &� �J8��i����h� �۵��`6�s��"KM�mI�u��m M���$�ְ�� �l      7�|�     sm�6�  m�6����� �`�j���*�햪�ڨ	A�!��d�9LA����.���@4(t�v6�Kh 9'h��Y�V/Y(�    qU	h
���(
��h �c��h�:I@I��ҷ`� m� �6^[�Y���e�u��6���m��T�  e���mH�V�� I�m�k�\d$�4� ��e�d̀ ڶ��҉���� � 9�!%���'�U��R�T��Ā66�:޶�� ���� $  � l��mյ���I��V�m��
��	V�aZ�[���V�a�   pM� �j���ZZ�j�����>�߄��mBRڕWe���n���- ޭ9����Y��M�UcB���URuӍ%��ɐ[@ kE�`t�� ��-��&ԫ�Yi�-U.��]�[@۫n�c,��`   vۯJ�kZ@��]�g6��&���	~n��e�-�M��p    �gH��*��l`MR�aYYZ�bKm��sm�_��m� �k�Bj�U�9��lK $���)�!
�PM���� � �n� m�^�8 -KQ��[L��R��嚶�<�O,S�����PI6[d����il.[�[@6ٶ�����Ce���Z��{B� �Iî�����km���)��U.�-|Q} ��m�Hm�;l[NR�hH���ml� [@͔^vh� CgR =��q՝r@�k �[tŷ`h�n@�X` �uԠ-�m��2�m�d�kn &�6�pV� �`:A�l�k�`H�z���A 0m��qr����ȁU��-��m��Z�Z�pUҭJ���4�6�-���@��zj�J	 ,X�mpH��s9UJ:C�WT�e�$&ک�T���U\���M�)�����IXCga�c�UV���sT4�t@UԼ�J�F�y�Um�Rڐ8h�3�Ž���e��	 ��m&�]�	��9��@`��i� 6�*Z�����`t�m�6�N]Zj6�$��EPh��=J��s�T�Ӳ�TI�` �$�4�n|��    l��     <]6���`  ��m �U�`A���
��� ��     9�l��  мV�l ��O���u��[&�X����k�����r[��$�H�c �d��7i+sm�"�mr޶�nY�` $ kXm��
ڪ�u$��  ��$� ��v��08U*�,�媗�5MT�� �Y)5�A�-m��S����Z �Kn[@ l���� l�V�[U+*�5c!]��sb�p���+ �M�$ v�&� =oP/[�����u���Y�-�])i'ZlH�m�oeUT�@��*�WU[j��e�	i6 �6n� Z` �jU��MJ�E�]�\F٦�  6ۀ��Æ�I�l�i�[V��>  �m�md`�k��:I� �Ysm�-6];;]$���l  �[�[@[@�` ��-�Ԁ�Iy���:��^���~����-�m"�#m�����m�I�k��  m���k�  	$ 6ۀ��`�  H p ��$	$ [BM�l	m�FK�}��>� �l  m�H 6�pm�m�m��`���km�`   ����hm�D�    ��8m� p��h����m$��ܰ��-���  ��z�b�  ��
����DP�À۵��4����T��Wf�n�������[�����"��n�[@FE�vݪ��UVV��VM1���V��"Ll�t�J�)<��WU�u��N�I妷69!�� ���V��U���^i6mz��]skapl��� [��-�Fݛn�� -mҭ���5R�iy溕�]`
��"8U涺��eUSSTY�T�ͦ�Y*)�;5[�`�C�6����m�&�:U�;2�*��C����c[H�eY������M�*K� �^�l6ۉ �[w9:�[@	  So�86�6�YF�F�u$!K�*d�m�UV��� -�ց��m $�p$-�t�涀�	E�Sv�@@@R�@U,�G���6Z��  p �h �m���m��õ�Jm��Z�6�p$m��i6UJ�R��@UJ��=�[4��K@6� � 8�>�l�+�@ʵJ��uUHJ��P6�z��\6�I6�Y����jD�m�   �lm�ى6Ͷj��Z�Rvj�.!ZtJ���UUU*�TZ�� &ٷ �  ��[Z� m�E�ŲP6�Z� ���v��n$N�඀���6�   ޜ0 �jۀ�[.[@0��S[�i�&�n�m��p   l �d��	,�� p�nnScZ�� � �Ҷ�5��-�    �cm� I�[s  ��h7m��Y�p�H��Z+j��� 6�@  h��ڶp�ͳl 6�`Kl�.��[J�	6�#tv�o�_�� ��ڐ	     �m�[@�
@@�tUO$a����R��L �`   m"���  -�    F� m�      l	� $-�  7n�vӥ�N����v� 8 m��  �        �m m m�e��ր 	��`kzE�r���-�ݶM���@UU@JH
�m�59�%��t[@ s�J��v���  6�t��2�UJ��*U�WZ�g;Y+ � �  ��;J�vؑ��m5  ��@R����    �b@     V�l	kV���m��p�8j�@[V�-� $m�"��ۖ���dM0m %���d�  9J$ ���m� �`�� �]��l"�=��  m�  @pp$:ޡmAm�m � [\  ���a��H�  m�X�h-�Mm�[�     �   �p8m$�m6["�m��6��$rCm�-�       [@ k5  h 6��^�p���le��H ��   �c�Ͷڷ\;d�j��������Z����ـ�UBl�m� H �  ��9�����o�ݻc�5�$ ph  N|m��h����[j/	mY	(8�i� �!Ӧ�6ݤI$P嵷��q�  �iY�E�ovvZ�M@cMUU[�.�<��#�����3�V�sz�uؔ�Г��o/j���IE.�!r��U ��G�e�$'���sgp�5 �d�OQggguR��G�y�U��<�@Zhפ�ۇ[vٴ��f��[R-ɤE��&Ev"EJ���V��"��ݰ��i�  p��h >��t� pe6 ���l   	���*�
��ʰR�!4�  � ڶ�8�K��x���.��m(M�3m� ��` m��  �m��lq�mm�������� z�m�@9mp    m��m�6H�6�l�a� ��L�[s3332�_������E������?�QP�� �$P�"�X$D��U~�(hT\@ �U	�&E�I �$XI�*� :�� �#ĀUM(mTL
�>��P ����|���qA�P:��x�T[�X��HB��+Dv�B 4�� ҿ('�S�C����
�I`@� �����E�� �P�l Ҁ��T�= �� 	�h(�ϟ�<y�N� tP�TF ��(�P�#�Dv���viTS��'�����D�~����@�lA1E���@�TT>Ut �D���P�����A?�EAU���?�DX,P�F#_w���ֿ���   �        �l  k           m� -�k.�rU�Pl�Tݩ�m$��,ڙP\��k˛8^C�\�Kծ݂4fxS�MT$�(90ݬ�iV�
۝�.4�Z�-Eu{m�݂汉�g6�i��((��� �ە܇cN�!2�4� Z,��:y]���3�V�O��A�@y��ke@dt�[v�2��y����U��@YZ�H{;n�)T��t�B�t��r���A؇��Q\9�%��Ymr�jX*��iV�ݰ!�*�YRy��'��I;<ե��0852��ݰ*����ci
 ��"�iwnzZ��X���=PKl��`v�-qm��gM���:C��Y�ɤU�U����$�f�\dT���6�ʌݥ^�,bR���e�/FØV�GH9��D���Q����]lrLN��2K�Z\i���vUv���/m��������	���9q�4���Y$ ݙZq�N�Lݵ7]�;K8%��v�qے{!;�#��c�n�fwAb��j���6FKm��h��K�	��m���38��F�N̮ґ�wM�Ʀ��	K���nI`Bvd"7McJ���� ��!�W�Y�c�8���xl;l�Z�d��n\��q�b,��4�T˳3�젎�[�b��c�k���X�4��rm;!f�*�5��\�4� �x[A����on'U@)-*�UJ���Y2=`���qL,x +�C8D�h��J'nN���\b8*U�T�� %[u�0�m��/E��B��@©z�g�b�b�;`R�*�@f+��lUT��p���]@U�^w1�[!��`v��ש�V��9�0�z��p��N��-�]����;U���[�����=k�	n@)Ր�g��e�s,�t���٥@��F�ʖ��m$�i,��NՆa�I4p���{�wJ� ��'�P�&{���}�����������  �l�j���Sf�@N�ckd�v�N^�l��Uƌ���t�6�1y��N�,�4۵͹^��l��K3�4�bN��Ғ�:j*�Sr�k2�Y�9��y���vMiBҁb���SՋ�t������S�ݖ�t�L`��*ݲ���2�����ݡ�����j.{FN�S*�����՞�i'��A'[c[��������N�'�{ew.�`\��c����&�������h[�D��4j���f��'{��$�H���7�O�}� �Bz&�X�'��m9ı,_�g��j�&f�E�5�ț�bX�%�ﻛNC�@�MD�>��J��bX�'��m9ı,K���D�Kı/�Ӡ���UW*������
HRB��["n%�bX���y��Kı/�ܩ��%�b^~����Kİo�>�e�SW
\��[�aq,K���ͧ"X�%�{�s"n%�bX����m9ı �?}s���X�%�ο?R��c�[�w�{��7������D�Kı/���r%�bX����Sq,K���{ͧ"X�%��w����Q�v��#[p1�����:�8�BP)�ќ��"��ݠ5
Ӣ�M55�n�"n%�bX����m9ı,O�\쩸�%�b~���ӑ,KĿw]ʛ�bX�'�}�j���.�jY�fm9ı,O�w["nC�'�t*��2%����M�"X�%�{�s"n%�bX����m9ı,�^����ѭY�d���%�b~����r%�bX���̉��%�b_�w���Kı;�u�&�X�%�~;�L&D�k&�e��iȖ%�b^��ț�bX�%��{�ND�,K�{��7ı,O�w}�ND�,K=�����
jdƖ����7���{����r%�bX�����ț�bX�'﻾ͧ"X�%�~���7ĳ�ow�������=����;wVx�ĺl��ml��f
���Ų�/JA�5�]��SkYMf����r%�bX���l���%�b~����r%�bX�ﻙq,KĿ��siȖ%�`���s,���R�ֲ]k��bX�'﻾ͧ"X�%�~���7ı,K���6��bX�'��["n�ؖ%�{�����'3d��������oq���V�%�b_�w���K��b��$D����Ț��w��7ı,O���6��bX�{������F{9�k{���{��"_�w���Kı?w��q,K���wٴ�Kı/�w2&�X�%���Xo��f\%�WVɭfm9ı,O��D�Kı?}��m9ı,K��̉��%�b_�w���K�7���ݿ;���VQ��f+��a��Gg\\X�cf�"�Md1Fժ2>����N1�.Ja�M�˘D�Kı>���Kı/�w2&�X�%�}��ӑ,K����dMı,K�w��	�\5�Z2�ɴ�Kı/�w2&�X�%�}��ӑ,K����dMı,K���fӑ,K����~@�v�v�����7���{�����|��bX�'��["n%� %����iȖ%�b_��dMı,K��ΝԗZ�k)��k36��bX�'��["n%�bX����6��bX�%���D�K���O�<�G����fӑ,K���]M\)r�0��7ı,O�w�6��bX�%���D�Kı/���r%�bX���l���%�by�=�[�T೉&ȺҢ:y+0�\p�b�V���\��s�k�>��wwr�����-�kXm?D�,K��̉��%�b_�w���Kı?w�����D�K�����"X�%�~�{W.f����u�q,KĿ��siȖ%�b~�u�&�X�%�����ӑ,KĿ}�ț�bX�'�}�R�֬���j�Y�fm9ı,O��D�Kı?}���r%�bX�k��n%�bX����m9ı,�^�����֮\�&�X�
�b~����Kı>���D�Kı/���r%�bX���l���%�o�~�I3����s4]k�u�@��s ��� �(��K�"�.��ݫ� H   I��Nf,��0���v|��ݬ����j�n�҅�`}w.�)�/mlfy�b���cnqg��n�u���d�[&갧i��F$ѧZ�]6@�#���BL�s�)��4kWn���1�>Q�+{4�,�������}����6�08j Ḧ���	��cc&.y����<gGG��7\��/��ܶ^Ѣ��m�6��۰��dݴ����&��\��E�*m���7Z
�s=A�&ҘH�"n? z��4[w4kx�IDB_Hl����vU3jj�wJ���6�g�
&M}ذ/���u�ʇ;�jb��s4�d�K`�1��GL��,����m�&$�r�^�{�����	Q�����X�٪�u76�J*f��ylӦ06H�����Il�?;���[�[������L(Ӛ��Q���n�V�c�\KY�f��;�)8�Mb�X��3�w�|�����IlӦ0>ғ�D��j�����`�x��!r���"*�5�X�}x�x�TD$� �=nL&1�2C@�ֽ ��h��h�S@�=Ipq&ҘK��*��9%<�� ��ŀ?kŀj�^�}���`&Ҙ�Y�M��X�I$���_��� ?7x��\� �ۓ]��P�������|�O�n.�֎=��2�h��e����k��`N��ˤ��&06H�x�����ۘL���9u�g�$���7��`�l�i;C�.nɚ
��殰�]�m��R�Q�"(^C �J�]�����;{��r�%��h�`���@��s@�빠r�^�}m��<�ZDH�&��,�`wtt���[ ��$t��;�\���SMbɓ�`<��̱�DZ�j�/V��ûfj��for��h�)���
�{7��<�ȓ��*�����@��4���$�S	pn= �Ɍ	; �����l��R��m)�őH��=m��;��h�נ[f����o��D�M�h<�Jwu��-���w�)BBQ.���}�V7#i��F�h^�@>��ޔ�;��h,�[nI�Œ�F��+�no2�e�jL�����գѺgcy\c����:���t3��??&0$����S��;�v��D�*�swx{l��(V��}� ��~�@>���_��&I�c"̦wGL]%�I1��GLkݖb�<��$�h�נ�������_�@�:�c�6��G�^[ �&0$�wGL�K`Ow����ޞ�������?� �6�  �Eyk�d�Zu�l9!�4���F�*��n��K���eے�b��Mas�b��[��Zٸ�͚3OdػX�7���ƌ�kZ�8���}�q��F�d�W%/jR��f�4;+67\�dE]oY텶�\��l!�uٳ]/&'���l���-�'9O=c�@k��=;��:;];��Ҽ��N|H�J��GM*��]Fet�`�Ӈ���a�b��y����v�p��f�1G�3�m)�ő8������4�w4
�W����y$��N	8h�:`E:[ �&0$� �Yw�E�MU�3j�`^�����
D�s�0o�`���f�����`d���`N���l��WZb$�D6a��)�~������:y�`�w�	�f]]YAB�D���]9�.�Iq�3F�]vT�E�gU.{��'�"X<��H�&�$��^����[ �&06H�ml�����Lpo"Nf�˭{��nͅv��]��]���u�$�S	j$��wL`l��^�K`E�*��S�$x'&��n��u��9u�@>�@�x���S(� ���׋ �"!�<�^��,6��{���߿���qU���m��j�쮪�I�y5�B�b�I�|�L�3ѪQe"i�S#s>�������=m�5��s@=���)���8���$t��tt���[������`�#�h��hw]�>�����4d �E ł��F)$�`0!�@�,$H$cĈ�D5I�LAo� T���8 E7 D$H*�-!i�����D�,Ql�HZ$��Ab��B���)JA�!P�D"�"� B"��]�$J�J� ��n�0�P(/�M�Z���X�����;��5��kh
' �`�`�`�{��f�A B����I��M[��3	�C30؃� � ؊`�����<����u�{[T�lllo��ٱ�A����{�6 �6667�z{��.��5�b�ֳf�A����ｭ�<��667�{�؃� �(�`�`����y��mD�A�B��o��V�k.�$�0�%�wV�q\����YS��m�W��>��v睪�)��`P�C,�������~���}�����rI�����
�[��{[��I)��:��j�mU\�SsWx�v-�� �*��O��훜}}����'Q	}!�Ӧ�©T܄�ՖUZ��%>o�X��<�^��, �Ҷ����%2)3@�ֽ��z��I9�������`0BD�#�`(>�ٜ7$����s&\�5�K3�W��=�1���0=� �ռ[m����?�V����CX��۔��Sۦ�9z�M

`��smUȬWB��R��(�̒I�}�w4��h�נ�1�Pı,Feb��ox�|a�	L�}Հ�_BI}!�݋�Q3��h�R&իUAe]��˫:"!)��������w��<���I$�=���c�6��&�I�z��٘����7��`k�`:Ӭ����*�S�&(ܚ����e4]r�	?������������~?� ]6   `�λ�Im�m�qӮ!xr\���sA�i�-t��.љ1�pU�&69u�YJ����)�k�9��{V.
�em�}�_!� ܡDCۊ���K�?|_w�HXR�Ka9��\=�gY���M�ݴ��ه#����&���rmZ�ٺ�Y��c Bx7��mL�G����f����৅���ڗti���-���i��g�U�nJe���ꇳ�!MCK�e��K\,q7]�yE{���Q�5%������@��+�wY�z۹�z�����(�I�@���`�1��GLt�0�]Wb�A&�)1�����h��hu��-uנ}�n�D�0Q�L��0=� ����`�1��B�(�D�6"G3@����k�� �u����s�bmǍ��1��һ��UD���� =v��o��ң�p<'R��Y��r	��L�9������{u���/�I%�_�}�M��L�.j��� =��-*�	(JH�J*j̟{�ٹ'���M�ˮW��?+�W��cD�LQ�4��0=� ��ҥ�����+�&,Q8A���e4]r� �u����׫I���"����.�-�{zcd���`v�D>c���kdl����VuS��V�u���9�qB�B�������DVU���+����$t���t��ҥ�;��+���<Cd�M����u��9u���u�ݎ�"Q)�L&�.������6u�XZ�J�Q�@��s@=�I���"<�9����u��loL`l��oGLg���cS�p�#��@���������`:Ӭ�yUUt��)m��)�ݦ�[��g�ȷ�)��\���V �24��G64LQ���@��s@����J��&�����Wf
�%���z:~�UT�˥;`zf��n�{:֓q�!�Hґ��9t�loL`l��oGLk�UȢ�m���<�@/��������r
� %E��krN���d�ԗD�4�����,b!Cݿg�r����hvt�)I���1G*/64�#T����g�^y�a�P�d;O\�H����Jb��H�h��h�T��0$� ����(�W���A9�W�����ޔ�/u��=��b�LJa$S"S#�/�ŀ7��*"!)��l���`u9`��1G�A���)�_YM��^�{���v��,Q(%x0'tt��uK`M��N�0$�~  �h  
�V�/$^�M���t�8䱞��I)uӲŃ�h�������Y��AX�L���\��MIlm�X*86�����km����4)wv�iK��!$]��s�3x v�6���k�3�6��펬uF��ZQUyN	g���'�#]QƞjkEq��cs�M�x̗smt3�_K�tL�a5]n�T�`ں�ogg�Jl�^%�wE���](u;��]d�[���,k��ªI`Yte�Ff����y����X{l��)(I}A��, �Dꮹ��*��Wjf���orQ	L����}� r�:�=�����#�����ޔ�/u��*�����hv:�D�)0LR)�GL�T��0�UUR���V�	�hl�9�W�������`u��7�[2��U�D��x�\3G1�a����z烣���<�����EƎ-���b�LJa#�D�G�_[��[ҚW���g!��y%�V��َ:%]�O�`<�V}�s~���Ą�$݀�J	8`��`^�XrJg��,���u+i��l�1�3@��W�_uŀ7���Q
{_|��ʺ���6��LI�z�]�ޔ�/��h^��vY[ncn?��Ѧ8;��n0�\�v�[Q�췒�v4KO�CZ�v�&������-�M���U�@�빠}̨�J%1I�b�Hh��gD%2t�]Xk�X{l�{-&	�hl�9�W�� ��x
""�ـ=׋ ��<�nI�f��G	2= ��h���{��U�@��UQ��h���qI4[w4.�^�_u�v;cm��d�gG���!g���#1s@��m=�v�	h��7aL��puhAkg�[i����wGL]*[ �&06H�z��6�Q�FI&h��z}l�=m��/u���e��b�f91'���1��GL	�09t�lL��1F��f��n�{��}~��nL�c > %	$` A�,�P
��X �$F1�>v���ߟ�nh��~"Q)�L#��^��˥K`M�遲GLmL���������Gl�z3-�DZ�l�'#�d�aݩ7��_}��v�km��6.��dˬ7 r�u`��`m�����C��,ɾ�&�RZ.n�f�� ��r���M��Xk�Xδ� s�.�f���7VZ�j���,�^,9D%2����@�����v�ɂ�I�`��`:Ӭ�^,Q
w��X��6�Q�FI&h��z�<X�x��x�^��$�	RJ�����E�v�0�����$���0�	k`�V��:1j���$� ��Ą���C�J���1HB,P��`�EH�Y�1.
�tS� � b���FaT��1"E�H�XX&�A,�"�4�E! �*B$GB�.$Ą*�EP�� 4Ҏ�0�X��A�`��E�% ���h�:�d$ �`X,H�$�!@ЊA`D���"�kw�    ��        �m�  �             m{M������[���P	tJdB����
ge�U]H� սWF2�K"��ݻk9���Gm��PN� ��6�m�$�]�W9��Q&s3�J�5��o����Ɵm̂�*.�6��V+nWg�Mh�T�vs��pK 6d�QȏN���f�Y�k�ػk�̪gCK+�%v�jڤ ��#�k˳���CS��Q�^5�P$N1l�æ't���t����Z�M/���mpS�%���s�1X|盐���+:聹vu��,�W�屡���[�X� �;r��	Z5"��v3��csU���gce�`��L�H[%�'-������d"b�֣�^)��iXz�i�V�h�)ulܙi���B
l���&�g�iM͢���>�i#i٭g����;s��C�۴$����mr-M�:gL��ת76;t��L 5),m*]5��[��j�eW�)�6����Wu
�x�����Z�b&Pl�p� ��;vl۱��SQ�cuhܺ�v\��|�[��gcZ�ZBwaE\Z��c�Fev��ۍ�g�j�T{W[]���T6$���ڕI�r:bک�HH]u��I5d�5��R��]�lv�;0F��C�>������3�m���&7c�6
6qv8�k���T�9�7�q�1rl��[�LC�:�+�V�t[PR�J��ҏl�UJ�UA�s\v�G�ҩ��t����X͏q�� #SIp �E.�*�]��G��qtX��K;��y��4�����*�R�(��2�#���3ή����m�7���
�mgm/%�vڒ� 6���L���]�9ݪlX���:sā�C�� EqtA�h�f�]m9n��6�n��%VvZ�v.�ZTj��R�P  T=�ghUH~�C�˖��UB*ڠ�<�� C��o�"m�� /7����� ��  k.�s\��9���(<��]�V��z����Dt������r��yd�/���v�fn^Ll�gk�3�������nnn�;�5��0�Zۇo1��+�e�I,�����Lusz�wJm����t\�m���{z�X@tq&�,4��gn@��c.�0��M�M�ۜ�s�=�:��`�]M����%�e���\�S���.��U��N.�6��y΄��]�b,GӃ�:�E�kHo+�{:�.�M+�.nK�EWjf���݋ �o}�s@��+�;�.�c�#�7fSd��z:`r�R�z:`}̨�J%18	����/��h�T�ގ�$t�=�,�e0�]�+�`r�R�z:`l��oG���V�X�0�F�S#�/��h��h�w4]r��X�cR�݇��w`Ԉ�԰��J�%��@<�Sf�YNFP4i�a�������0&�t��ҥ�&�t��԰ʺ-����� ��T(�B_�I"�$(P�	$+���Հ=�f��, ��x�j5�$d�f�z�Y�{� ������ �B�f,FX��Į�1����GLwGLf[4��Y1��0ndru��wGLeI�	�:`��K���9��xMӋ�Lv��4ř�su:�W�rű����R����!p�57}��ʓdt��� ݩq"`�S$�'3@=r٠_[��wW� {�r�=ΜSs*iZ.n�U+��;{�`���ˢt�(��� w���h{*��6���w[����� �Rc�::�<�%�,3& �M��;�2 }��4���u��Ymm��jO梌Cm!��Y쮪�Y��k���g�N��z^q:�A��ͧ���l�27 ��f�z���������eL$�c�'�F�0;�t��2eI�����F�p��w[��^����������H�Jbp%Z��f y�� z�,B��o {�]H�0R�r�����u���)���q���ĩf�Օ�Z{ju�#����ݻk���}���ϛVQx�58����O/U��~�~���m����/YM ��f�WUcm&�"#����;���/YM ��f�z����]��ɂ�I�h���l�1�:GL�0ur�X��!�E2�@=r٠w[��w[��z�M �Iv�@�F9x��;�ŀn�� �v� �M� $$�",�$��bS����� m   ;��ً"�-��A'�Ĝ�X�v\e6�;�J#C�Tq�q�Zs	��hV���cvH��Z���>�FK���Ii��/^�8J�y��@��d�{���q;I�Ãc\�4��4�]q�-i����!Oa��wL�㔤su��%^�W���n�;�1kA{w;mE�d� `/X��gy�K�ݗ�];
h���{��PJ��N}�kg[V7N۔���ۧ��^��B��Kpnm��
ڶ���]&�Ӝ��w�c���X��`�n�D%�}ذueG�$Ҙ��H�h�S@=r٠w[��w[���-0x)�ee�eI��0;�t��2���[�%���)7�M��������h�[4]�VF�i�!H�nf��n��e4�-�u�����mɓ�#�����L���B���-�VT�ɘf���=�z�q�s;V�.�,��nf��e4�-�u��u���g*�j!�E2�@=q��$�*���`��`nٜ�L�iV�&L�F9x��-��s@�s@�������6LM���*�`���<ݳ <�w���w� ��D�&���#��Z���BS����;�b�7[ŀ�GsUWIͱ���o%Q)���l�|����K�t�Vf��D:��.��t��m���u�X�x�7l�>�h��ʚV�f��R��u�Y�!(Q27݋@�ߧ�@=r٠r��m��A1H��`����s���n���h/�6@Y�'��hmI�	::`l� �W(��ve&���IŠ�h���=zS@��Z쵥�,@�dȤf)#mp&VuS�g7g��]&s`&06����N�&Fb�<rh���=zS@��Z��f����{0��1��nf���&��0ړtt����R$Ҙ�Bb�Hh��@;�l�-빠z���{ʪ�0x)�dr\�tBP��z�� �}� ��fD$����}8�ӧ�ʚV�f��R���x�=�`ֹ��n����~~�m˔;l��/=6���vV�l�o<U�M��b�k��<[R��;�	/�`�&0$���������p�-}V�w�٠[�s@��M ���I��bl�O� �1�'GL��`I} �%p�&F#�<rh���=zS@��Z��f����{0��1��nf��Қ����[4z�}$�����8 �` 
���[](�����<;��I�j4:�j
�Zɸ�T�mu�t&�FO��W��c�B�-�m�`�q�]�M˙|vȭj�J��c2��d�8hxu�ٯN�7L�ȶ#�%'����x���盳��Řx��Ӽ]��4��RT�<b"<�v�ӱ"Y;m���@��܍d�=���X��m�r�nzD+�J.4�6G��www?u|i�!��ex��a���-���6�7l8nf�!����c')`�\��b�}s��;jL`I��gd4�E�&1�#�- �e�@�����0$�������0UveD���I4z�h�)�Z�� �e�@��
��Ca�R73@��F��0ړtt����ul�,�����k����޻��Jh���r�i|�,J#���|���V�bҲ�X�t�;]��.<`P.��#d����8� ���M޻��Jh��@:���&F`یYwxz�g�$�EQ����O� 7ˬ�>�\{&(��LCp��}zS@��&�]1�'GL��Pĭ,���C@��Z�γ@�����M ��d��9�drE���	::`zvA�%�LоJ^V]�sۭS��F��b:�^.�:9�+��J덛�S��A�z2F��
��>�޼X�m�u�z"!} �S���+�#ka1)���>�)�Z������;�)�yx9��`�jf��>u�p�s��$�	T""$`�"2�ˢ0H���I�����#��D�&��R0a �*��|+ c �)@��H�,E$AFE 1$ |@���` Z� ؿ�U:��6(�D@����""�BP�QX�,3����f y�V�&6�j$��;����Қץ4���XV�3���f&od��`z_D���{����߿~���h7gٞl�[2R�f6㮥�u��݆f`�f)V��q�f�Y�ncr��~4���>�@�����U�I�1���H�4_T���tt��� �jKU�]
c�6G$Z{�@����n�k����Y0X�DJH�)�gGL�0$������� ��t����LJD�s4�w4_U�z�i䭻��$��lm���Fx��	�k�QsY,�t���`KG�ͱ9^��X���֫-�����~c����/y$���I%�'��I!w
Z�-�j5?�pZ�K�%��Jۺ�K�߳�J�(�$���´L��)����{�%$lI.�=^�IIy�Iz�}�Iy�$���)�np5$�t��y$���i$�VH�䒒6�K�ګȓJcq�JI3�J�(�I-��/y$���I%�'��I"�~����"Ŋ�`(B.O��  �  Y��	]v��p��mX�tfݶ�$8�]�g��\i�^۴��c���az񳭝����>��یg7��⬭��m7q=hĪܙu��uN���D��ڔʗ9������G��ٶ��2�l���a�%�P�ͫ�tx;k��d��6z�5�M�����Q����v?�N����6�h�C��p��~n�wwqt��l����`:��v��Xn�k�� �u�';�I��}�-Y�rđ7GMһ:m���$����RF������$��QjI/��/�)���"RF�H��$���I%�'��I)/ �I-��/y$���X�H%"r8�K�߳�JK�&�Ked��I)#`�Iz�:�x�0_�HG3�J�(�$��KW�$��t5$�u�g�$��ʴȞF6��Rx&�Ked��I)#`�IwI��䒵�-I%^^��$��Eك����M���B֌��],i��k��\V���+�xFɓ#1�#O#��Jۺ�K�߳�J�(�$��KW�$��)rLmA6�����ə��o���@�BQ�u// �I.����RF�����LVLR!�II&}�IZ�����j�䒶�����<<���<�0l���4��w�"m$���I%�ΛI.�8Z�K��!�0X�DJD�H��$���I%�'��I)/ �I-��/x ����U�5�8����fl �hVf�XGB�R������yc#�c���8z�P�IRIw[�}�IZ�����j�䒶���[�`����W��R^A4�[+$^�II�K�O��H^�ZdO#����Ԓ^����-����&�؋A����g{Ü��l�5$��%�*�2df4�I�$�tlI.�=^�I-���Il��{�%_GrL��L�7RIw[�}�[#����Y"��K�6$���G�6y�z�{�5��A�"�ӢcQ���r�
�c=L���i��.ua�2��fW��Kdx4�[+$^�IwF�������<<�d��9��q��KҲE�$�tlI.�=^�I-���I}���6���H�I�$�u�I%�'��I%�<I-��/y$��,���O$�rH����~�}�I.��a�$�VH�䒪���r��I%����`����g�$���I%����%�wCRIw[�}�IU��m�1���^�d���粺�M&�狩��]�qL�A2C*;N�%:k| ��~~�$�tlI.�=^�I-���I-�ҭ�&F1$��K������^�a�$�rZ��$��.I���Fp��$���>�$���jI/\���I.��K�ڕ"M)��7�,����Il��Ked��I.��4�]���|�G����<�0O9I%��E�$�tlI.�=^�I-���V�����w~�???� ?���m� �W��L,Ӯ�v��q,Ⳏ�֤@7��r\�ݱ˪m�$��Q�����]"KI:�9�tT,��M�`��ڻ��l��s����n�hwkr�:k���
���a�D��d�0�`r�z΄cb����aν��n�^{O�%Nq;&�\�q�@����v
�jzwj8t�D7m��r��N99�܋�q!2��c�.3.�
��6�0�:L��v�7�}����r���㞵�R�ا)v9dbY�Vf/rII�`�IwI���Il��K�%��H�e.�5��P�I��IwI���Il��Ked��I.��K��Ԉx�0_�HG3�IzǃI%��E�$�tlI.�=^�I
�m���$j)�Ԓ^�-_|�]Ѱi$���{�$�G�I$���J]�&F1HђE��%�wCRIw[�}�I-���Il����U~����/Yv�,yy���y�Gd���ۧ��^��Þ%�76��+jۥQn�Q��-�� ��{�$�G�I%�����K�6$��9�`�S����L��^�a����U~�_�ĺVO/y$��`�Iv����H��ѓ���	�G!�$�ru_y$��`�Iv����Il��Kս=bj`񸈔�dq}�Iw]�Ԓ]�~�y$���i/��w�S�/y$��������2[�5��&������[o�����$�������$��ߛn#m��-��)�$�03P�֮F�[\�:��y��jW�.�{��}�q}�"k��n�?�Iw�<I.�N�IwF����'��I!^���0��E#r�K����(���[��ə����}��ϩ��:"�m%�*���2dc#�5�|�V�ݓv�w���\T_�s2���&�����7�� ���S�ӱq��m����*���/������2ffwZ�}���IBIR���5$��??�iLn&�"I3�KnGcI%����O���
O�06H�����ߐ��-u�9�m�u�%5��m�]s��7�/�\�R�=������{�:�λ<M��MAuu�;�+�`n�X�x��uz���c��H���׋?�"�UC���,g��`�[0��K�F�dD&9&h��h.�XrJ&[�|`o�`Jju�%MIaQsw7V�:Q3���|���׋�!B���{[ŀ9m�T�]���������ճ �G���k�ŀwY�w��K\X�652dII��1�&VuS�g7g�Y�Y{q`6
��t�H$%�&F28�Y!�}�w4u���u��I}!���ϕ���]7U����=���Q	)��}x|���י�}��$4�7O!� ����V�:Dϛ�X>�X�KZ��H�Uh�Auw��w�g��X�x�?BJg���[ݔMM�����n�fwGL�0wL`l��`u>��T4�l$�v�H�)!$�0&��Cm����I�N�/ ?��?E*@���	]�!)�I��Ҩj��&�(ҜB����P�Do*�`�A -Q�����D� �> "p�`)�7@�CBG����     m�        'l  ��             ��/b]�պN���cr-,Yغ�&�ivZ��s���z�W0n�+��6�^��N���F' ��Z��i���n���i��ی�Jnɳ$�m��jq��*�\8h�V7i	��f��sm�]x�G$�L�P�t���1�ۉP�u�h�*h'�E��ݽ��@p��ؘw�����+�%�q���ۇm�k�j�vo9UL��s��)2mm��zv_IF�vY�ivG�sٶj��D�XB��Z���l-���S�n�v�m˦Mص�]��-a8��wgt;;�i��V�Y���n��橶��ͧv�[WV���6U�˰ԯ4�,k�	�vL���*K;(���4�94<��˲���źv6I��\�X� ��ƕ�F��99��h�[.�4�Zݫv����OQ��Us��b�@.y��H�҃�::�):g̜�Ug��SS,�d[�C.��b�exLSGjn���+Df.�Y��S�k��Vi��P.�m�b3�Gh����yz�<��G�`��֖l�5Kb 6�Ӻ��5��P1�X*��N�U���3&9����P2��u�2<b��� @.�dVyb�p�W]�s���Zb4�)��;p˚�H\�mk@W[r�����C��l�	K&��i^O5U4�km�U73��%P�g\��lq�`Uj��j��kn$���+`6�
C�ڨ z���8۴郝�HR���o*�vѷJ� =�m�pUU^U�-��U�.壝��/F�W������h@T�U*�*Ҭ�Mj<�OS�UR�2��uq��کs��+j^d�ڠ#v�d��ĬY�a÷m5O&����cse����e���;۵W����؍�S��9vـ��U�S�ļ�7IUC6��fx�;;��]nv�ʪdtUT�j�&h���b�)�T��)��?�@�C���z����33 �   i�e̹1�\s�'fDr�.�i��A�V:4��\�'tU��h�e�����m�˷TE'bg.�;T&�al\��C�r�*�lZ�\�(��B��kSd����ӹ�:�s�l�k��(��'9�u��؜��+=�su�T�u�v�l��j�,����W#�2���H�atf�5�q��G�'��Hqm2��1��W<%ӜW�\�p9�[\�s�kn�vJ�o}���ySuJ�ԫV]v�wv, ��ͫgDG�_b�=)�|\��������遲VA�����n���H��e��L#	��آs4�W���ŀn�� �u��7T�(� F8�md���u��=��hw]��rS@=z�H�F�nD�SzGLwGL�Y�������Ͽ@���<��"�,�E�5�e�u�e�۞���n��!��ڈ�T8Xq��ej�f^W��>t�ޕ�`{�:`oH� �R֨�R&�Z&���`֭�����B��%	}�/=� �7� �u��P�DL�M��T�*��]M��+� �>t�ޑ����zVA���Tu7T��J�e�����N�����)�}�w4�vs�!�����e�S���zVA���遽#����P�C�ְ���q�Q ���"HYz��Ƶ09uvp���̨�s�5Z+�`oJ�0=�07�u�� �>���~�Ѧ� F8�S$4��恽#������� ���˳,.�5WS7k ��� �u���"�(��+5�0k�XΔ�sD�3j�榢�`rID���`�0�^,����y�0x)�`��rf��rA���遲GL�`l��P���ue;fڗ[I��1�u��͓�ù*�ټ��^K�I�+����M��&�06H��2�Y�W�5��Y2�4[w4�)�{�Jh��h ��TCM1�D�&h� �ޕ�`l��zGL�]i*Lq�d���)�z۹�{[Ł*9(QQ�}� k�|������q�L��=m��=m��;����ճ �KԹ�UU�U�	��r��*)*$0�\�ml��2�ח��M*[��C,��D�#�M�)3�;��ۚ��h�%4u����[Ҙ�M�$�X��3�I)��W�����f�|�r	���	�$s4뒚����0=�0=[a҅�]]^VZ̻��ގ�$t���t��)�}��]j7��Y2$�4[u`{^,u�f����)$�(dB��G��8 �@  ���d�von���������Z{dבֲtO.�[GV9�a�'�hm؂����N�t��2�9-����:��YvI��N�s�7T:���Q���ԁLm���Q��a�<�vY�e�M�G��ӣ�ڽ��m���Ƕá���4dN��؉X����7�f:��m�j:���I�v��bg��,�ݹ{e�O�{�=����Mm�뭇��:�]X!���[WY���kq�;q��&g����ț�}^ehwL`wJ�0=�06H��մ-R�WR�����7Z�gDD��}� ��ŀ{]��gZ���.�1�2C@��w4[w4�f${��w\��w7����$���}�ۚ��4뒚�빠}�+u�)���2I��@�)�}����=ZU�ldPn`��!��� ��2�E��\8�g��w����d9�-�����\ȚTM���k�|`{^,��/�	B��_�@=�����X�L�H�����d��[��ҲVԉ���,�	�I������^��rS@��w4��er1����	�L`yoK`wJ�0=�06H�&X�a1�Ƣ�qǠw\��>�]������@�/Vۏ�Gcf�B��:m����s����`.��}Lsqv4I9��� F8�S$4��s@�[��|���뒚���0��UrM��=���Q�ON���W�����IB�<�uWUTͪ�������zu�`�[0�I)��DBJ=	*ʭy�z���t�Ʉ�Lp�$�@�jـ}�x�6�`r������˖�cǊdjD�Hh�]��n����@�\����m�B�Pݕŭ��m
���*��ه�ql�mA�y⠰� �Q�Na�!2I3@�[��|�k�=�%4{���;9��h�Ad�7k �|�g%&�W����orJ"d�e<h�Ss5wXO�>�07�t���-�ou��Q6H�8����s@�[��r���rW�(EB ���3�rC���$#Da����4u��˭z�䦁�빠�䫏�A�Ƥ<5j0�b�Ea�Dƣ��b�\�lg��*n�����!r»������~?`ޕ�`ott�ޑ�i|J�(ĳ�H�u�M��s@�s@�u��J(����C�T�M�����v`�b�7[Ň%�ϥ�V����=��V���2�4�w4�[�ͫf(��:�|�H�]wT4ѓAcRf���^��rS@�u��7[ŀ>I(I.쾻�����������  �ۭ�1�����򽍻p� �`;Q�f����,6܁웞�Tٶu����%�sz���ne���m�X��̠ݹ���ֹb����	���6¨Jٮ��T"m�H�r���YD,���4@�����[� uuA{�S��Z�j����2�ڙ�]v�P��ڦ���t=�<�p�ǋ��COd�5q?���~�V�6�n��	�nm���uV�Mʚ�[z�n9.�E8�k �, 䶝��-~J�3@��g�{��t���٠��\�6H�8����VtL��b�>��<ڶ`�i����f6�JL�;����٠zܔ�=�w4�ʝhCJcq6�G3@:I����:`wH�4�%2a1�M�9�䦁�������s@.{�U� ����8�G5�bU���7;�?�����vtr�:�3i\�%���<x�F�M��u��4�w0��_�ID}!����5j��)MZ�-Uݬu�Y{�,I-If�34�d���빠|��u�ƚ2c�J��Xۯ�ճ�L��ŀ7ݙ�Uy��(
a1��5&h�%4�^,u�X���� 7�Ur����F8�S$4����n��u��=nJh����b�O&�(��䝭5�����g�%�E�7gslָVշJ��K��$�mĔ������}�w4[����s@����x)���!Xۯ~P�L�ܯ���,u�X���Ʉ�6dRf��rS@�ﻳs��(�!]hD�"'6� ~��e%�!,����S���X2$��P�H�`� Ĉ�:E�"A��#*���+4������X "$	 ��@S@Ȑ�IZ���"I �C�H�A�� � �b���1`�Z]h�!��R$RQ����M`!*hU$H�@��с0`��H�*J HA!�Gm�@�HAӭ�c�ca�X�Ted	��$�D�!"1I6����Z�Oʨ��t�(����
m��B �*�?)�W���5����;�]� �<��Ǐ�ԉ���=�07�t��tt�ޕ�`z��$�)MZ�-Uݬ��,�G���u���}�w4�[�����Ǔ�;I,Ɏ{y�
^M#�`�]�x�t˶y��V8��Gli�&<q8)3@���h뒌wGL�0"�uwV�,�*�/��e07�d�:`{�:`;����F8�28����ף����J���l]0A�eUU����5�ŀn�f�V���P�R<�X�C���b;}٠{�'��4�7lD�f����Z� �o�^,�BJ9�Ϸ�+r�4��n���F��m�mq=�Kwܼ�r�2�=�]Yʮ��k6&�n�ߕw��<�ŀk׋ �v� �ˎcǊdjF�8�[w4�0=�0:U�LV�"J���*�2�::`{�:`{�d�:�(4ѓ2893@���h�Y����GL�L������nT�ݬ�jـ~������k}� �u��:$���뻻Wwwwwwe�m� m�;l�d�&��C�R���;GP��A��U3���������/8�u���d��յ�к㕱���!gN�3�ӻp��@���㪞��ʼԉE�v������N�	vi�=�����Ĺ�[�X�nwD@뙞!ɛ��%y����"�t�m͏q�5�l�@�:��Nݨݗ����=@�.�՗*�����>C�MH�WV�]r&Va�l9�MR��}>�Lű^_n�u$�m��c�a2C�u�ۚ����u��>뒚�� �@���IKX�^,�׋ �Z�`n�Y��P�?���?��cQ4�I�~����>�Y����GL	�Ĭ2�U�3TIuV�:'ϖq�y�ŀ{u���f�}�{.\s<S#RcY!�zۋ �o�_ 7�x�ճ �7UM�;�L��w"K�*���A��^m1�N9��>�N��z��5�ݳ�9�}$�����&07�d$t�'J�Z���V�Que]� �n�b-%J)qer�Ӏ{��`����we��	�2�b��f0:U�L�:g�O�Θ��M �Ȩ��F8�#�@�o�^, �n�9N�Y� =�ȸ0�#1�Rf��s@;���䦁�s@��J��$�ō�<m8����9j�`�m�tv��]v;��^�,�(ܲ��<)�D��I&h]k�=�%46�w���`�3��&�Y3T]�e�7�d�:`oH遫����q�x�L�H���n���<����Ҳ��!�uw�2���X:��X���ճ ������j4dǌ�L�<�נ{Z�`��`��`���OU���8�xwWg���Ō6��33hqOGI�n,���.\����A���b�rG!O���g�zGL�05t��4�Tel�#s�!�{�����G_߷4W��{�Jhpta Fcn]MU���,ӭ�
g_+� �ݙ�}J�x[�D�ń�f��ֽ	��ٹ'�ݛ����,ੂ'�I$�$�s���>���ʋE�j�f�����=�[0�-}�/��݋ ��u�z�䫘�0b�J219!���LGWnuc�6GB��ֲ�z�@�<�����7sT����,��, ���?$���+�`w�&�U�Z��.�`��`�w�{Z�`��͈䒪��cM��� w�ߦ��������?u��]�̙�c��@�jـn�� �oBJ&w�� 8?~F~l�#s�!�w[��w[�����䦁޷d�$�I$�M�  fY6�k��ָ�\��s�y�`��x���N�|z�Qy-p��v虵��֖Gk��>�t�ˮ@��5k���u:�e��]��N��4\�X��[I�N�c����Xj7..<��c���V.�w$kӪ�O�bc`t.ݙ�6{v1[u�IdA����d��5�5J��H[m�N�-�ٌ�n]I.h�t��5�k5�f�.�	�)���B`)W3[=iԡH�4��"�Lj�ߩBSf^+����U\�v��ذ�٠zܔ�;���>��^Ƣi࣒f�z�4[��u��kx���;�ڮTZ(�Ws4���� ��|`����S-�b��������6�Bm]M��+��Q�!Ww��Xw�ذ7l�<ڶ`�G&YJ��L��$������h�%4�w4�퍶 ƐF�r73I�z�t34��U�>������ls�f�f��w��?pY�����Rg�w���zܔ�;���;���*�N�$�Lx�q8hm[3�S#}ذ��`nـ�[#�$�!�w[��w[��z�M�䦀x�\���f6�v�?(�P�$��wߌ���^�f�n��u:��5O#p�<ݳ �	G�J;�/����X��`ÿ��?g�ko�j^�ڢ��s�G\!�vv���g]�\N�U�:E�v��\�t�����Y�����Ӳl�4�ge��ƁL�H�� ����$�L���{{�`�[0/1ɖ<l�L��)&�ץ4�n��?���P�b&�)�b;@���U T-*�R)�_ ��P�_+�`�� m:jfʚ��]^+���GL�Y��:S@��<t��a1�8�h����P�B�o�_������,�O]+W���W�7\l,4�k�.�k����7X���\ˣ�ƓX��F��9��nɌ	��`{du�UW�}�s��<w��L$�7#NM��4�n�}���{��=�U�1Lj'4�����7� ~U�p脦M�׀~�?�L��b��"OQ9��>s�����ف�,J!*�P�"v��4᝟��S25#YZ�u��Jh޶h��� ���ݵ�^ŭ�,��T�2=j��}�����U�ݬ��ˮ�Z����`�n��Z�"����~���%���'�p��l�/��� ��� ���興�:u�)]w!tWK�3u\�0ޘ����u��A�ղ0�r@�Z�K�z��|`��x�BSڭ����/Ʉ��nF���Jh{����rI��w7$Ã�N"�(�`�Q�UaA"�	�%L\  L
@����4�T�,c4F���B�C`h��@d@�%��X� ]����=׺^�������     �        N6�  m�            ���ݭ���mUWOm�-4�L��]�$ m��)v^��yU�k+U�D���X�J/lX�� Gl�oUӗ�{v�9ظ�\�*�MLn�m�eA7ayKd�!��㶐IIcx�����S�R��BL�̰=���*�؎{[rmT����b`�g� ����*�%eQ��ٗT�{s\p���RM�eeW������8^����Y�x�3��
,O���mT̻y�u*v�$r���g�y�5p2�]�e��#p�&�d���.��':V�wVҙ����[g���f��<�up=*+H][�y��6�sljU��Jp��j�k���b���rgcf�A�&�E��Zɹ��	�E��F��܏B�Sf�H:4���xQ�(ݶ��v����m���{e���I t<E�Uʶ�J���b},q����@��qb�&S�l��nʯtl�]R��UL��t�S�as���v{h�V�y�j�W(	;M� �yz��G�Ƀ�L[�Z��ϭ�E�@Zسۧ����%��x����uk/Yۆ��9'����:ס�E���@2�lke�Y�ge�G�V�6۴.�Q��\[��e�`��V�'\YW�Ŷ�`(���0���	�,I�u˺�-��d��],˦q��*���O'Ugf. ����clC��hkX�n$m��86�]f��֖k61�ج��Jd�R*�Wm�ت��.�̱�l�p�i6(&�t�n�m�^q��/Z�n8'6v%��������iV���RV�UJ��FUݎ6�ݫj�Uzܥ]5Lkd (�qK�sc&M�oiy��˶�ڰ���NLm���`ݣ�Ij��Kմ�wK�;/X˷G�Լ�r�ܧ`�-uNtb�F��s�Pn�B^��5355�r٨]RMO�� *�P�C@�?!��#��`��B�:G�Ƞt�w���{�{������  �   �Itj�[��K0��  �������/`'m��k	]��͵�D.9��5��h�Xp��]�m��զH�ᬭ箎�]���B�K�N�Mk8ֳ�zvڔ����u�;��{��ם�ݷ<�/��v�kt��-7c��g@c�;Fp5�=ssU]��3���ۓ扗�r��S�ؽ�l��b�`���au?�{��s���?��f�s Q�����p�Vv�3���͕���l멹NR�냌��1Lj&�,�8P;��h��� ���/�;]�>sttU��m]�ң.�j�&��{ �����P�d5w*�U!6����U� {_^7�oGL	�}ka��!"�@��M ��f�}����	L�_^ {�W)�*jnQJ˥3V`��0&��Lw�0&�A���ww��N�rλI��H8��2&�����g]<�q�t�&��}�;�b�s�
]��v�}8����m��_Hn�ŀ���~l�#�&G�}�f�3�(� �A�D���!�%��	)����ΰz���d<w�k�a F3�nM���y{��;��� ������b�j&�*�����z[���`�c�o��h�U���PS$I����>�@=�f���M ��4�R�ۍ�r��������
3QU�K�W���㝾��t�ɫ��^�W��ܗ&�����m�����`zvA�zI��YWB!�lq��H�$�:���{���d��{�����\��_�� yL��O���rO�񝛔 � @S��fN޳@��M地�b0��D��V�U� <���m�.�����_�͑�c�	L��^�@�Қ.��{%4�ե�ő�$X�t��[vE�4�Y��z�Yl�i�9њӔ�m�@�l$�cr
I�[Қ��xz��ė��u�u3�҂��j&�)#��˺���M ��4zS@��ɄJd�Lr9�oVA�zI�	; �7�c �:���L�)$y!�u�@��4���BDDB�z����5�Uj��$D�h���{����M ����[��lF8a1�6�/*����k6��*=])���ɺЩ]=��dͻ5�B���0;j�&�?�A�Y��<��3��L&<Q$9&����s��y�^�w� {u�~�2�LS�$���߿M�Қ�3;��4���{��a F3����>�`���7ʵ��L���@��*��1Lj!�$���h�!B���O�{� �� �Q������ޝ���?��� �[~6�  ��W�&iۢt3�<��Tˑ.��@kk������"�3�<��.7����lu�
�����nn5�	�n�Ù���ͤgV0�DAXg�jg�ظѳ�dF��'���s�9�k{:6�kj���&�Ŭ�n�ӹ��l��qD���M��5��v����CӍ�[�x��H\�uͩ��]�k܋�w{��{�ۋP��@������[�EN�H�m��mٻ+#E/Yص��p��0�L�)�q�������������Hl�u`��ujej�f�0�1����%�=Kz[��*651d�H��h{�4+ְ��|�_V =� ��YRR����^S��;j�&�&0��%>�`�p.됛E�Ss2U��)���?�
���t������C�H�s+[u����Va���#�S/M(���&�c�
p�rn�NӚ�Ȥz޶hyڴ׬�fg�-�- �\��	1�܌nI�}]�u%�!BPD*��}xR�� o����Ƞ1F(��8�׬�;����S#���=��8۷U.*��ͩ�ڒM�U��f��v�׮�}��X�%��"N3�@;���"����7�b�7Uk���+n�����uu��s��cY�8ղ�j��\�ݛΘ����sMa5�ם�T} ��::`wU�L�L`;��T�����wx��Y�(��DUʻ��?߯ >m����n�&ЭR��]Z�7Uk� �7xZ���A��� 1rw~�nI���7$�A�ê.�誻��us��(��^�^ {�� �׋ �U�p�\�vE܌nI�[f���s@���hz٠z�%1��F�cg�m���9j�`:m��v)�����n���LmN���w{����4�cxd�O�����ݏ����@>���蚿�b�L�)����7Uk��t(��P>�wu�ݵ�(���rU��M������ o��`�cgGL꾉����xZ��V���������(IUo�߯ ��,uV���QP��QJ*�n��wF����)&�z��v>�@7�� |ۼ�D$��}S=S*�UJ#����^�m��͡Xz:�b�y^���'f�7V�-�ʢ����,�a�&��f��Uߧ 7�� |ۼ�^, �h�ղ0�rAL�- �[4�l�=w�n��9��D�{F����.�*�2����}�06tt���l�@�ir((��#�@=z�uV���w��")�wu�n槡LQ)�%1�$�v>�@;�� ��4^���?���I&I$�I$�  �^���j[�%f��3l��!������k�j͟l�m�[j�968e�:z�-Ŵ4�k�m����k�f��sn���r��J�K�&ʮ�-M^�E��p��h�"�08�nj{k��%]&]Ԅ�v9�q�qg�ѡ�t'k�%S{�t&tv��jd�<����Z[��v��r}��]�.p���ϫ���v�������_|78���BD�,6YR�ԕ��3�s�8�݁��v�r]��Ncx)�&�18����@>���^/���A�O� ռt�eMM�WB�X�1�zI��0;��&�&0��A�Ƀ�Bc�@=z��V�ÔDB��^ {�� �G$�܄a�A���v>�@/����h�@8.��Dcr%28����?��BP�~�~ �����Z���~~~*ʖ�D��8�%kA�����=52���kn�V�	���.մ�cr1�&�}m�{��;��Z}l�=p�1kcxH���f�]+@("��v(PD %��5O� ;{� n��<�j�J%2D�8���~������ �٠^빠��q9��R�3�C�D%3��x��x�x��78��.ljb�̑E$�m���Z}l�-��6�F�(bմ��F^�	L��/U֧�y�ݹt�clgF��9����WV�ҴM��U7w��,�v� ��h���P�DѓA����[�ՠ�� �٠=׋9(�GGU\ԗD��M��� �� m��-J�(�����5
������!����lP���B %�l	E
�D)���	�v~�*�$�(�G�(M%w{�� ڦ� <��["��f7#�h����M�M�B��ou��a�Q9D���iɠ^빠[�ՠ�� �����������l����h���v����\݇[(e�B �.������n�L��]w3j�j�xߕ~�8 ���m�������� 4?��R�m]��Ц�pl��$��:`IW"`mmp\�4�ő�$�m�@��S@��@>��@3��`��!�]�~S���O� >�w�脔ϛɠ|��[D�y��ݏ���l���@��S@��ն��D@.���z�p3vMKZ��J�k�M��O��h4b��zXM9h.+}������`�cw��� ���vb�F3���4�l�ؑ��ۚ�g�@/����1F&#�@���� �=�c ����\��S$Jcp�;��4�[4�l�/u�����ks!�����
!O���u���f䟁B��EG�0u��fa� ր  n.\�l���ӵd,�n99[,u�O+�y�\9�����wێ�v:r�ܔ���|���9���k���)Ӭ�Ibӌ��ؚ�6��Ӵ��ւ��L���At��݃r�a�W��m�2=�zpy�g���*��om;; k�]�24����Sl�t<��>&�Y2�tQ:���u�od[�p+mЦ5��jd�[��_� ������?��U� �{��Sp�Fj�1���*x\�<N��N�Gp玧v���dK��Աfg�>�����`wWd�L`�[�1��
&1�4�w4��M ��h�٠|�؈� <�MI3@�Δ��f�}m��P��n6�br528��٠[f�{��ݏ����VȢ#������h��h��� ��h}�J����%�,�	H�4C	۷Ea�����^zl*��[su6S�Ѯ�������2'&�{��ݏ���f�}m���w���S$Jcq�3@�5�n�Q�`�R ֡6L`�1�����꒳)]%yX\՗*n� 7�� |ۼ?B�3��,�w��=�๰i��&2DI&�}$��GL꾉�{��^�Q�6�`�c�@�u��;��Z�[4�l�;�n�ܓ�HL0Nb��s:�[vWMO Ҷ��m�t�U�]�&֌�"#iLAc�f�ݏ���٠[f��빠�
�V�iF'#S%\����DB��wu��b�7UkZ�vul�"1�܌NI�[f����ٹ� H � �g�5����f����@b��Ba�94wGL꾉�{���&0=;s�S$Jc#s4�}V�}�� ��4w]������n&�lR�h����ETa�ܯ�}��q��Wg��nW��L�Ĝ�D�)�;���4�l�=�w4�}V���R�`�SLd$���&07�:`wU�L�&0
���1��
&1�4w]��U�u�@>����I[J`�����$��o� <�� >m��H�j�DR��Q�;���'O�3�殪f蚻��us�kw��
'����,uV��7V���,�Wsu�l���G�-��Κv8R9�l�"�l�v���F�ͷ�����Кs�k�W�m����GL꾉�{���%�@1Lj!?�����ݏ���٠[f���;�LQ)�%1�$��n��8��xrJ"d�w^��, �;-�1<ĪNb�h�l���@�u��;��Z�Ԩ�4�œ.K�� ��x%���/�mS����������w~���  �   �i{h^l�˪�Όs�������Z���uF{CΎ,���8e���3sx^�9Ք#��^�zv�[J��v[ �md����/\YF1fʝ#۩��"�r��kdGV�sc�C����r���X\S
lR%d�Gl��m���Skjf⛳gtr�v�;B��p6���qq��\����\�s����د�4 �B�8 f�޳Zֲh��n�F��]ף��"�����6��]����ɺЩ,Jd�'�468�Ci�4���ݏ���٠[f��;�h���RY*��`S��?%	%2}׀߿M��s@:���T�b�nE2' �I�vL`ott��[%�o"�Ț#�ɂ�h�l�=�w4)�u��$�&|�� z>��(�U7"���^c�����-�zI�v٠}s�bm�x<q5�#��Lp�.�-:q#�_�o���n�H����ڹ�r����Jd�LmI&|b�ߞ�}�� ����yd�{훒O�����˗X�yl�L~���L`ott��S��=��Tlj ��I$���@�uՇ%
L���pϺ��uT��*�&�WUuw��JJ[}��;�>� ��4�٠|�U��ئ4A29�� ���1����mH��2���]:����[*ˎt����6�Wh�"����C�������^�����Jd�|�߿M ���;��\���@�P�dQ����I4���{q`��8���	%'��I� yBl�94[�s@�U���S M���Q>?~��~��'w��z�Xa1D�H���f�n>�@>�w��P�B�7�, �r}E��)�b�3�@;��oY�z۹�[���>�v��k$bƆC�.�`�r�ƷW#��Y5`�m�5�f�ٮ0p�g�sD�MD�ē�@-�4[w4q�Z�l�gvX�68Ģ��^��,脡D�ܩ��}׀��bK��m�1�	���-��ht��$��:`��X�ŖU]̫Ww8	(�o�����m�?�� �Q�L����ﵩ��nFE$�z�ޔ�-��h�f���+m̒D�6�s"�L�d9�ncQا���a����͛�{���"���0�@��4q�Z ޻�	%�����_+.I��Ws7���4q�ZoY����)���VL%2LQ�b�h�f�7���"�s�0�O� լre�4L'�$�z�ޔ�-�j�z� ���X�651(���{l�T��m� 6��%?�#C�#ˮ���iD"6��"@_�j'��B�b�ec�$$H�H��R7t��eZ*AғD��!�B$B0O�&�n 2p����T�,H5���!4IU��ی[�4��	��#"�0b0`�Q""B �B��6�4aP�p4�� �)"Db�
� ��RF�]�](l9�NM ?0 И��)"�?M��fffffff`  �         ��   �`             kG�©��n1<�WN�-���9�	�Z��TW9��M�W��YچM���m����Ә����W��f(��-�8{j�q�]0��H�,�������cvrb��Uei���;眝�;N�,E2W��=93^1��aV�s�5��=�=��r�m8��%is���W3�&-$����A��T�q�i�Á�J�6�N}����٫���Zm,9�;%]�M��BL�;6�s��+�m�6� 8�l��T�Y����\�,m���� [es�[�"n*�q��E�o�]a��6E�]�V���m��H{v��!'-+�D�B�>�u�]#��ڗ&���j��5�G��W����1-�3�]W0��s��v]=�s��
�gP.@=[V�:F�����ԟi��A���t���{li��WGPgm M+�ŰM&X��;m[�T��#ST�/.)�gikz�\ڹCp2	��"�6-lN�)�1���m=%����S���`�P�t����J�J`�-EIif�5�a��!f�[&R�p��XGX��i-�R��F ���&��j��:nj��*��Xݢ�U�;S;�s�E.�6e�8��m�2�T�b(+�Rٜ�-/;t�x5��dM�ͯAc��]���EU�Ȁ������wGM.�m#m���-��V��a�nm6y�=m,���(1 =��\�
���U*�WR�C�p�j
�[���\�q�k��Ӎ�ֶUek�����p����1���`i5�@%Nwk����ovBm��� �ڀx�K��k9�t[��㝤�b�X�z8(�����Y��v�<���v�]�>���~x6��Z[�,
N����q���T�7S��6��V۶x�U]G6�Y��W4[sE��Dx�J��¡( lTM��i�>
=���u���  ��� *��c�RU5�*,2�n9Ѻ'N�k e�pq�lQ��h�i���b�	��vi@5����W������Dld���1[E�Ӷ[q�Xz�F��꧲@�����W�JgnZ���v�Q�[�ցM$u��մa��p�����lʯ�����O6�y����u�	u�t���y^��j�l����O9z�M~�{�}�w|���䫌<�s�=��F�W #16�^��u�b���m�N��=�\�}����Z�1��ƈ,���?���- �٠�4l��\�/�R6�cr%���p��?�$�D�ww^��� �;V���3�3࿛"��f7#r����ݶa�"&{�wN {�� ��ʀ"������;�S@�s�6��P�&}�׀n��XZ�&��Jjj��uV��?%	O��� �w�wt���ϒ�xĘ�0��Ѷ��Ce�U%���uf��)7`nz^�u�؋��0x��1G�Š[f�}z���4�>�@��Tlh�O�#�wx��y*"�������� z���ͻ��B���n��tԕEM�l�B���>�} ���Lܓ��m�]�K�W
\�����ʧ�sYߧ 7�~� ��}�� ��تFҌnA#�@;�� ����Jh�}V�V{�mǒF�nC	�rTt�R�e�cf�ft�ե��0����uk0�r6E�nF'$��Y�w[��o�k�_H�׀o;�� .mL�*�ř��0;j�&�L`�1���X�
d���rf����h�����%"� ��# D(�AB�
l�yx��, �7G4Z)LիE�ښ���
������}��0;j�&�x�xZ�e��qI4��h���;��� �l�-��6�$80x��	Lx0҈�����Mu����Cclg��'f�5����m󲖲��Zfx��:`v��Lt��>�f�򸒮�'�LX�LRf�ޫ��1�zt��0�'�Y��܆�"��� ����w4�>�@=C�dQ���crM ���x��s�)B��L(�P�YϺ��j�rsjf�T������ �*�9�HRB���
HSĿ��fӑ,K��G��}�5d���t���\{7j���jζ�v6X�T�˹����A::�q7]X�ߩ��bX��;��Kı/{�fӑ,KĿ��fӑ,K�����"X�%�~'{=u0�-�e�ˬ�ND�,K���m9�c���b_����ND�,K����6��bX�'~���9ı,O�ǧ��M]Y��Yu����Kı/�wٴ�Kı>���iȖ?D�Ow=�v��bX�%����iȖ%�b_�-�Ԛ���\������Kı>���iȖ%�bw��ӑ,KĽ｛ND�,K��}�ND�,K��[{�d�SW
\���6��bX�'~���9ı,��ٴ�Kı/�wٴ�Kı>���iȖ%�biD_���ff������l   ���K����8��t�9gZ�s)����q'�m�8�:�ݯG+uیi=�r��etin���ѝ@�j�16�Udx��W79.�خ-,��X��PHX�֖'yc�fU���b8{d�]�F�G�qy��x���<sxV�Ś��0d��c�F�K#�v��Iъ9皮�[R��4,�W��,։�����ER�mP��oZֳE��{0p苲��]Uk�ɧ5��Ÿ-ez��2^��IڛZ�bt�~�Ȗ%�b_}���ND�,K��}�ND�,K�{�6��bX�'~���9=���oq�����tF��Zr����ı,K���m9ı,O��p�r%�bX��;��Kı/{�fӑ,K���ޭ�Ԓe��&�L����Kı>���iȖ%�bw��ӑ,KĽ｛ND�,K��}�ND�,K�{7���fMY���6��bX�'~���9ı,K��ٴ�Kı/�wٴ�K��>���iȖ%�b_���]L&�u�5r�.ӑ,KĽ｛ND�,K��}�ND�,K�{�6��bX�'~�������oq���?e^�umc��It<YQ���v[r�N�����G+���vq�3&��p��.�36��bX�%���6��bX�'���m9ı,N����r%�bX����iȖ%�b_�%�Ԛ���\������Kı>�}�i��(��2&D�?��ܻND�,K���ٴ�Kı/�wٴ�Kı?k����%��-ԗ0�r%�bX��;��Kı/{�fӑ,KĿ��fӑ,K�����"�oq�����~��9kv�G����bX�%�}��r%�bX�����r%�bX�{���Kı;�w�i�����?�4F��Zr�����ı,K���m9ı,O��p�r%�bX��;��Kı/{�fӓ�oq�����_;5>Sp]nܖ<[m�Xi�%�/\�l*b����zW�W\\�F��.�5�e�ͧ"X�%����ND�,K�g}v��bX�%�}��r%�bX�����r%�bX��ٿd&%�2h����iȖ%�bw��ӑ,KĽ｛ND�,K��}�ND�,K�{�6��bX�%������h�Xa3W.��9ı,K��ٴ�Kı/�wٴ�K�Y`�A@���Sf�n'����m9ı,O��]�"X�%����.]kV�1�]ffm9İlK���m9ı,Ow���Kı;�w�iȖ%�b_w�ͧ"X�%�~���=�kSW	r��fӑ,K��}�ND�,K�g}v��bX�%�}��r%�bX����iȖ%�b{��浦m˛��8�棫cMKC���-p6�t[K�^z5΄�ڪp��خ�9ı,Ow=��Kı/��fӑ,Kľ｛ND�,K���o����{��7��ߟ��(Nj;j�iȖ%�b_w�ͧ"X�%�}�{6��bX�'��p�r%�bX��{�iȖ%�b_�'}�L�\԰ֳ5.k3iȖ%�b_w�ͧ"X�%�����"X%�b{��]�"X�%�}�{6��bX�'���l�f\-�WE��fӑ,K��{�ND�,K��z�9ı,K���m9İ181�)���=�{6��bX�'�zo�	��p̚�Yu�m9ı,Ow=��Kı/��fӑ,Kľ｛ND�,K���m9ı,O�_?���w�
�;'-�/,������5�zS����漣�Z�<���.���wwOk�����eə�v�D�,K����ͧ"X�%�}���ND�,K���6��bX�'����r%�bX�:�ӗ.��p�jd�ffӑ,Kľ��ͧ"X�%����6��bX�'����r%�bX��{ٴ�Kı/�{g�&�5p�)�s36��bX�'�w~�ND�,K����9�ı/���r%�bX��{ٴ�Kı?k��{3R�j�K��f�&ӑ,K��s��ND�,K���ͧ"X�%�}���ND�,K﻿M�"X�%�};��nf�njkY��32�9ı,K��{6��bX�%�}��r%�bX�w���r%�bX��{�iȖ%�bT)�'w���=�����    M��[۵�[����H�������D�	ك+��tg�:C��g��ɶ泼	�Qy��HpjX��M�U���:;P�란k<��Q�����In\��\9uAx������R\��x�P����o$���d{)�2l�c#\�sY�ݢ���&ܛ�'T���9N(���p�ک-��%�+���=�{?��������w�w��C�nQ�%�5/P\�gM;V�R�h���:4�%�vx�'S.5k�f�f��,KĿ���fӑ,K�����ND�,K��z�9ı,K��{6��bX�'��ݞ�V̸[���5�ͧ"X�%����6��bX�'����r%�bX����m9ı,K��ٴ�ı?w�~�L.K�d՚��fӑ,K��s޻ND�,K���ͧ"X�%�}�{6��bX�'�ﹴ�Kı/O^�SS	���,��˴�Kı/��ٴ�Kı/��fӑ,K����6��bX��O�o���9ı,N���.]kV�0�ɬ�ͧ"X�%�}�{6��bX� /�ﹴ�Kı=���ӑ,KĿ��fӑ,KĈ�ݿ��}���"q.�9��;k��,�z��LY1ZV���a�#�֮fpI�>�}��$�w�w�bH��ϻ�M��Kľ｛ND�,K��_{3R�j�K��\�m9ı,Ow=��? �P���D�K��m9ı,K��ٴ�Kı>����r�bX�%��ﭹsR榵�	33.ӑ,KĿ���iȖ%�b_��iȖ%�b}���iȖ%�bw��ӑ,KĽ�l�֦\.j�Z�-�ͧ"X�%�{�ͧ"X�%��{�M�"X�%�߳޻ND�,K�｛ND�,K��wg��f\-�WE˙�ND�,K��~�ND�,KQ���]�"X�%�w�ͧ"X�%�~�}�ND�,K�N��@z�f�fR\�.j���qqc�X�s��"���:�0W<����ud�5��O�,K��s���9ı,K���m9ı,K����r%�bX�}��m9ı,K����S	���,�33.ӑ,KĿ���iȖ%�b_��fӑ,K���ߦӑ,K����]� 
�bX�|{�.��p�jd�ffӑ,KĿ{�ͧ"X�%����6��c@��? |DaE�0�� <|�l�h�B;�A(��`�`Á
D�I(��HB��h!�*D�(d����> |���b@�V)��
B��b��A�	D��4#BM! ���鈌 ��iH4P!D���`DX�Dh�Б2�@@iD$��|ڰ"�D! ��X@$dD�X�H0B$HD�0� FF��*��))��)$!�
��4���?��ED�TH`�"��"m�蛉ϳ]�"X�%�~��ͧ"X�%�~>����kF��2浙��Kı=�{�ӑ,K����]�"X�%�}�{6��bX�%���m9ı,O�����Ժ��R�%�6��bX�'���6��bX�  �w�ͧ"X�%�w�ͧ"X�%����6���oq�߿�����%V�d��f�Y���r�/i��S"���P�ю���F��չ��fB[��iȖ%�b_w�ͧ"X�%�w�ͧ"X�%����ND�,K��~�ND�,K�>���2�sV��e����Kı/��ٴ�Kı>���iȖ%�b}���iȖ%�b^��ͧ" �bX��w�g�[2�n�.\��r%�bX�{���Kı>�w��Kı/{�fӑ,KĿ��fӑ,K����^f���%�-˘m9ı,O���m9ı,K��ٴ�Kı/��ٴ�K�逎��D��ND�,K�O{Ʀp�L�&fM�"X�%�{�{6��bX� #w�ͧ"X�%����ND�,K��~�ND�,K�I����a�Z[MkT��O]eD��-&e�ƛ$�N�FT�e�vٽX��8w3�.�T.�Ϫ�����7���{����ͧ"X�%����ND�,K��~�ND�,K���m9ı,K���}�5�\5�e5sZ��r%�bX�{���Q[ı>�w��Kı/{�fӑ,KĿ��fӑ?�P5^w�����������q�w����,K����ӑ,KĽ｛ND�,K�｛ND�,K�{�6��bX�%������չ��fB[��iȖ%�b^��ͧ"X�%�w�ͧ"X�%����ND�,�B*&�w����r%�bX���Կ��˅�Z�Y��fӑ,KĿ��fӑ,K�����"X�%��{�M�"X�%�{�{6��bX�'��{�߳33333333h  ��e�F���碇�g�عQ�%�`7��4�(s����f��՝�R��<�xw[�m�����6�-�n� �n�9��]\<Ұ��;x��>�b�+n�b������j�lX�nP5�grf㶆p�Y6�[��]�N�wX(�U8�l�i�J�K������9E�'��#�v��<����*w6�5�]���������?��U/lX�aI4��f���g0j������:�d�6j������~{�w���{���?�p�r%�bX�w���r%�bX����iȖ%�b_���iȖ%�b~�w�:��fI�In\�iȖ%�b}���iȨؖ%�{�{6��bX�%��{6��bX�'���m9ı,K�;��Mᬗ$��6��bX�%�}��r%�bX��}��r%���5Q;����iȖ%�bw����r%�bX���zr�ֵn.�Nffm9ı,K���m9ı,O��p�r%�bX�w���r%�b�b^��ͧ"X�����?8�vT�Y䖾�7��������"X�%��{�M�"X�%�{�{6��bX�%��{6��b�ow��_����K�nH��d��
5he��OlPr=-�!�5�+Ik��]5-�[�a��Kı>�w��Kı/{�fӑ,KĿ��fӑ,K�����"X�%�{>=�.f�njkY���d�r%�bX����i�x� � *�T8 /?D�,K���6��bX�'}�p�r%�HRB���
HRB�鮎���ޭu��s3iȖ%�b_���iȖ%�b{�ߦӑ,K���ߦӑ,Kľ�}�ND�,K���l�f\-�ZԹs3iȖ%�b{�ߦӑ,K��}�ND�,K���m9ı,K��ٴ�Kı?w�םYr\3$Ѣ��d�r%�bX���iȖ%�b%����r%�bX����iȖ%�b{�o�iȖ%�bt��~�F�-�nκ�9��Ա�DQ�:�aLݣ��v�ݳ[t��c��s��ͧ������,Kľ�}�ND�,K���m9ı,O}��m9ı,Ow���Kı:w�ח.��p�u�s33iȖ%�b_w�ͧ"X�%�ｿM�"X�%����6��bX�%�{��r X�%�|�ΞԗZ�]k4j浙��Kı>���iȖ%�b{���"X�T:lP4n&�\｛ND�,K���m9ı,O���ײK���.]k%��iȖ%�b{���"X�%�{���ND�,K���m9ı,O��p�r%�bX��Y�Yr��Mfe!na��Kı/{�fӑ,K���ٴ�Kı>���iȖ%�b{���"X�%��ﵭk5��v+tcZkj'Q���bbB:gjq����M�gcy\����
�.���AW����bX�%�}��r%�bX�{���Kı?{���Kı/{�fӑ,K����oƵf\-�ZԦ\��r%�bX���iȖ%�b~�}�iȖ%�b_w�ͧ"X�%�{�}�N@ı?w�םYr\3$Ѣ�a��Kı?{���Kı/��fӑ,KĽ��ͧ"X�%����6��bX�%����0�-�Y.Lֵ�ӑ,Kľ｛ND�,K���6��bX�'��p�r%�`hZ��D|�����ND�,K��g�.]kV�2�4�ffӑ,KĽ��ͧ"X�%��������ı,O����iȖ%�b_{�ͧ"X�%�������Wic�9^�Emϩ8�����zy����G9z����b�N�����.5�ѫ��fӑ,K���ߦӑ,K�����ӑ,Kľ�}�ND�,K���6��bX�'�x��j˩��.]k,�d�r%�bX���p�r%�bX���iȖ%�b^��fӑ,K�����ӑT�,K���ڗ3Z�55���5�6��bX�%���m9ı,K߻��r%�bX�����r%�bX���p�r%�bX��{Z׳Z�tf�l��e���r%�bX��wٴ�Kı=����Kı?{���K��f�k���ͧ"X�%���z��5�2�n֥˙�ND�,K�{~�ND�,K �{�6��bX�%�{��r%�bX����r%�bX�w���w��;���?�� -� ��K2Y��a]s����јtݹ�c��]�(���[�]=��ѱJ:QYj�4u���v���pp7;`b�n2���wN����ҧ��kQS�ニ��Kc��XD�2�^t%�:�/St-��=q9��qO4c�R�zy^+7Z9-a�I�>�v�� �۲p��6;X��g=YӺUf��sq��2�|
��u�/5o5�fjML�au.���q�tݦ��Vc(�܉�gU.�+Z����m��YrS�4h��2�=ı,O���M�"X�%�~�}�ND�,K���͇�(��MD�,O����iȖ%�b^����&E�k&h�s&ӑ,KĿw�ͧ"X�%�}�fӑ,K���ߦӑ,K���w��lK����^\�֭�e�i��ͧ"X�%�}�fӑ,K���ߦӑ,����w���ND�,K�{�ٴ�Kı/�x������Y�W5�ͧ"X�%�ｿM�"X�%�����iȖ%�b_w�ͧ"X�%�}�fӑ,K�����Yu5p�˭e�̛ND�,K��ߦӑ,K�R���m9ı,K���6��bX�'���6��bX�'�ﵭk4Mk2�����3a�쮪��p�k��\Y�Xd��s$�c�Ѯ)�(Nj;K[�w�{��7�����iȖ%�b_�wٴ�Kı?w;�� ��j%�b}�o�m9ı�{����W��J�_{���oq�Ŀ��i�|&DC�� vȜ�bk��]�"X�%��}�M�"X�%�w�ͧ"X�%���z��Y�pֵ.\��r%�bX�����r%�bX�����r%���b_w�ͧ"X�%�~�}�ND�,K�r���%0�&�̺ɴ�Kı?w=��Kı/��fӑ,KĿw�ͧ"X�%�ｿM�"X�%�~;�x�	��5�4d�˴�Kı/��fӑ,KĿw�ͧ"X�%�ｿM�"X�%����]�"X�%�|{ڷ�2�]ú,�Ņ�k6Tj�i�b�MX-���vT��n7Hβw��޽Q��Z蹼�r%�bX���ٴ�Kı?w=��Kı?}��m9ı,K�{��r%�bX���<{R]j�u�ѫ��fӑ,K���ߦӑ,K���w��Kı/��fӑ,KĿ��iȖ%�b~פ�,���R�ֲ۬6��bX�'﻿M�"X�%�}���ND�᠟��12H�$bA�J�K�O�"A2'�_��m9ı,O}��ND�,K=�������9��-o����7���%���m9ı,K���6��bX�'��p�r%�`MD�����r%��oq��E�i����h*�����%�b_�wٴ�Kı=���ӑ,K���w��Kı/���iȖ{��7�����?Z��C���[u����nP��OG7f^��B��
�nm��T�tO����Y�f�f\-�ZԹs3iȖ%�b{���"X�%�����iȖ%�b_}�fӑ,KĿ��iȖ%�b~�_>���ѣY��ND�,K��ߦӐ���j%�����ND�,K��fӑ,K��{�ND�,K�w��&E�k&h�s&ӑ,Kľ��ͧ"X�%�}�fӑ,��������"X�%��}���Kı>><o�n�n3Y�Lֳ6��bX��%��}�ND�,K��m9ı,O�w~�ND�,
� �>2&����6��bX�%����������Y�Y��fm9ı,Ow���Kı?}�siȖ%�b_}�fӑ,KĿ��iȖ%�b{��浭U�.�:"0����yv�
jZ7'VT���u��+�>Y�0<��F�B��}�,K���}ͧ"X�%�}�{6��bX�%��}�D�,K��}�ND�,K��j\�j���k-����r%�bX����iȖ%�b_�wٴ�Kı>����r%�bX��ﹴ�O�T�K�����f�]ud��e���r%�bX����6��bX�'��p�r%�bX��ﹴ�Kı/ou�/�RB���xQ<����3j���36��bX�#b{���"X�%�����ND�,K���m9İ?�I�����ͧ"X�%�������%0�5f����ӑ,K���}ͧ"X�%�7���bH$����pI���͉ �'�"����"�����*��PUh����*
����*���*����EB*�B  B(�A@
	T"���B( @ b
1Pb��	E�P�BAa	�B D(@�Eb �
1B" T"�1B( @��T *�B�E�� T �D � �! `AP�@,AP�B�"@�D�@�E@�@ ��@�E@*B  T  �Q��W��*
����*�PUh����EAU�aW�T_�PU�EAU��W�B*
�� _��

��PVI��G��N�Sl��@�����d/���2��U��u) i�`4 �*���v�m@`�{� :P(%D#�J *Q �*�@
R�)@ � (+g��D`>�|x  �s�r�GAMdo��}�v�vh�l���do�{      �� ����{�9�t=����P�����T46���A����ztkC��5����3��A&AO���}���^�4�k 7����H�l��Ç� ��F��������\��|.��t�A�����

� ��
y�'�AN�7�����G��X44}�:;�н�N�=�=47��$ h�<(:=h/{�C���A�����Q��Yɯ���\+��N�A��p둬�
��B   P !�$�MCS�b  �hhLE?��J�I��2��4 �a4db'�UJjji�F	���� 0� �S�j�	M*�4     HHe"MLM2=h�!�OS5=�ST�&��`      J{��?T~q�������̥~� 4�'�� X����Q�������l_���[ռY�l��6�	�7���s:����ٍ�,�>�(r?*�}zʿ�}>���������"�c��p6�pnA� l�@�T@���"�����@o���f�|�3� Ȣ�Ȣ� ��EC�-����m�@f�e�.��9ww��e������ͬ����{�ڻ����
���9�9���{���ۻ����������{��s������̻�ݾ���{�훻�www�wwwwwwwww�7ww.��Wwwwwwwww��wv���}wf�����������{�����www��ř����}=����^�Z_����������>k���aq��7UR�j�驃W=��G�w��ײo4��8w��K;CǍ҄��'�R���u�O<�z�FF�^:RJiI����o�s����@��;7����gb���{;�(�aY�fۏVc���5�&���
Y��yg�6w��T.xv��2%�H���m���I�Xbh���Q.L].��ٚ��C��N:�����s��y�K�If�)In�e�Ąh��YY�Ӣ�'��8��xx#�֝�Wq�p�b�FA^ӧ���-�!հ�V�^s8���l[Y��,#�227f��mki��-�-�a���([HU����DHB*�M'oiښ||-�!
�aK
U�:{{�An:;0),�6�c���HPX����Wfh�E�[�����Qf�h��%Q��a-%fh���Z0��&�F���;H�E��Y���HU�����(��YA*�%V^:;@�ޱ��S�uz�;:/���<��B�9u��rpY�,��;0�5ca�Z��PB���L�$H�
*�04B�cK(��/;N��u<�-h�u�8<<y	y4�����K댺$�=����n���G5����tZ�C�8s�'j�-�g�^��sܞU@��	���$�0�Wlg}}����4�:]u^vJ/(�����t�(�8�0 Sy0֘U�CF��w։W����H@����5�YI�L�
0��
 @�"PGhx� �����[{|�@J;��ﳣA�0�0��,��B�h�BŘ+@�J-!j�D�:#���Qf"@��-��m�"����čXb)�E�:�^k��lk
aM$��X�щ�a$�+2�u�٭gi
�4��LaNA&�5�3Z�u�z/"��N���BZ�i1�c���u���-"Yu+��h��xE��:��� �1H0��IwM�0�Z,'Z�j�z0�Є�)ѭ�ִ$���xy�arx���V�:5���1|9��B��C�%啲�uxy�tB���#xe:$zaA#%�:V[�F�$bPb�Sy���Z�%^h&k�'�T�,�X��,��g&�e��MAtj����'U�H����1 �%��Mdk��6��)K)e]�ꦼ,L#W���!����5��W |u��q�� �Sm���H-hh'�hG��jo{{�	����
���uk��ӡ������5��F�� ��"o������@v64����l�88�3{�u݂�4
@���r�/{z�n��G1����l
X�d��$i	��D��e�E�IV��S�.:��r�ӛ",�C���m���!�ɠi�n�0k�)�ǭT;�޸^�o�mƃ��K�Μ���[�ی������Q4$i��%:�Jq P6�I�ILB�U"]���^�!W0*�r��%1�tj�æV��B�b:J��h�U�=1��������}��$oV��-d(�ѓ�qEu߇s�w��h�Ӎ	��a��%���Y/u��T���a;ʰ��a���4^��h����W���B��&擫nj��9]",��¼�e������Z�z���Q����-n��gY����2k[sY�lAi��f����r+�nuy{���U�C�����c��Q��;:�#���t��	Ǝ;m	m���ᠱ�L�m��h������8Zg3�i��c��㤀D�qt��abA�����C
�th�A��Rw��=}CjPY� �is]�޼�����@�A(���f�:��E�:,��-�a��՗�F��%U掎���G 5�,Ņ�+�i�ގ�F�@
:��BNc���t�`ڲ�ǭHnw�Kx�(2�hCf�/)ͰiG]g��Kγ\��i�f��[+��1-[�&1﹉���i���:����ޒ���Z��$#R�����l|:��������/�����g�}vV�E��YU��$t}���������$�I$�      ��    m       6�	� m�l              ��                                                 :ɤ�oJZ�Cfy+`��w�����8qM�p�m;8��vŵ��a�A��nt�e���RT~*�ʩY9�p�\sv��Vm��I�A'�@���ljޮH�m�6��IkT�[h�&�sk5kr-6���km� m�  l��94�, p��v=`Uj�Wvc�$U���6��q��   �  m�m�zW��^8��N ���-�$m���z�IĀXGe͖մ�`$UmUmVҭ+���Q���]T�eyVs$�R�� �ۜ� H-��R�A�ij�8�hi\�U���o����i�[v�hmqÃ�A+6�l9n��&�L��t�*�S!=<F�U:]�7�*�r���q@U6  X
���˵���IA�mmP%�p��@��X.{v��l%������N�q�9c�'�"Nm�u�NX �6�v�m���PЄn
9�%PUU ��k�k�#n����`i��B�öU��cb���xr�h�Ŵ lO��  �. d�U�C�����]����m������q��ހ7i6�� $m�p �6�l @�	-�n �u�knp���� �	 $�<��"Kh-���!���� ����� m�m��pn��ח� յ�ۀ	8�m -�UT���g�U�@UW��   4������z�[F��� :�f�ڀ_-X�U���g���m�[s�y�Ĳ��U�׷�U�<�iM<�lv�\1;��]�v�YvZE��%��u��kjB@Am�o	n   �  ٳl$�I�q�� 	m ,�vKҗM�`,��޲{���� $C�l C��,���ŵ �譶��Am��*:�u�Pʂ�1�y�#��J=�@#mz[.$r@ ��yP�6�mH��R�� Hm���z�[6-�I  ��m�  E�Z^l�d��r*մ�{8.
��nl]e�-�� ��Z�����a�.#mf����
kt�N� !��l�T8b���mp˷��L	   Zˣ'D�mAC��Xɵ��RF8��[@[KgS![4��J\֒m�����L�:��ۮ��[x��@��   MKNsm�6l�/]{]n���88-��p�dI�e���[�`�kX�o ���<����P���%� ���mRli�	 j� પ�Z�`9c����F� p�$:ս�E� �9��ٮһ&v9��5�@t���$m[5�V� m�� �_o{��Mmm m����V��U%U�o�`�kѠ�]v��m��o 8Ht�H�iX��6@������m[@�
�R�T�2�UWP�v�wm�M����]g�o@q�m -���e  �am�t��Z��b�T���h�	�ض� m� �-����|(U�X��R�>25@  okw�ŭ�[q p e�6݀ ��[@ �.�m����W�� �nm� /Zݼ�[d�l��Hu�#	9�I�6Z     5�6٭�@ $  $  -��$m   � ���m�l���Y}O69m[M�-�$ �H� �`�$2�T#���IR\&���<kpn�  ��[@�&ꭁ 6Ͱ	6�zSa�' 5UUTd�`8-��m� m�m� ��^��l �`$�	�lh:-�  [@  hH   ��` 4P �� 	�� �  �mm�    '%( 	 �6�-6K��  ���I�U^CT�Kۯ�J�'���@dg`*����ɍ�9H�V�'Kv�)\  ol��r�m��H�[�U�5nE���  ���%�bCv�� !�` l� �m,[�m��ZHҫ��͜�d���J���c���W�&n�y�U٪ f�D���:PH*�d|���!��Km��2e�v��Q�7n^�y�������s��0q�f�n]�C+3$�eIy��H
�� �z�D�T���_����ۈ�(!�%�R�Ʃ˚�)n\�\��DP�����s�n�+S\�-�,�n�tY2���A=�_�v"��(���m�&b6c��o6��'�yY�y�p<lc�3+�h`*iJ � :���AmAM>�� ��B(��ҥi4+�C}��� J�O;Q6Øx6�8u��;g�&@�H'�	�O �7�D6��G�3�{1mcw�ʰz��{ax��sf��mf�Ԉ��m�MlD� AmTҭ��Aoq�� mPڈC� �!4t(�x����u��<Lw� x^�o|������
��������r*�����򪪪��*���������*��dUUU2<����������*���������*�*�������*   o������ @�� +���jO�{�����g�w}�9[�D�H`�rI;J�ı��R��B��W��=��Л�]#��v{��1�'���  m[6Z  �         Ӳg�S���j���c���X(2ـ�6�x��U�݄�-�КՔݻJ��U�;�9�}��v��d�]�`6�w�Ȳ�Κ�#��ȅm�3�\v��U��`Ņѵ�m�� ����кL�J˱����d탪�u;T@�Շg�(������l�8N�G�]�:^����-�,�n3g�Z�i���4�b�՜Ө���]^=Qpt���-#���+,��Q=S���T�A�[yˠ�{��]7������s�-���S6Y�3=	y�w,UV��2�1���&z���t6�na66BYzJu��Cq�����D�W$	���e��n�WXiI`�ݷPt�;���f�[d�lHm�l���%6i�2�;]u8���i�َ��چ���
��$$:uq�[��N�e^�5Mʇ"��#'@��M�Jen��Y�*�p%sGB%�qD�`STK}��z��YM��ݖ���W�D0(�ZiS�CO�x�`(x���t�w)�YW��fl �\ܽ��.��NX�l������v֢�k��%���k�d��r���ڃ'W���9�G������cY��K�N�Ѭ��������ns,e�U���}�;y9�i9=1��--��Sk��@�e2>\�*�����3���>��Ъ�3:ƿ�eޑl���냼��X�e�=�c
-Uݰ;ޱdv]NtX��N��m��u����2����ݰ.��`Z��B{�3���td��R��q!�(�@j�pq��X����̍�o{�kD��1�`! @�P�  ����c�G���&��\T��b��^����a��,�Z�v��O,�t�d�JCy�s\u��������3e�m�q�Hh�h�jF �R�n-3wn�ݺ��cdk�$I@╫�+����V�˷�@��l��ܠ�uwn��r(����j��n����]�FdiG�wn�އVi]����@��
B�Kh�$oV�
�2�"l����s�Ϛ�i]�wl����Q=t�4��5v���w�E0b5��9�:�uf�XZ�,��7���[�Q=�4�*:8���5c�@�u�w+���.ͺ��Ͼ���Qkt3�\-Ѻ��e��ٮ�V�k��s�����]��owQF�5��5�rUطBq";����ҍ]��y�Vi�\=�
J:�ۮWo���Pgw��$��"��<X�X/\�@^s�Q��vkl|�nw�:SIK�ӧ��<|{� �0 ��<Rup��\�GC���\{[#V�ukμ��5�+�+���(vY2�q�B���r�m��;Vpt����P�nR��g
.�&/e 7��� \u��6e+�Q�ܰ\�#��!#f'$�I�"�1*��uB��0*��]�]���ԓ.�M�{�=�D��������k͜3*�����`��Z���w��&�w�5YS+	������w��.��j=u7�VV]�a2�{�]w݂�~X.�.nk[�n]pM�Y���ϪN�D�(d�2�iFuT*��\����Z�v��쬹�.��w����A-�)�Iof�G}�c��s��	vL��.�-u�X���s~Z�z�y�]ɕ=
,�^�G���_^��^@]���RL����v��]��K1�
�V�́�L���[��v�W�a����c�5����]�v��7j;��5�{��ɆT���9H�ߖ���3@κ�[�r8�������T+|� V���ȥoV�y��Ys2�ViG~n�{��Iw{��oee̹u���`��
�n�j;7����>obU�%dhݐd���LQ��,� I��VhUi��
������\��T��d���]�/9݂�)�"�º�I��Z�9`�y݂���`�߆�ʬ+*�w�,��݊i<���X/}u�نV+H���_V��$��.�ݨ����SL�d�˦�]�i���8��������ôNs�799�q������PN�ی��Fj�Uݰ��o�P^@{��,z��J�Ys�Y`�ߖ���G{ݠn)::���VI�z���j;�����c�M��W�ު]ɕz�]ڝ�s��k��SW�ɕ����� 77_|F�-K3��IaC,��[��h�Ym6"�{p^3�WLm$#�W��z^8C;7O�^�܆���Y�Ks��y��v�ǆj�(A�+3�.%Mxx�r��{�pd����-q��A!Q���F�^�։1�V��]���w`�����.w��̪²�z����/pw�Q��`�k���&aYZE�E���(�{�]o�Q���.s.�@]��Q�}�.��x�����yrfUV^�w�ڥ���,}�-�v��S��%�d	dR�V�8��e�gT+�SIFc-FV��\4*�۪wl}N��®L��.�D{R�/��G{��w�-M�r��5r�L��9j=�ݫQs��w�+]I2�ViG~n�|���wk{��N�܆eV5�`����[ݨ�{�K��rrz�^�ۘX(D�l�k�1A��Fe.c$6�,���ֺ��y�X.��Q�}wXe̻�u��T�מX/9�E�@/��W�3.�/J;���<�/pT5����3�w9�����9����u�9(�A � �V�j�҄�f�*U���N�+h$���ҏ�
�N(���)���V���Yl��vL�%��ڳ��"Q_�H�'�����N��t@ �����V"�N('�/۾���qB��_�ZIO^�Ys.]e�j=��ȇ�
�7�Zd��9h�W����®N���r!�=F���y�Z��sv���L�)��el�e2� �	�_`ܛ�Ù�.�$*�I��=�����ymSf���]�w��e2�L�S)��2�L���e2�L�I��eL��?�e2�L�I��e2�L�S)��2�L�S)��e2��׾ݲ�L�V�e2�L�I��e2�L�S)��2�L�V�����L�S)�e2�L�S)��e2L�S)���L�S)�8�)��e2�L�S)�e2�L�S)��e2L�S)�Ϟ>9��]�˿>YL�S)�e2�L�S)��e2L�V�e2�L���gϟ;v�e2�L���e2�&S)��e2�L�S$�e2�L����S)��d�L�S)��e2�L��e2�L�S)��g�8�e2�L�S)��d�L���e2�L�S$�e2�L����e2�L�I��el��nL�S)��L�S)����S)��e��Ͼ]��v�t��e2�L�V��L�I��e2�L�S)��2�E52�����S)��d�L�S)��e2�L�)��e2�L�S)���)��e2�L�S)�e2�S)��e2�L�)��e3����e2�L�I��e2�L�S)��[)��e2�L�S)�>�]�e2�L�S)��e2L���e2�L�S)�e2�L�x��{��]��y��e2�L��e2�L�S)��d�L�S)��e2�L��L�S)��e2�L�)��e2�L�S)�el�S)�y��l�S)��2�L�S)���L�I��e2�L�S)�ϟ>v��e2�L�S)�SKmL�S)��e2���|��>�o��y�-��e2�w���L�S)��el�S)��e2�L�S)�ĊH$�H$�o~rh˙w��$�L�S)��e2�L�S)��e2�L�S)��g����e2�S)��e2�L�S)��e2�L�S+ebm�}��f��n�U�QWe�u.��&���uٍQ�x�Vi��;��S)���L�S)��e2�L�S)��e2�L�S)�>|�S)��g�q��52�L�S)��e2�L�S)��e��}w2�L�S)B�L�S)��e2�L�S)���L�S)�9�S)��e2�L�S)��e2�L�S)��e2�L�u��}��L�S)��e2�L�S)��e2�L�S)��e3�=�|�;u�W9�^L�S+e2�L�S)��e2�L�S)��e2�L�|���L�S)��e2�L�S+bA$D�yo|�#�r�y�U�&�ef��BD�A���r�r�y��N����1[ݼ�#�~Zs�oH<�<����fhG�圊��v�a�+1
f��f<� �<��H$�  �Nv��9zKc�u���[�ٹ:ge8���KnZ=Ė�������6z��_�i'E�cBP2�yK3ԈUmu�����ΤFv��,�]�y����>���-:��TJX\��6�d8Q~�o'n��zڼ���)��딣�r�s[��I3
�Ҏ�.�ը�{�^s�b�]sɆ�w�󔣚���P�9j<���s��/.V^�y�X/<��\��P^r��.O7ʬ/.XX/9�Q�"�1U
���*���h6�d1d�J�#�*wDY
�U��k�h�(�k��99�Z{��S׮Z�S�W���L��v���z�\�`�k�j>���@��b��I�UY�D���X/��b�">�/9@���eV�`����"H�R�9��y��*L²����QMuJ;��{��wߞ����C2��q\6]�]l)G6�f�1�ղs��^rq�́C���j�n����&iG�r�z��Q���Qq'��V�(��^s���W�4�5�<EC+�|�P�{l�*����@�1M
����Ρ��!��Ώ1���eJ�CZ۬ �3�ϓ���E[fQYe�n�d��f�]�噕@r�����]b�����.%f84s1���C3s{]6�@��Y���uwlo{V ���.��z۫�c�n�1�x�Ơq����ηޱ����$۳H4�l�F9��\��eф׵u�2P8�Q���5��f:����(�F(�0��<
�c�]���6�(��Y�w�u��0�u�bR�u����*�U%�%)Dfc5v�ݺ��,��6��� tɥ�-MnѦu�ǳ]��^*�8%CgnR%5cQ�[r2������f��p�@���x��B�ڂ́��RՖ���7\�J�����M���_vm�;7�9�'x��s���9�ْ���,��l��w�����0)E�g�9�>�.�3�k|�3j��@�u��a�cY�q�4=��� 9v �Y�3�Ġq����c����h��-��M�h�gV��WNor�oo;q�`���R�.����n26br�R4�(�Fb��+3�*�b;Ht7v�� Qcْ��?x��(L3 �� ��J���`2�qW8�uv�t�ߠ���$f*�C��zu��OqV���Ċ!H�"��-�-�n|���z�
g1�43��}�j�S<������wy<(P;5�!�y�����3�lY�m|��B���u�y��8�l�+ذ�|u��r��n#���hfc���Yó�����r-ȭ��En��V�cFۆ�",H�
& �̝$�`\9��#{��Zohfc��cZ݈ ���1s����a�/X�.2D���[�z}O�ˬ��Yy.6&�{ 67���7��#IG]�~=5��k:��}B����[��7d`Q�M�If1��"��b�k[B��]۩|\E��������f���#���F-�:�zŚ�X{��X�FC���c���U{ޘG9�t 2�ǉ5�!������M߲~ִ��9�g_{����z�� "�0�a�Ѥ��#�R�����2#��g5�˗��kj,ss�q�7{-��8$�3����di�.�X�:�\4ĈEcă���$��Hac#��'F3�b�%�"�u�t�3��b�Yg��Zŵ���,k5�.cp#�N+.Nk�$7	y���'�\�љ�#;_��t�ۺw�vC   }����            6�zڕ���aF�M�Ȁf�CdD��ն��v�sn���-(%m�r��lڝ>����v�:�π-��&�ݰM�AV�s��&J��E]C��y�byu�A�v��N�����TC�n��6�2S[� [َ<�m4M��6uu)���lfШv5 Zu����a�m �ͧ���|�<j݊ت٪� d+T@93��W�(]�+� ���Ϯ-��B6��3,l
E�v%�Ӫ���^�X�̡mc�V��r��b���9�aNcf�c7��Z�rk��*��+pK6C V]����Ⱥ7n�n-Cޠ�Ԝ�fnJ����s�%�]Iz�t�;��F2���1�KP�n�јy���Ӝ6ɱ[o15��چ��/IpEmu�uqO<�[f�n[la�r��:%�ԤKH-F�n���VW/+s�] (�c���.�7��bS��N.�D2��	j�U�sJ��*����:_��S���D=
�H��k�;�Fw[�ɔ` ^���R��*FV�4uV��D�r�{l��F��ۥG�U `n{�oPy����+��6�%فD�uv���&i;r��i�M���6�-����;*��0�Z��w�c�I$ܗ
��<�:���Ζk���[�q�}$:��M�Bdf 9�&���Ő#�R4f��3r� f*g�h�ciGWvٜ\#�P�b�5�`^���3�4���6A���n����[(��7��������o� �ĄE�l�U�]Z�hƱ�g߿w�{�xp����x!�����Z��1͗� ��τ@�����>�:��5��HL����1s����z� ;�\;�w��#MM�ί��0����&�di1s���q:��\EǬ=$R#!��j��f!32Vo��Fb*9�d��uwo���;e����!��1��r��~�����{�c��*hz��{��f�n!:;b��s���uΝ��bR

'� ��1Ѧ%�f]��V�|���˻|# ��0�Bdf 3
�rT��0�%�E�F����Y��0a���
�1me� f!�:(
��R����8�>�������:��5gm��w3	���*��x�5P�D_�OL�Q�>#�C�ۯ{�a�Ά�Qf�fd�@31��� ༄D�q�v����u�n����[Mo�fi�'/ ��vBTh�b{uwn���������=}��Er�����-�q�:x�Ƙ���̭͇��M�+YDV�9�Tc���Ul��.����q�]���5/A�`���G����b�����fˀm�o�X��ZV�
�c����A�Ϻ���l�j�rk�3��[�S!�	I��"���^J��p|@�@3��d1�ܕwo�G�x�y{ν��^QD�SC{b��Ù���|�ʵ�=�9�:��z ;á�$M�u�w3�x^�IH�J�
Q@���MP�E����F�ǵ�ϖ�Ma�C3o[�8!���ʪ�T@��=���@�9�z���@{�M��{��'dt��[<�̑E���u���f�[��@��k���1���c�B��N��A��D�6�H�[iZ�;<�f�Z�[����>�z���\��Z��;m4��ϼ�7�^���A�sGE��s4o{��<�p�S��UM��5����q:��u���z�U�����P8�<G�s�fc��`M���M�����v��P������@Ll�]�7�Wv�55���(�9���j�+��Y�>��d1����u�]�.���d)E5Vk[B�v{~�٠U�9�s߾s*��P3��k|��{�C�_���=��(��$�K�
y�s�Հ��]V�&[��w�u���}�q��q:�fAMf!����7��-�5�!w��fc\�3&FL5����]۫5!�9
�f�ݺ�z�E����tq!@��   78�v�F��9�t�C+�:��p���[KWnd��#v�ru9�n�cg�P�\�̳1��)�f�������ݲc@j�	��M��X�δYX���n�s���&Rw1@���1�j�f�gHcM��{�u�^.�^��d�R�j�ֶ�ݺ��S3�������c��u3Y�b�6"b����a��CF���u�Wx��t�b�c��^�:W�*-��m�*.�]��@�4#P8�^5���y��cc|�3.L�9^ᴠF �A��Y��SY�̑��ƈ�z��]���ِ��i���5��f:�m^!J!5Vkh]۫�b|���$���A]�:	�ɿ}޶�J�5�!�m׽ￕB��Ƶ��#��{�u뻕��w�#0\n������ާ�Z�go��{��w��{��r�o�R	V�7%�$U�\�j-T�x�����m���m�il{	}��{NiŎM&ku��=wk�$¡T%G�����rӓY4<.\�D"H�ԓ�ɭl�CYm+H�L`�1��xO�Њ�:P��@�DA���z�꟒�{�x����=sV��u��F�qj�k[B��]���A��G㘆��8s1�#� 7�ޔM$$��!V-��k �)��͙[X".D����9v%x�b�1�m��̕dp�P��s|W��Rb���a�o�fc��bο����ei���������~-��YZ*���ow��|�{��{�Vj���V䄄m@!5��Q�ⶶ�u$=8�]ۮ�^9��owx�1@�ݑ��Lk1���0s�X �FL#�1s����}�������Y��yn��m�v̆2ʎ�� �Y���ޕ�  к*�T��O�����$�I*��n��f�k�r��r:˃���B���z'r;�[��̡�<z+�b�6A��rT���7�*�u���0bݲV��)i��Z�T3�L+��R��OW68]r&�~�I�%���!_�y�E��i����8�S?e[ނ�(�p�7�=�u���$���ƛ(i��޶����vv8"����w�uf����a�LaE*�߁'����Z��#Q��ox�f:��3 �0��fS��Q�1/l^��,�Ѽ(�HɅ����"��Y�w��!r#4.��|�U��{�^5�v���Y�d1��zWH����Y�+�d)E/b��P�C�T{�zB9��4�ZG�|������4���{�K���QF���KMv�v0���}�����n��b��X�#%]�J��9����ΣP8�6k[_�ʡd�P��`�',(��Wպ�:��rd�Y�Mm�ݺ�\���H\Q�N���o���k"	���� �	[��:���ƻzµKQ�JF�3<5w��f?|��d)����Ad�W�u���ƛ+H������}�ҼkX<N�x��Q�����:���@�K~\��`b0���u�,�.�ַ쾦����(D������G!u	��F�F%�8�4��31�u���PA#&�Bkn��՚}��!r#4.����Vj�{n�P��n�����C�+7�x��!�a�oL]۫ж>=u*�I$�U�[	'''�'�����e�*�W*���Fyr�c���m��p�wl&��xspW@�̳l�:^8���m��,�
"�$��yzv]�2�.�9a�$�����1۶���=20�gj��l��]����zvK[L���M�mB�z�c@�u�m�)vi��QvD��]v/i�ϖ;����}#c3Ga(Zx�UQ�`�5���0��wn�j��u�w��&(Z�>#|C3���s9�2j�Cz۫�l�4�{2$!��J!Q�f(�B���m�d��8�#631���ܬ:��s����cee��/��z ���9f���Q!}��/�2�P�ֶ�w_m���Ͻ�6V�#�@ }�9�:��ĺ�)a�þ��Qhfc�?�U����^�0�<�J%"AR�ᆚ����X��9$�M���u�Y�]ۭk�6!�S�Ug(P��
��3` K��PHc3%j�𣙮����G�����V\�ԛ��fHL��PC���]��Y�3˴d1����cU
�a8Q1ff�'t$��Y�v �:�c]H�)*���T�9�rrW��ֻ�'
$��I��	7w!$��]ě+H�%��UT4(
�u�	?}��'�h��蓙��o�!�EP�l��p�Iz��8Z*)ݢz �@�+3ZԒnT�rT��`���՞�_Y$����@�z$�(��*�R�d�̐��������;�w2e͍�aڙ�U*F��]s���T�҉9�sZ$�d�UU�x�I;�vZ��9ܓ���Sg��M�2I�V+kK8�ʑ6�z$�ސ�zQ�*�	I��1#��FB�Q�P�	x�I�D�̐�UA{��$���dI�R�;1#���7!'�􄓅]Y�o$��[�w��{Ξ���{��w`���E�B�Ġ��Z�p��96���Zl�,[e�����Y��'8s�ss��s�TL�M*�5����r����ǀzA�K)��妺���vl}_=��??  � $�            T����έ��٦�v{!�1�S��캁�`)C�J�\����ܴ��kv{:�u�z�naY�m� �6���\�c&h�1�hxۋ��	��(*���ӬY�0)c
�R���^�����gI!��Pl,����AcL�f�Bq=�қ���`t07<q�ʹy�iyo<y2�Z\)l˵t�
���5A�nX��&/EY�*kg����]�lU���[���1�A;�#4��ڍq���6ɭ^��JvD�\k��mZy�����7h�Ћj�$��b�+�,h�YVˁ�@���@���+ �X,x�g��4�I�k��b�.n�:(��*T�K@7-��LM�P	:�M���
����g�ܗE��n��5��h�,NZ	�ym��U�9�L�$����Y(��H0rUNC�Z�1k��]������2���-��Ж�tn ��h�ˍmK.;���ߺ�J�$gڮe�IY!R��Ѣ��e�z����P���'?9'�N1�DT>@�*'�*%���G�DP��>(5[匏����{}�8  ݳ�Y�k�pJ��U6�Mխn�c�ْ흹�����AYs9*�93�K��9Pe��bd�&y׍�ݣ�rۆ����#�^�U,�īq���۰��I�$�;�+n��2�f��U��Tъ����9q���h����P=���'P �8Q&f�p�b��'3$$�:h��s2L H���E�=N�'es2BK��h��c�Ј�H�D� XY'[䄜̐� ��Z��ϻ��PN�����~��(��;�[�d�[��ڧ	G6f���e�9�޽��mU��߿~�eNI���"s;4�
Z i�l�p�(v�Ф(P�A-���>�$$�ݐ�u�Ϯ�M��}�I�D�o�t}�:�u�l"�q?�@�� ���������tb���u���f:�9�0�c�
^�-�ڶ���ݶX4���1a5��� އ��'�.�"-�5^55�31���N��Ќ���9�:��=qV�b�AD=
�q��I��d�������U��5�^�]��J(���ۮ���w��y���Ԃ%���X3=��ݡ��nڇCDH��5l�������ǽ�Wj����q��9�:�Ug�(U Gf`|CC3w���ݸA�mD"����V�]���"����ُ��N{�L�{BD�ػ��.��[٪�d�$	E��b���<݃���[���ִ#.Da��1��׼�0 f�d��'�wo�T< ��^��</�qڊ$����l�
�(����s���ein�5�m�Ìz������x�P(�fc��u�b�5+���Z�X��m�$� :�ӲN]u؛^��J��",�[d�kj	4mj!�iri��[2�+��\�pdZK�C��l�3� ���ŉ��1ўRX��=1�,��M�i��%j�=�s�st����\e3Ak�[]-HF\����9Ğ��p�Tnǽ�S�Y������o3��.7^��8k3��� ��`2���Z�ѼU���0�l�FUU��o��1Yi��2�SC3e ��Y��h�#qF��lN�zwn�A�ť�)Z :'�k
<5��@p{ν��Ϛ������Ü��������7��㭞�B#Y��{α���G�Å���fd��Xk����a��*٬�b��k}7��SG��6��A�U,r٥R�6$`Ƅ�H�5�,ַ�/v������"0�f< b��~#^U��Q�}�d1������!�]�c� ��	u�1��IE$>�k3���^��{����ein�5�m��uv�Yݮ��،ѕK
RͲ���Ս4��	!l�P(�]��]�՚�Å��.��
]���{Φg��(N�l�V�ݺ��9b"��ꬁ5�.��i� <�9�c�@�F̶>��]��^#�{Gލ��&LA#�wWgu�L%�.(̑�j��f:��8Ff1�J��QGY��xE�b�߈�s����Z[�޶�$}�ҳg��P(����'y�Y�}T(W=��,š����	�Wv�� �|��R0 ^���$�K8�T����3�p�v�T��P��[���v(�4h���ݮQb3�j�z�Xl���&���Qc7��z��hc86簘�U����j�ԏ�I;�t�!ҳ^�K`1��`+[�B�Yn�m�:�kb�.7Y�:�澄�c�
ᾜ�Dj��( F��31�b�k܁@�F��5�:�L�4�{VLf6�л�\꫈z�~����+�"�QױV�fcf��A/�}��>�W���K��ܰ�r8N��?kz3Q��{ʵ�1=�W{b{|	0�5w���*�� Я����m׺���v{��11hn�2U��T�Y��]�E��bxk3���=o�+�̙�f�G�J�߆�^���u����!BB�*2�
Dӌ�`�ζ]�\�����\5�Vf1���b�4�vɌ�Қv�U
�;aVfn�W�(��:ͪ�C�U]�5����w��9�ps��{���?�h�?UB�*���,����TSV�a���T���笑e�M2�W:�Vg)��̫n���SIk-�ŔKV�Z�i�Cn�*���9�JJi��XD����E������y�S���
P7-)7���-��SKoA���9�O0xS����� r��vt��<�7"<��N���s��<<<�)u����tg��`ݷ�I'X
���X"��A���~
�J��0�y�ٽ�������˩Z����
���9�1�y����#6�l��j��t �]��y��^4�
��
DCWZĜF�6�{h�{x-$�
M���/��Ug
���;TE�㈙�Vg]pջb��UP������f���]�;f�f!%��F��,��,9�=àP;:L���9S�6�r�#�Uf��b'v�L4K�ap���x�Uv�*�2����Q�h�Z���Y��I��ݺ�in���U I��ǽ�Y�23Oa&F��o�0`@��F���b5�f:�UYB�Q��!��(�����?P �^�����+�Y�������J���v.`2:M��w��A\f�c8����av�d�w=�r��[b��g!ۖ�d�i8�5�zvÝTd��S��+xz�m��v��7c�J۠]q��pg�Rk�s�#ޮ��`ftn�F�p��U�}����N��}E.���<5��� �Fb�rJBMffM�ΧY���*���T ^:[������p��x�^1�J��QF<*���!��Y�Ƴ^���\i����^��{����1�ZX������p@\`��ƓD�h�Ί�dl��Jӟ~��:�f*�*虁�1��v���B�U?B�C1W�#��'��2��[#(@��A����[�d*4,�o�fcuB�%�kY�b%!$l�c�v�wa��f`HS&�(H�-���`.�`�G\��Ɲ5��.��:�π ��p�����QNJ�U�Y�b��UQ�~�H�3���z���(Wι���)��G���u��8k�0>1Mp���5j�j�1Ǵ�~���-Q�lcZ<�] ��Q��oZ1� �J�U�Y��9w%owޣ!P��g �:�sf/�z�"1Ĝ$�{�s�c� ����M,ֱ�m)�
��W��:�|@U@����׾1D�2:��8ff�������~���0S�n�;U�ڈb1$l�ʟ�h����x����?}��D{�{H-�$�. FϽ���R�������2��Uf��u�]� �F�]�٫�b��k]�!P��S[b��]���O;y�v��~o���  ����a�.�밨v�Լչ��7\tS��T.�h{cvF˰��åm3��T�hU�^��w�cE��cnnԄl\CC�¦X�ε�h��s�����*K��j�uls-�`�8
U09jBc�1��1�q�\uf��v�f0Қv]>u՚���+0��FG�C��@��c����>��4T[�޶�f:�C�q�&�Q���7�:�Uf��n1NB�RB����P�p��ۅ�
�̘ogϟ7=��f����l@Ă50���!�^�����Z�b2�3Uf���ݱ�v���p��LB?
���>�nW��Ɩ^��m)�wods��Իc|;�m��I��3�����If{\IsX����;J�j�ػ�W���+An��������9�B3��6\F�1�o�~��h( � ��*Ѭ�>aƢ����z��v�� �F���?z����y�??6�O=~Q�!��K�Q�-��k͢��.PR�y���}z�]��@��7��F8��^1��9���� Og<�f6�����WT(�f1��w���FGY��k3�Р*�TwޛDz�����OOu�k|���\�sϧ�]�����30�)e�̚jV�NC$l��D�.#Y�Ʒ�WyT(:�]�g��Z���Cv�fc�P ��	�5+0 ��Mfc|u��Lf2��B� �o��������޳��M@��5�:�C"�_�C�@�TחI'��~�����z;����{ޓP�M�8�(����r�����f���O�	Б���+��`$f�#�bP"$D� �"���3�T��ǃ����4�i4:'9�g��̸�#��-d9�q�-��3��l�[&��v�k�Π�����t�zwۜ�$��#a��m�.u7�|�����  m� -�            S�Y��g��[��BpV��lϳ�We����)=%�����D�[�	{u7\g[��\���a�jr�@M��,�r
ꬁ�����.ڧT��-u���¡�Q���:@�(]*�[v���`R]X# 0��7GF;J�\m�RřE%�m��*U �Pm�<�U ,�az@,��.�sj���SMN��f�P��3u�U�n,h�6�P�s�ձ�:�*�k*��x��v.v�m�3n<�ٌ)��tu��*���Ķ�fѩ;(�Kmg<N��m�i�$��i���֚ݭ��h�ܮ�xB�]�H�ݣ�N�l��L�ک���9��az.ȸ��[����.���X���j�����
��Y+����jx���AĐq�+#p\����H4��5R��	�F���.'�V%^��+��t�+b����m(gv3��8�qt*Ɏs���˺���'��"��ްAbொ�P)]'��Jv���t�_{�Er������vvt�h��ca����r:�}5Yn݌rU�4��\`�=�G�]��w\[�lp!@��Co\��iӸu4&5�j�"s�L�&��]�1���h;-�����I�<��۲�b!bl�u�Hl���Q9M����gc��:�����  C��Ş-�
h�^򭚻�.�<� ;9��K񍤎��ő�m��ސ�����)�&�cz�7he
���4x��E�����Vj�m�Y[H�8R0����8nq	�-�mgy�t-Mĕ���Y�]۩��Ɍ�I��?��;'X��<���(o;�$�5��7�:�Uf�ޭ�l%4.��:���Pfc�#X�ZSR����|9�����0S)$8`Q�a	���p�f:c+��~ͿO|�Խ����o�}��]�ȗ��L%��~�<�Y"fXk�f�j-Î���C`US���Z�$$�J�G#�rýsɘ$
)Wj�j����PW��W;��1��|k[���1�SD7�!BF�1�WGGֈ4���#�]���zq(!��c[�9���8p�5�g|�f6��߇���U��1�b�-�
�z��p����c��k�>��in�5�m��c��@~��!�5ƺaDE�y��������=�<��h.Յv+�]6�^�"F%B��cQ�`w�u��p�n�H$
)Y�����0g2~Hs��"�3ۢjko�(�ޕ�!&�(����Ʒ�Wh`��� &[�c2�/G9�}�ݼ�9�=�Kj��	��}RK�M~Q� ��XK��i�nְ.�SQ�콹n� �f���l�@��
���6�u��n:�B��=�maK��7 ���;n�W��"s
���n8]�+ָ�c��P\G�&'' �.N�1����۞u�b���!N����I���l��{�31�o���+Ku�[����^�a�3o��D�c��G1V�L��Z��Ude�,e��HR�l��ػ�=�>|��%�rV]k��ip�4���j�iX=���ϟ7��CZ�@c�6����<�]f*�K/X�f6�׎f>�WڪC-W5�kJ��I�빎�fc��Y���	@P��z�>$�v	��B3�9�#p%A�$=�/^�d筹���p�a���c�㫵Vk�,7�cQhffH ]��Ff05���(�v�l�����w<٩�7�}#|�P%SCb��S{��똆�V���l�Wv��(pv�^��5uZ�^�@��14�0����!
85� ��Ho����ݪj6
3���uY5���X��)5f-��fc��(Uus����$�����~��\���S">�����v��G�{�$`2*��H�h��1��31��XC9���mxcP����it::�7�P�ݶ�� �9�$0���k3�̕��+����57�.��f?�@US�;�Lq6a���k|u�*�J��Q5Jh]ۮuU��@P9� �+��0��u��qW33���?nw�{9�ϛ+r����3����� +*��k��X
��s5	����0�5�kID�X�C�3ZM�L^k��1�F��fw��-m�g��lu�g�#"�ۅ\n7]�3�$+s:������w�����`4!Ժ�8X\�Xddl���&�m�n���B�����}� ^!;�1�Ǉ���Xk�07�c���uެ�	:�Y���g��b���e�wl]ۭ����Ȓ��Uڬ@o��Y�#����qFC
JIJC$݇.������4F`z�F���:���E�w{ډ��SB�����C�T �*ѭ{��� �^��!I��3���1���g����%ilr���\���f Ƚ=��1��9�:���.>���j�̬Z�m����rpURoA=�-��u����l��H�*�B6j��^��
j��Ȓ��V��:�^���'�w��{����~����׷���KVr*U�E=G�AX�VB0��-�K.Y7T].q�Ƹ2�q�'�$�ٮw}i�t�)I l�1ֲН����A
%%�Af�G��1,a.� �%Y*�jc�é����������}�]��Tgz�.c�1w1�o��fq�( pֳ7�Q��f:�UY�Ï�B���D��M�@vI����.`���Md)5{ʷ�Y����V���^��ϘQ���_�Ǽ�����!��S#Wv�w�����u�ǴLj-��
�����}���~-�}�Ej�*ZUB# C�D�^�`Bz�і\�ec��|xk3y�*Y�0(Y���MB�@F�^u$���6Q��$�YkoF��^�c{��̑&5��k|u�UY���Q�Jh]���&����-"8#Ԅf!�f31���2�������������6*�����ώ��y�~��}:_�  цq�%�f��{����tIa<��[�zͳ�����[g���1��Z�����n�Л{eu���ДNj5�%'&���,�<6gc,`g�T�N䶝�ν�!1ĸv"֓��JY���t�F8�UWs�2~߷�=:���Mq���&5�9���	�`fc��3�Vg��n��\�vܑ(���<F��=�:���6�2D�5�3��e��V�mq�7�@�-©�@����F�*#2[���:��_mԵ�-Aj:�_��
����� lY��c��W��������o�P��y�b��q���fc�]��\���2(�.��z��\��s�p��e�i(�4
�R3���Z�Tr���+��f��(U
����!�Z�!L�����
#|���{�k�2D���]�����v�
(�z��@�I(�=�u:���UG3�xZ�"�u��;5wl]���
;��h��}ѩ���u�!�/5�%��+Ku�[���ﾕ��#7��`�f1����hq���&E�ݺ�Vqa�DfiЗ�CEA���ᡙ��{����9F�[�޻w�w[��W%VhYZ�໷R�p�{.!%Tl�]<\�g]���ꁄ�c[㫴,��v�E��
h]ۮu ]��sx�j�Qֱ����{����o�~��M�����9���E�q�0�y�J�A���*��zE|��` ]۪c�:���5��n���pw^��	<���=�7Y�j��D�3h[�i�:0���{��On9��C�^hy�:�M�MJ�Ҫׁ�qT���:�~��$���Qu'�ګ�+���Go%�jSl�ɍEc�?:�P��wlp��b8c*'_�OH��9�����!L�d	��wn�З��d�4a��c{㫴0᧚�0'Jhf,5Ϊ�WvŊ�ӷm�rvJ�^ga��pU���$JB����[#f1��#��=q���[��c����e����"�1���;κ�U�a�/��Z���\�"�`j�b8`1J�U�Wv�ݺ�l�}s��ӵp�d�ʚ�##nHQpE!L�5Vjkl]��D��3$I�@��5�:�dJ�l��I,�'9�<�u�1D��"�A:�T�0�FF���������P�f:����1������[���f!���R�5nu��=�����=l$bG �7")�`�,s|uv��8�e��B��w�Y32CY��$0�f.�3#v�Z�R�-� k[L]���  )��s�q�"N=�5�:�*�h|D��bD$�0
P��h���.�����J�.m�����u΄6sj���Zݖ�)&䫵[5wl]۫��e��mi���o�{�u��#7��`�j��y�Y��N��`��&5�r�Uڬ#�3��ۍ~�o|�{�����3���y*y�m�%��6R��#j6v�a��� � �@����T��*��I���%�I[Z�r�m|6	js������  �[@            �$r%��_������jͣMi��)tIi��f��
�M�V�.�v�v�y���ۊ�m����6�����{r$i�F�{4�Ld:��eCn��,l���mAq�m�yU!���3�G!v`�D��펔!�86*;-Xf�gXk�X�b��5��D�Ƭ�6�m3�Hƅ&E��,0��=*�ԭJ�9��O����9�ڽ.�JG]�VE��cZՊE�;�ٺ���%�<���].w���J;���EU�����(�n.��P���m;r�N�C)2�{9�֌�s�]�lF�����εqg��@+t�l"�3n��K�-��R]�6�g*�%�;CP�nb��,�n�;`�!���U0b�]r4�u����k�y�;�@6�%����V�
��$$8�H�ͻa��b��m��S����f�S\1ڊ��ɡU`v��u�����]0�u�V[Q�d�ʨ��j�B.�S�H hA<�=-��B�j��.Ȟ�����fd��  �Mt�n�6&��\ŌlTuc��t�X���4 ��8�$CͲ2.C
q��b��f,���c�l�
����oo����y���}��%-m�.�b�RX�eM;4��!��d��ei��0ٙ\�߮oz%�l��E��|�f��c��f���R���55�.����@�9�Z�$�4s2o�t  Y��Ғ��\i)�{λj���%��jB�Q�����^�����꽰}w?{�JP�K��<� ����P6���|kZ�}󫰃"���a��]���U@U� �ݦ����� �|<���š�c��!�wl�ْPx�����f:֮�T�1в�ػ�Wh1Z��,0��gK�i:�o�٣Ga��v���hYC��q���^:�P�ݱ�5��!A5��C��ؠ�@a�~w��~�n�Z_p|@��X���1E�q�0�.:�|'�d���p���Ż�m8A�cJ�ˊm3��f�}��s׻0�wl�ْR���@U�=�1�yֵ�t�"�� M틻uv����!��>�	�rμ��Cת=�8*$\<���=���QJhz��:�����l�Lٴ����e�[q�حG�&�
�$���1�g�`��Y��}�4��{5��
Bs��������!��I�d5��&��F *���-�p�Z���X��`_v�E*���]��̕���0��I$�I$�UUy��Ɣ�p1��7:��eؽgjt�TEx��/-�
.����i�]2se/4���E7&�f����ڀ��ѭ�69�ˠ\�Σ[.����B�)�9��I'9;�#a�$��(�dGRM4�4e�� QN�Holfc��5||b8�p���5�:��@�T�Ӹ�������uΞ�dv�7�*8�j:����1�����쁦���olfc����;m��ۮ��c.A/p�.\9$���&	�j�o���Ő-�p�ѓB�����������8Fo�q��V���]�wn���J��Z@Z�vło�gv�r4�Wlk|䫻�$���ʹml��*M�r�7(̐419rH�24���̕۶0����(؉���8ivŋ�W���Li������`�UT@UyiF�3lB3���	�k1����̶& 2k�0��]ۮ��YCVġΛ�&m�2�����U%����E��q7f(�Uݱ��b���-��* Qj������W}cu[6_r8�F�vƷ�W}aZox�25.�ts���<���z}��hPֺ�Vjkׂ�$���8@Wl]�u�@�g�� x���3n7�׮
�o4��_��m��?|�|�}��� G�}pl����bHg^�v�����3{�}dƌ�̷]�]���W�Y��s��H1��u5w�2���ŋ�W}};��*��:F��C[O�I$�  4��S^Kt�%��<u�:�ҷ n�-�Ԕ��1��(im��T�U�(����F�S���D����z��{V�g�,1	�p�Ʌ�rC���6��5^��TU�^�����]utZ�;�3��m(0R���P�5&��z�N;�1����w@�M㈸�e�p�^J��`��=�
C����;��c3f�s����������>2����[��������a�0��d�$�#q���7��sT�t��TQ�f*�8��]^�n)Wv�+�  P�	d�cY���+|̆2d
-��ǳ2s-��{R2� ^�s���Őu�qE��u�� [�\:��,�U!�1�l� �V�FHK��JB�Q��XΠc��5���e�����X��W}b|�E�L]�9�1��s�֤�g9��9�s���9�c��ޛXN-���d�����m��Bs,�m7vw�����%�3�7�p�4['5��&8s��J�Y��iD"�J��X#6�$�8������5�4i���<�sV��A3�c�hF�J/�l�i5e�ֶ�Y�HDVPq�
t�6��QiR�W��Z�-��56�I�E�¨U?}��Y��<@~�W�y	����c�v�ݿ�����tYi��fK���;���Q���V�}$�y�߿w����)b�cþu�e���;��1�\e)��{һv�Ɩcһ�c��s-��y�{ݞ�t�a��3;��~��2�zOu�K[c3]��l
�Ϣ�,�N��\��Ӆ�v�0� n4�Ɉ���fu՚�cOh�ʏB��g��uf�ަUty���&�V�'�p�����J�^[� Qj����6�1�ݱ��c�Fن��ƷǄf[�5�,h4I��C��  5דZ�jΖ�E�+���0B≰3�a�f�X�[ʨX76`n^�"ݪf�������c��&����+�o&� 6��뛳)�Q����mua�q[��Ns��{��G���Q�ݻufv�{���u,�g+��]w�u�l��5j�L�4�uwo�t��c3f��}M3��<|i���fu�E�Ɉ���1w�Ԭ�b"���Oh�ҏB��w�b�
�Mݹ#I�ӭļ��Ղ����nۆ%q��1J�����p-�ʚ�t�Lx]V���; �{Q4���,�9o3�h_9�5�q��v@w�[��ʏ^=�u۷��ŝCGY��
틻~#�P�<����(��쩖�����5��ſ��ZM='�����?~���lh��b-�LY�s|uw܃+X6������]�_���t����z�W�4���FV�s�쎚nػ�SW}1� QhY���.�9��0��B[P�%7�81���р�̺�U���k�uw�,�!�QQ�]��n�a/1�b�&	IGY��
틻u{��q���Oc{c3�T(� �Un� %ޘ�wl��h���]���&~^��Ws5�`�]�hH����	""�&4f�ݿwla������1A�3��F31���Ld��B�[P�d�VƆ�#Q���w޺̶0��Y�!q��ݺ�z��
�UB��n���I*���0Ȗ4�v��,�t����`�Q�8iT.��6A&!f",U	��۱7g���W=)F#��k��]a�ML�XL�h����%5G.�#.�4�%����^\#b������&�$˼�ـ�T��2�0�уs�n��feހ�I�����2�-���0���31��X�_9L ���]��5����Lh��h����2nnV��b�19Z�c�Z@<�31��<�a� �^���5�m��[:�3I�2��[cٙ+2����VT̺ʨ뜿�к($A�`%(� @�	���=C^�����}�p�\M8�=�:�n�x��bb�	J<#3t��c3^�s�l='��K{,fc�����d>�YfBb0 a����xj�*0�����s|u����[���L�wo��Xig5�����&V;�v��V
�A�E˽ٽ�nl�~^\��ej���ػ�,���ھE���5��3���u��7�i��L�P(Cq'D9.h��򎍭r�T3�Y�gϖ�	�]Y�;lKW`�#)GWv놕�vv��ޣ-��^�-m�f:���E��Q�� y�w�u�׆�����E�lq��C3w�cy�v��}ٵ��)F�,*�m�P � ��0A)Y�놱�x 4=�:�s��2��*��c3fu��;QF�#���o�u��="-ڌ��SB��s�uf����0H�i��31���#����տ�?��I!	�$�$ ��*� �����h� ~ϰ�RW��u�����\�חp$�DTlƬ��caM�7��j��!"*(�@R��jj����.���^<9�RQaKKk
��\2�U&��*������hZ����4I*��Jɭ[Y��f��4i��y�sc7U��[[@�[B�-&�@��t��qAL�+C ���ͥ�mM�YF�@�[ln�fr��m���ڶ���7���\��U�9��X�6q��b��2�`�R�Q�b6_�Ҟ������� ���Y~�ο|��� PO�������)p��(%���(=�������&3�� ���?�쎣��k�Ge9�@����T@���~������D �$<�T@�
F����~���?H�4��\�qT�������>��~$#� ğ֢� o�G�>�o���:B�F�>�����񸄌d~�t�
�����u����*"}g��}T2uG�ԒB����,�gB"��
�RA$E6Ɖ��mL�6�2�m��e6̦6�`I�چmM�ձ�)���V�*YY��Ʀ6�c����m���ʵj���b����m�j���lj�6�m�l
2��(�VV͵m�4�X+l��f�6�[2�
���6��1�b�eb���fVڨH�Y��U�0�mLe�
ٕ�k�9�ɶ�+
қM�Ֆb�ԣ,Ĭ!+5�����g~�O��fg�q�/�����I��������j����}��>���������σ۰�=�����?��A�������1ED ��I�Ak��C�:���ܸO�/���������X{'�q���r|��������������HH6�7��a'��G���槏���,~c�?+~nͳ���߿�>sA��?}U'�ћP����=��@ ��c�p�?��A@
HBӯ���S��A&������ʎ��<ޠ}���v����gB* Q�����}B* ��g��~_s�PS�o������W���Ū�����}��� ~����������~`O������#>z?�����'�g�����> >�}à>:4�?{��A���X�z��l7�����9�m�O3�>#�q��E'�؁S������?O�yA(���F���:��_��{"$Q ?���p��@O�Q������T@���[����S�_�����i�'Ї��3|�}���rE8P���q�